magic
tech sky130A
magscale 1 2
timestamp 1607327525
<< checkpaint >>
rect -3932 -3932 43584 45728
<< locali >>
rect 28917 28951 28951 29257
rect 29285 28407 29319 28577
rect 31953 23103 31987 23273
rect 5089 21879 5123 22049
rect 5181 21879 5215 21981
rect 5825 20247 5859 20417
rect 17233 19159 17267 19261
rect 17325 19227 17359 19329
rect 17601 19159 17635 19465
rect 29377 18615 29411 18853
rect 8493 18139 8527 18241
rect 17601 18071 17635 18173
rect 14289 16983 14323 17085
rect 15669 16983 15703 17085
rect 11345 15895 11379 15997
rect 11621 14807 11655 14909
rect 12081 14807 12115 14977
rect 13277 13787 13311 13957
rect 23397 13379 23431 13481
rect 23397 13175 23431 13345
rect 18429 12223 18463 12393
rect 19533 12291 19567 12393
rect 24777 12291 24811 12393
rect 17233 9367 17267 9469
<< viali >>
rect 3801 39049 3835 39083
rect 8769 39049 8803 39083
rect 9597 39049 9631 39083
rect 11437 39049 11471 39083
rect 26617 39049 26651 39083
rect 6653 38981 6687 39015
rect 12817 38981 12851 39015
rect 4353 38913 4387 38947
rect 7481 38913 7515 38947
rect 10149 38913 10183 38947
rect 13553 38913 13587 38947
rect 15301 38913 15335 38947
rect 15761 38913 15795 38947
rect 4077 38845 4111 38879
rect 6285 38845 6319 38879
rect 7205 38845 7239 38879
rect 9873 38845 9907 38879
rect 13461 38845 13495 38879
rect 14289 38845 14323 38879
rect 14381 38845 14415 38879
rect 15485 38845 15519 38879
rect 27077 38845 27111 38879
rect 27353 38845 27387 38879
rect 5733 38777 5767 38811
rect 28733 38777 28767 38811
rect 3433 38709 3467 38743
rect 13277 38709 13311 38743
rect 17049 38709 17083 38743
rect 26249 38709 26283 38743
rect 13645 38505 13679 38539
rect 3157 38437 3191 38471
rect 5733 38369 5767 38403
rect 13369 38369 13403 38403
rect 17509 38369 17543 38403
rect 23213 38369 23247 38403
rect 26801 38369 26835 38403
rect 29837 38369 29871 38403
rect 32413 38369 32447 38403
rect 1501 38301 1535 38335
rect 1777 38301 1811 38335
rect 5457 38301 5491 38335
rect 7113 38301 7147 38335
rect 11713 38301 11747 38335
rect 11989 38301 12023 38335
rect 17233 38301 17267 38335
rect 22937 38301 22971 38335
rect 26525 38301 26559 38335
rect 29561 38301 29595 38335
rect 32137 38301 32171 38335
rect 7389 38165 7423 38199
rect 9873 38165 9907 38199
rect 15485 38165 15519 38199
rect 18613 38165 18647 38199
rect 19441 38165 19475 38199
rect 24317 38165 24351 38199
rect 27905 38165 27939 38199
rect 30941 38165 30975 38199
rect 33517 38165 33551 38199
rect 1961 37961 1995 37995
rect 5549 37961 5583 37995
rect 7205 37961 7239 37995
rect 11897 37961 11931 37995
rect 23029 37961 23063 37995
rect 27629 37961 27663 37995
rect 29561 37961 29595 37995
rect 30021 37961 30055 37995
rect 31401 37961 31435 37995
rect 32045 37961 32079 37995
rect 5825 37825 5859 37859
rect 7665 37825 7699 37859
rect 11161 37825 11195 37859
rect 19257 37825 19291 37859
rect 19625 37825 19659 37859
rect 26157 37825 26191 37859
rect 26525 37825 26559 37859
rect 32413 37825 32447 37859
rect 35725 37825 35759 37859
rect 36093 37825 36127 37859
rect 7389 37757 7423 37791
rect 10793 37757 10827 37791
rect 17325 37757 17359 37791
rect 19349 37757 19383 37791
rect 26249 37757 26283 37791
rect 32321 37757 32355 37791
rect 33149 37757 33183 37791
rect 33241 37757 33275 37791
rect 35817 37757 35851 37791
rect 9045 37689 9079 37723
rect 10609 37689 10643 37723
rect 1685 37621 1719 37655
rect 10425 37621 10459 37655
rect 11437 37621 11471 37655
rect 12173 37621 12207 37655
rect 17693 37621 17727 37655
rect 20729 37621 20763 37655
rect 23397 37621 23431 37655
rect 25697 37621 25731 37655
rect 31769 37621 31803 37655
rect 37197 37621 37231 37655
rect 26801 37417 26835 37451
rect 35173 37417 35207 37451
rect 32781 37349 32815 37383
rect 5641 37281 5675 37315
rect 5917 37281 5951 37315
rect 9689 37281 9723 37315
rect 9965 37281 9999 37315
rect 12449 37281 12483 37315
rect 15577 37281 15611 37315
rect 16957 37281 16991 37315
rect 18613 37281 18647 37315
rect 26249 37281 26283 37315
rect 32413 37281 32447 37315
rect 34069 37281 34103 37315
rect 35817 37281 35851 37315
rect 12173 37213 12207 37247
rect 15301 37213 15335 37247
rect 18337 37213 18371 37247
rect 33793 37213 33827 37247
rect 7021 37077 7055 37111
rect 11253 37077 11287 37111
rect 13553 37077 13587 37111
rect 19717 37077 19751 37111
rect 1685 36873 1719 36907
rect 2329 36873 2363 36907
rect 5733 36873 5767 36907
rect 9781 36873 9815 36907
rect 10057 36873 10091 36907
rect 12173 36873 12207 36907
rect 12633 36873 12667 36907
rect 15393 36873 15427 36907
rect 18429 36873 18463 36907
rect 26893 36873 26927 36907
rect 33885 36873 33919 36907
rect 34253 36873 34287 36907
rect 35173 36873 35207 36907
rect 6009 36737 6043 36771
rect 19073 36737 19107 36771
rect 19441 36737 19475 36771
rect 25145 36737 25179 36771
rect 25605 36737 25639 36771
rect 35817 36737 35851 36771
rect 1409 36669 1443 36703
rect 1593 36669 1627 36703
rect 19165 36669 19199 36703
rect 25329 36669 25363 36703
rect 35725 36669 35759 36703
rect 36415 36669 36449 36703
rect 36553 36669 36587 36703
rect 20821 36601 20855 36635
rect 15761 36533 15795 36567
rect 35449 36533 35483 36567
rect 10425 36329 10459 36363
rect 5181 36193 5215 36227
rect 10609 36193 10643 36227
rect 16405 36193 16439 36227
rect 4905 36125 4939 36159
rect 16681 36125 16715 36159
rect 18061 36125 18095 36159
rect 1685 35989 1719 36023
rect 6469 35989 6503 36023
rect 18337 35989 18371 36023
rect 19165 35989 19199 36023
rect 25329 35989 25363 36023
rect 35633 35989 35667 36023
rect 4997 35785 5031 35819
rect 5365 35785 5399 35819
rect 10517 35785 10551 35819
rect 24961 35785 24995 35819
rect 25421 35649 25455 35683
rect 35725 35649 35759 35683
rect 36093 35649 36127 35683
rect 18061 35581 18095 35615
rect 18337 35581 18371 35615
rect 25145 35581 25179 35615
rect 35817 35581 35851 35615
rect 17785 35513 17819 35547
rect 19717 35513 19751 35547
rect 26801 35513 26835 35547
rect 16405 35445 16439 35479
rect 16865 35445 16899 35479
rect 37197 35445 37231 35479
rect 11713 35241 11747 35275
rect 29377 35241 29411 35275
rect 7297 35105 7331 35139
rect 11897 35105 11931 35139
rect 14197 35105 14231 35139
rect 7021 35037 7055 35071
rect 8585 34901 8619 34935
rect 14013 34901 14047 34935
rect 14749 34901 14783 34935
rect 18153 34901 18187 34935
rect 24041 34901 24075 34935
rect 25145 34901 25179 34935
rect 35909 34901 35943 34935
rect 7021 34697 7055 34731
rect 7389 34697 7423 34731
rect 11805 34697 11839 34731
rect 14013 34697 14047 34731
rect 25881 34697 25915 34731
rect 37381 34697 37415 34731
rect 30665 34629 30699 34663
rect 14749 34561 14783 34595
rect 19717 34561 19751 34595
rect 20085 34561 20119 34595
rect 21189 34561 21223 34595
rect 26341 34561 26375 34595
rect 26709 34561 26743 34595
rect 29101 34561 29135 34595
rect 29561 34561 29595 34595
rect 35725 34561 35759 34595
rect 36093 34561 36127 34595
rect 15025 34493 15059 34527
rect 19809 34493 19843 34527
rect 24593 34493 24627 34527
rect 26433 34493 26467 34527
rect 29285 34493 29319 34527
rect 35817 34493 35851 34527
rect 14565 34425 14599 34459
rect 16129 34357 16163 34391
rect 24409 34357 24443 34391
rect 27813 34357 27847 34391
rect 15117 34153 15151 34187
rect 15761 34153 15795 34187
rect 27261 34153 27295 34187
rect 27813 34153 27847 34187
rect 9965 34017 9999 34051
rect 16129 34017 16163 34051
rect 16497 34017 16531 34051
rect 16681 34017 16715 34051
rect 17969 34017 18003 34051
rect 21925 34017 21959 34051
rect 22477 34017 22511 34051
rect 23489 34017 23523 34051
rect 24317 34017 24351 34051
rect 24501 34017 24535 34051
rect 27445 34017 27479 34051
rect 30021 34017 30055 34051
rect 30297 34017 30331 34051
rect 9689 33949 9723 33983
rect 15945 33949 15979 33983
rect 17693 33949 17727 33983
rect 19809 33949 19843 33983
rect 21741 33949 21775 33983
rect 24041 33949 24075 33983
rect 29653 33949 29687 33983
rect 30389 33949 30423 33983
rect 22385 33881 22419 33915
rect 11253 33813 11287 33847
rect 16957 33813 16991 33847
rect 19073 33813 19107 33847
rect 20361 33813 20395 33847
rect 25421 33813 25455 33847
rect 28089 33813 28123 33847
rect 29377 33813 29411 33847
rect 35909 33813 35943 33847
rect 9781 33609 9815 33643
rect 10057 33609 10091 33643
rect 14473 33609 14507 33643
rect 16221 33609 16255 33643
rect 17785 33609 17819 33643
rect 22201 33609 22235 33643
rect 24317 33609 24351 33643
rect 26709 33609 26743 33643
rect 22477 33541 22511 33575
rect 16681 33473 16715 33507
rect 20269 33473 20303 33507
rect 20453 33473 20487 33507
rect 20545 33473 20579 33507
rect 25513 33473 25547 33507
rect 27445 33473 27479 33507
rect 14841 33405 14875 33439
rect 16589 33405 16623 33439
rect 16957 33405 16991 33439
rect 17141 33405 17175 33439
rect 21281 33405 21315 33439
rect 21373 33405 21407 33439
rect 25421 33405 25455 33439
rect 26249 33405 26283 33439
rect 26341 33405 26375 33439
rect 27353 33405 27387 33439
rect 28181 33405 28215 33439
rect 28273 33405 28307 33439
rect 29929 33405 29963 33439
rect 30297 33405 30331 33439
rect 23857 33337 23891 33371
rect 24869 33337 24903 33371
rect 29101 33337 29135 33371
rect 30021 33337 30055 33371
rect 15209 33269 15243 33303
rect 15577 33269 15611 33303
rect 18245 33269 18279 33303
rect 19073 33269 19107 33303
rect 21833 33269 21867 33303
rect 23489 33269 23523 33303
rect 25237 33269 25271 33303
rect 27169 33269 27203 33303
rect 28641 33269 28675 33303
rect 10885 33065 10919 33099
rect 15117 33065 15151 33099
rect 17141 33065 17175 33099
rect 20453 33065 20487 33099
rect 24961 33065 24995 33099
rect 28273 33065 28307 33099
rect 29929 33065 29963 33099
rect 15577 32997 15611 33031
rect 19993 32997 20027 33031
rect 29561 32997 29595 33031
rect 30205 32997 30239 33031
rect 6285 32929 6319 32963
rect 11069 32929 11103 32963
rect 16037 32929 16071 32963
rect 24961 32929 24995 32963
rect 25421 32929 25455 32963
rect 26525 32929 26559 32963
rect 26985 32929 27019 32963
rect 27353 32929 27387 32963
rect 28365 32929 28399 32963
rect 28917 32929 28951 32963
rect 30113 32929 30147 32963
rect 31033 32929 31067 32963
rect 6009 32861 6043 32895
rect 12633 32861 12667 32895
rect 12909 32861 12943 32895
rect 15761 32861 15795 32895
rect 18337 32861 18371 32895
rect 18613 32861 18647 32895
rect 21649 32861 21683 32895
rect 21925 32861 21959 32895
rect 27445 32861 27479 32895
rect 28825 32861 28859 32895
rect 30757 32861 30791 32895
rect 31217 32861 31251 32895
rect 7573 32725 7607 32759
rect 14013 32725 14047 32759
rect 23213 32725 23247 32759
rect 27813 32725 27847 32759
rect 6009 32521 6043 32555
rect 6377 32521 6411 32555
rect 12265 32521 12299 32555
rect 16681 32521 16715 32555
rect 18245 32521 18279 32555
rect 18981 32521 19015 32555
rect 21741 32521 21775 32555
rect 25329 32521 25363 32555
rect 25881 32521 25915 32555
rect 28641 32521 28675 32555
rect 29653 32521 29687 32555
rect 30021 32521 30055 32555
rect 31585 32521 31619 32555
rect 15669 32453 15703 32487
rect 17785 32453 17819 32487
rect 27629 32453 27663 32487
rect 29009 32453 29043 32487
rect 13553 32385 13587 32419
rect 19349 32385 19383 32419
rect 23765 32385 23799 32419
rect 14013 32317 14047 32351
rect 14197 32317 14231 32351
rect 14381 32317 14415 32351
rect 14933 32317 14967 32351
rect 15853 32317 15887 32351
rect 16037 32317 16071 32351
rect 16221 32317 16255 32351
rect 18061 32317 18095 32351
rect 19073 32317 19107 32351
rect 23489 32317 23523 32351
rect 24409 32317 24443 32351
rect 26249 32317 26283 32351
rect 27813 32317 27847 32351
rect 28181 32317 28215 32351
rect 28273 32317 28307 32351
rect 30297 32317 30331 32351
rect 15209 32249 15243 32283
rect 18521 32249 18555 32283
rect 26617 32249 26651 32283
rect 27261 32249 27295 32283
rect 30941 32249 30975 32283
rect 10977 32181 11011 32215
rect 12725 32181 12759 32215
rect 13001 32181 13035 32215
rect 13369 32181 13403 32215
rect 20453 32181 20487 32215
rect 22017 32181 22051 32215
rect 24961 32181 24995 32215
rect 31309 32181 31343 32215
rect 13645 31977 13679 32011
rect 16129 31977 16163 32011
rect 18613 31977 18647 32011
rect 19165 31977 19199 32011
rect 19625 31977 19659 32011
rect 26341 31977 26375 32011
rect 28089 31977 28123 32011
rect 30297 31977 30331 32011
rect 14381 31909 14415 31943
rect 15761 31909 15795 31943
rect 16589 31909 16623 31943
rect 24409 31909 24443 31943
rect 26893 31909 26927 31943
rect 27261 31909 27295 31943
rect 13921 31841 13955 31875
rect 17049 31841 17083 31875
rect 17233 31841 17267 31875
rect 17417 31841 17451 31875
rect 18429 31841 18463 31875
rect 19441 31841 19475 31875
rect 24685 31841 24719 31875
rect 25421 31841 25455 31875
rect 25513 31841 25547 31875
rect 26709 31841 26743 31875
rect 26801 31841 26835 31875
rect 27905 31841 27939 31875
rect 28273 31841 28307 31875
rect 28825 31841 28859 31875
rect 29009 31841 29043 31875
rect 29193 31841 29227 31875
rect 29837 31841 29871 31875
rect 30573 31841 30607 31875
rect 13829 31773 13863 31807
rect 19993 31773 20027 31807
rect 24593 31773 24627 31807
rect 26525 31773 26559 31807
rect 28365 31773 28399 31807
rect 3249 31637 3283 31671
rect 12909 31637 12943 31671
rect 23673 31637 23707 31671
rect 25881 31637 25915 31671
rect 27537 31637 27571 31671
rect 30941 31637 30975 31671
rect 10885 31433 10919 31467
rect 16129 31433 16163 31467
rect 16865 31433 16899 31467
rect 23121 31433 23155 31467
rect 28641 31433 28675 31467
rect 30665 31433 30699 31467
rect 35633 31433 35667 31467
rect 3065 31365 3099 31399
rect 16405 31365 16439 31399
rect 18245 31365 18279 31399
rect 3157 31297 3191 31331
rect 3893 31297 3927 31331
rect 4077 31297 4111 31331
rect 12909 31297 12943 31331
rect 15761 31297 15795 31331
rect 19901 31297 19935 31331
rect 23857 31297 23891 31331
rect 25513 31297 25547 31331
rect 25605 31297 25639 31331
rect 27905 31297 27939 31331
rect 30021 31297 30055 31331
rect 30941 31297 30975 31331
rect 32137 31297 32171 31331
rect 36093 31297 36127 31331
rect 3801 31229 3835 31263
rect 4169 31229 4203 31263
rect 10517 31229 10551 31263
rect 13185 31229 13219 31263
rect 16589 31229 16623 31263
rect 16681 31229 16715 31263
rect 18061 31229 18095 31263
rect 18889 31229 18923 31263
rect 19257 31229 19291 31263
rect 19625 31229 19659 31263
rect 23765 31229 23799 31263
rect 24593 31229 24627 31263
rect 24685 31229 24719 31263
rect 25789 31229 25823 31263
rect 26341 31229 26375 31263
rect 29561 31229 29595 31263
rect 29745 31229 29779 31263
rect 31677 31229 31711 31263
rect 31953 31229 31987 31263
rect 35817 31229 35851 31263
rect 14565 31161 14599 31195
rect 17417 31161 17451 31195
rect 25973 31161 26007 31195
rect 27169 31161 27203 31195
rect 27537 31161 27571 31195
rect 29101 31161 29135 31195
rect 31125 31161 31159 31195
rect 2697 31093 2731 31127
rect 10333 31093 10367 31127
rect 12817 31093 12851 31127
rect 18613 31093 18647 31127
rect 19073 31093 19107 31127
rect 21005 31093 21039 31127
rect 23489 31093 23523 31127
rect 25053 31093 25087 31127
rect 25881 31093 25915 31127
rect 26617 31093 26651 31127
rect 26985 31093 27019 31127
rect 27353 31093 27387 31127
rect 27445 31093 27479 31127
rect 28181 31093 28215 31127
rect 37381 31093 37415 31127
rect 3249 30889 3283 30923
rect 13921 30889 13955 30923
rect 14289 30889 14323 30923
rect 16681 30889 16715 30923
rect 17233 30889 17267 30923
rect 19441 30889 19475 30923
rect 19901 30889 19935 30923
rect 23765 30889 23799 30923
rect 24593 30889 24627 30923
rect 26341 30889 26375 30923
rect 28733 30889 28767 30923
rect 29745 30889 29779 30923
rect 35909 30889 35943 30923
rect 13093 30821 13127 30855
rect 25237 30821 25271 30855
rect 27353 30821 27387 30855
rect 27445 30821 27479 30855
rect 28457 30821 28491 30855
rect 11989 30753 12023 30787
rect 13185 30753 13219 30787
rect 18521 30753 18555 30787
rect 18705 30753 18739 30787
rect 18889 30753 18923 30787
rect 20269 30753 20303 30787
rect 21373 30753 21407 30787
rect 23029 30753 23063 30787
rect 25053 30753 25087 30787
rect 25145 30753 25179 30787
rect 27261 30753 27295 30787
rect 30021 30753 30055 30787
rect 30757 30753 30791 30787
rect 31217 30753 31251 30787
rect 31493 30753 31527 30787
rect 12081 30685 12115 30719
rect 15301 30685 15335 30719
rect 15577 30685 15611 30719
rect 21649 30685 21683 30719
rect 24869 30685 24903 30719
rect 25605 30685 25639 30719
rect 27077 30685 27111 30719
rect 27813 30685 27847 30719
rect 18337 30617 18371 30651
rect 6929 30549 6963 30583
rect 10425 30549 10459 30583
rect 12541 30549 12575 30583
rect 12909 30549 12943 30583
rect 13369 30549 13403 30583
rect 24133 30549 24167 30583
rect 25973 30549 26007 30583
rect 26709 30549 26743 30583
rect 29285 30549 29319 30583
rect 14013 30345 14047 30379
rect 14565 30345 14599 30379
rect 16037 30345 16071 30379
rect 17785 30345 17819 30379
rect 18337 30345 18371 30379
rect 21373 30345 21407 30379
rect 28273 30345 28307 30379
rect 31769 30345 31803 30379
rect 4537 30277 4571 30311
rect 9229 30277 9263 30311
rect 10425 30277 10459 30311
rect 11897 30277 11931 30311
rect 12541 30277 12575 30311
rect 13921 30277 13955 30311
rect 26801 30277 26835 30311
rect 28825 30277 28859 30311
rect 35725 30277 35759 30311
rect 3065 30209 3099 30243
rect 7849 30209 7883 30243
rect 10241 30209 10275 30243
rect 13461 30209 13495 30243
rect 15301 30209 15335 30243
rect 18061 30209 18095 30243
rect 18889 30209 18923 30243
rect 19441 30209 19475 30243
rect 21097 30209 21131 30243
rect 24593 30209 24627 30243
rect 24961 30209 24995 30243
rect 25973 30209 26007 30243
rect 26985 30209 27019 30243
rect 28641 30209 28675 30243
rect 29377 30209 29411 30243
rect 30297 30209 30331 30243
rect 32321 30209 32355 30243
rect 36093 30209 36127 30243
rect 2697 30141 2731 30175
rect 3157 30141 3191 30175
rect 3433 30141 3467 30175
rect 7389 30141 7423 30175
rect 7665 30141 7699 30175
rect 8861 30141 8895 30175
rect 10425 30141 10459 30175
rect 10977 30141 11011 30175
rect 11069 30141 11103 30175
rect 12449 30141 12483 30175
rect 12725 30141 12759 30175
rect 14197 30141 14231 30175
rect 14749 30141 14783 30175
rect 14841 30141 14875 30175
rect 18153 30141 18187 30175
rect 19717 30141 19751 30175
rect 21925 30141 21959 30175
rect 22293 30141 22327 30175
rect 22569 30141 22603 30175
rect 25513 30141 25547 30175
rect 25881 30141 25915 30175
rect 27813 30141 27847 30175
rect 27951 30141 27985 30175
rect 29009 30141 29043 30175
rect 30205 30141 30239 30175
rect 32137 30141 32171 30175
rect 32781 30141 32815 30175
rect 33057 30141 33091 30175
rect 35817 30141 35851 30175
rect 6837 30073 6871 30107
rect 9873 30073 9907 30107
rect 13185 30073 13219 30107
rect 15577 30073 15611 30107
rect 25053 30073 25087 30107
rect 27077 30073 27111 30107
rect 29469 30073 29503 30107
rect 31033 30073 31067 30107
rect 33333 30073 33367 30107
rect 6653 30005 6687 30039
rect 8677 30005 8711 30039
rect 12173 30005 12207 30039
rect 17509 30005 17543 30039
rect 19349 30005 19383 30039
rect 22293 30005 22327 30039
rect 23489 30005 23523 30039
rect 24133 30005 24167 30039
rect 26433 30005 26467 30039
rect 30757 30005 30791 30039
rect 37381 30005 37415 30039
rect 3433 29801 3467 29835
rect 6929 29801 6963 29835
rect 12541 29801 12575 29835
rect 12817 29801 12851 29835
rect 14105 29801 14139 29835
rect 15485 29801 15519 29835
rect 17601 29801 17635 29835
rect 18245 29801 18279 29835
rect 18521 29801 18555 29835
rect 19165 29801 19199 29835
rect 21373 29801 21407 29835
rect 22109 29801 22143 29835
rect 23765 29801 23799 29835
rect 24225 29801 24259 29835
rect 27813 29801 27847 29835
rect 28273 29801 28307 29835
rect 29745 29801 29779 29835
rect 32321 29801 32355 29835
rect 13001 29733 13035 29767
rect 1685 29665 1719 29699
rect 7573 29665 7607 29699
rect 7941 29665 7975 29699
rect 10149 29665 10183 29699
rect 11437 29665 11471 29699
rect 11713 29665 11747 29699
rect 13645 29665 13679 29699
rect 16497 29665 16531 29699
rect 19901 29665 19935 29699
rect 22569 29665 22603 29699
rect 23305 29665 23339 29699
rect 25237 29665 25271 29699
rect 26525 29665 26559 29699
rect 28273 29665 28307 29699
rect 28457 29665 28491 29699
rect 28825 29665 28859 29699
rect 30021 29665 30055 29699
rect 30481 29665 30515 29699
rect 34897 29665 34931 29699
rect 1409 29597 1443 29631
rect 7205 29597 7239 29631
rect 10057 29597 10091 29631
rect 10609 29597 10643 29631
rect 11897 29597 11931 29631
rect 16221 29597 16255 29631
rect 19993 29597 20027 29631
rect 22477 29597 22511 29631
rect 23397 29597 23431 29631
rect 24409 29597 24443 29631
rect 24501 29597 24535 29631
rect 25329 29597 25363 29631
rect 29929 29597 29963 29631
rect 30757 29597 30791 29631
rect 34069 29597 34103 29631
rect 34161 29597 34195 29631
rect 34989 29597 35023 29631
rect 7849 29529 7883 29563
rect 10885 29529 10919 29563
rect 11529 29529 11563 29563
rect 25789 29529 25823 29563
rect 27445 29529 27479 29563
rect 2789 29461 2823 29495
rect 8585 29461 8619 29495
rect 20453 29461 20487 29495
rect 26157 29461 26191 29495
rect 26709 29461 26743 29495
rect 27077 29461 27111 29495
rect 29469 29461 29503 29495
rect 31217 29461 31251 29495
rect 35449 29461 35483 29495
rect 35909 29461 35943 29495
rect 1685 29257 1719 29291
rect 4905 29257 4939 29291
rect 7849 29257 7883 29291
rect 10149 29257 10183 29291
rect 11253 29257 11287 29291
rect 12173 29257 12207 29291
rect 13277 29257 13311 29291
rect 15209 29257 15243 29291
rect 16313 29257 16347 29291
rect 22109 29257 22143 29291
rect 22845 29257 22879 29291
rect 23489 29257 23523 29291
rect 27997 29257 28031 29291
rect 28917 29257 28951 29291
rect 33701 29257 33735 29291
rect 33977 29257 34011 29291
rect 34345 29257 34379 29291
rect 36553 29257 36587 29291
rect 11529 29189 11563 29223
rect 21189 29189 21223 29223
rect 24777 29189 24811 29223
rect 27629 29189 27663 29223
rect 2053 29121 2087 29155
rect 3341 29121 3375 29155
rect 8493 29121 8527 29155
rect 13737 29121 13771 29155
rect 18797 29121 18831 29155
rect 19625 29121 19659 29155
rect 20269 29121 20303 29155
rect 24041 29121 24075 29155
rect 26985 29121 27019 29155
rect 3617 29053 3651 29087
rect 8585 29053 8619 29087
rect 8861 29053 8895 29087
rect 11345 29053 11379 29087
rect 12817 29053 12851 29087
rect 13829 29053 13863 29087
rect 14105 29053 14139 29087
rect 18889 29053 18923 29087
rect 20361 29053 20395 29087
rect 20913 29053 20947 29087
rect 21281 29053 21315 29087
rect 24869 29053 24903 29087
rect 25605 29053 25639 29087
rect 25973 29053 26007 29087
rect 26433 29053 26467 29087
rect 27445 29053 27479 29087
rect 3157 28985 3191 29019
rect 7113 28985 7147 29019
rect 7481 28985 7515 29019
rect 10517 28985 10551 29019
rect 11897 28985 11931 29019
rect 12725 28985 12759 29019
rect 18705 28985 18739 29019
rect 19349 28985 19383 29019
rect 24409 28985 24443 29019
rect 25053 28985 25087 29019
rect 25237 28985 25271 29019
rect 26249 28985 26283 29019
rect 27261 28985 27295 29019
rect 28733 28985 28767 29019
rect 30573 29189 30607 29223
rect 30941 29189 30975 29223
rect 29285 29121 29319 29155
rect 30297 29121 30331 29155
rect 31309 29121 31343 29155
rect 35449 29121 35483 29155
rect 29101 29053 29135 29087
rect 29837 29053 29871 29087
rect 30113 29053 30147 29087
rect 31217 29053 31251 29087
rect 32045 29053 32079 29087
rect 32137 29053 32171 29087
rect 35173 29053 35207 29087
rect 13001 28917 13035 28951
rect 16681 28917 16715 28951
rect 22477 28917 22511 28951
rect 25145 28917 25179 28951
rect 26617 28917 26651 28951
rect 28917 28917 28951 28951
rect 4905 28713 4939 28747
rect 11529 28713 11563 28747
rect 13461 28713 13495 28747
rect 16681 28713 16715 28747
rect 19349 28713 19383 28747
rect 20361 28713 20395 28747
rect 26249 28713 26283 28747
rect 28089 28713 28123 28747
rect 35265 28713 35299 28747
rect 26893 28645 26927 28679
rect 30757 28645 30791 28679
rect 1777 28577 1811 28611
rect 4721 28577 4755 28611
rect 6653 28577 6687 28611
rect 7021 28577 7055 28611
rect 8677 28577 8711 28611
rect 10609 28577 10643 28611
rect 10977 28577 11011 28611
rect 12909 28577 12943 28611
rect 13829 28577 13863 28611
rect 15577 28577 15611 28611
rect 22201 28577 22235 28611
rect 22937 28577 22971 28611
rect 24409 28577 24443 28611
rect 24961 28577 24995 28611
rect 25329 28577 25363 28611
rect 25421 28577 25455 28611
rect 26709 28577 26743 28611
rect 26801 28577 26835 28611
rect 28641 28577 28675 28611
rect 28825 28577 28859 28611
rect 29009 28577 29043 28611
rect 29285 28577 29319 28611
rect 30297 28577 30331 28611
rect 30481 28577 30515 28611
rect 33793 28577 33827 28611
rect 34161 28577 34195 28611
rect 1501 28509 1535 28543
rect 6745 28509 6779 28543
rect 7113 28509 7147 28543
rect 8033 28509 8067 28543
rect 11069 28509 11103 28543
rect 13001 28509 13035 28543
rect 14381 28509 14415 28543
rect 15301 28509 15335 28543
rect 17785 28509 17819 28543
rect 18061 28509 18095 28543
rect 22109 28509 22143 28543
rect 23029 28509 23063 28543
rect 23765 28509 23799 28543
rect 24501 28509 24535 28543
rect 26525 28509 26559 28543
rect 27261 28509 27295 28543
rect 10425 28441 10459 28475
rect 28457 28441 28491 28475
rect 33701 28509 33735 28543
rect 34253 28509 34287 28543
rect 32781 28441 32815 28475
rect 3065 28373 3099 28407
rect 6101 28373 6135 28407
rect 9137 28373 9171 28407
rect 14013 28373 14047 28407
rect 19809 28373 19843 28407
rect 27537 28373 27571 28407
rect 29285 28373 29319 28407
rect 29561 28373 29595 28407
rect 29929 28373 29963 28407
rect 31217 28373 31251 28407
rect 33241 28373 33275 28407
rect 35817 28373 35851 28407
rect 1593 28169 1627 28203
rect 2053 28169 2087 28203
rect 4721 28169 4755 28203
rect 6469 28169 6503 28203
rect 7389 28169 7423 28203
rect 10609 28169 10643 28203
rect 11253 28169 11287 28203
rect 11805 28169 11839 28203
rect 23121 28169 23155 28203
rect 24777 28169 24811 28203
rect 28181 28169 28215 28203
rect 28641 28169 28675 28203
rect 31677 28169 31711 28203
rect 32505 28169 32539 28203
rect 34529 28169 34563 28203
rect 5733 28101 5767 28135
rect 8309 28101 8343 28135
rect 10241 28101 10275 28135
rect 18613 28101 18647 28135
rect 19073 28101 19107 28135
rect 28917 28101 28951 28135
rect 30297 28101 30331 28135
rect 31309 28101 31343 28135
rect 8953 28033 8987 28067
rect 13553 28033 13587 28067
rect 14381 28033 14415 28067
rect 20913 28033 20947 28067
rect 22753 28033 22787 28067
rect 33425 28033 33459 28067
rect 34069 28033 34103 28067
rect 35725 28033 35759 28067
rect 36093 28033 36127 28067
rect 6101 27965 6135 27999
rect 7481 27965 7515 27999
rect 8861 27965 8895 27999
rect 9689 27965 9723 27999
rect 9781 27965 9815 27999
rect 13277 27965 13311 27999
rect 13461 27965 13495 27999
rect 14289 27965 14323 27999
rect 18337 27965 18371 27999
rect 19257 27965 19291 27999
rect 19441 27965 19475 27999
rect 19625 27965 19659 27999
rect 20545 27965 20579 27999
rect 21557 27965 21591 27999
rect 21833 27965 21867 27999
rect 22017 27965 22051 27999
rect 23949 27965 23983 27999
rect 24225 27965 24259 27999
rect 25329 27965 25363 27999
rect 25789 27965 25823 27999
rect 27353 27965 27387 27999
rect 27445 27965 27479 27999
rect 29101 27965 29135 27999
rect 29929 27965 29963 27999
rect 30481 27965 30515 27999
rect 30665 27965 30699 27999
rect 30849 27965 30883 27999
rect 32689 27965 32723 27999
rect 33149 27965 33183 27999
rect 35817 27965 35851 27999
rect 12725 27897 12759 27931
rect 17785 27897 17819 27931
rect 20085 27897 20119 27931
rect 21005 27897 21039 27931
rect 23489 27897 23523 27931
rect 25237 27897 25271 27931
rect 27169 27897 27203 27931
rect 27537 27897 27571 27931
rect 27905 27897 27939 27931
rect 29561 27897 29595 27931
rect 5365 27829 5399 27863
rect 7665 27829 7699 27863
rect 8585 27829 8619 27863
rect 10977 27829 11011 27863
rect 15393 27829 15427 27863
rect 15761 27829 15795 27863
rect 17509 27829 17543 27863
rect 22293 27829 22327 27863
rect 23765 27829 23799 27863
rect 25421 27829 25455 27863
rect 26525 27829 26559 27863
rect 26985 27829 27019 27863
rect 33701 27829 33735 27863
rect 37381 27829 37415 27863
rect 7481 27625 7515 27659
rect 8861 27625 8895 27659
rect 14197 27625 14231 27659
rect 21097 27625 21131 27659
rect 21557 27625 21591 27659
rect 22109 27625 22143 27659
rect 27721 27625 27755 27659
rect 29653 27625 29687 27659
rect 8585 27557 8619 27591
rect 11713 27557 11747 27591
rect 11805 27557 11839 27591
rect 12541 27557 12575 27591
rect 13829 27557 13863 27591
rect 23949 27557 23983 27591
rect 25973 27557 26007 27591
rect 29285 27557 29319 27591
rect 32689 27557 32723 27591
rect 1685 27489 1719 27523
rect 5733 27489 5767 27523
rect 6009 27489 6043 27523
rect 6653 27489 6687 27523
rect 6837 27489 6871 27523
rect 8033 27489 8067 27523
rect 8217 27489 8251 27523
rect 11069 27489 11103 27523
rect 13369 27489 13403 27523
rect 15301 27489 15335 27523
rect 16589 27489 16623 27523
rect 18797 27489 18831 27523
rect 22845 27489 22879 27523
rect 23857 27489 23891 27523
rect 24685 27489 24719 27523
rect 26893 27489 26927 27523
rect 27997 27489 28031 27523
rect 28825 27489 28859 27523
rect 31125 27489 31159 27523
rect 32137 27489 32171 27523
rect 32321 27489 32355 27523
rect 33517 27489 33551 27523
rect 34529 27489 34563 27523
rect 35817 27489 35851 27523
rect 36645 27489 36679 27523
rect 1409 27421 1443 27455
rect 3065 27421 3099 27455
rect 5549 27421 5583 27455
rect 12173 27421 12207 27455
rect 16313 27421 16347 27455
rect 22201 27421 22235 27455
rect 23673 27421 23707 27455
rect 24777 27421 24811 27455
rect 28089 27421 28123 27455
rect 28917 27421 28951 27455
rect 31217 27421 31251 27455
rect 35909 27421 35943 27455
rect 36737 27421 36771 27455
rect 5181 27353 5215 27387
rect 9965 27353 9999 27387
rect 18981 27353 19015 27387
rect 26341 27353 26375 27387
rect 27077 27353 27111 27387
rect 34713 27353 34747 27387
rect 3433 27285 3467 27319
rect 4997 27285 5031 27319
rect 7941 27285 7975 27319
rect 9321 27285 9355 27319
rect 10333 27285 10367 27319
rect 10793 27285 10827 27319
rect 11943 27285 11977 27319
rect 12081 27285 12115 27319
rect 13553 27285 13587 27319
rect 15485 27285 15519 27319
rect 17693 27285 17727 27319
rect 19349 27285 19383 27319
rect 25421 27285 25455 27319
rect 26709 27285 26743 27319
rect 27445 27285 27479 27319
rect 30205 27285 30239 27319
rect 31493 27285 31527 27319
rect 33149 27285 33183 27319
rect 33701 27285 33735 27319
rect 34989 27285 35023 27319
rect 2053 27081 2087 27115
rect 4537 27081 4571 27115
rect 5273 27081 5307 27115
rect 6009 27081 6043 27115
rect 7113 27081 7147 27115
rect 11897 27081 11931 27115
rect 13369 27081 13403 27115
rect 21005 27081 21039 27115
rect 22845 27081 22879 27115
rect 23489 27081 23523 27115
rect 25973 27081 26007 27115
rect 27905 27081 27939 27115
rect 28365 27081 28399 27115
rect 30205 27081 30239 27115
rect 31861 27081 31895 27115
rect 33977 27081 34011 27115
rect 36277 27081 36311 27115
rect 6285 27013 6319 27047
rect 8125 27013 8159 27047
rect 8585 27013 8619 27047
rect 12633 27013 12667 27047
rect 28733 27013 28767 27047
rect 30021 27013 30055 27047
rect 3433 26945 3467 26979
rect 21465 26945 21499 26979
rect 23765 26945 23799 26979
rect 25053 26945 25087 26979
rect 26341 26945 26375 26979
rect 30849 26945 30883 26979
rect 31217 26945 31251 26979
rect 34713 26945 34747 26979
rect 3249 26877 3283 26911
rect 3525 26877 3559 26911
rect 4077 26877 4111 26911
rect 4261 26877 4295 26911
rect 6837 26877 6871 26911
rect 6929 26877 6963 26911
rect 8493 26877 8527 26911
rect 8861 26877 8895 26911
rect 9137 26877 9171 26911
rect 10333 26877 10367 26911
rect 10701 26877 10735 26911
rect 11161 26877 11195 26911
rect 12449 26877 12483 26911
rect 14013 26877 14047 26911
rect 14473 26877 14507 26911
rect 16037 26877 16071 26911
rect 16129 26877 16163 26911
rect 16865 26877 16899 26911
rect 18521 26877 18555 26911
rect 19533 26877 19567 26911
rect 19717 26877 19751 26911
rect 19901 26877 19935 26911
rect 22017 26877 22051 26911
rect 22293 26877 22327 26911
rect 22477 26877 22511 26911
rect 24593 26877 24627 26911
rect 24685 26877 24719 26911
rect 26249 26877 26283 26911
rect 26801 26877 26835 26911
rect 26985 26877 27019 26911
rect 27169 26877 27203 26911
rect 28181 26877 28215 26911
rect 29653 26877 29687 26911
rect 30757 26877 30791 26911
rect 31125 26877 31159 26911
rect 32413 26877 32447 26911
rect 32505 26877 32539 26911
rect 33793 26877 33827 26911
rect 34897 26877 34931 26911
rect 35173 26877 35207 26911
rect 2881 26809 2915 26843
rect 5641 26809 5675 26843
rect 9689 26809 9723 26843
rect 11437 26809 11471 26843
rect 14841 26809 14875 26843
rect 15301 26809 15335 26843
rect 16589 26809 16623 26843
rect 17325 26809 17359 26843
rect 19073 26809 19107 26843
rect 21373 26809 21407 26843
rect 23857 26809 23891 26843
rect 25605 26809 25639 26843
rect 32965 26809 32999 26843
rect 33609 26809 33643 26843
rect 1593 26741 1627 26775
rect 7665 26741 7699 26775
rect 10149 26741 10183 26775
rect 12173 26741 12207 26775
rect 12909 26741 12943 26775
rect 15853 26741 15887 26775
rect 18797 26741 18831 26775
rect 26065 26741 26099 26775
rect 32229 26741 32263 26775
rect 34345 26741 34379 26775
rect 36921 26741 36955 26775
rect 1685 26537 1719 26571
rect 3341 26537 3375 26571
rect 4537 26537 4571 26571
rect 6193 26537 6227 26571
rect 8033 26537 8067 26571
rect 14289 26537 14323 26571
rect 16405 26537 16439 26571
rect 16865 26537 16899 26571
rect 24041 26537 24075 26571
rect 24409 26537 24443 26571
rect 25973 26537 26007 26571
rect 27997 26537 28031 26571
rect 31953 26537 31987 26571
rect 34713 26537 34747 26571
rect 35725 26537 35759 26571
rect 36093 26537 36127 26571
rect 9689 26469 9723 26503
rect 16957 26469 16991 26503
rect 19993 26469 20027 26503
rect 23765 26469 23799 26503
rect 26249 26469 26283 26503
rect 28273 26469 28307 26503
rect 29101 26469 29135 26503
rect 32873 26469 32907 26503
rect 4905 26401 4939 26435
rect 5273 26401 5307 26435
rect 6469 26401 6503 26435
rect 6653 26401 6687 26435
rect 7021 26401 7055 26435
rect 7481 26401 7515 26435
rect 10149 26401 10183 26435
rect 10517 26401 10551 26435
rect 10609 26401 10643 26435
rect 12265 26401 12299 26435
rect 12449 26401 12483 26435
rect 12725 26401 12759 26435
rect 14105 26401 14139 26435
rect 15301 26401 15335 26435
rect 17601 26401 17635 26435
rect 17969 26401 18003 26435
rect 18153 26401 18187 26435
rect 19533 26401 19567 26435
rect 21097 26401 21131 26435
rect 21465 26401 21499 26435
rect 21833 26401 21867 26435
rect 27445 26401 27479 26435
rect 27537 26401 27571 26435
rect 29745 26401 29779 26435
rect 29837 26401 29871 26435
rect 30113 26401 30147 26435
rect 30297 26401 30331 26435
rect 31309 26401 31343 26435
rect 33057 26401 33091 26435
rect 33701 26401 33735 26435
rect 34529 26401 34563 26435
rect 34989 26401 35023 26435
rect 5549 26333 5583 26367
rect 9137 26333 9171 26367
rect 11805 26333 11839 26367
rect 13001 26333 13035 26367
rect 13185 26333 13219 26367
rect 17417 26333 17451 26367
rect 19441 26333 19475 26367
rect 26617 26333 26651 26367
rect 26709 26333 26743 26367
rect 4997 26265 5031 26299
rect 7481 26265 7515 26299
rect 8401 26265 8435 26299
rect 8769 26265 8803 26299
rect 11345 26265 11379 26299
rect 13553 26265 13587 26299
rect 15485 26265 15519 26299
rect 19165 26265 19199 26299
rect 21741 26265 21775 26299
rect 29009 26265 29043 26299
rect 32505 26265 32539 26299
rect 10977 26197 11011 26231
rect 15761 26197 15795 26231
rect 18429 26197 18463 26231
rect 22385 26197 22419 26231
rect 30665 26197 30699 26231
rect 30941 26197 30975 26231
rect 31125 26197 31159 26231
rect 2789 25993 2823 26027
rect 4997 25993 5031 26027
rect 8953 25993 8987 26027
rect 11805 25993 11839 26027
rect 13829 25993 13863 26027
rect 15301 25993 15335 26027
rect 17049 25993 17083 26027
rect 17693 25993 17727 26027
rect 19625 25993 19659 26027
rect 21005 25993 21039 26027
rect 21373 25993 21407 26027
rect 21741 25993 21775 26027
rect 22477 25993 22511 26027
rect 26065 25993 26099 26027
rect 26525 25993 26559 26027
rect 27813 25993 27847 26027
rect 29561 25993 29595 26027
rect 30113 25993 30147 26027
rect 30941 25993 30975 26027
rect 34529 25993 34563 26027
rect 37381 25993 37415 26027
rect 10425 25925 10459 25959
rect 12633 25925 12667 25959
rect 17417 25925 17451 25959
rect 26801 25925 26835 25959
rect 29101 25925 29135 25959
rect 1409 25857 1443 25891
rect 4629 25857 4663 25891
rect 6837 25857 6871 25891
rect 7849 25857 7883 25891
rect 8677 25857 8711 25891
rect 10241 25857 10275 25891
rect 10885 25857 10919 25891
rect 14197 25857 14231 25891
rect 16405 25857 16439 25891
rect 18521 25857 18555 25891
rect 23489 25857 23523 25891
rect 30665 25857 30699 25891
rect 35725 25857 35759 25891
rect 1685 25789 1719 25823
rect 3801 25789 3835 25823
rect 4537 25789 4571 25823
rect 5917 25789 5951 25823
rect 7389 25789 7423 25823
rect 7665 25789 7699 25823
rect 8769 25789 8803 25823
rect 10977 25789 11011 25823
rect 11345 25789 11379 25823
rect 11529 25789 11563 25823
rect 12265 25789 12299 25823
rect 14381 25789 14415 25823
rect 14841 25789 14875 25823
rect 15945 25789 15979 25823
rect 16221 25789 16255 25823
rect 18245 25789 18279 25823
rect 22661 25789 22695 25823
rect 23673 25789 23707 25823
rect 23949 25789 23983 25823
rect 26617 25789 26651 25823
rect 27077 25789 27111 25823
rect 27629 25789 27663 25823
rect 29285 25789 29319 25823
rect 29377 25789 29411 25823
rect 30757 25789 30791 25823
rect 31493 25789 31527 25823
rect 31953 25789 31987 25823
rect 32873 25789 32907 25823
rect 33241 25789 33275 25823
rect 33333 25789 33367 25823
rect 33701 25789 33735 25823
rect 35817 25789 35851 25823
rect 36093 25789 36127 25823
rect 13001 25721 13035 25755
rect 15393 25721 15427 25755
rect 30573 25721 30607 25755
rect 32413 25721 32447 25755
rect 5273 25653 5307 25687
rect 6193 25653 6227 25687
rect 6561 25653 6595 25687
rect 8217 25653 8251 25687
rect 8585 25653 8619 25687
rect 9781 25653 9815 25687
rect 13369 25653 13403 25687
rect 14565 25653 14599 25687
rect 20269 25653 20303 25687
rect 25053 25653 25087 25687
rect 28181 25653 28215 25687
rect 28733 25653 28767 25687
rect 32321 25653 32355 25687
rect 6193 25449 6227 25483
rect 9965 25449 9999 25483
rect 12081 25449 12115 25483
rect 12541 25449 12575 25483
rect 14381 25449 14415 25483
rect 15485 25449 15519 25483
rect 18337 25449 18371 25483
rect 19441 25449 19475 25483
rect 21189 25449 21223 25483
rect 23673 25449 23707 25483
rect 29009 25449 29043 25483
rect 30205 25449 30239 25483
rect 30941 25449 30975 25483
rect 31861 25449 31895 25483
rect 33701 25449 33735 25483
rect 35817 25449 35851 25483
rect 7205 25381 7239 25415
rect 8953 25381 8987 25415
rect 10425 25381 10459 25415
rect 16681 25381 16715 25415
rect 27261 25381 27295 25415
rect 29837 25381 29871 25415
rect 32689 25381 32723 25415
rect 4353 25313 4387 25347
rect 4629 25313 4663 25347
rect 5181 25313 5215 25347
rect 7665 25313 7699 25347
rect 7849 25313 7883 25347
rect 8125 25313 8159 25347
rect 8677 25313 8711 25347
rect 11253 25313 11287 25347
rect 11621 25313 11655 25347
rect 12633 25313 12667 25347
rect 13185 25313 13219 25347
rect 13369 25313 13403 25347
rect 13553 25313 13587 25347
rect 14105 25313 14139 25347
rect 17141 25313 17175 25347
rect 17509 25313 17543 25347
rect 21557 25313 21591 25347
rect 21925 25313 21959 25347
rect 25421 25313 25455 25347
rect 28089 25313 28123 25347
rect 29285 25313 29319 25347
rect 29377 25313 29411 25347
rect 30665 25313 30699 25347
rect 30849 25313 30883 25347
rect 32229 25313 32263 25347
rect 33517 25313 33551 25347
rect 5273 25245 5307 25279
rect 8309 25245 8343 25279
rect 11345 25245 11379 25279
rect 11713 25245 11747 25279
rect 13737 25245 13771 25279
rect 15945 25245 15979 25279
rect 17601 25245 17635 25279
rect 21373 25245 21407 25279
rect 21833 25245 21867 25279
rect 27813 25245 27847 25279
rect 28273 25245 28307 25279
rect 29101 25245 29135 25279
rect 31493 25245 31527 25279
rect 32137 25245 32171 25279
rect 4721 25177 4755 25211
rect 10701 25177 10735 25211
rect 15117 25177 15151 25211
rect 25053 25177 25087 25211
rect 1685 25109 1719 25143
rect 6469 25109 6503 25143
rect 6929 25109 6963 25143
rect 9505 25109 9539 25143
rect 16221 25109 16255 25143
rect 25605 25109 25639 25143
rect 26801 25109 26835 25143
rect 27077 25109 27111 25143
rect 30573 25109 30607 25143
rect 10793 24905 10827 24939
rect 13921 24905 13955 24939
rect 17233 24905 17267 24939
rect 17509 24905 17543 24939
rect 26985 24905 27019 24939
rect 29101 24905 29135 24939
rect 8217 24837 8251 24871
rect 12541 24837 12575 24871
rect 27721 24837 27755 24871
rect 32781 24837 32815 24871
rect 4261 24769 4295 24803
rect 4629 24769 4663 24803
rect 5273 24769 5307 24803
rect 5825 24769 5859 24803
rect 8769 24769 8803 24803
rect 11805 24769 11839 24803
rect 13553 24769 13587 24803
rect 14289 24769 14323 24803
rect 15301 24769 15335 24803
rect 16221 24769 16255 24803
rect 19809 24769 19843 24803
rect 20177 24769 20211 24803
rect 21557 24769 21591 24803
rect 22201 24769 22235 24803
rect 24869 24769 24903 24803
rect 27261 24769 27295 24803
rect 29745 24769 29779 24803
rect 31217 24769 31251 24803
rect 35725 24769 35759 24803
rect 36093 24769 36127 24803
rect 3433 24701 3467 24735
rect 4169 24701 4203 24735
rect 5365 24701 5399 24735
rect 6101 24701 6135 24735
rect 7113 24701 7147 24735
rect 7573 24701 7607 24735
rect 9413 24701 9447 24735
rect 9689 24701 9723 24735
rect 9781 24701 9815 24735
rect 10057 24701 10091 24735
rect 10425 24701 10459 24735
rect 11345 24701 11379 24735
rect 13093 24701 13127 24735
rect 13185 24701 13219 24735
rect 13461 24701 13495 24735
rect 14473 24701 14507 24735
rect 14933 24701 14967 24735
rect 16313 24701 16347 24735
rect 16681 24701 16715 24735
rect 16865 24701 16899 24735
rect 19901 24701 19935 24735
rect 24961 24701 24995 24735
rect 25329 24701 25363 24735
rect 25697 24701 25731 24735
rect 26249 24701 26283 24735
rect 27629 24701 27663 24735
rect 27905 24701 27939 24735
rect 29285 24701 29319 24735
rect 30113 24701 30147 24735
rect 30573 24701 30607 24735
rect 31493 24701 31527 24735
rect 31677 24701 31711 24735
rect 32597 24701 32631 24735
rect 35817 24701 35851 24735
rect 6837 24633 6871 24667
rect 7205 24633 7239 24667
rect 8953 24633 8987 24667
rect 11161 24633 11195 24667
rect 26157 24633 26191 24667
rect 28365 24633 28399 24667
rect 30665 24633 30699 24667
rect 5089 24565 5123 24599
rect 6653 24565 6687 24599
rect 7021 24565 7055 24599
rect 7849 24565 7883 24599
rect 11529 24565 11563 24599
rect 12265 24565 12299 24599
rect 14657 24565 14691 24599
rect 15945 24565 15979 24599
rect 21833 24565 21867 24599
rect 24409 24565 24443 24599
rect 28641 24565 28675 24599
rect 29469 24565 29503 24599
rect 32229 24565 32263 24599
rect 33517 24565 33551 24599
rect 37197 24565 37231 24599
rect 2973 24361 3007 24395
rect 3525 24361 3559 24395
rect 7757 24361 7791 24395
rect 16681 24361 16715 24395
rect 17049 24361 17083 24395
rect 21189 24361 21223 24395
rect 24041 24361 24075 24395
rect 25053 24361 25087 24395
rect 28273 24361 28307 24395
rect 31217 24361 31251 24395
rect 31493 24361 31527 24395
rect 32321 24361 32355 24395
rect 32597 24361 32631 24395
rect 32965 24361 32999 24395
rect 35817 24361 35851 24395
rect 4353 24293 4387 24327
rect 9689 24293 9723 24327
rect 11805 24293 11839 24327
rect 14657 24293 14691 24327
rect 15301 24293 15335 24327
rect 17325 24293 17359 24327
rect 25973 24293 26007 24327
rect 26893 24293 26927 24327
rect 1409 24225 1443 24259
rect 4997 24225 5031 24259
rect 5365 24225 5399 24259
rect 6193 24225 6227 24259
rect 6377 24225 6411 24259
rect 7113 24225 7147 24259
rect 7389 24225 7423 24259
rect 7573 24225 7607 24259
rect 8217 24225 8251 24259
rect 10241 24225 10275 24259
rect 10333 24225 10367 24259
rect 10517 24225 10551 24259
rect 12541 24225 12575 24259
rect 13921 24225 13955 24259
rect 16129 24225 16163 24259
rect 17877 24225 17911 24259
rect 22661 24225 22695 24259
rect 25421 24225 25455 24259
rect 27261 24225 27295 24259
rect 28457 24225 28491 24259
rect 28733 24225 28767 24259
rect 30021 24225 30055 24259
rect 31033 24225 31067 24259
rect 32137 24225 32171 24259
rect 1685 24157 1719 24191
rect 4905 24157 4939 24191
rect 5457 24157 5491 24191
rect 8953 24157 8987 24191
rect 10885 24157 10919 24191
rect 11069 24157 11103 24191
rect 12449 24157 12483 24191
rect 13001 24157 13035 24191
rect 13829 24157 13863 24191
rect 14381 24157 14415 24191
rect 15853 24157 15887 24191
rect 16313 24157 16347 24191
rect 17601 24157 17635 24191
rect 21465 24157 21499 24191
rect 22937 24157 22971 24191
rect 28549 24157 28583 24191
rect 29193 24157 29227 24191
rect 5825 24089 5859 24123
rect 9321 24089 9355 24123
rect 12357 24089 12391 24123
rect 13737 24089 13771 24123
rect 15117 24089 15151 24123
rect 20637 24089 20671 24123
rect 25605 24089 25639 24123
rect 30205 24089 30239 24123
rect 3893 24021 3927 24055
rect 8677 24021 8711 24055
rect 11529 24021 11563 24055
rect 13369 24021 13403 24055
rect 18981 24021 19015 24055
rect 19993 24021 20027 24055
rect 27905 24021 27939 24055
rect 29561 24021 29595 24055
rect 30757 24021 30791 24055
rect 1593 23817 1627 23851
rect 3801 23817 3835 23851
rect 5181 23817 5215 23851
rect 5917 23817 5951 23851
rect 9781 23817 9815 23851
rect 10149 23817 10183 23851
rect 12173 23817 12207 23851
rect 12725 23817 12759 23851
rect 15301 23817 15335 23851
rect 17417 23817 17451 23851
rect 18889 23817 18923 23851
rect 20361 23817 20395 23851
rect 23121 23817 23155 23851
rect 25881 23817 25915 23851
rect 27169 23817 27203 23851
rect 28641 23817 28675 23851
rect 30389 23817 30423 23851
rect 1961 23749 1995 23783
rect 2329 23749 2363 23783
rect 4905 23749 4939 23783
rect 14381 23749 14415 23783
rect 24869 23749 24903 23783
rect 25237 23749 25271 23783
rect 27721 23749 27755 23783
rect 3433 23681 3467 23715
rect 6837 23681 6871 23715
rect 7573 23681 7607 23715
rect 11529 23681 11563 23715
rect 17141 23681 17175 23715
rect 17785 23681 17819 23715
rect 18521 23681 18555 23715
rect 21465 23681 21499 23715
rect 29101 23681 29135 23715
rect 30113 23681 30147 23715
rect 31125 23681 31159 23715
rect 35725 23681 35759 23715
rect 36093 23681 36127 23715
rect 5733 23613 5767 23647
rect 6193 23613 6227 23647
rect 6653 23613 6687 23647
rect 7113 23613 7147 23647
rect 8861 23613 8895 23647
rect 10701 23613 10735 23647
rect 10793 23613 10827 23647
rect 11069 23613 11103 23647
rect 13553 23613 13587 23647
rect 13645 23613 13679 23647
rect 13921 23613 13955 23647
rect 14013 23613 14047 23647
rect 15117 23613 15151 23647
rect 15577 23613 15611 23647
rect 16681 23613 16715 23647
rect 16957 23613 16991 23647
rect 18613 23613 18647 23647
rect 18705 23613 18739 23647
rect 21005 23613 21039 23647
rect 21189 23613 21223 23647
rect 21557 23613 21591 23647
rect 25053 23613 25087 23647
rect 26157 23613 26191 23647
rect 27445 23613 27479 23647
rect 27629 23613 27663 23647
rect 27905 23613 27939 23647
rect 29561 23613 29595 23647
rect 29653 23613 29687 23647
rect 30849 23613 30883 23647
rect 31493 23613 31527 23647
rect 31769 23613 31803 23647
rect 35817 23613 35851 23647
rect 3065 23545 3099 23579
rect 4537 23545 4571 23579
rect 5641 23545 5675 23579
rect 7205 23545 7239 23579
rect 8585 23545 8619 23579
rect 8953 23545 8987 23579
rect 9321 23545 9355 23579
rect 10977 23545 11011 23579
rect 12909 23545 12943 23579
rect 15025 23545 15059 23579
rect 16129 23545 16163 23579
rect 19441 23545 19475 23579
rect 19993 23545 20027 23579
rect 22753 23545 22787 23579
rect 26801 23545 26835 23579
rect 28365 23545 28399 23579
rect 32045 23545 32079 23579
rect 4169 23477 4203 23511
rect 7021 23477 7055 23511
rect 8033 23477 8067 23511
rect 8401 23477 8435 23511
rect 8769 23477 8803 23511
rect 11805 23477 11839 23511
rect 16037 23477 16071 23511
rect 20821 23477 20855 23511
rect 25513 23477 25547 23511
rect 32413 23477 32447 23511
rect 37381 23477 37415 23511
rect 3893 23273 3927 23307
rect 6101 23273 6135 23307
rect 6469 23273 6503 23307
rect 9045 23273 9079 23307
rect 9873 23273 9907 23307
rect 10149 23273 10183 23307
rect 10517 23273 10551 23307
rect 14657 23273 14691 23307
rect 15669 23273 15703 23307
rect 16865 23273 16899 23307
rect 17693 23273 17727 23307
rect 21097 23273 21131 23307
rect 23857 23273 23891 23307
rect 25605 23273 25639 23307
rect 26249 23273 26283 23307
rect 27629 23273 27663 23307
rect 27997 23273 28031 23307
rect 28365 23273 28399 23307
rect 29837 23273 29871 23307
rect 31033 23273 31067 23307
rect 31401 23273 31435 23307
rect 31769 23273 31803 23307
rect 31953 23273 31987 23307
rect 35817 23273 35851 23307
rect 6285 23205 6319 23239
rect 6653 23205 6687 23239
rect 7021 23205 7055 23239
rect 8401 23205 8435 23239
rect 12081 23205 12115 23239
rect 12909 23205 12943 23239
rect 17969 23205 18003 23239
rect 26525 23205 26559 23239
rect 1501 23137 1535 23171
rect 4261 23137 4295 23171
rect 4813 23137 4847 23171
rect 4997 23137 5031 23171
rect 6561 23137 6595 23171
rect 8217 23137 8251 23171
rect 8309 23137 8343 23171
rect 9689 23137 9723 23171
rect 11529 23137 11563 23171
rect 11621 23137 11655 23171
rect 13369 23137 13403 23171
rect 13553 23137 13587 23171
rect 13829 23137 13863 23171
rect 15117 23137 15151 23171
rect 16037 23137 16071 23171
rect 16405 23137 16439 23171
rect 18889 23137 18923 23171
rect 19073 23137 19107 23171
rect 19257 23137 19291 23171
rect 20913 23137 20947 23171
rect 21373 23137 21407 23171
rect 22753 23137 22787 23171
rect 25421 23137 25455 23171
rect 29101 23137 29135 23171
rect 29377 23137 29411 23171
rect 29561 23137 29595 23171
rect 32321 23137 32355 23171
rect 33057 23137 33091 23171
rect 1777 23069 1811 23103
rect 4169 23069 4203 23103
rect 7665 23069 7699 23103
rect 8033 23069 8067 23103
rect 8769 23069 8803 23103
rect 14197 23069 14231 23103
rect 14289 23069 14323 23103
rect 15853 23069 15887 23103
rect 16313 23069 16347 23103
rect 17233 23069 17267 23103
rect 22477 23069 22511 23103
rect 26893 23069 26927 23103
rect 28549 23069 28583 23103
rect 31953 23069 31987 23103
rect 32229 23069 32263 23103
rect 33149 23069 33183 23103
rect 5181 23001 5215 23035
rect 10885 23001 10919 23035
rect 18705 23001 18739 23035
rect 26801 23001 26835 23035
rect 3065 22933 3099 22967
rect 3525 22933 3559 22967
rect 5733 22933 5767 22967
rect 7297 22933 7331 22967
rect 9413 22933 9447 22967
rect 11345 22933 11379 22967
rect 12449 22933 12483 22967
rect 12817 22933 12851 22967
rect 20545 22933 20579 22967
rect 25973 22933 26007 22967
rect 26663 22933 26697 22967
rect 27169 22933 27203 22967
rect 30297 22933 30331 22967
rect 1685 22729 1719 22763
rect 4169 22729 4203 22763
rect 4537 22729 4571 22763
rect 5181 22729 5215 22763
rect 10590 22729 10624 22763
rect 11069 22729 11103 22763
rect 12265 22729 12299 22763
rect 13645 22729 13679 22763
rect 15945 22729 15979 22763
rect 17417 22729 17451 22763
rect 18245 22729 18279 22763
rect 18613 22729 18647 22763
rect 19257 22729 19291 22763
rect 19625 22729 19659 22763
rect 19993 22729 20027 22763
rect 21557 22729 21591 22763
rect 22569 22729 22603 22763
rect 22937 22729 22971 22763
rect 25881 22729 25915 22763
rect 26985 22729 27019 22763
rect 28641 22729 28675 22763
rect 32137 22729 32171 22763
rect 32505 22729 32539 22763
rect 8309 22661 8343 22695
rect 8677 22661 8711 22695
rect 9873 22661 9907 22695
rect 10701 22661 10735 22695
rect 11437 22661 11471 22695
rect 13093 22661 13127 22695
rect 13323 22661 13357 22695
rect 26157 22661 26191 22695
rect 27169 22661 27203 22695
rect 28917 22661 28951 22695
rect 29469 22661 29503 22695
rect 32965 22661 32999 22695
rect 2145 22593 2179 22627
rect 3341 22593 3375 22627
rect 8861 22593 8895 22627
rect 10793 22593 10827 22627
rect 12725 22593 12759 22627
rect 13553 22593 13587 22627
rect 14289 22593 14323 22627
rect 16681 22593 16715 22627
rect 17141 22593 17175 22627
rect 18889 22593 18923 22627
rect 20184 22593 20218 22627
rect 25513 22593 25547 22627
rect 28089 22593 28123 22627
rect 35725 22593 35759 22627
rect 37289 22593 37323 22627
rect 2513 22525 2547 22559
rect 3249 22525 3283 22559
rect 3617 22525 3651 22559
rect 3801 22525 3835 22559
rect 4905 22525 4939 22559
rect 4997 22525 5031 22559
rect 5733 22525 5767 22559
rect 7481 22525 7515 22559
rect 9045 22525 9079 22559
rect 13415 22525 13449 22559
rect 14657 22525 14691 22559
rect 14749 22525 14783 22559
rect 14841 22525 14875 22559
rect 15577 22525 15611 22559
rect 16957 22525 16991 22559
rect 18061 22525 18095 22559
rect 20453 22525 20487 22559
rect 24685 22525 24719 22559
rect 25421 22525 25455 22559
rect 27077 22525 27111 22559
rect 27353 22525 27387 22559
rect 27813 22525 27847 22559
rect 29285 22525 29319 22559
rect 30113 22525 30147 22559
rect 30389 22525 30423 22559
rect 35817 22525 35851 22559
rect 36093 22525 36127 22559
rect 2605 22457 2639 22491
rect 7297 22457 7331 22491
rect 7665 22457 7699 22491
rect 8033 22457 8067 22491
rect 9229 22457 9263 22491
rect 9597 22457 9631 22491
rect 10425 22457 10459 22491
rect 11897 22457 11931 22491
rect 13185 22457 13219 22491
rect 15301 22457 15335 22491
rect 16129 22457 16163 22491
rect 17785 22457 17819 22491
rect 26617 22457 26651 22491
rect 29745 22457 29779 22491
rect 31033 22457 31067 22491
rect 6377 22389 6411 22423
rect 7205 22389 7239 22423
rect 7573 22389 7607 22423
rect 9137 22389 9171 22423
rect 10241 22389 10275 22423
rect 3065 22185 3099 22219
rect 3893 22185 3927 22219
rect 5365 22185 5399 22219
rect 5733 22185 5767 22219
rect 6469 22185 6503 22219
rect 8769 22185 8803 22219
rect 9045 22185 9079 22219
rect 9413 22185 9447 22219
rect 9965 22185 9999 22219
rect 15853 22185 15887 22219
rect 16221 22185 16255 22219
rect 19533 22185 19567 22219
rect 20177 22185 20211 22219
rect 26341 22185 26375 22219
rect 35817 22185 35851 22219
rect 5825 22117 5859 22151
rect 8033 22117 8067 22151
rect 10057 22117 10091 22151
rect 10701 22117 10735 22151
rect 12541 22117 12575 22151
rect 15577 22117 15611 22151
rect 2697 22049 2731 22083
rect 4445 22049 4479 22083
rect 4997 22049 5031 22083
rect 5089 22049 5123 22083
rect 5457 22049 5491 22083
rect 5641 22049 5675 22083
rect 7021 22049 7055 22083
rect 7168 22049 7202 22083
rect 8585 22049 8619 22083
rect 9873 22049 9907 22083
rect 11069 22049 11103 22083
rect 11253 22049 11287 22083
rect 11437 22049 11471 22083
rect 12633 22049 12667 22083
rect 12817 22049 12851 22083
rect 13921 22049 13955 22083
rect 14657 22049 14691 22083
rect 16773 22049 16807 22083
rect 17141 22049 17175 22083
rect 18981 22049 19015 22083
rect 21281 22049 21315 22083
rect 22097 22049 22131 22083
rect 23673 22049 23707 22083
rect 24041 22049 24075 22083
rect 27353 22049 27387 22083
rect 28825 22049 28859 22083
rect 30481 22049 30515 22083
rect 31033 22049 31067 22083
rect 32689 22049 32723 22083
rect 1685 21981 1719 22015
rect 4353 21981 4387 22015
rect 4629 21913 4663 21947
rect 2053 21845 2087 21879
rect 3525 21845 3559 21879
rect 5089 21845 5123 21879
rect 5181 21981 5215 22015
rect 6193 21981 6227 22015
rect 7389 21981 7423 22015
rect 7665 21981 7699 22015
rect 9689 21981 9723 22015
rect 10425 21981 10459 22015
rect 12081 21981 12115 22015
rect 14289 21981 14323 22015
rect 16589 21981 16623 22015
rect 17049 21981 17083 22015
rect 18153 21981 18187 22015
rect 18705 21981 18739 22015
rect 19165 21981 19199 22015
rect 21373 21981 21407 22015
rect 22201 21981 22235 22015
rect 23305 21981 23339 22015
rect 26525 21981 26559 22015
rect 27077 21981 27111 22015
rect 27537 21981 27571 22015
rect 30297 21981 30331 22015
rect 30941 21981 30975 22015
rect 32965 21981 32999 22015
rect 17601 21913 17635 21947
rect 23949 21913 23983 21947
rect 5181 21845 5215 21879
rect 6929 21845 6963 21879
rect 7297 21845 7331 21879
rect 8493 21845 8527 21879
rect 11529 21845 11563 21879
rect 12909 21845 12943 21879
rect 13553 21845 13587 21879
rect 15025 21845 15059 21879
rect 17969 21845 18003 21879
rect 25697 21845 25731 21879
rect 28641 21845 28675 21879
rect 31585 21845 31619 21879
rect 34069 21845 34103 21879
rect 4077 21641 4111 21675
rect 5549 21641 5583 21675
rect 5917 21641 5951 21675
rect 9413 21641 9447 21675
rect 9762 21641 9796 21675
rect 10241 21641 10275 21675
rect 11989 21641 12023 21675
rect 16221 21641 16255 21675
rect 17785 21641 17819 21675
rect 20177 21641 20211 21675
rect 21189 21641 21223 21675
rect 27077 21641 27111 21675
rect 28549 21641 28583 21675
rect 32781 21641 32815 21675
rect 33057 21641 33091 21675
rect 35265 21641 35299 21675
rect 37197 21641 37231 21675
rect 1869 21573 1903 21607
rect 5181 21573 5215 21607
rect 9137 21573 9171 21607
rect 9873 21573 9907 21607
rect 11069 21573 11103 21607
rect 13369 21573 13403 21607
rect 20821 21573 20855 21607
rect 24501 21573 24535 21607
rect 26525 21573 26559 21607
rect 28181 21573 28215 21607
rect 30205 21573 30239 21607
rect 30481 21573 30515 21607
rect 1961 21505 1995 21539
rect 2697 21505 2731 21539
rect 4813 21505 4847 21539
rect 6653 21505 6687 21539
rect 6837 21505 6871 21539
rect 9965 21505 9999 21539
rect 14105 21505 14139 21539
rect 15945 21505 15979 21539
rect 18705 21505 18739 21539
rect 23489 21505 23523 21539
rect 23857 21505 23891 21539
rect 28825 21505 28859 21539
rect 32413 21505 32447 21539
rect 36093 21505 36127 21539
rect 2605 21437 2639 21471
rect 2973 21437 3007 21471
rect 3065 21437 3099 21471
rect 4261 21437 4295 21471
rect 5733 21437 5767 21471
rect 6193 21437 6227 21471
rect 7021 21437 7055 21471
rect 8585 21437 8619 21471
rect 9597 21437 9631 21471
rect 10609 21437 10643 21471
rect 11161 21437 11195 21471
rect 12541 21437 12575 21471
rect 13553 21437 13587 21471
rect 13645 21437 13679 21471
rect 14841 21437 14875 21471
rect 15485 21437 15519 21471
rect 15761 21437 15795 21471
rect 16589 21437 16623 21471
rect 18797 21437 18831 21471
rect 19073 21437 19107 21471
rect 21649 21437 21683 21471
rect 24041 21437 24075 21471
rect 24501 21437 24535 21471
rect 25513 21437 25547 21471
rect 25605 21437 25639 21471
rect 25973 21437 26007 21471
rect 26433 21437 26467 21471
rect 27997 21437 28031 21471
rect 29285 21437 29319 21471
rect 30297 21437 30331 21471
rect 30757 21437 30791 21471
rect 31217 21437 31251 21471
rect 31401 21437 31435 21471
rect 31677 21437 31711 21471
rect 32137 21437 32171 21471
rect 35725 21437 35759 21471
rect 35817 21437 35851 21471
rect 3433 21369 3467 21403
rect 7113 21369 7147 21403
rect 7205 21369 7239 21403
rect 7573 21369 7607 21403
rect 7941 21369 7975 21403
rect 14933 21369 14967 21403
rect 21281 21369 21315 21403
rect 4445 21301 4479 21335
rect 8401 21301 8435 21335
rect 8769 21301 8803 21335
rect 11345 21301 11379 21335
rect 11621 21301 11655 21335
rect 12725 21301 12759 21335
rect 13093 21301 13127 21335
rect 14381 21301 14415 21335
rect 16957 21301 16991 21335
rect 17325 21301 17359 21335
rect 18245 21301 18279 21335
rect 22385 21301 22419 21335
rect 22661 21301 22695 21335
rect 23121 21301 23155 21335
rect 27353 21301 27387 21335
rect 27721 21301 27755 21335
rect 29469 21301 29503 21335
rect 29837 21301 29871 21335
rect 3893 21097 3927 21131
rect 4353 21097 4387 21131
rect 6009 21097 6043 21131
rect 6929 21097 6963 21131
rect 7297 21097 7331 21131
rect 9137 21097 9171 21131
rect 9965 21097 9999 21131
rect 10701 21097 10735 21131
rect 12633 21097 12667 21131
rect 15485 21097 15519 21131
rect 16129 21097 16163 21131
rect 16865 21097 16899 21131
rect 24041 21097 24075 21131
rect 25697 21097 25731 21131
rect 26709 21097 26743 21131
rect 30205 21097 30239 21131
rect 36277 21097 36311 21131
rect 3157 21029 3191 21063
rect 7481 21029 7515 21063
rect 9873 21029 9907 21063
rect 10057 21029 10091 21063
rect 10425 21029 10459 21063
rect 14657 21029 14691 21063
rect 24225 21029 24259 21063
rect 27629 21029 27663 21063
rect 33333 21029 33367 21063
rect 1777 20961 1811 20995
rect 4813 20961 4847 20995
rect 5549 20961 5583 20995
rect 5641 20961 5675 20995
rect 6193 20961 6227 20995
rect 7389 20961 7423 20995
rect 11253 20961 11287 20995
rect 11437 20961 11471 20995
rect 13921 20961 13955 20995
rect 14197 20961 14231 20995
rect 15301 20961 15335 20995
rect 17233 20961 17267 20995
rect 17601 20961 17635 20995
rect 17785 20961 17819 20995
rect 18613 20961 18647 20995
rect 20453 20961 20487 20995
rect 22661 20961 22695 20995
rect 23121 20961 23155 20995
rect 25053 20961 25087 20995
rect 26525 20961 26559 20995
rect 28457 20961 28491 20995
rect 28917 20961 28951 20995
rect 29469 20961 29503 20995
rect 30297 20961 30331 20995
rect 32597 20961 32631 20995
rect 33057 20961 33091 20995
rect 34897 20961 34931 20995
rect 1501 20893 1535 20927
rect 7113 20893 7147 20927
rect 7849 20893 7883 20927
rect 9689 20893 9723 20927
rect 12265 20893 12299 20927
rect 13369 20893 13403 20927
rect 14381 20893 14415 20927
rect 17049 20893 17083 20927
rect 21649 20893 21683 20927
rect 22385 20893 22419 20927
rect 23673 20893 23707 20927
rect 24777 20893 24811 20927
rect 25237 20893 25271 20927
rect 28181 20893 28215 20927
rect 32321 20893 32355 20927
rect 35173 20893 35207 20927
rect 4721 20825 4755 20859
rect 20637 20825 20671 20859
rect 23121 20825 23155 20859
rect 27169 20825 27203 20859
rect 29009 20825 29043 20859
rect 8125 20757 8159 20791
rect 8861 20757 8895 20791
rect 11069 20757 11103 20791
rect 13277 20757 13311 20791
rect 15025 20757 15059 20791
rect 15853 20757 15887 20791
rect 18245 20757 18279 20791
rect 20085 20757 20119 20791
rect 21281 20757 21315 20791
rect 25973 20757 26007 20791
rect 27905 20757 27939 20791
rect 30481 20757 30515 20791
rect 30849 20757 30883 20791
rect 31309 20757 31343 20791
rect 31769 20757 31803 20791
rect 4629 20553 4663 20587
rect 5273 20553 5307 20587
rect 6009 20553 6043 20587
rect 6653 20553 6687 20587
rect 7113 20553 7147 20587
rect 9873 20553 9907 20587
rect 10498 20553 10532 20587
rect 12633 20553 12667 20587
rect 13093 20553 13127 20587
rect 17049 20553 17083 20587
rect 17417 20553 17451 20587
rect 18981 20553 19015 20587
rect 22385 20553 22419 20587
rect 24685 20553 24719 20587
rect 26525 20553 26559 20587
rect 28457 20553 28491 20587
rect 29009 20553 29043 20587
rect 30665 20553 30699 20587
rect 35449 20553 35483 20587
rect 4353 20485 4387 20519
rect 8677 20485 8711 20519
rect 10609 20485 10643 20519
rect 10793 20485 10827 20519
rect 11437 20485 11471 20519
rect 11805 20485 11839 20519
rect 13461 20485 13495 20519
rect 14473 20485 14507 20519
rect 15669 20485 15703 20519
rect 16773 20485 16807 20519
rect 25973 20485 26007 20519
rect 30113 20485 30147 20519
rect 32045 20485 32079 20519
rect 2421 20417 2455 20451
rect 3157 20417 3191 20451
rect 3341 20417 3375 20451
rect 5825 20417 5859 20451
rect 7941 20417 7975 20451
rect 8769 20417 8803 20451
rect 10149 20417 10183 20451
rect 10701 20417 10735 20451
rect 17785 20417 17819 20451
rect 19441 20417 19475 20451
rect 26985 20417 27019 20451
rect 3065 20349 3099 20383
rect 3433 20349 3467 20383
rect 4445 20349 4479 20383
rect 5457 20349 5491 20383
rect 1961 20281 1995 20315
rect 7389 20349 7423 20383
rect 7481 20349 7515 20383
rect 8953 20349 8987 20383
rect 9505 20349 9539 20383
rect 10333 20349 10367 20383
rect 13645 20349 13679 20383
rect 13829 20349 13863 20383
rect 14013 20349 14047 20383
rect 15853 20349 15887 20383
rect 16037 20349 16071 20383
rect 16221 20349 16255 20383
rect 19165 20349 19199 20383
rect 25053 20349 25087 20383
rect 25145 20349 25179 20383
rect 25697 20349 25731 20383
rect 25973 20349 26007 20383
rect 27629 20349 27663 20383
rect 27905 20349 27939 20383
rect 28089 20349 28123 20383
rect 29377 20349 29411 20383
rect 29653 20349 29687 20383
rect 30113 20349 30147 20383
rect 31217 20349 31251 20383
rect 31585 20349 31619 20383
rect 32137 20349 32171 20383
rect 7205 20281 7239 20315
rect 7565 20281 7599 20315
rect 9137 20281 9171 20315
rect 12081 20281 12115 20315
rect 14933 20281 14967 20315
rect 20821 20281 20855 20315
rect 23029 20281 23063 20315
rect 23949 20281 23983 20315
rect 27077 20281 27111 20315
rect 32965 20281 32999 20315
rect 2329 20213 2363 20247
rect 3985 20213 4019 20247
rect 4905 20213 4939 20247
rect 5641 20213 5675 20247
rect 5825 20213 5859 20247
rect 8217 20213 8251 20247
rect 9045 20213 9079 20247
rect 15301 20213 15335 20247
rect 18337 20213 18371 20247
rect 18613 20213 18647 20247
rect 21097 20213 21131 20247
rect 22661 20213 22695 20247
rect 24317 20213 24351 20247
rect 31125 20213 31159 20247
rect 32597 20213 32631 20247
rect 35173 20213 35207 20247
rect 1961 20009 1995 20043
rect 2513 20009 2547 20043
rect 3525 20009 3559 20043
rect 4629 20009 4663 20043
rect 4905 20009 4939 20043
rect 6193 20009 6227 20043
rect 7113 20009 7147 20043
rect 7481 20009 7515 20043
rect 8309 20009 8343 20043
rect 9413 20009 9447 20043
rect 10609 20009 10643 20043
rect 13645 20009 13679 20043
rect 19165 20009 19199 20043
rect 25237 20009 25271 20043
rect 26341 20009 26375 20043
rect 27629 20009 27663 20043
rect 29009 20009 29043 20043
rect 31493 20009 31527 20043
rect 1685 19941 1719 19975
rect 2881 19941 2915 19975
rect 5273 19941 5307 19975
rect 6837 19941 6871 19975
rect 7665 19941 7699 19975
rect 11621 19941 11655 19975
rect 15853 19941 15887 19975
rect 25881 19941 25915 19975
rect 34253 19941 34287 19975
rect 4721 19873 4755 19907
rect 5733 19873 5767 19907
rect 6009 19873 6043 19907
rect 7573 19873 7607 19907
rect 9965 19873 9999 19907
rect 12449 19873 12483 19907
rect 13921 19873 13955 19907
rect 15393 19873 15427 19907
rect 16957 19873 16991 19907
rect 17049 19873 17083 19907
rect 17417 19873 17451 19907
rect 17509 19873 17543 19907
rect 22109 19873 22143 19907
rect 22385 19873 22419 19907
rect 24041 19873 24075 19907
rect 24409 19873 24443 19907
rect 25421 19873 25455 19907
rect 27813 19873 27847 19907
rect 28365 19873 28399 19907
rect 28549 19873 28583 19907
rect 29745 19873 29779 19907
rect 30113 19873 30147 19907
rect 30297 19873 30331 19907
rect 33149 19873 33183 19907
rect 33517 19873 33551 19907
rect 33977 19873 34011 19907
rect 35909 19873 35943 19907
rect 7297 19805 7331 19839
rect 8033 19805 8067 19839
rect 10333 19805 10367 19839
rect 11345 19805 11379 19839
rect 12173 19805 12207 19839
rect 12633 19805 12667 19839
rect 13829 19805 13863 19839
rect 15301 19805 15335 19839
rect 21741 19805 21775 19839
rect 23673 19805 23707 19839
rect 32413 19805 32447 19839
rect 35081 19805 35115 19839
rect 35633 19805 35667 19839
rect 36093 19805 36127 19839
rect 5825 19737 5859 19771
rect 10241 19737 10275 19771
rect 15117 19737 15151 19771
rect 16589 19737 16623 19771
rect 17877 19737 17911 19771
rect 22385 19737 22419 19771
rect 24317 19737 24351 19771
rect 25605 19737 25639 19771
rect 30297 19737 30331 19771
rect 3893 19669 3927 19703
rect 5641 19669 5675 19703
rect 8861 19669 8895 19703
rect 10103 19669 10137 19703
rect 11069 19669 11103 19703
rect 13185 19669 13219 19703
rect 14105 19669 14139 19703
rect 14657 19669 14691 19703
rect 16221 19669 16255 19703
rect 18429 19669 18463 19703
rect 19809 19669 19843 19703
rect 26801 19669 26835 19703
rect 27077 19669 27111 19703
rect 29377 19669 29411 19703
rect 31125 19669 31159 19703
rect 33057 19669 33091 19703
rect 1869 19465 1903 19499
rect 3709 19465 3743 19499
rect 7849 19465 7883 19499
rect 8953 19465 8987 19499
rect 10149 19465 10183 19499
rect 13093 19465 13127 19499
rect 17509 19465 17543 19499
rect 17601 19465 17635 19499
rect 21741 19465 21775 19499
rect 23949 19465 23983 19499
rect 2329 19329 2363 19363
rect 4721 19329 4755 19363
rect 5917 19329 5951 19363
rect 7573 19329 7607 19363
rect 9137 19329 9171 19363
rect 11529 19329 11563 19363
rect 16129 19329 16163 19363
rect 17325 19329 17359 19363
rect 2605 19261 2639 19295
rect 4353 19261 4387 19295
rect 6285 19261 6319 19295
rect 6837 19261 6871 19295
rect 9321 19261 9355 19295
rect 10793 19261 10827 19295
rect 12265 19261 12299 19295
rect 12817 19261 12851 19295
rect 12909 19261 12943 19295
rect 14197 19261 14231 19295
rect 14289 19261 14323 19295
rect 14749 19261 14783 19295
rect 16681 19261 16715 19295
rect 16957 19261 16991 19295
rect 17141 19261 17175 19295
rect 17233 19261 17267 19295
rect 2237 19193 2271 19227
rect 5181 19193 5215 19227
rect 5457 19193 5491 19227
rect 5549 19193 5583 19227
rect 7205 19193 7239 19227
rect 8309 19193 8343 19227
rect 9505 19193 9539 19227
rect 9873 19193 9907 19227
rect 11161 19193 11195 19227
rect 11897 19193 11931 19227
rect 12725 19193 12759 19227
rect 15025 19193 15059 19227
rect 17325 19193 17359 19227
rect 5089 19125 5123 19159
rect 5365 19125 5399 19159
rect 6653 19125 6687 19159
rect 7021 19125 7055 19159
rect 7113 19125 7147 19159
rect 8585 19125 8619 19159
rect 9413 19125 9447 19159
rect 10701 19125 10735 19159
rect 10977 19125 11011 19159
rect 11069 19125 11103 19159
rect 13829 19125 13863 19159
rect 15485 19125 15519 19159
rect 16037 19125 16071 19159
rect 17233 19125 17267 19159
rect 23489 19397 23523 19431
rect 24501 19397 24535 19431
rect 26157 19397 26191 19431
rect 17785 19329 17819 19363
rect 19717 19329 19751 19363
rect 26801 19329 26835 19363
rect 30297 19329 30331 19363
rect 32045 19329 32079 19363
rect 32965 19329 32999 19363
rect 19993 19261 20027 19295
rect 24317 19261 24351 19295
rect 25145 19261 25179 19295
rect 25329 19261 25363 19295
rect 25697 19261 25731 19295
rect 26157 19261 26191 19295
rect 27169 19261 27203 19295
rect 27537 19261 27571 19295
rect 28089 19261 28123 19295
rect 28273 19261 28307 19295
rect 29285 19261 29319 19295
rect 29561 19261 29595 19295
rect 31033 19261 31067 19295
rect 31585 19261 31619 19295
rect 31861 19261 31895 19295
rect 33517 19261 33551 19295
rect 33793 19261 33827 19295
rect 33977 19261 34011 19295
rect 34253 19261 34287 19295
rect 35449 19261 35483 19295
rect 19625 19193 19659 19227
rect 21373 19193 21407 19227
rect 24869 19193 24903 19227
rect 29101 19193 29135 19227
rect 29481 19193 29515 19227
rect 30021 19193 30055 19227
rect 34621 19193 34655 19227
rect 35817 19193 35851 19227
rect 17601 19125 17635 19159
rect 18245 19125 18279 19159
rect 18613 19125 18647 19159
rect 22109 19125 22143 19159
rect 22477 19125 22511 19159
rect 23121 19125 23155 19159
rect 27353 19125 27387 19159
rect 28641 19125 28675 19159
rect 30941 19125 30975 19159
rect 32505 19125 32539 19159
rect 32781 19125 32815 19159
rect 35081 19125 35115 19159
rect 3525 18921 3559 18955
rect 4905 18921 4939 18955
rect 6193 18921 6227 18955
rect 6469 18921 6503 18955
rect 6837 18921 6871 18955
rect 8769 18921 8803 18955
rect 11713 18921 11747 18955
rect 13461 18921 13495 18955
rect 14657 18921 14691 18955
rect 16221 18921 16255 18955
rect 17233 18921 17267 18955
rect 18521 18921 18555 18955
rect 18889 18921 18923 18955
rect 22569 18921 22603 18955
rect 24501 18921 24535 18955
rect 25053 18921 25087 18955
rect 26985 18921 27019 18955
rect 28273 18921 28307 18955
rect 30021 18921 30055 18955
rect 30297 18921 30331 18955
rect 31401 18921 31435 18955
rect 32873 18921 32907 18955
rect 5181 18853 5215 18887
rect 7849 18853 7883 18887
rect 10333 18853 10367 18887
rect 10425 18853 10459 18887
rect 10793 18853 10827 18887
rect 15945 18853 15979 18887
rect 23029 18853 23063 18887
rect 25973 18853 26007 18887
rect 27813 18853 27847 18887
rect 29377 18853 29411 18887
rect 34069 18853 34103 18887
rect 1685 18785 1719 18819
rect 5641 18785 5675 18819
rect 6653 18785 6687 18819
rect 7665 18785 7699 18819
rect 7941 18785 7975 18819
rect 10241 18785 10275 18819
rect 12265 18785 12299 18819
rect 12449 18785 12483 18819
rect 12817 18785 12851 18819
rect 14197 18785 14231 18819
rect 16129 18785 16163 18819
rect 17325 18785 17359 18819
rect 17417 18785 17451 18819
rect 18705 18785 18739 18819
rect 23673 18785 23707 18819
rect 24041 18785 24075 18819
rect 25145 18785 25179 18819
rect 26801 18785 26835 18819
rect 28181 18785 28215 18819
rect 29009 18785 29043 18819
rect 1409 18717 1443 18751
rect 10057 18717 10091 18751
rect 23305 18717 23339 18751
rect 29101 18717 29135 18751
rect 4445 18649 4479 18683
rect 5825 18649 5859 18683
rect 9873 18649 9907 18683
rect 12817 18649 12851 18683
rect 15025 18649 15059 18683
rect 16865 18649 16899 18683
rect 23949 18649 23983 18683
rect 25329 18649 25363 18683
rect 25697 18649 25731 18683
rect 33517 18785 33551 18819
rect 33793 18785 33827 18819
rect 33057 18717 33091 18751
rect 2789 18581 2823 18615
rect 3801 18581 3835 18615
rect 7297 18581 7331 18615
rect 8125 18581 8159 18615
rect 9137 18581 9171 18615
rect 11161 18581 11195 18615
rect 13737 18581 13771 18615
rect 14381 18581 14415 18615
rect 15577 18581 15611 18615
rect 17601 18581 17635 18615
rect 18245 18581 18279 18615
rect 19717 18581 19751 18615
rect 27445 18581 27479 18615
rect 29377 18581 29411 18615
rect 29653 18581 29687 18615
rect 30665 18581 30699 18615
rect 31033 18581 31067 18615
rect 1685 18377 1719 18411
rect 1961 18377 1995 18411
rect 4169 18377 4203 18411
rect 4905 18377 4939 18411
rect 5273 18377 5307 18411
rect 5641 18377 5675 18411
rect 5917 18377 5951 18411
rect 8677 18377 8711 18411
rect 10701 18377 10735 18411
rect 15669 18377 15703 18411
rect 23213 18377 23247 18411
rect 23949 18377 23983 18411
rect 24317 18377 24351 18411
rect 28733 18377 28767 18411
rect 29837 18377 29871 18411
rect 13185 18309 13219 18343
rect 16405 18309 16439 18343
rect 19073 18309 19107 18343
rect 22293 18309 22327 18343
rect 32045 18309 32079 18343
rect 32689 18309 32723 18343
rect 33701 18309 33735 18343
rect 7113 18241 7147 18275
rect 8493 18241 8527 18275
rect 8861 18241 8895 18275
rect 9597 18241 9631 18275
rect 11345 18241 11379 18275
rect 12081 18241 12115 18275
rect 16589 18241 16623 18275
rect 19717 18241 19751 18275
rect 25973 18241 26007 18275
rect 28089 18241 28123 18275
rect 30113 18241 30147 18275
rect 31125 18241 31159 18275
rect 31401 18241 31435 18275
rect 5733 18173 5767 18207
rect 6653 18173 6687 18207
rect 7205 18173 7239 18207
rect 7389 18173 7423 18207
rect 9137 18173 9171 18207
rect 10425 18173 10459 18207
rect 10517 18173 10551 18207
rect 11621 18173 11655 18207
rect 13553 18173 13587 18207
rect 13921 18173 13955 18207
rect 14105 18173 14139 18207
rect 14749 18173 14783 18207
rect 14841 18173 14875 18207
rect 16681 18173 16715 18207
rect 17601 18173 17635 18207
rect 17785 18173 17819 18207
rect 18153 18173 18187 18207
rect 19993 18173 20027 18207
rect 22385 18173 22419 18207
rect 24133 18173 24167 18207
rect 25053 18173 25087 18207
rect 25145 18173 25179 18207
rect 25697 18173 25731 18207
rect 26065 18173 26099 18207
rect 27353 18173 27387 18207
rect 28365 18173 28399 18207
rect 29285 18173 29319 18207
rect 31585 18173 31619 18207
rect 32045 18173 32079 18207
rect 7573 18105 7607 18139
rect 7941 18105 7975 18139
rect 8401 18105 8435 18139
rect 8493 18105 8527 18139
rect 9229 18105 9263 18139
rect 10149 18105 10183 18139
rect 13277 18105 13311 18139
rect 17141 18105 17175 18139
rect 17509 18105 17543 18139
rect 18061 18105 18095 18139
rect 21373 18105 21407 18139
rect 27261 18105 27295 18139
rect 27721 18105 27755 18139
rect 30757 18105 30791 18139
rect 33057 18105 33091 18139
rect 4537 18037 4571 18071
rect 6193 18037 6227 18071
rect 7481 18037 7515 18071
rect 9045 18037 9079 18071
rect 12817 18037 12851 18071
rect 16037 18037 16071 18071
rect 17601 18037 17635 18071
rect 19533 18037 19567 18071
rect 22569 18037 22603 18071
rect 24685 18037 24719 18071
rect 26893 18037 26927 18071
rect 27537 18037 27571 18071
rect 27629 18037 27663 18071
rect 29469 18037 29503 18071
rect 33333 18037 33367 18071
rect 1869 17833 1903 17867
rect 4629 17833 4663 17867
rect 5181 17833 5215 17867
rect 7205 17833 7239 17867
rect 7665 17833 7699 17867
rect 8677 17833 8711 17867
rect 11529 17833 11563 17867
rect 12357 17833 12391 17867
rect 12725 17833 12759 17867
rect 15485 17833 15519 17867
rect 18061 17833 18095 17867
rect 18429 17833 18463 17867
rect 20637 17833 20671 17867
rect 21557 17833 21591 17867
rect 23949 17833 23983 17867
rect 26709 17833 26743 17867
rect 30849 17833 30883 17867
rect 1961 17765 1995 17799
rect 4997 17765 5031 17799
rect 10701 17765 10735 17799
rect 11621 17765 11655 17799
rect 11989 17765 12023 17799
rect 13645 17765 13679 17799
rect 22569 17765 22603 17799
rect 24409 17765 24443 17799
rect 30389 17765 30423 17799
rect 2421 17697 2455 17731
rect 2605 17697 2639 17731
rect 2973 17697 3007 17731
rect 5365 17697 5399 17731
rect 5549 17697 5583 17731
rect 5917 17697 5951 17731
rect 7021 17697 7055 17731
rect 8033 17697 8067 17731
rect 9505 17697 9539 17731
rect 9689 17697 9723 17731
rect 9965 17697 9999 17731
rect 11253 17697 11287 17731
rect 11437 17697 11471 17731
rect 13185 17697 13219 17731
rect 16129 17697 16163 17731
rect 16497 17697 16531 17731
rect 16681 17697 16715 17731
rect 17325 17697 17359 17731
rect 17785 17697 17819 17731
rect 19441 17697 19475 17731
rect 22109 17697 22143 17731
rect 23121 17697 23155 17731
rect 23397 17697 23431 17731
rect 23581 17697 23615 17731
rect 25237 17697 25271 17731
rect 26525 17697 26559 17731
rect 27997 17697 28031 17731
rect 28181 17697 28215 17731
rect 28273 17697 28307 17731
rect 29561 17697 29595 17731
rect 30665 17697 30699 17731
rect 32413 17697 32447 17731
rect 32873 17697 32907 17731
rect 33333 17697 33367 17731
rect 34529 17697 34563 17731
rect 34805 17697 34839 17731
rect 35265 17697 35299 17731
rect 35541 17697 35575 17731
rect 2881 17629 2915 17663
rect 6469 17629 6503 17663
rect 8401 17629 8435 17663
rect 10425 17629 10459 17663
rect 13093 17629 13127 17663
rect 14657 17629 14691 17663
rect 15853 17629 15887 17663
rect 18797 17629 18831 17663
rect 24961 17629 24995 17663
rect 25421 17629 25455 17663
rect 27445 17629 27479 17663
rect 30021 17629 30055 17663
rect 32689 17629 32723 17663
rect 33609 17629 33643 17663
rect 8309 17561 8343 17595
rect 9781 17561 9815 17595
rect 11161 17561 11195 17595
rect 22477 17561 22511 17595
rect 24225 17561 24259 17595
rect 26341 17561 26375 17595
rect 3893 17493 3927 17527
rect 6929 17493 6963 17527
rect 8171 17493 8205 17527
rect 9045 17493 9079 17527
rect 14289 17493 14323 17527
rect 15025 17493 15059 17527
rect 19901 17493 19935 17527
rect 20177 17493 20211 17527
rect 25973 17493 26007 17527
rect 27077 17493 27111 17527
rect 27721 17493 27755 17527
rect 28457 17493 28491 17527
rect 29377 17493 29411 17527
rect 29745 17493 29779 17527
rect 31217 17493 31251 17527
rect 31585 17493 31619 17527
rect 2053 17289 2087 17323
rect 3525 17289 3559 17323
rect 4445 17289 4479 17323
rect 5641 17289 5675 17323
rect 8125 17289 8159 17323
rect 8769 17289 8803 17323
rect 9137 17289 9171 17323
rect 12725 17289 12759 17323
rect 14197 17289 14231 17323
rect 15301 17289 15335 17323
rect 16681 17289 16715 17323
rect 17601 17289 17635 17323
rect 18245 17289 18279 17323
rect 18889 17289 18923 17323
rect 20269 17289 20303 17323
rect 22937 17289 22971 17323
rect 26157 17289 26191 17323
rect 26525 17289 26559 17323
rect 28641 17289 28675 17323
rect 30297 17289 30331 17323
rect 30665 17289 30699 17323
rect 32597 17289 32631 17323
rect 35081 17289 35115 17323
rect 5181 17221 5215 17255
rect 16313 17221 16347 17255
rect 19257 17221 19291 17255
rect 19901 17221 19935 17255
rect 22293 17221 22327 17255
rect 25789 17221 25823 17255
rect 26019 17221 26053 17255
rect 2421 17153 2455 17187
rect 5365 17153 5399 17187
rect 6285 17153 6319 17187
rect 7021 17153 7055 17187
rect 9505 17153 9539 17187
rect 16405 17153 16439 17187
rect 26249 17153 26283 17187
rect 28365 17153 28399 17187
rect 30021 17153 30055 17187
rect 31125 17153 31159 17187
rect 33977 17153 34011 17187
rect 34621 17153 34655 17187
rect 2145 17085 2179 17119
rect 5457 17085 5491 17119
rect 7205 17085 7239 17119
rect 8585 17085 8619 17119
rect 9689 17085 9723 17119
rect 10241 17085 10275 17119
rect 10517 17085 10551 17119
rect 12449 17085 12483 17119
rect 12582 17085 12616 17119
rect 14013 17085 14047 17119
rect 14289 17085 14323 17119
rect 14841 17085 14875 17119
rect 15025 17085 15059 17119
rect 15117 17085 15151 17119
rect 15669 17085 15703 17119
rect 16497 17085 16531 17119
rect 18061 17085 18095 17119
rect 19073 17085 19107 17119
rect 20085 17085 20119 17119
rect 20545 17085 20579 17119
rect 21465 17085 21499 17119
rect 21925 17085 21959 17119
rect 22293 17085 22327 17119
rect 24225 17085 24259 17119
rect 25881 17085 25915 17119
rect 27905 17085 27939 17119
rect 29561 17085 29595 17119
rect 31677 17085 31711 17119
rect 31953 17085 31987 17119
rect 32137 17085 32171 17119
rect 33517 17085 33551 17119
rect 33793 17085 33827 17119
rect 1685 17017 1719 17051
rect 4813 17017 4847 17051
rect 7297 17017 7331 17051
rect 7389 17017 7423 17051
rect 7757 17017 7791 17051
rect 8493 17017 8527 17051
rect 12265 17017 12299 17051
rect 13369 17017 13403 17051
rect 19533 17017 19567 17051
rect 21005 17017 21039 17051
rect 27629 17017 27663 17051
rect 27997 17017 28031 17051
rect 29101 17017 29135 17051
rect 29285 17017 29319 17051
rect 29653 17017 29687 17051
rect 32965 17017 32999 17051
rect 34253 17017 34287 17051
rect 6653 16949 6687 16983
rect 9781 16949 9815 16983
rect 11345 16949 11379 16983
rect 11621 16949 11655 16983
rect 13645 16949 13679 16983
rect 14289 16949 14323 16983
rect 14565 16949 14599 16983
rect 15669 16949 15703 16983
rect 15945 16949 15979 16983
rect 17233 16949 17267 16983
rect 18521 16949 18555 16983
rect 21373 16949 21407 16983
rect 23213 16949 23247 16983
rect 24133 16949 24167 16983
rect 24409 16949 24443 16983
rect 24869 16949 24903 16983
rect 25329 16949 25363 16983
rect 26893 16949 26927 16983
rect 27537 16949 27571 16983
rect 27813 16949 27847 16983
rect 29469 16949 29503 16983
rect 1685 16745 1719 16779
rect 2053 16745 2087 16779
rect 2421 16745 2455 16779
rect 2697 16745 2731 16779
rect 3157 16745 3191 16779
rect 3525 16745 3559 16779
rect 4445 16745 4479 16779
rect 6837 16745 6871 16779
rect 7113 16745 7147 16779
rect 9413 16745 9447 16779
rect 9965 16745 9999 16779
rect 11805 16745 11839 16779
rect 13369 16745 13403 16779
rect 14105 16745 14139 16779
rect 14749 16745 14783 16779
rect 16037 16745 16071 16779
rect 16497 16745 16531 16779
rect 18429 16745 18463 16779
rect 20729 16745 20763 16779
rect 25421 16745 25455 16779
rect 26341 16745 26375 16779
rect 27721 16745 27755 16779
rect 29837 16745 29871 16779
rect 31309 16745 31343 16779
rect 31585 16745 31619 16779
rect 32873 16745 32907 16779
rect 34805 16745 34839 16779
rect 6193 16677 6227 16711
rect 6561 16677 6595 16711
rect 7481 16677 7515 16711
rect 7757 16677 7791 16711
rect 8033 16677 8067 16711
rect 8125 16677 8159 16711
rect 10241 16677 10275 16711
rect 11161 16677 11195 16711
rect 13093 16677 13127 16711
rect 17141 16677 17175 16711
rect 19441 16677 19475 16711
rect 19809 16677 19843 16711
rect 20361 16677 20395 16711
rect 22937 16677 22971 16711
rect 26525 16677 26559 16711
rect 27261 16677 27295 16711
rect 29193 16677 29227 16711
rect 30297 16677 30331 16711
rect 34529 16677 34563 16711
rect 3893 16609 3927 16643
rect 4905 16609 4939 16643
rect 4997 16609 5031 16643
rect 5181 16609 5215 16643
rect 5365 16609 5399 16643
rect 5641 16609 5675 16643
rect 6653 16609 6687 16643
rect 7941 16609 7975 16643
rect 8493 16609 8527 16643
rect 9781 16609 9815 16643
rect 10977 16609 11011 16643
rect 11069 16609 11103 16643
rect 12265 16609 12299 16643
rect 12541 16609 12575 16643
rect 12633 16609 12667 16643
rect 13737 16609 13771 16643
rect 13921 16609 13955 16643
rect 14381 16609 14415 16643
rect 15577 16609 15611 16643
rect 16681 16609 16715 16643
rect 17417 16609 17451 16643
rect 18613 16609 18647 16643
rect 18797 16609 18831 16643
rect 21557 16609 21591 16643
rect 21925 16609 21959 16643
rect 22385 16609 22419 16643
rect 22753 16609 22787 16643
rect 23765 16609 23799 16643
rect 24317 16609 24351 16643
rect 24777 16609 24811 16643
rect 29009 16609 29043 16643
rect 29101 16609 29135 16643
rect 30573 16609 30607 16643
rect 30757 16609 30791 16643
rect 32413 16609 32447 16643
rect 33517 16609 33551 16643
rect 33793 16609 33827 16643
rect 10793 16541 10827 16575
rect 11529 16541 11563 16575
rect 16589 16541 16623 16575
rect 19165 16541 19199 16575
rect 21373 16541 21407 16575
rect 21833 16541 21867 16575
rect 23489 16541 23523 16575
rect 23949 16541 23983 16575
rect 25145 16541 25179 16575
rect 26893 16541 26927 16575
rect 28825 16541 28859 16575
rect 29561 16541 29595 16575
rect 33057 16541 33091 16575
rect 34069 16541 34103 16575
rect 12357 16473 12391 16507
rect 26801 16473 26835 16507
rect 9045 16405 9079 16439
rect 10609 16405 10643 16439
rect 15761 16405 15795 16439
rect 18061 16405 18095 16439
rect 21189 16405 21223 16439
rect 24685 16405 24719 16439
rect 24915 16405 24949 16439
rect 25053 16405 25087 16439
rect 25881 16405 25915 16439
rect 26663 16405 26697 16439
rect 28089 16405 28123 16439
rect 28641 16405 28675 16439
rect 30941 16405 30975 16439
rect 3525 16201 3559 16235
rect 4813 16201 4847 16235
rect 6285 16201 6319 16235
rect 6653 16201 6687 16235
rect 8309 16201 8343 16235
rect 10977 16201 11011 16235
rect 11253 16201 11287 16235
rect 14289 16201 14323 16235
rect 16681 16201 16715 16235
rect 17049 16201 17083 16235
rect 19901 16201 19935 16235
rect 21373 16201 21407 16235
rect 23029 16201 23063 16235
rect 25237 16201 25271 16235
rect 26617 16201 26651 16235
rect 28641 16201 28675 16235
rect 29101 16201 29135 16235
rect 30849 16201 30883 16235
rect 33977 16201 34011 16235
rect 4629 16133 4663 16167
rect 7941 16133 7975 16167
rect 13553 16133 13587 16167
rect 16221 16133 16255 16167
rect 17417 16133 17451 16167
rect 22385 16133 22419 16167
rect 25053 16133 25087 16167
rect 26506 16133 26540 16167
rect 26801 16133 26835 16167
rect 30573 16133 30607 16167
rect 1409 16065 1443 16099
rect 1685 16065 1719 16099
rect 3893 16065 3927 16099
rect 5273 16065 5307 16099
rect 7573 16065 7607 16099
rect 10241 16065 10275 16099
rect 21005 16065 21039 16099
rect 21741 16065 21775 16099
rect 24685 16065 24719 16099
rect 25145 16065 25179 16099
rect 25789 16065 25823 16099
rect 26709 16065 26743 16099
rect 30205 16065 30239 16099
rect 32229 16065 32263 16099
rect 5365 15997 5399 16031
rect 5733 15997 5767 16031
rect 5917 15997 5951 16031
rect 6837 15997 6871 16031
rect 7113 15997 7147 16031
rect 8677 15997 8711 16031
rect 8861 15997 8895 16031
rect 9229 15997 9263 16031
rect 9781 15997 9815 16031
rect 10149 15997 10183 16031
rect 11069 15997 11103 16031
rect 11345 15997 11379 16031
rect 12633 15997 12667 16031
rect 13921 15997 13955 16031
rect 14013 15997 14047 16031
rect 14197 15997 14231 16031
rect 16037 15997 16071 16031
rect 18337 15997 18371 16031
rect 19625 15997 19659 16031
rect 19717 15997 19751 16031
rect 21925 15997 21959 16031
rect 22477 15997 22511 16031
rect 23673 15997 23707 16031
rect 24924 15997 24958 16031
rect 27353 15997 27387 16031
rect 28181 15997 28215 16031
rect 29745 15997 29779 16031
rect 30297 15997 30331 16031
rect 31861 15997 31895 16031
rect 32873 15997 32907 16031
rect 33149 15997 33183 16031
rect 33333 15997 33367 16031
rect 34897 15997 34931 16031
rect 35357 15997 35391 16031
rect 3065 15929 3099 15963
rect 4261 15929 4295 15963
rect 7205 15929 7239 15963
rect 12173 15929 12207 15963
rect 12449 15929 12483 15963
rect 12817 15929 12851 15963
rect 13185 15929 13219 15963
rect 15669 15929 15703 15963
rect 18061 15929 18095 15963
rect 18429 15929 18463 15963
rect 18797 15929 18831 15963
rect 24777 15929 24811 15963
rect 26341 15929 26375 15963
rect 31217 15929 31251 15963
rect 32321 15929 32355 15963
rect 33609 15929 33643 15963
rect 7021 15861 7055 15895
rect 10609 15861 10643 15895
rect 11345 15861 11379 15895
rect 11621 15861 11655 15895
rect 12725 15861 12759 15895
rect 14841 15861 14875 15895
rect 15209 15861 15243 15895
rect 17785 15861 17819 15895
rect 18245 15861 18279 15895
rect 19073 15861 19107 15895
rect 19533 15861 19567 15895
rect 20453 15861 20487 15895
rect 23489 15861 23523 15895
rect 23857 15861 23891 15895
rect 24317 15861 24351 15895
rect 26249 15861 26283 15895
rect 28089 15861 28123 15895
rect 28365 15861 28399 15895
rect 35081 15861 35115 15895
rect 1685 15657 1719 15691
rect 4445 15657 4479 15691
rect 5457 15657 5491 15691
rect 7389 15657 7423 15691
rect 7849 15657 7883 15691
rect 8585 15657 8619 15691
rect 10793 15657 10827 15691
rect 13001 15657 13035 15691
rect 16129 15657 16163 15691
rect 16681 15657 16715 15691
rect 18705 15657 18739 15691
rect 19165 15657 19199 15691
rect 20361 15657 20395 15691
rect 20729 15657 20763 15691
rect 22017 15657 22051 15691
rect 22385 15657 22419 15691
rect 23029 15657 23063 15691
rect 24869 15657 24903 15691
rect 26249 15657 26283 15691
rect 27169 15657 27203 15691
rect 27905 15657 27939 15691
rect 28549 15657 28583 15691
rect 31217 15657 31251 15691
rect 32229 15657 32263 15691
rect 33241 15657 33275 15691
rect 5641 15589 5675 15623
rect 11253 15589 11287 15623
rect 11621 15589 11655 15623
rect 12541 15589 12575 15623
rect 16497 15589 16531 15623
rect 16865 15589 16899 15623
rect 19257 15589 19291 15623
rect 21097 15589 21131 15623
rect 22661 15589 22695 15623
rect 23397 15589 23431 15623
rect 23857 15589 23891 15623
rect 25973 15589 26007 15623
rect 26525 15589 26559 15623
rect 28641 15589 28675 15623
rect 29009 15589 29043 15623
rect 29377 15589 29411 15623
rect 30205 15589 30239 15623
rect 4629 15521 4663 15555
rect 6101 15521 6135 15555
rect 6285 15521 6319 15555
rect 6469 15521 6503 15555
rect 7113 15521 7147 15555
rect 7941 15521 7975 15555
rect 9689 15521 9723 15555
rect 11069 15521 11103 15555
rect 11161 15521 11195 15555
rect 13185 15521 13219 15555
rect 13645 15521 13679 15555
rect 13737 15521 13771 15555
rect 14289 15521 14323 15555
rect 15301 15521 15335 15555
rect 16773 15521 16807 15555
rect 19073 15521 19107 15555
rect 21833 15521 21867 15555
rect 22845 15521 22879 15555
rect 24004 15521 24038 15555
rect 25421 15521 25455 15555
rect 26672 15521 26706 15555
rect 28457 15521 28491 15555
rect 30021 15521 30055 15555
rect 30113 15521 30147 15555
rect 32137 15521 32171 15555
rect 32597 15521 32631 15555
rect 34437 15521 34471 15555
rect 34805 15521 34839 15555
rect 3525 15453 3559 15487
rect 6745 15453 6779 15487
rect 8309 15453 8343 15487
rect 10885 15453 10919 15487
rect 17233 15453 17267 15487
rect 18889 15453 18923 15487
rect 19625 15453 19659 15487
rect 24225 15453 24259 15487
rect 25329 15453 25363 15487
rect 26893 15453 26927 15487
rect 28273 15453 28307 15487
rect 29837 15453 29871 15487
rect 30573 15453 30607 15487
rect 30849 15453 30883 15487
rect 34161 15453 34195 15487
rect 3157 15385 3191 15419
rect 4813 15385 4847 15419
rect 8217 15385 8251 15419
rect 9873 15385 9907 15419
rect 15485 15385 15519 15419
rect 17785 15385 17819 15419
rect 21741 15385 21775 15419
rect 24317 15385 24351 15419
rect 25605 15385 25639 15419
rect 34805 15385 34839 15419
rect 3893 15317 3927 15351
rect 5181 15317 5215 15351
rect 8079 15317 8113 15351
rect 8953 15317 8987 15351
rect 9321 15317 9355 15351
rect 10241 15317 10275 15351
rect 12173 15317 12207 15351
rect 14749 15317 14783 15351
rect 15117 15317 15151 15351
rect 18061 15317 18095 15351
rect 19901 15317 19935 15351
rect 23765 15317 23799 15351
rect 24133 15317 24167 15351
rect 26801 15317 26835 15351
rect 27629 15317 27663 15351
rect 29745 15317 29779 15351
rect 2973 15113 3007 15147
rect 5733 15113 5767 15147
rect 8493 15113 8527 15147
rect 10958 15113 10992 15147
rect 11069 15113 11103 15147
rect 11805 15113 11839 15147
rect 13461 15113 13495 15147
rect 13829 15113 13863 15147
rect 14381 15113 14415 15147
rect 16589 15113 16623 15147
rect 17601 15113 17635 15147
rect 18613 15113 18647 15147
rect 21189 15113 21223 15147
rect 23121 15113 23155 15147
rect 23489 15113 23523 15147
rect 24317 15113 24351 15147
rect 24501 15113 24535 15147
rect 26111 15113 26145 15147
rect 27353 15113 27387 15147
rect 28273 15113 28307 15147
rect 28641 15113 28675 15147
rect 29469 15113 29503 15147
rect 30757 15113 30791 15147
rect 31953 15113 31987 15147
rect 32413 15113 32447 15147
rect 33793 15113 33827 15147
rect 34253 15113 34287 15147
rect 34621 15113 34655 15147
rect 7665 15045 7699 15079
rect 9965 15045 9999 15079
rect 11253 15045 11287 15079
rect 22477 15045 22511 15079
rect 26249 15045 26283 15079
rect 26985 15045 27019 15079
rect 27721 15045 27755 15079
rect 35081 15045 35115 15079
rect 1409 14977 1443 15011
rect 1685 14977 1719 15011
rect 7757 14977 7791 15011
rect 7849 14977 7883 15011
rect 8861 14977 8895 15011
rect 11161 14977 11195 15011
rect 12081 14977 12115 15011
rect 12449 14977 12483 15011
rect 13185 14977 13219 15011
rect 14565 14977 14599 15011
rect 18484 14977 18518 15011
rect 18705 14977 18739 15011
rect 19073 14977 19107 15011
rect 24409 14977 24443 15011
rect 26341 14977 26375 15011
rect 30573 14977 30607 15011
rect 33057 14977 33091 15011
rect 3801 14909 3835 14943
rect 4353 14909 4387 14943
rect 4537 14909 4571 14943
rect 4905 14909 4939 14943
rect 5089 14909 5123 14943
rect 7536 14909 7570 14943
rect 9689 14909 9723 14943
rect 10793 14909 10827 14943
rect 11621 14909 11655 14943
rect 7389 14841 7423 14875
rect 8953 14841 8987 14875
rect 9321 14841 9355 14875
rect 3433 14773 3467 14807
rect 3985 14773 4019 14807
rect 6009 14773 6043 14807
rect 6469 14773 6503 14807
rect 7205 14773 7239 14807
rect 9137 14773 9171 14807
rect 9229 14773 9263 14807
rect 10701 14773 10735 14807
rect 11621 14773 11655 14807
rect 12725 14909 12759 14943
rect 14473 14909 14507 14943
rect 15209 14909 15243 14943
rect 15301 14909 15335 14943
rect 15669 14909 15703 14943
rect 16773 14909 16807 14943
rect 17233 14909 17267 14943
rect 18337 14909 18371 14943
rect 19717 14909 19751 14943
rect 20177 14909 20211 14943
rect 21649 14909 21683 14943
rect 22201 14909 22235 14943
rect 22569 14909 22603 14943
rect 24041 14909 24075 14943
rect 24188 14909 24222 14943
rect 25145 14909 25179 14943
rect 25973 14909 26007 14943
rect 27537 14909 27571 14943
rect 29929 14909 29963 14943
rect 30481 14909 30515 14943
rect 31033 14909 31067 14943
rect 33333 14909 33367 14943
rect 33517 14909 33551 14943
rect 12817 14841 12851 14875
rect 19901 14841 19935 14875
rect 26709 14841 26743 14875
rect 31401 14841 31435 14875
rect 32505 14841 32539 14875
rect 12081 14773 12115 14807
rect 12173 14773 12207 14807
rect 12633 14773 12667 14807
rect 16957 14773 16991 14807
rect 19349 14773 19383 14807
rect 21557 14773 21591 14807
rect 23949 14773 23983 14807
rect 25513 14773 25547 14807
rect 25881 14773 25915 14807
rect 29009 14773 29043 14807
rect 1961 14569 1995 14603
rect 3525 14569 3559 14603
rect 3893 14569 3927 14603
rect 4353 14569 4387 14603
rect 5365 14569 5399 14603
rect 6101 14569 6135 14603
rect 7481 14569 7515 14603
rect 10977 14569 11011 14603
rect 11713 14569 11747 14603
rect 13369 14569 13403 14603
rect 14197 14569 14231 14603
rect 17509 14569 17543 14603
rect 17785 14569 17819 14603
rect 18705 14569 18739 14603
rect 19073 14569 19107 14603
rect 20545 14569 20579 14603
rect 21649 14569 21683 14603
rect 22109 14569 22143 14603
rect 22753 14569 22787 14603
rect 26985 14569 27019 14603
rect 27353 14569 27387 14603
rect 27905 14569 27939 14603
rect 29929 14569 29963 14603
rect 30389 14569 30423 14603
rect 32321 14569 32355 14603
rect 33057 14569 33091 14603
rect 3157 14501 3191 14535
rect 7113 14501 7147 14535
rect 8309 14501 8343 14535
rect 9965 14501 9999 14535
rect 10333 14501 10367 14535
rect 10701 14501 10735 14535
rect 13461 14501 13495 14535
rect 13829 14501 13863 14535
rect 15577 14501 15611 14535
rect 16313 14501 16347 14535
rect 16681 14501 16715 14535
rect 17877 14501 17911 14535
rect 17969 14501 18003 14535
rect 18337 14501 18371 14535
rect 19533 14501 19567 14535
rect 19901 14501 19935 14535
rect 26065 14501 26099 14535
rect 31493 14501 31527 14535
rect 4169 14433 4203 14467
rect 6469 14433 6503 14467
rect 7849 14433 7883 14467
rect 7941 14433 7975 14467
rect 8125 14433 8159 14467
rect 8217 14433 8251 14467
rect 10149 14433 10183 14467
rect 10241 14433 10275 14467
rect 11897 14433 11931 14467
rect 12909 14433 12943 14467
rect 13277 14433 13311 14467
rect 15117 14433 15151 14467
rect 16129 14433 16163 14467
rect 16221 14433 16255 14467
rect 19349 14433 19383 14467
rect 19441 14433 19475 14467
rect 20913 14433 20947 14467
rect 21925 14433 21959 14467
rect 22937 14433 22971 14467
rect 23949 14433 23983 14467
rect 24096 14433 24130 14467
rect 26525 14433 26559 14467
rect 28641 14433 28675 14467
rect 28733 14433 28767 14467
rect 30113 14433 30147 14467
rect 30941 14433 30975 14467
rect 31125 14433 31159 14467
rect 32137 14433 32171 14467
rect 33793 14433 33827 14467
rect 34253 14433 34287 14467
rect 8677 14365 8711 14399
rect 13093 14365 13127 14399
rect 15945 14365 15979 14399
rect 17601 14365 17635 14399
rect 19165 14365 19199 14399
rect 23489 14365 23523 14399
rect 24317 14365 24351 14399
rect 25697 14365 25731 14399
rect 29193 14365 29227 14399
rect 33609 14365 33643 14399
rect 4721 14297 4755 14331
rect 6653 14297 6687 14331
rect 9321 14297 9355 14331
rect 14473 14297 14507 14331
rect 20177 14297 20211 14331
rect 21097 14297 21131 14331
rect 22477 14297 22511 14331
rect 24409 14297 24443 14331
rect 28273 14297 28307 14331
rect 29469 14297 29503 14331
rect 34253 14297 34287 14331
rect 1593 14229 1627 14263
rect 5733 14229 5767 14263
rect 8953 14229 8987 14263
rect 11345 14229 11379 14263
rect 12081 14229 12115 14263
rect 12541 14229 12575 14263
rect 17049 14229 17083 14263
rect 23121 14229 23155 14263
rect 23857 14229 23891 14263
rect 24225 14229 24259 14263
rect 25329 14229 25363 14263
rect 26709 14229 26743 14263
rect 28457 14229 28491 14263
rect 31953 14229 31987 14263
rect 32597 14229 32631 14263
rect 2697 14025 2731 14059
rect 4629 14025 4663 14059
rect 5273 14025 5307 14059
rect 5641 14025 5675 14059
rect 7113 14025 7147 14059
rect 7757 14025 7791 14059
rect 9597 14025 9631 14059
rect 12265 14025 12299 14059
rect 15393 14025 15427 14059
rect 15945 14025 15979 14059
rect 16570 14025 16604 14059
rect 18429 14025 18463 14059
rect 18889 14025 18923 14059
rect 19257 14025 19291 14059
rect 19993 14025 20027 14059
rect 20361 14025 20395 14059
rect 21005 14025 21039 14059
rect 23121 14025 23155 14059
rect 24041 14025 24075 14059
rect 25513 14025 25547 14059
rect 26138 14025 26172 14059
rect 26617 14025 26651 14059
rect 26985 14025 27019 14059
rect 27721 14025 27755 14059
rect 28457 14025 28491 14059
rect 30665 14025 30699 14059
rect 32229 14025 32263 14059
rect 34529 14025 34563 14059
rect 5917 13957 5951 13991
rect 13277 13957 13311 13991
rect 16681 13957 16715 13991
rect 19146 13957 19180 13991
rect 22385 13957 22419 13991
rect 25881 13957 25915 13991
rect 26249 13957 26283 13991
rect 30297 13957 30331 13991
rect 3157 13889 3191 13923
rect 9229 13889 9263 13923
rect 10793 13889 10827 13923
rect 13185 13889 13219 13923
rect 3249 13821 3283 13855
rect 3525 13821 3559 13855
rect 5733 13821 5767 13855
rect 6285 13821 6319 13855
rect 6653 13821 6687 13855
rect 6837 13821 6871 13855
rect 6929 13821 6963 13855
rect 8401 13821 8435 13855
rect 8769 13821 8803 13855
rect 11805 13821 11839 13855
rect 12633 13821 12667 13855
rect 13645 13889 13679 13923
rect 14749 13889 14783 13923
rect 16773 13889 16807 13923
rect 16865 13889 16899 13923
rect 19349 13889 19383 13923
rect 26341 13889 26375 13923
rect 31493 13889 31527 13923
rect 34161 13889 34195 13923
rect 13921 13821 13955 13855
rect 15209 13821 15243 13855
rect 16405 13821 16439 13855
rect 18981 13821 19015 13855
rect 19717 13821 19751 13855
rect 20545 13821 20579 13855
rect 21649 13821 21683 13855
rect 21925 13821 21959 13855
rect 22477 13821 22511 13855
rect 24409 13821 24443 13855
rect 24501 13821 24535 13855
rect 25973 13821 26007 13855
rect 27445 13821 27479 13855
rect 27537 13821 27571 13855
rect 28181 13821 28215 13855
rect 29285 13821 29319 13855
rect 29469 13821 29503 13855
rect 29561 13821 29595 13855
rect 30941 13821 30975 13855
rect 31769 13821 31803 13855
rect 31953 13821 31987 13855
rect 32689 13821 32723 13855
rect 32781 13821 32815 13855
rect 33149 13821 33183 13855
rect 33609 13821 33643 13855
rect 33885 13821 33919 13855
rect 8493 13753 8527 13787
rect 8861 13753 8895 13787
rect 10057 13753 10091 13787
rect 10425 13753 10459 13787
rect 13277 13753 13311 13787
rect 13553 13753 13587 13787
rect 14013 13753 14047 13787
rect 14381 13753 14415 13787
rect 15117 13753 15151 13787
rect 29009 13753 29043 13787
rect 29653 13753 29687 13787
rect 30021 13753 30055 13787
rect 8677 13685 8711 13719
rect 9873 13685 9907 13719
rect 10241 13685 10275 13719
rect 10333 13685 10367 13719
rect 11161 13685 11195 13719
rect 11529 13685 11563 13719
rect 12817 13685 12851 13719
rect 13829 13685 13863 13719
rect 17693 13685 17727 13719
rect 20729 13685 20763 13719
rect 21465 13685 21499 13719
rect 23489 13685 23523 13719
rect 5273 13481 5307 13515
rect 5641 13481 5675 13515
rect 7481 13481 7515 13515
rect 8217 13481 8251 13515
rect 9505 13481 9539 13515
rect 10517 13481 10551 13515
rect 11069 13481 11103 13515
rect 13921 13481 13955 13515
rect 14381 13481 14415 13515
rect 14749 13481 14783 13515
rect 16497 13481 16531 13515
rect 18153 13481 18187 13515
rect 19073 13481 19107 13515
rect 19901 13481 19935 13515
rect 20729 13481 20763 13515
rect 21189 13481 21223 13515
rect 22845 13481 22879 13515
rect 23213 13481 23247 13515
rect 23397 13481 23431 13515
rect 23581 13481 23615 13515
rect 24685 13481 24719 13515
rect 25053 13481 25087 13515
rect 25421 13481 25455 13515
rect 25973 13481 26007 13515
rect 26709 13481 26743 13515
rect 27629 13481 27663 13515
rect 29285 13481 29319 13515
rect 30849 13481 30883 13515
rect 31585 13481 31619 13515
rect 32229 13481 32263 13515
rect 33149 13481 33183 13515
rect 33609 13481 33643 13515
rect 33885 13481 33919 13515
rect 3065 13413 3099 13447
rect 7021 13413 7055 13447
rect 8401 13413 8435 13447
rect 10885 13413 10919 13447
rect 11253 13413 11287 13447
rect 15945 13413 15979 13447
rect 16589 13413 16623 13447
rect 16681 13413 16715 13447
rect 18245 13413 18279 13447
rect 18613 13413 18647 13447
rect 28917 13413 28951 13447
rect 1409 13345 1443 13379
rect 5641 13345 5675 13379
rect 6193 13345 6227 13379
rect 6377 13345 6411 13379
rect 7941 13345 7975 13379
rect 8309 13345 8343 13379
rect 9689 13345 9723 13379
rect 11161 13345 11195 13379
rect 12725 13345 12759 13379
rect 12909 13345 12943 13379
rect 13277 13345 13311 13379
rect 15301 13345 15335 13379
rect 16313 13345 16347 13379
rect 17417 13345 17451 13379
rect 18061 13345 18095 13379
rect 19441 13345 19475 13379
rect 20269 13345 20303 13379
rect 21465 13345 21499 13379
rect 22385 13345 22419 13379
rect 22661 13345 22695 13379
rect 23397 13345 23431 13379
rect 23673 13345 23707 13379
rect 23820 13345 23854 13379
rect 25237 13345 25271 13379
rect 26525 13345 26559 13379
rect 26985 13345 27019 13379
rect 28365 13345 28399 13379
rect 28457 13345 28491 13379
rect 29745 13345 29779 13379
rect 30021 13345 30055 13379
rect 32413 13345 32447 13379
rect 32597 13345 32631 13379
rect 1685 13277 1719 13311
rect 8033 13277 8067 13311
rect 8769 13277 8803 13311
rect 11621 13277 11655 13311
rect 11897 13277 11931 13311
rect 17049 13277 17083 13311
rect 17877 13277 17911 13311
rect 4353 13209 4387 13243
rect 9137 13209 9171 13243
rect 13277 13209 13311 13243
rect 15485 13209 15519 13243
rect 19625 13209 19659 13243
rect 24041 13277 24075 13311
rect 28181 13277 28215 13311
rect 30481 13277 30515 13311
rect 31125 13277 31159 13311
rect 24133 13209 24167 13243
rect 27997 13209 28031 13243
rect 29837 13209 29871 13243
rect 4905 13141 4939 13175
rect 9873 13141 9907 13175
rect 10241 13141 10275 13175
rect 12265 13141 12299 13175
rect 15117 13141 15151 13175
rect 17693 13141 17727 13175
rect 22017 13141 22051 13175
rect 23397 13141 23431 13175
rect 23949 13141 23983 13175
rect 31861 13141 31895 13175
rect 1593 12937 1627 12971
rect 5089 12937 5123 12971
rect 8125 12937 8159 12971
rect 10701 12937 10735 12971
rect 10958 12937 10992 12971
rect 11805 12937 11839 12971
rect 12265 12937 12299 12971
rect 12909 12937 12943 12971
rect 16221 12937 16255 12971
rect 17325 12937 17359 12971
rect 18981 12937 19015 12971
rect 19717 12937 19751 12971
rect 20085 12937 20119 12971
rect 21097 12937 21131 12971
rect 23121 12937 23155 12971
rect 24133 12937 24167 12971
rect 25237 12937 25271 12971
rect 26230 12937 26264 12971
rect 27537 12937 27571 12971
rect 29009 12937 29043 12971
rect 30205 12937 30239 12971
rect 30573 12937 30607 12971
rect 32505 12937 32539 12971
rect 32873 12937 32907 12971
rect 5457 12869 5491 12903
rect 5825 12869 5859 12903
rect 9873 12869 9907 12903
rect 10333 12869 10367 12903
rect 11069 12869 11103 12903
rect 11253 12869 11287 12903
rect 13553 12869 13587 12903
rect 16083 12869 16117 12903
rect 22477 12869 22511 12903
rect 24022 12869 24056 12903
rect 24869 12869 24903 12903
rect 26341 12869 26375 12903
rect 31401 12869 31435 12903
rect 1961 12801 1995 12835
rect 6653 12801 6687 12835
rect 6929 12801 6963 12835
rect 11161 12801 11195 12835
rect 13921 12801 13955 12835
rect 16313 12801 16347 12835
rect 17785 12801 17819 12835
rect 19073 12801 19107 12835
rect 19349 12801 19383 12835
rect 24225 12801 24259 12835
rect 25973 12801 26007 12835
rect 26433 12801 26467 12835
rect 27629 12801 27663 12835
rect 28641 12801 28675 12835
rect 29929 12801 29963 12835
rect 31033 12801 31067 12835
rect 35725 12801 35759 12835
rect 37289 12801 37323 12835
rect 6285 12733 6319 12767
rect 7113 12733 7147 12767
rect 7665 12733 7699 12767
rect 8493 12733 8527 12767
rect 8953 12733 8987 12767
rect 9505 12733 9539 12767
rect 9781 12733 9815 12767
rect 10793 12733 10827 12767
rect 12449 12733 12483 12767
rect 13645 12733 13679 12767
rect 14013 12733 14047 12767
rect 14565 12733 14599 12767
rect 14933 12733 14967 12767
rect 15853 12733 15887 12767
rect 15945 12733 15979 12767
rect 17049 12733 17083 12767
rect 18705 12733 18739 12767
rect 18852 12733 18886 12767
rect 20453 12733 20487 12767
rect 21557 12733 21591 12767
rect 21833 12733 21867 12767
rect 22109 12733 22143 12767
rect 22569 12733 22603 12767
rect 23857 12733 23891 12767
rect 26065 12733 26099 12767
rect 27905 12733 27939 12767
rect 29561 12733 29595 12767
rect 31125 12733 31159 12767
rect 31677 12733 31711 12767
rect 31953 12733 31987 12767
rect 35817 12733 35851 12767
rect 36093 12733 36127 12767
rect 7297 12665 7331 12699
rect 20269 12665 20303 12699
rect 20821 12665 20855 12699
rect 26801 12665 26835 12699
rect 27169 12665 27203 12699
rect 27813 12665 27847 12699
rect 27997 12665 28031 12699
rect 28365 12665 28399 12699
rect 29377 12665 29411 12699
rect 7205 12597 7239 12631
rect 12633 12597 12667 12631
rect 15393 12597 15427 12631
rect 16589 12597 16623 12631
rect 18613 12597 18647 12631
rect 23397 12597 23431 12631
rect 24501 12597 24535 12631
rect 5273 12393 5307 12427
rect 5733 12393 5767 12427
rect 7757 12393 7791 12427
rect 8033 12393 8067 12427
rect 8677 12393 8711 12427
rect 9045 12393 9079 12427
rect 9873 12393 9907 12427
rect 11621 12393 11655 12427
rect 11897 12393 11931 12427
rect 12633 12393 12667 12427
rect 14381 12393 14415 12427
rect 14841 12393 14875 12427
rect 18153 12393 18187 12427
rect 18429 12393 18463 12427
rect 6377 12325 6411 12359
rect 10609 12325 10643 12359
rect 11253 12325 11287 12359
rect 13277 12325 13311 12359
rect 14105 12325 14139 12359
rect 1777 12257 1811 12291
rect 3157 12257 3191 12291
rect 4169 12257 4203 12291
rect 5917 12257 5951 12291
rect 6193 12257 6227 12291
rect 6837 12257 6871 12291
rect 7205 12257 7239 12291
rect 8217 12257 8251 12291
rect 9689 12257 9723 12291
rect 10793 12257 10827 12291
rect 12081 12257 12115 12291
rect 14197 12257 14231 12291
rect 15301 12257 15335 12291
rect 16589 12257 16623 12291
rect 17325 12257 17359 12291
rect 17693 12257 17727 12291
rect 19533 12393 19567 12427
rect 20269 12393 20303 12427
rect 21097 12393 21131 12427
rect 22109 12393 22143 12427
rect 22937 12393 22971 12427
rect 23581 12393 23615 12427
rect 24685 12393 24719 12427
rect 24777 12393 24811 12427
rect 26709 12393 26743 12427
rect 27721 12393 27755 12427
rect 28273 12393 28307 12427
rect 28825 12393 28859 12427
rect 29469 12393 29503 12427
rect 30481 12393 30515 12427
rect 30849 12393 30883 12427
rect 31217 12393 31251 12427
rect 21741 12325 21775 12359
rect 24317 12325 24351 12359
rect 19257 12257 19291 12291
rect 19533 12257 19567 12291
rect 20913 12257 20947 12291
rect 22385 12257 22419 12291
rect 23397 12257 23431 12291
rect 24777 12257 24811 12291
rect 24869 12257 24903 12291
rect 25605 12257 25639 12291
rect 27077 12257 27111 12291
rect 28641 12257 28675 12291
rect 29653 12257 29687 12291
rect 31033 12257 31067 12291
rect 32781 12257 32815 12291
rect 1501 12189 1535 12223
rect 7297 12189 7331 12223
rect 10701 12189 10735 12223
rect 16681 12189 16715 12223
rect 17141 12189 17175 12223
rect 17601 12189 17635 12223
rect 18429 12189 18463 12223
rect 18613 12189 18647 12223
rect 18705 12189 18739 12223
rect 25237 12189 25271 12223
rect 27445 12189 27479 12223
rect 4353 12121 4387 12155
rect 8401 12121 8435 12155
rect 10241 12121 10275 12155
rect 12265 12121 12299 12155
rect 13645 12121 13679 12155
rect 25145 12121 25179 12155
rect 29837 12121 29871 12155
rect 30205 12121 30239 12155
rect 4629 12053 4663 12087
rect 5641 12053 5675 12087
rect 9413 12053 9447 12087
rect 13001 12053 13035 12087
rect 15485 12053 15519 12087
rect 16037 12053 16071 12087
rect 16405 12053 16439 12087
rect 19717 12053 19751 12087
rect 20637 12053 20671 12087
rect 22569 12053 22603 12087
rect 23857 12053 23891 12087
rect 25034 12053 25068 12087
rect 26065 12053 26099 12087
rect 27215 12053 27249 12087
rect 27353 12053 27387 12087
rect 31493 12053 31527 12087
rect 32413 12053 32447 12087
rect 35817 12053 35851 12087
rect 6009 11849 6043 11883
rect 7297 11849 7331 11883
rect 8217 11849 8251 11883
rect 9597 11849 9631 11883
rect 11897 11849 11931 11883
rect 14289 11849 14323 11883
rect 16773 11849 16807 11883
rect 17509 11849 17543 11883
rect 19073 11849 19107 11883
rect 19533 11849 19567 11883
rect 20913 11849 20947 11883
rect 23489 11849 23523 11883
rect 24041 11849 24075 11883
rect 24961 11849 24995 11883
rect 27261 11849 27295 11883
rect 27721 11849 27755 11883
rect 27997 11849 28031 11883
rect 28641 11849 28675 11883
rect 29653 11849 29687 11883
rect 31953 11849 31987 11883
rect 32873 11849 32907 11883
rect 37381 11849 37415 11883
rect 5641 11781 5675 11815
rect 11529 11781 11563 11815
rect 14657 11781 14691 11815
rect 17141 11781 17175 11815
rect 23121 11781 23155 11815
rect 31125 11781 31159 11815
rect 3341 11713 3375 11747
rect 3709 11713 3743 11747
rect 8677 11713 8711 11747
rect 9229 11713 9263 11747
rect 12265 11713 12299 11747
rect 14749 11713 14783 11747
rect 19901 11713 19935 11747
rect 22569 11713 22603 11747
rect 26985 11713 27019 11747
rect 31677 11713 31711 11747
rect 32505 11713 32539 11747
rect 35725 11713 35759 11747
rect 3433 11645 3467 11679
rect 6653 11645 6687 11679
rect 7481 11645 7515 11679
rect 8769 11645 8803 11679
rect 9965 11645 9999 11679
rect 10701 11645 10735 11679
rect 12541 11645 12575 11679
rect 13093 11645 13127 11679
rect 13277 11645 13311 11679
rect 13737 11645 13771 11679
rect 14933 11645 14967 11679
rect 15393 11645 15427 11679
rect 15485 11645 15519 11679
rect 16957 11645 16991 11679
rect 18153 11645 18187 11679
rect 20545 11645 20579 11679
rect 21557 11645 21591 11679
rect 21833 11645 21867 11679
rect 22017 11645 22051 11679
rect 22477 11645 22511 11679
rect 24409 11645 24443 11679
rect 25697 11645 25731 11679
rect 26157 11645 26191 11679
rect 26709 11645 26743 11679
rect 27813 11645 27847 11679
rect 28273 11645 28307 11679
rect 30757 11645 30791 11679
rect 31769 11645 31803 11679
rect 35817 11645 35851 11679
rect 36093 11645 36127 11679
rect 5089 11577 5123 11611
rect 6377 11577 6411 11611
rect 7941 11577 7975 11611
rect 10057 11577 10091 11611
rect 16037 11577 16071 11611
rect 18061 11577 18095 11611
rect 31493 11577 31527 11611
rect 1593 11509 1627 11543
rect 1961 11509 1995 11543
rect 6469 11509 6503 11543
rect 11161 11509 11195 11543
rect 12541 11509 12575 11543
rect 17785 11509 17819 11543
rect 25237 11509 25271 11543
rect 30389 11509 30423 11543
rect 6009 11305 6043 11339
rect 7665 11305 7699 11339
rect 9413 11305 9447 11339
rect 9965 11305 9999 11339
rect 13001 11305 13035 11339
rect 14749 11305 14783 11339
rect 16497 11305 16531 11339
rect 17049 11305 17083 11339
rect 18521 11305 18555 11339
rect 18889 11305 18923 11339
rect 19257 11305 19291 11339
rect 19993 11305 20027 11339
rect 20361 11305 20395 11339
rect 20637 11305 20671 11339
rect 21741 11305 21775 11339
rect 22109 11305 22143 11339
rect 23673 11305 23707 11339
rect 24041 11305 24075 11339
rect 26801 11305 26835 11339
rect 3065 11237 3099 11271
rect 6101 11237 6135 11271
rect 8677 11237 8711 11271
rect 12173 11237 12207 11271
rect 17417 11237 17451 11271
rect 17509 11237 17543 11271
rect 19625 11237 19659 11271
rect 25237 11237 25271 11271
rect 29929 11237 29963 11271
rect 1409 11169 1443 11203
rect 4721 11169 4755 11203
rect 5089 11169 5123 11203
rect 5273 11169 5307 11203
rect 6745 11169 6779 11203
rect 7113 11169 7147 11203
rect 8217 11169 8251 11203
rect 10885 11169 10919 11203
rect 11069 11169 11103 11203
rect 11621 11169 11655 11203
rect 11805 11169 11839 11203
rect 13645 11169 13679 11203
rect 13921 11169 13955 11203
rect 15485 11169 15519 11203
rect 15577 11169 15611 11203
rect 16037 11169 16071 11203
rect 16221 11169 16255 11203
rect 17601 11169 17635 11203
rect 19073 11169 19107 11203
rect 23489 11169 23523 11203
rect 24869 11169 24903 11203
rect 26617 11169 26651 11203
rect 28549 11169 28583 11203
rect 30665 11169 30699 11203
rect 30757 11169 30791 11203
rect 31033 11169 31067 11203
rect 31125 11169 31159 11203
rect 1685 11101 1719 11135
rect 4169 11101 4203 11135
rect 4629 11101 4663 11135
rect 6561 11101 6595 11135
rect 7021 11101 7055 11135
rect 7941 11101 7975 11135
rect 8125 11101 8159 11135
rect 10793 11101 10827 11135
rect 13185 11101 13219 11135
rect 27077 11101 27111 11135
rect 30021 11101 30055 11135
rect 3525 11033 3559 11067
rect 5549 11033 5583 11067
rect 12633 11033 12667 11067
rect 13921 11033 13955 11067
rect 25605 11033 25639 11067
rect 26157 11033 26191 11067
rect 27537 11033 27571 11067
rect 28917 11033 28951 11067
rect 9045 10965 9079 10999
rect 10241 10965 10275 10999
rect 35817 10965 35851 10999
rect 3709 10761 3743 10795
rect 4537 10761 4571 10795
rect 8217 10761 8251 10795
rect 8493 10761 8527 10795
rect 10517 10761 10551 10795
rect 13185 10761 13219 10795
rect 13921 10761 13955 10795
rect 14657 10761 14691 10795
rect 15301 10761 15335 10795
rect 15761 10761 15795 10795
rect 16129 10761 16163 10795
rect 19349 10761 19383 10795
rect 20085 10761 20119 10795
rect 23949 10761 23983 10795
rect 25329 10761 25363 10795
rect 25697 10761 25731 10795
rect 28089 10761 28123 10795
rect 28641 10761 28675 10795
rect 29653 10761 29687 10795
rect 4169 10693 4203 10727
rect 9873 10693 9907 10727
rect 12817 10693 12851 10727
rect 16681 10693 16715 10727
rect 24317 10693 24351 10727
rect 30113 10693 30147 10727
rect 14381 10625 14415 10659
rect 26617 10625 26651 10659
rect 30757 10625 30791 10659
rect 31309 10625 31343 10659
rect 4813 10557 4847 10591
rect 5825 10557 5859 10591
rect 8677 10557 8711 10591
rect 8769 10557 8803 10591
rect 8953 10557 8987 10591
rect 9413 10557 9447 10591
rect 9505 10557 9539 10591
rect 12265 10557 12299 10591
rect 13001 10557 13035 10591
rect 14473 10557 14507 10591
rect 14933 10557 14967 10591
rect 16313 10557 16347 10591
rect 17877 10557 17911 10591
rect 18429 10557 18463 10591
rect 19901 10557 19935 10591
rect 20361 10557 20395 10591
rect 24133 10557 24167 10591
rect 24593 10557 24627 10591
rect 24961 10557 24995 10591
rect 25145 10557 25179 10591
rect 26709 10557 26743 10591
rect 26985 10557 27019 10591
rect 30849 10557 30883 10591
rect 31217 10557 31251 10591
rect 5457 10489 5491 10523
rect 10977 10489 11011 10523
rect 18337 10489 18371 10523
rect 30205 10489 30239 10523
rect 1593 10421 1627 10455
rect 1961 10421 1995 10455
rect 4629 10421 4663 10455
rect 6193 10421 6227 10455
rect 6561 10421 6595 10455
rect 7849 10421 7883 10455
rect 11345 10421 11379 10455
rect 11713 10421 11747 10455
rect 17417 10421 17451 10455
rect 26157 10421 26191 10455
rect 31677 10421 31711 10455
rect 4353 10217 4387 10251
rect 6837 10217 6871 10251
rect 8493 10217 8527 10251
rect 9137 10217 9171 10251
rect 11989 10217 12023 10251
rect 12449 10217 12483 10251
rect 13185 10217 13219 10251
rect 14841 10217 14875 10251
rect 16589 10217 16623 10251
rect 17693 10217 17727 10251
rect 19165 10217 19199 10251
rect 19533 10217 19567 10251
rect 21741 10217 21775 10251
rect 25605 10217 25639 10251
rect 26985 10217 27019 10251
rect 27997 10217 28031 10251
rect 30205 10217 30239 10251
rect 30665 10217 30699 10251
rect 30941 10217 30975 10251
rect 36553 10217 36587 10251
rect 4721 10149 4755 10183
rect 12817 10149 12851 10183
rect 15853 10149 15887 10183
rect 16221 10149 16255 10183
rect 23949 10149 23983 10183
rect 5549 10081 5583 10115
rect 8585 10081 8619 10115
rect 11437 10081 11471 10115
rect 13461 10081 13495 10115
rect 15301 10081 15335 10115
rect 16957 10081 16991 10115
rect 17969 10081 18003 10115
rect 18981 10081 19015 10115
rect 21925 10081 21959 10115
rect 22569 10081 22603 10115
rect 25421 10081 25455 10115
rect 26801 10081 26835 10115
rect 27813 10081 27847 10115
rect 29929 10081 29963 10115
rect 35449 10081 35483 10115
rect 5273 10013 5307 10047
rect 7389 10013 7423 10047
rect 11713 10013 11747 10047
rect 13369 10013 13403 10047
rect 13921 10013 13955 10047
rect 22293 10013 22327 10047
rect 35173 10013 35207 10047
rect 8769 9945 8803 9979
rect 17141 9945 17175 9979
rect 7757 9877 7791 9911
rect 9505 9877 9539 9911
rect 14289 9877 14323 9911
rect 15485 9877 15519 9911
rect 18153 9877 18187 9911
rect 18797 9877 18831 9911
rect 19809 9877 19843 9911
rect 27353 9877 27387 9911
rect 11069 9673 11103 9707
rect 12633 9673 12667 9707
rect 13461 9673 13495 9707
rect 15393 9673 15427 9707
rect 17509 9673 17543 9707
rect 18337 9673 18371 9707
rect 18889 9673 18923 9707
rect 21833 9673 21867 9707
rect 26801 9673 26835 9707
rect 27813 9673 27847 9707
rect 5365 9605 5399 9639
rect 7205 9605 7239 9639
rect 11989 9605 12023 9639
rect 16497 9605 16531 9639
rect 25789 9605 25823 9639
rect 35265 9605 35299 9639
rect 1869 9537 1903 9571
rect 3341 9537 3375 9571
rect 6653 9537 6687 9571
rect 8033 9537 8067 9571
rect 8217 9537 8251 9571
rect 13829 9537 13863 9571
rect 24317 9537 24351 9571
rect 35541 9537 35575 9571
rect 1961 9469 1995 9503
rect 2237 9469 2271 9503
rect 5733 9469 5767 9503
rect 7941 9469 7975 9503
rect 8309 9469 8343 9503
rect 8861 9469 8895 9503
rect 13921 9469 13955 9503
rect 14381 9469 14415 9503
rect 14473 9469 14507 9503
rect 15945 9469 15979 9503
rect 16957 9469 16991 9503
rect 17233 9469 17267 9503
rect 19441 9469 19475 9503
rect 19625 9469 19659 9503
rect 19947 9469 19981 9503
rect 20177 9469 20211 9503
rect 23489 9469 23523 9503
rect 24409 9469 24443 9503
rect 24685 9469 24719 9503
rect 7297 9401 7331 9435
rect 15025 9401 15059 9435
rect 20453 9401 20487 9435
rect 13001 9333 13035 9367
rect 16129 9333 16163 9367
rect 17141 9333 17175 9367
rect 17233 9333 17267 9367
rect 17877 9333 17911 9367
rect 19257 9333 19291 9367
rect 22293 9333 22327 9367
rect 22661 9333 22695 9367
rect 23305 9333 23339 9367
rect 23857 9333 23891 9367
rect 1961 9129 1995 9163
rect 8493 9129 8527 9163
rect 10057 9129 10091 9163
rect 12633 9129 12667 9163
rect 13921 9129 13955 9163
rect 24501 9129 24535 9163
rect 25973 9129 26007 9163
rect 14657 9061 14691 9095
rect 19993 9061 20027 9095
rect 25513 9061 25547 9095
rect 6101 8993 6135 9027
rect 7389 8993 7423 9027
rect 9873 8993 9907 9027
rect 10333 8993 10367 9027
rect 10885 8993 10919 9027
rect 11069 8993 11103 9027
rect 11621 8993 11655 9027
rect 11805 8993 11839 9027
rect 13185 8993 13219 9027
rect 15485 8993 15519 9027
rect 16037 8993 16071 9027
rect 16221 8993 16255 9027
rect 18337 8993 18371 9027
rect 18613 8993 18647 9027
rect 26157 8993 26191 9027
rect 7113 8925 7147 8959
rect 13093 8925 13127 8959
rect 15301 8925 15335 8959
rect 6285 8857 6319 8891
rect 9137 8789 9171 8823
rect 12081 8789 12115 8823
rect 13369 8789 13403 8823
rect 14381 8789 14415 8823
rect 16497 8789 16531 8823
rect 6101 8585 6135 8619
rect 7481 8585 7515 8619
rect 10609 8585 10643 8619
rect 11621 8585 11655 8619
rect 12817 8585 12851 8619
rect 13185 8585 13219 8619
rect 14933 8585 14967 8619
rect 15393 8585 15427 8619
rect 15669 8585 15703 8619
rect 18245 8585 18279 8619
rect 18521 8585 18555 8619
rect 18889 8585 18923 8619
rect 26065 8585 26099 8619
rect 7205 8517 7239 8551
rect 8861 8517 8895 8551
rect 10977 8517 11011 8551
rect 17877 8517 17911 8551
rect 8493 8449 8527 8483
rect 9689 8449 9723 8483
rect 11253 8449 11287 8483
rect 14197 8449 14231 8483
rect 15945 8449 15979 8483
rect 16405 8449 16439 8483
rect 16865 8449 16899 8483
rect 17417 8449 17451 8483
rect 9597 8381 9631 8415
rect 9965 8381 9999 8415
rect 10149 8381 10183 8415
rect 13737 8381 13771 8415
rect 14105 8381 14139 8415
rect 16589 8381 16623 8415
rect 16957 8381 16991 8415
rect 18061 8381 18095 8415
rect 8953 8313 8987 8347
rect 13277 8313 13311 8347
rect 14657 8313 14691 8347
rect 12173 8245 12207 8279
rect 9045 8041 9079 8075
rect 11069 8041 11103 8075
rect 13553 8041 13587 8075
rect 13829 8041 13863 8075
rect 15117 8041 15151 8075
rect 16681 8041 16715 8075
rect 20269 8041 20303 8075
rect 12633 7905 12667 7939
rect 13001 7905 13035 7939
rect 13093 7905 13127 7939
rect 15577 7905 15611 7939
rect 18061 7905 18095 7939
rect 21557 7905 21591 7939
rect 21925 7905 21959 7939
rect 23121 7905 23155 7939
rect 9689 7837 9723 7871
rect 9965 7837 9999 7871
rect 12173 7837 12207 7871
rect 15301 7837 15335 7871
rect 17785 7837 17819 7871
rect 21373 7837 21407 7871
rect 21833 7837 21867 7871
rect 19349 7701 19383 7735
rect 21189 7701 21223 7735
rect 22937 7701 22971 7735
rect 8493 7497 8527 7531
rect 9505 7497 9539 7531
rect 10149 7497 10183 7531
rect 11897 7497 11931 7531
rect 15025 7497 15059 7531
rect 15393 7497 15427 7531
rect 16313 7497 16347 7531
rect 17877 7497 17911 7531
rect 20085 7497 20119 7531
rect 21741 7497 21775 7531
rect 23029 7497 23063 7531
rect 12173 7429 12207 7463
rect 16037 7429 16071 7463
rect 10885 7361 10919 7395
rect 11253 7361 11287 7395
rect 13185 7361 13219 7395
rect 20453 7361 20487 7395
rect 22109 7361 22143 7395
rect 8861 7293 8895 7327
rect 10977 7293 11011 7327
rect 11345 7293 11379 7327
rect 12909 7293 12943 7327
rect 18337 7293 18371 7327
rect 20177 7293 20211 7327
rect 9873 7225 9907 7259
rect 12725 7225 12759 7259
rect 8677 7157 8711 7191
rect 10425 7157 10459 7191
rect 14289 7157 14323 7191
rect 10425 6953 10459 6987
rect 13001 6953 13035 6987
rect 20269 6953 20303 6987
rect 21097 6953 21131 6987
rect 21557 6953 21591 6987
rect 9505 6817 9539 6851
rect 10057 6817 10091 6851
rect 13737 6817 13771 6851
rect 14105 6817 14139 6851
rect 16773 6817 16807 6851
rect 17141 6817 17175 6851
rect 17233 6817 17267 6851
rect 19165 6817 19199 6851
rect 19533 6817 19567 6851
rect 27353 6817 27387 6851
rect 28733 6817 28767 6851
rect 10517 6749 10551 6783
rect 10793 6749 10827 6783
rect 11897 6749 11931 6783
rect 13093 6749 13127 6783
rect 13829 6749 13863 6783
rect 14013 6749 14047 6783
rect 16129 6749 16163 6783
rect 16681 6749 16715 6783
rect 19073 6749 19107 6783
rect 19441 6749 19475 6783
rect 22201 6749 22235 6783
rect 22477 6749 22511 6783
rect 23581 6749 23615 6783
rect 27077 6749 27111 6783
rect 14933 6681 14967 6715
rect 12541 6613 12575 6647
rect 14565 6613 14599 6647
rect 18797 6613 18831 6647
rect 10057 6409 10091 6443
rect 10609 6409 10643 6443
rect 12265 6409 12299 6443
rect 12817 6409 12851 6443
rect 13921 6409 13955 6443
rect 16589 6409 16623 6443
rect 17877 6409 17911 6443
rect 20453 6409 20487 6443
rect 22569 6409 22603 6443
rect 27445 6409 27479 6443
rect 7665 6341 7699 6375
rect 11253 6341 11287 6375
rect 15853 6341 15887 6375
rect 18521 6341 18555 6375
rect 15025 6273 15059 6307
rect 16221 6273 16255 6307
rect 18981 6273 19015 6307
rect 7849 6205 7883 6239
rect 8217 6205 8251 6239
rect 10241 6205 10275 6239
rect 10885 6205 10919 6239
rect 13553 6205 13587 6239
rect 14565 6205 14599 6239
rect 14749 6205 14783 6239
rect 15117 6205 15151 6239
rect 19073 6205 19107 6239
rect 19349 6205 19383 6239
rect 13185 6137 13219 6171
rect 22293 6137 22327 6171
rect 14381 6069 14415 6103
rect 16957 6069 16991 6103
rect 27077 6069 27111 6103
rect 14289 5865 14323 5899
rect 14749 5865 14783 5899
rect 17049 5865 17083 5899
rect 18889 5865 18923 5899
rect 18613 5797 18647 5831
rect 13001 5729 13035 5763
rect 15945 5729 15979 5763
rect 23673 5729 23707 5763
rect 12725 5661 12759 5695
rect 15669 5661 15703 5695
rect 19257 5525 19291 5559
rect 23489 5525 23523 5559
rect 10425 5321 10459 5355
rect 12817 5321 12851 5355
rect 16037 5321 16071 5355
rect 23857 5321 23891 5355
rect 13093 5253 13127 5287
rect 15761 5253 15795 5287
rect 8769 5185 8803 5219
rect 8861 5117 8895 5151
rect 9137 5117 9171 5151
rect 21833 5117 21867 5151
rect 22201 5117 22235 5151
rect 25605 5117 25639 5151
rect 25881 5117 25915 5151
rect 21649 4981 21683 5015
rect 25421 4981 25455 5015
rect 8861 4777 8895 4811
rect 12173 4777 12207 4811
rect 33517 4777 33551 4811
rect 19441 4709 19475 4743
rect 28181 4709 28215 4743
rect 10793 4641 10827 4675
rect 17785 4641 17819 4675
rect 32413 4641 32447 4675
rect 11069 4573 11103 4607
rect 18061 4573 18095 4607
rect 26525 4573 26559 4607
rect 26801 4573 26835 4607
rect 32137 4573 32171 4607
rect 9965 4233 9999 4267
rect 11253 4233 11287 4267
rect 18245 4233 18279 4267
rect 27353 4233 27387 4267
rect 8401 4097 8435 4131
rect 19073 4097 19107 4131
rect 19441 4097 19475 4131
rect 20821 4097 20855 4131
rect 25329 4097 25363 4131
rect 26893 4097 26927 4131
rect 8677 4029 8711 4063
rect 17877 4029 17911 4063
rect 19165 4029 19199 4063
rect 25421 4029 25455 4063
rect 25697 4029 25731 4063
rect 10793 3961 10827 3995
rect 32229 3961 32263 3995
rect 8309 3893 8343 3927
rect 32505 3893 32539 3927
rect 8401 3689 8435 3723
rect 11529 3689 11563 3723
rect 19165 3689 19199 3723
rect 24685 3689 24719 3723
rect 33517 3689 33551 3723
rect 16957 3621 16991 3655
rect 1777 3553 1811 3587
rect 4353 3553 4387 3587
rect 10149 3553 10183 3587
rect 15301 3553 15335 3587
rect 23397 3553 23431 3587
rect 1501 3485 1535 3519
rect 3157 3485 3191 3519
rect 4077 3485 4111 3519
rect 10425 3485 10459 3519
rect 15577 3485 15611 3519
rect 23121 3485 23155 3519
rect 32137 3485 32171 3519
rect 32413 3485 32447 3519
rect 5457 3349 5491 3383
rect 19993 3349 20027 3383
rect 25513 3349 25547 3383
rect 26801 3349 26835 3383
rect 35817 3349 35851 3383
rect 1961 3145 1995 3179
rect 4169 3145 4203 3179
rect 10057 3145 10091 3179
rect 10793 3145 10827 3179
rect 15301 3145 15335 3179
rect 16957 3145 16991 3179
rect 21281 3145 21315 3179
rect 23857 3145 23891 3179
rect 24593 3145 24627 3179
rect 26341 3145 26375 3179
rect 29101 3145 29135 3179
rect 33149 3145 33183 3179
rect 37381 3145 37415 3179
rect 1685 3077 1719 3111
rect 23213 3077 23247 3111
rect 8401 3009 8435 3043
rect 8769 3009 8803 3043
rect 14565 3009 14599 3043
rect 15393 3009 15427 3043
rect 15669 3009 15703 3043
rect 19809 3009 19843 3043
rect 25053 3009 25087 3043
rect 29285 3009 29319 3043
rect 31677 3009 31711 3043
rect 32045 3009 32079 3043
rect 8493 2941 8527 2975
rect 10517 2941 10551 2975
rect 14933 2941 14967 2975
rect 19901 2941 19935 2975
rect 20177 2941 20211 2975
rect 24777 2941 24811 2975
rect 29561 2941 29595 2975
rect 31217 2941 31251 2975
rect 31769 2941 31803 2975
rect 35817 2941 35851 2975
rect 36093 2941 36127 2975
rect 30941 2873 30975 2907
rect 4445 2805 4479 2839
rect 35633 2805 35667 2839
rect 3433 2601 3467 2635
rect 8493 2601 8527 2635
rect 11437 2601 11471 2635
rect 12449 2601 12483 2635
rect 15761 2601 15795 2635
rect 17785 2601 17819 2635
rect 22845 2601 22879 2635
rect 29377 2601 29411 2635
rect 31861 2601 31895 2635
rect 35173 2601 35207 2635
rect 6009 2533 6043 2567
rect 11989 2533 12023 2567
rect 28825 2533 28859 2567
rect 4629 2465 4663 2499
rect 9597 2465 9631 2499
rect 10333 2465 10367 2499
rect 13185 2465 13219 2499
rect 18613 2465 18647 2499
rect 21005 2465 21039 2499
rect 21741 2465 21775 2499
rect 26709 2465 26743 2499
rect 34897 2465 34931 2499
rect 35449 2465 35483 2499
rect 4353 2397 4387 2431
rect 9229 2397 9263 2431
rect 10057 2397 10091 2431
rect 12909 2397 12943 2431
rect 14565 2397 14599 2431
rect 18337 2397 18371 2431
rect 20637 2397 20671 2431
rect 21465 2397 21499 2431
rect 24869 2397 24903 2431
rect 26341 2397 26375 2431
rect 27169 2397 27203 2431
rect 27445 2397 27479 2431
rect 35725 2397 35759 2431
rect 18061 2329 18095 2363
rect 3801 2261 3835 2295
rect 19901 2261 19935 2295
rect 32229 2261 32263 2295
rect 36829 2261 36863 2295
<< metal1 >>
rect 3418 40196 3424 40248
rect 3476 40236 3482 40248
rect 7006 40236 7012 40248
rect 3476 40208 7012 40236
rect 3476 40196 3482 40208
rect 7006 40196 7012 40208
rect 7064 40196 7070 40248
rect 2958 40128 2964 40180
rect 3016 40168 3022 40180
rect 19150 40168 19156 40180
rect 3016 40140 19156 40168
rect 3016 40128 3022 40140
rect 19150 40128 19156 40140
rect 19208 40128 19214 40180
rect 3234 40060 3240 40112
rect 3292 40100 3298 40112
rect 20070 40100 20076 40112
rect 3292 40072 20076 40100
rect 3292 40060 3298 40072
rect 20070 40060 20076 40072
rect 20128 40060 20134 40112
rect 26878 40060 26884 40112
rect 26936 40100 26942 40112
rect 35250 40100 35256 40112
rect 26936 40072 35256 40100
rect 26936 40060 26942 40072
rect 35250 40060 35256 40072
rect 35308 40060 35314 40112
rect 15746 39380 15752 39432
rect 15804 39420 15810 39432
rect 33594 39420 33600 39432
rect 15804 39392 33600 39420
rect 15804 39380 15810 39392
rect 33594 39380 33600 39392
rect 33652 39380 33658 39432
rect 4154 39312 4160 39364
rect 4212 39352 4218 39364
rect 5166 39352 5172 39364
rect 4212 39324 5172 39352
rect 4212 39312 4218 39324
rect 5166 39312 5172 39324
rect 5224 39312 5230 39364
rect 8846 39312 8852 39364
rect 8904 39352 8910 39364
rect 22922 39352 22928 39364
rect 8904 39324 22928 39352
rect 8904 39312 8910 39324
rect 22922 39312 22928 39324
rect 22980 39312 22986 39364
rect 11422 39244 11428 39296
rect 11480 39284 11486 39296
rect 34514 39284 34520 39296
rect 11480 39256 34520 39284
rect 11480 39244 11486 39256
rect 34514 39244 34520 39256
rect 34572 39244 34578 39296
rect 1104 39194 38548 39216
rect 1104 39142 4246 39194
rect 4298 39142 4310 39194
rect 4362 39142 4374 39194
rect 4426 39142 4438 39194
rect 4490 39142 34966 39194
rect 35018 39142 35030 39194
rect 35082 39142 35094 39194
rect 35146 39142 35158 39194
rect 35210 39142 38548 39194
rect 1104 39120 38548 39142
rect 2774 39040 2780 39092
rect 2832 39080 2838 39092
rect 3789 39083 3847 39089
rect 3789 39080 3801 39083
rect 2832 39052 3801 39080
rect 2832 39040 2838 39052
rect 3789 39049 3801 39052
rect 3835 39049 3847 39083
rect 3789 39043 3847 39049
rect 8757 39083 8815 39089
rect 8757 39049 8769 39083
rect 8803 39080 8815 39083
rect 8846 39080 8852 39092
rect 8803 39052 8852 39080
rect 8803 39049 8815 39052
rect 8757 39043 8815 39049
rect 3804 38944 3832 39043
rect 8846 39040 8852 39052
rect 8904 39040 8910 39092
rect 9585 39083 9643 39089
rect 9585 39049 9597 39083
rect 9631 39080 9643 39083
rect 9674 39080 9680 39092
rect 9631 39052 9680 39080
rect 9631 39049 9643 39052
rect 9585 39043 9643 39049
rect 9674 39040 9680 39052
rect 9732 39040 9738 39092
rect 11422 39080 11428 39092
rect 11383 39052 11428 39080
rect 11422 39040 11428 39052
rect 11480 39040 11486 39092
rect 26234 39040 26240 39092
rect 26292 39080 26298 39092
rect 26605 39083 26663 39089
rect 26605 39080 26617 39083
rect 26292 39052 26617 39080
rect 26292 39040 26298 39052
rect 26605 39049 26617 39052
rect 26651 39080 26663 39083
rect 27338 39080 27344 39092
rect 26651 39052 27344 39080
rect 26651 39049 26663 39052
rect 26605 39043 26663 39049
rect 27338 39040 27344 39052
rect 27396 39040 27402 39092
rect 6454 38972 6460 39024
rect 6512 39012 6518 39024
rect 6641 39015 6699 39021
rect 6641 39012 6653 39015
rect 6512 38984 6653 39012
rect 6512 38972 6518 38984
rect 6641 38981 6653 38984
rect 6687 38981 6699 39015
rect 6641 38975 6699 38981
rect 4341 38947 4399 38953
rect 4341 38944 4353 38947
rect 3804 38916 4353 38944
rect 4341 38913 4353 38916
rect 4387 38913 4399 38947
rect 6656 38944 6684 38975
rect 7469 38947 7527 38953
rect 7469 38944 7481 38947
rect 6656 38916 7481 38944
rect 4341 38907 4399 38913
rect 7469 38913 7481 38916
rect 7515 38913 7527 38947
rect 9692 38944 9720 39040
rect 12805 39015 12863 39021
rect 12805 38981 12817 39015
rect 12851 39012 12863 39015
rect 12851 38984 14412 39012
rect 12851 38981 12863 38984
rect 12805 38975 12863 38981
rect 10137 38947 10195 38953
rect 10137 38944 10149 38947
rect 9692 38916 10149 38944
rect 7469 38907 7527 38913
rect 10137 38913 10149 38916
rect 10183 38913 10195 38947
rect 10137 38907 10195 38913
rect 12894 38904 12900 38956
rect 12952 38944 12958 38956
rect 13541 38947 13599 38953
rect 13541 38944 13553 38947
rect 12952 38916 13553 38944
rect 12952 38904 12958 38916
rect 13541 38913 13553 38916
rect 13587 38913 13599 38947
rect 13541 38907 13599 38913
rect 14384 38888 14412 38984
rect 19978 38972 19984 39024
rect 20036 39012 20042 39024
rect 20036 38984 26924 39012
rect 20036 38972 20042 38984
rect 15289 38947 15347 38953
rect 15289 38913 15301 38947
rect 15335 38944 15347 38947
rect 15746 38944 15752 38956
rect 15335 38916 15752 38944
rect 15335 38913 15347 38916
rect 15289 38907 15347 38913
rect 15746 38904 15752 38916
rect 15804 38904 15810 38956
rect 26896 38944 26924 38984
rect 35250 38944 35256 38956
rect 26896 38916 35256 38944
rect 35250 38904 35256 38916
rect 35308 38904 35314 38956
rect 4065 38879 4123 38885
rect 4065 38876 4077 38879
rect 3436 38848 4077 38876
rect 2774 38700 2780 38752
rect 2832 38740 2838 38752
rect 3436 38749 3464 38848
rect 4065 38845 4077 38848
rect 4111 38876 4123 38879
rect 5442 38876 5448 38888
rect 4111 38848 5448 38876
rect 4111 38845 4123 38848
rect 4065 38839 4123 38845
rect 5442 38836 5448 38848
rect 5500 38876 5506 38888
rect 6273 38879 6331 38885
rect 6273 38876 6285 38879
rect 5500 38848 6285 38876
rect 5500 38836 5506 38848
rect 6273 38845 6285 38848
rect 6319 38876 6331 38879
rect 7193 38879 7251 38885
rect 7193 38876 7205 38879
rect 6319 38848 7205 38876
rect 6319 38845 6331 38848
rect 6273 38839 6331 38845
rect 7193 38845 7205 38848
rect 7239 38845 7251 38879
rect 7193 38839 7251 38845
rect 7300 38848 9628 38876
rect 5721 38811 5779 38817
rect 5721 38777 5733 38811
rect 5767 38808 5779 38811
rect 7300 38808 7328 38848
rect 5767 38780 7328 38808
rect 9600 38808 9628 38848
rect 9674 38836 9680 38888
rect 9732 38876 9738 38888
rect 9861 38879 9919 38885
rect 9861 38876 9873 38879
rect 9732 38848 9873 38876
rect 9732 38836 9738 38848
rect 9861 38845 9873 38848
rect 9907 38845 9919 38879
rect 13354 38876 13360 38888
rect 9861 38839 9919 38845
rect 9968 38848 13360 38876
rect 9968 38808 9996 38848
rect 13354 38836 13360 38848
rect 13412 38836 13418 38888
rect 13449 38879 13507 38885
rect 13449 38845 13461 38879
rect 13495 38845 13507 38879
rect 13449 38839 13507 38845
rect 9600 38780 9996 38808
rect 5767 38777 5779 38780
rect 5721 38771 5779 38777
rect 3421 38743 3479 38749
rect 3421 38740 3433 38743
rect 2832 38712 3433 38740
rect 2832 38700 2838 38712
rect 3421 38709 3433 38712
rect 3467 38709 3479 38743
rect 3421 38703 3479 38709
rect 13265 38743 13323 38749
rect 13265 38709 13277 38743
rect 13311 38740 13323 38743
rect 13464 38740 13492 38839
rect 13630 38836 13636 38888
rect 13688 38876 13694 38888
rect 14277 38879 14335 38885
rect 14277 38876 14289 38879
rect 13688 38848 14289 38876
rect 13688 38836 13694 38848
rect 14277 38845 14289 38848
rect 14323 38845 14335 38879
rect 14277 38839 14335 38845
rect 14366 38836 14372 38888
rect 14424 38876 14430 38888
rect 15473 38879 15531 38885
rect 14424 38848 14469 38876
rect 14424 38836 14430 38848
rect 15473 38845 15485 38879
rect 15519 38845 15531 38879
rect 27065 38879 27123 38885
rect 27065 38876 27077 38879
rect 15473 38839 15531 38845
rect 26252 38848 27077 38876
rect 15286 38768 15292 38820
rect 15344 38808 15350 38820
rect 15488 38808 15516 38839
rect 26142 38808 26148 38820
rect 15344 38780 15516 38808
rect 16408 38780 26148 38808
rect 15344 38768 15350 38780
rect 16408 38740 16436 38780
rect 26142 38768 26148 38780
rect 26200 38768 26206 38820
rect 13311 38712 16436 38740
rect 17037 38743 17095 38749
rect 13311 38709 13323 38712
rect 13265 38703 13323 38709
rect 17037 38709 17049 38743
rect 17083 38740 17095 38743
rect 17862 38740 17868 38752
rect 17083 38712 17868 38740
rect 17083 38709 17095 38712
rect 17037 38703 17095 38709
rect 17862 38700 17868 38712
rect 17920 38700 17926 38752
rect 26050 38700 26056 38752
rect 26108 38740 26114 38752
rect 26252 38749 26280 38848
rect 27065 38845 27077 38848
rect 27111 38845 27123 38879
rect 27338 38876 27344 38888
rect 27299 38848 27344 38876
rect 27065 38839 27123 38845
rect 27338 38836 27344 38848
rect 27396 38836 27402 38888
rect 28718 38808 28724 38820
rect 28679 38780 28724 38808
rect 28718 38768 28724 38780
rect 28776 38768 28782 38820
rect 26237 38743 26295 38749
rect 26237 38740 26249 38743
rect 26108 38712 26249 38740
rect 26108 38700 26114 38712
rect 26237 38709 26249 38712
rect 26283 38709 26295 38743
rect 26237 38703 26295 38709
rect 1104 38650 38548 38672
rect 1104 38598 19606 38650
rect 19658 38598 19670 38650
rect 19722 38598 19734 38650
rect 19786 38598 19798 38650
rect 19850 38598 38548 38650
rect 1104 38576 38548 38598
rect 5534 38496 5540 38548
rect 5592 38536 5598 38548
rect 6730 38536 6736 38548
rect 5592 38508 6736 38536
rect 5592 38496 5598 38508
rect 6730 38496 6736 38508
rect 6788 38496 6794 38548
rect 13354 38496 13360 38548
rect 13412 38536 13418 38548
rect 13630 38536 13636 38548
rect 13412 38508 13636 38536
rect 13412 38496 13418 38508
rect 13630 38496 13636 38508
rect 13688 38496 13694 38548
rect 19426 38496 19432 38548
rect 19484 38536 19490 38548
rect 24578 38536 24584 38548
rect 19484 38508 24584 38536
rect 19484 38496 19490 38508
rect 24578 38496 24584 38508
rect 24636 38496 24642 38548
rect 31478 38496 31484 38548
rect 31536 38536 31542 38548
rect 37734 38536 37740 38548
rect 31536 38508 37740 38536
rect 31536 38496 31542 38508
rect 37734 38496 37740 38508
rect 37792 38496 37798 38548
rect 14 38428 20 38480
rect 72 38468 78 38480
rect 474 38468 480 38480
rect 72 38440 480 38468
rect 72 38428 78 38440
rect 474 38428 480 38440
rect 532 38428 538 38480
rect 3145 38471 3203 38477
rect 3145 38437 3157 38471
rect 3191 38468 3203 38471
rect 3694 38468 3700 38480
rect 3191 38440 3700 38468
rect 3191 38437 3203 38440
rect 3145 38431 3203 38437
rect 3694 38428 3700 38440
rect 3752 38428 3758 38480
rect 4614 38360 4620 38412
rect 4672 38400 4678 38412
rect 5534 38400 5540 38412
rect 4672 38372 5540 38400
rect 4672 38360 4678 38372
rect 5534 38360 5540 38372
rect 5592 38400 5598 38412
rect 5721 38403 5779 38409
rect 5721 38400 5733 38403
rect 5592 38372 5733 38400
rect 5592 38360 5598 38372
rect 5721 38369 5733 38372
rect 5767 38369 5779 38403
rect 13354 38400 13360 38412
rect 13315 38372 13360 38400
rect 5721 38363 5779 38369
rect 13354 38360 13360 38372
rect 13412 38360 13418 38412
rect 17310 38360 17316 38412
rect 17368 38400 17374 38412
rect 17497 38403 17555 38409
rect 17497 38400 17509 38403
rect 17368 38372 17509 38400
rect 17368 38360 17374 38372
rect 17497 38369 17509 38372
rect 17543 38369 17555 38403
rect 23198 38400 23204 38412
rect 23159 38372 23204 38400
rect 17497 38363 17555 38369
rect 23198 38360 23204 38372
rect 23256 38360 23262 38412
rect 26786 38400 26792 38412
rect 26747 38372 26792 38400
rect 26786 38360 26792 38372
rect 26844 38360 26850 38412
rect 29454 38360 29460 38412
rect 29512 38400 29518 38412
rect 29825 38403 29883 38409
rect 29825 38400 29837 38403
rect 29512 38372 29837 38400
rect 29512 38360 29518 38372
rect 29825 38369 29837 38372
rect 29871 38369 29883 38403
rect 29825 38363 29883 38369
rect 31754 38360 31760 38412
rect 31812 38400 31818 38412
rect 32401 38403 32459 38409
rect 32401 38400 32413 38403
rect 31812 38372 32413 38400
rect 31812 38360 31818 38372
rect 32401 38369 32413 38372
rect 32447 38369 32459 38403
rect 32401 38363 32459 38369
rect 1486 38332 1492 38344
rect 1447 38304 1492 38332
rect 1486 38292 1492 38304
rect 1544 38292 1550 38344
rect 1670 38292 1676 38344
rect 1728 38332 1734 38344
rect 1765 38335 1823 38341
rect 1765 38332 1777 38335
rect 1728 38304 1777 38332
rect 1728 38292 1734 38304
rect 1765 38301 1777 38304
rect 1811 38301 1823 38335
rect 5442 38332 5448 38344
rect 5403 38304 5448 38332
rect 1765 38295 1823 38301
rect 5442 38292 5448 38304
rect 5500 38292 5506 38344
rect 7101 38335 7159 38341
rect 7101 38301 7113 38335
rect 7147 38332 7159 38335
rect 7650 38332 7656 38344
rect 7147 38304 7656 38332
rect 7147 38301 7159 38304
rect 7101 38295 7159 38301
rect 7650 38292 7656 38304
rect 7708 38292 7714 38344
rect 11698 38332 11704 38344
rect 9876 38304 11704 38332
rect 7374 38196 7380 38208
rect 7335 38168 7380 38196
rect 7374 38156 7380 38168
rect 7432 38156 7438 38208
rect 9674 38156 9680 38208
rect 9732 38196 9738 38208
rect 9876 38205 9904 38304
rect 11698 38292 11704 38304
rect 11756 38292 11762 38344
rect 11882 38292 11888 38344
rect 11940 38332 11946 38344
rect 11977 38335 12035 38341
rect 11977 38332 11989 38335
rect 11940 38304 11989 38332
rect 11940 38292 11946 38304
rect 11977 38301 11989 38304
rect 12023 38301 12035 38335
rect 17218 38332 17224 38344
rect 17179 38304 17224 38332
rect 11977 38295 12035 38301
rect 17218 38292 17224 38304
rect 17276 38292 17282 38344
rect 22925 38335 22983 38341
rect 22925 38301 22937 38335
rect 22971 38332 22983 38335
rect 23382 38332 23388 38344
rect 22971 38304 23388 38332
rect 22971 38301 22983 38304
rect 22925 38295 22983 38301
rect 23382 38292 23388 38304
rect 23440 38292 23446 38344
rect 26050 38292 26056 38344
rect 26108 38332 26114 38344
rect 26513 38335 26571 38341
rect 26513 38332 26525 38335
rect 26108 38304 26525 38332
rect 26108 38292 26114 38304
rect 26513 38301 26525 38304
rect 26559 38301 26571 38335
rect 26513 38295 26571 38301
rect 29549 38335 29607 38341
rect 29549 38301 29561 38335
rect 29595 38332 29607 38335
rect 30006 38332 30012 38344
rect 29595 38304 30012 38332
rect 29595 38301 29607 38304
rect 29549 38295 29607 38301
rect 30006 38292 30012 38304
rect 30064 38332 30070 38344
rect 32122 38332 32128 38344
rect 30064 38304 32128 38332
rect 30064 38292 30070 38304
rect 32122 38292 32128 38304
rect 32180 38292 32186 38344
rect 9861 38199 9919 38205
rect 9861 38196 9873 38199
rect 9732 38168 9873 38196
rect 9732 38156 9738 38168
rect 9861 38165 9873 38168
rect 9907 38165 9919 38199
rect 9861 38159 9919 38165
rect 15286 38156 15292 38208
rect 15344 38196 15350 38208
rect 15473 38199 15531 38205
rect 15473 38196 15485 38199
rect 15344 38168 15485 38196
rect 15344 38156 15350 38168
rect 15473 38165 15485 38168
rect 15519 38165 15531 38199
rect 15473 38159 15531 38165
rect 18230 38156 18236 38208
rect 18288 38196 18294 38208
rect 18601 38199 18659 38205
rect 18601 38196 18613 38199
rect 18288 38168 18613 38196
rect 18288 38156 18294 38168
rect 18601 38165 18613 38168
rect 18647 38165 18659 38199
rect 19426 38196 19432 38208
rect 19387 38168 19432 38196
rect 18601 38159 18659 38165
rect 19426 38156 19432 38168
rect 19484 38156 19490 38208
rect 24302 38196 24308 38208
rect 24263 38168 24308 38196
rect 24302 38156 24308 38168
rect 24360 38156 24366 38208
rect 27890 38196 27896 38208
rect 27851 38168 27896 38196
rect 27890 38156 27896 38168
rect 27948 38156 27954 38208
rect 30929 38199 30987 38205
rect 30929 38165 30941 38199
rect 30975 38196 30987 38199
rect 31018 38196 31024 38208
rect 30975 38168 31024 38196
rect 30975 38165 30987 38168
rect 30929 38159 30987 38165
rect 31018 38156 31024 38168
rect 31076 38156 31082 38208
rect 33226 38156 33232 38208
rect 33284 38196 33290 38208
rect 33505 38199 33563 38205
rect 33505 38196 33517 38199
rect 33284 38168 33517 38196
rect 33284 38156 33290 38168
rect 33505 38165 33517 38168
rect 33551 38165 33563 38199
rect 33505 38159 33563 38165
rect 1104 38106 38548 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 34966 38106
rect 35018 38054 35030 38106
rect 35082 38054 35094 38106
rect 35146 38054 35158 38106
rect 35210 38054 38548 38106
rect 1104 38032 38548 38054
rect 1486 37952 1492 38004
rect 1544 37992 1550 38004
rect 1949 37995 2007 38001
rect 1949 37992 1961 37995
rect 1544 37964 1961 37992
rect 1544 37952 1550 37964
rect 1949 37961 1961 37964
rect 1995 37992 2007 37995
rect 2682 37992 2688 38004
rect 1995 37964 2688 37992
rect 1995 37961 2007 37964
rect 1949 37955 2007 37961
rect 2682 37952 2688 37964
rect 2740 37952 2746 38004
rect 5534 37992 5540 38004
rect 5495 37964 5540 37992
rect 5534 37952 5540 37964
rect 5592 37952 5598 38004
rect 7006 37952 7012 38004
rect 7064 37992 7070 38004
rect 7193 37995 7251 38001
rect 7193 37992 7205 37995
rect 7064 37964 7205 37992
rect 7064 37952 7070 37964
rect 7193 37961 7205 37964
rect 7239 37961 7251 37995
rect 11882 37992 11888 38004
rect 11843 37964 11888 37992
rect 7193 37955 7251 37961
rect 5442 37816 5448 37868
rect 5500 37856 5506 37868
rect 5813 37859 5871 37865
rect 5813 37856 5825 37859
rect 5500 37828 5825 37856
rect 5500 37816 5506 37828
rect 5813 37825 5825 37828
rect 5859 37825 5871 37859
rect 7208 37856 7236 37955
rect 11882 37952 11888 37964
rect 11940 37952 11946 38004
rect 23017 37995 23075 38001
rect 23017 37961 23029 37995
rect 23063 37992 23075 37995
rect 23198 37992 23204 38004
rect 23063 37964 23204 37992
rect 23063 37961 23075 37964
rect 23017 37955 23075 37961
rect 23198 37952 23204 37964
rect 23256 37952 23262 38004
rect 25222 37952 25228 38004
rect 25280 37992 25286 38004
rect 27617 37995 27675 38001
rect 27617 37992 27629 37995
rect 25280 37964 27629 37992
rect 25280 37952 25286 37964
rect 27617 37961 27629 37964
rect 27663 37961 27675 37995
rect 27617 37955 27675 37961
rect 29454 37952 29460 38004
rect 29512 37992 29518 38004
rect 29549 37995 29607 38001
rect 29549 37992 29561 37995
rect 29512 37964 29561 37992
rect 29512 37952 29518 37964
rect 29549 37961 29561 37964
rect 29595 37961 29607 37995
rect 30006 37992 30012 38004
rect 29967 37964 30012 37992
rect 29549 37955 29607 37961
rect 30006 37952 30012 37964
rect 30064 37952 30070 38004
rect 31386 37992 31392 38004
rect 31347 37964 31392 37992
rect 31386 37952 31392 37964
rect 31444 37952 31450 38004
rect 31754 37952 31760 38004
rect 31812 37992 31818 38004
rect 32033 37995 32091 38001
rect 32033 37992 32045 37995
rect 31812 37964 32045 37992
rect 31812 37952 31818 37964
rect 32033 37961 32045 37964
rect 32079 37961 32091 37995
rect 32033 37955 32091 37961
rect 7653 37859 7711 37865
rect 7653 37856 7665 37859
rect 7208 37828 7665 37856
rect 5813 37819 5871 37825
rect 7653 37825 7665 37828
rect 7699 37825 7711 37859
rect 7653 37819 7711 37825
rect 11149 37859 11207 37865
rect 11149 37825 11161 37859
rect 11195 37856 11207 37859
rect 11900 37856 11928 37952
rect 33226 37884 33232 37936
rect 33284 37884 33290 37936
rect 11195 37828 11928 37856
rect 19245 37859 19303 37865
rect 11195 37825 11207 37828
rect 11149 37819 11207 37825
rect 19245 37825 19257 37859
rect 19291 37856 19303 37859
rect 19613 37859 19671 37865
rect 19613 37856 19625 37859
rect 19291 37828 19625 37856
rect 19291 37825 19303 37828
rect 19245 37819 19303 37825
rect 19613 37825 19625 37828
rect 19659 37856 19671 37859
rect 19978 37856 19984 37868
rect 19659 37828 19984 37856
rect 19659 37825 19671 37828
rect 19613 37819 19671 37825
rect 5828 37788 5856 37819
rect 19978 37816 19984 37828
rect 20036 37816 20042 37868
rect 26145 37859 26203 37865
rect 26145 37825 26157 37859
rect 26191 37856 26203 37859
rect 26513 37859 26571 37865
rect 26513 37856 26525 37859
rect 26191 37828 26525 37856
rect 26191 37825 26203 37828
rect 26145 37819 26203 37825
rect 26513 37825 26525 37828
rect 26559 37856 26571 37859
rect 26694 37856 26700 37868
rect 26559 37828 26700 37856
rect 26559 37825 26571 37828
rect 26513 37819 26571 37825
rect 26694 37816 26700 37828
rect 26752 37816 26758 37868
rect 32398 37856 32404 37868
rect 32359 37828 32404 37856
rect 32398 37816 32404 37828
rect 32456 37816 32462 37868
rect 33244 37856 33272 37884
rect 33152 37828 33272 37856
rect 35713 37859 35771 37865
rect 7374 37788 7380 37800
rect 5828 37760 7380 37788
rect 7374 37748 7380 37760
rect 7432 37748 7438 37800
rect 10781 37791 10839 37797
rect 10781 37757 10793 37791
rect 10827 37788 10839 37791
rect 17310 37788 17316 37800
rect 10827 37760 11008 37788
rect 17271 37760 17316 37788
rect 10827 37757 10839 37760
rect 10781 37751 10839 37757
rect 9030 37720 9036 37732
rect 8991 37692 9036 37720
rect 9030 37680 9036 37692
rect 9088 37680 9094 37732
rect 10597 37723 10655 37729
rect 10597 37720 10609 37723
rect 10428 37692 10609 37720
rect 10428 37664 10456 37692
rect 10597 37689 10609 37692
rect 10643 37689 10655 37723
rect 10597 37683 10655 37689
rect 10980 37664 11008 37760
rect 17310 37748 17316 37760
rect 17368 37748 17374 37800
rect 19337 37791 19395 37797
rect 19337 37788 19349 37791
rect 18156 37760 19349 37788
rect 18156 37664 18184 37760
rect 19337 37757 19349 37760
rect 19383 37788 19395 37791
rect 19426 37788 19432 37800
rect 19383 37760 19432 37788
rect 19383 37757 19395 37760
rect 19337 37751 19395 37757
rect 19426 37748 19432 37760
rect 19484 37748 19490 37800
rect 33152 37797 33180 37828
rect 35713 37825 35725 37859
rect 35759 37856 35771 37859
rect 36078 37856 36084 37868
rect 35759 37828 36084 37856
rect 35759 37825 35771 37828
rect 35713 37819 35771 37825
rect 36078 37816 36084 37828
rect 36136 37816 36142 37868
rect 26237 37791 26295 37797
rect 26237 37788 26249 37791
rect 26068 37760 26249 37788
rect 26068 37664 26096 37760
rect 26237 37757 26249 37760
rect 26283 37757 26295 37791
rect 32309 37791 32367 37797
rect 32309 37788 32321 37791
rect 26237 37751 26295 37757
rect 31864 37760 32321 37788
rect 31864 37664 31892 37760
rect 32309 37757 32321 37760
rect 32355 37757 32367 37791
rect 32309 37751 32367 37757
rect 33137 37791 33195 37797
rect 33137 37757 33149 37791
rect 33183 37757 33195 37791
rect 33137 37751 33195 37757
rect 33226 37748 33232 37800
rect 33284 37788 33290 37800
rect 35805 37791 35863 37797
rect 33284 37760 33329 37788
rect 33284 37748 33290 37760
rect 35805 37757 35817 37791
rect 35851 37757 35863 37791
rect 35805 37751 35863 37757
rect 35710 37680 35716 37732
rect 35768 37720 35774 37732
rect 35820 37720 35848 37751
rect 35768 37692 35848 37720
rect 35768 37680 35774 37692
rect 1670 37652 1676 37664
rect 1631 37624 1676 37652
rect 1670 37612 1676 37624
rect 1728 37612 1734 37664
rect 10410 37652 10416 37664
rect 10371 37624 10416 37652
rect 10410 37612 10416 37624
rect 10468 37612 10474 37664
rect 10962 37612 10968 37664
rect 11020 37652 11026 37664
rect 11425 37655 11483 37661
rect 11425 37652 11437 37655
rect 11020 37624 11437 37652
rect 11020 37612 11026 37624
rect 11425 37621 11437 37624
rect 11471 37621 11483 37655
rect 11425 37615 11483 37621
rect 11698 37612 11704 37664
rect 11756 37652 11762 37664
rect 12158 37652 12164 37664
rect 11756 37624 12164 37652
rect 11756 37612 11762 37624
rect 12158 37612 12164 37624
rect 12216 37612 12222 37664
rect 17218 37612 17224 37664
rect 17276 37652 17282 37664
rect 17681 37655 17739 37661
rect 17681 37652 17693 37655
rect 17276 37624 17693 37652
rect 17276 37612 17282 37624
rect 17681 37621 17693 37624
rect 17727 37652 17739 37655
rect 18138 37652 18144 37664
rect 17727 37624 18144 37652
rect 17727 37621 17739 37624
rect 17681 37615 17739 37621
rect 18138 37612 18144 37624
rect 18196 37612 18202 37664
rect 20714 37652 20720 37664
rect 20675 37624 20720 37652
rect 20714 37612 20720 37624
rect 20772 37612 20778 37664
rect 23382 37652 23388 37664
rect 23295 37624 23388 37652
rect 23382 37612 23388 37624
rect 23440 37652 23446 37664
rect 25685 37655 25743 37661
rect 25685 37652 25697 37655
rect 23440 37624 25697 37652
rect 23440 37612 23446 37624
rect 25685 37621 25697 37624
rect 25731 37652 25743 37655
rect 26050 37652 26056 37664
rect 25731 37624 26056 37652
rect 25731 37621 25743 37624
rect 25685 37615 25743 37621
rect 26050 37612 26056 37624
rect 26108 37612 26114 37664
rect 31757 37655 31815 37661
rect 31757 37621 31769 37655
rect 31803 37652 31815 37655
rect 31846 37652 31852 37664
rect 31803 37624 31852 37652
rect 31803 37621 31815 37624
rect 31757 37615 31815 37621
rect 31846 37612 31852 37624
rect 31904 37612 31910 37664
rect 36538 37612 36544 37664
rect 36596 37652 36602 37664
rect 37185 37655 37243 37661
rect 37185 37652 37197 37655
rect 36596 37624 37197 37652
rect 36596 37612 36602 37624
rect 37185 37621 37197 37624
rect 37231 37621 37243 37655
rect 37185 37615 37243 37621
rect 1104 37562 38548 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 38548 37562
rect 1104 37488 38548 37510
rect 1578 37408 1584 37460
rect 1636 37448 1642 37460
rect 2314 37448 2320 37460
rect 1636 37420 2320 37448
rect 1636 37408 1642 37420
rect 2314 37408 2320 37420
rect 2372 37408 2378 37460
rect 26786 37448 26792 37460
rect 26747 37420 26792 37448
rect 26786 37408 26792 37420
rect 26844 37408 26850 37460
rect 34790 37408 34796 37460
rect 34848 37448 34854 37460
rect 35161 37451 35219 37457
rect 35161 37448 35173 37451
rect 34848 37420 35173 37448
rect 34848 37408 34854 37420
rect 35161 37417 35173 37420
rect 35207 37417 35219 37451
rect 35161 37411 35219 37417
rect 32122 37340 32128 37392
rect 32180 37380 32186 37392
rect 32769 37383 32827 37389
rect 32769 37380 32781 37383
rect 32180 37352 32781 37380
rect 32180 37340 32186 37352
rect 32769 37349 32781 37352
rect 32815 37380 32827 37383
rect 32815 37352 33824 37380
rect 32815 37349 32827 37352
rect 32769 37343 32827 37349
rect 5442 37272 5448 37324
rect 5500 37312 5506 37324
rect 5629 37315 5687 37321
rect 5629 37312 5641 37315
rect 5500 37284 5641 37312
rect 5500 37272 5506 37284
rect 5629 37281 5641 37284
rect 5675 37281 5687 37315
rect 5629 37275 5687 37281
rect 5905 37315 5963 37321
rect 5905 37281 5917 37315
rect 5951 37312 5963 37315
rect 5994 37312 6000 37324
rect 5951 37284 6000 37312
rect 5951 37281 5963 37284
rect 5905 37275 5963 37281
rect 5994 37272 6000 37284
rect 6052 37272 6058 37324
rect 9674 37312 9680 37324
rect 9635 37284 9680 37312
rect 9674 37272 9680 37284
rect 9732 37272 9738 37324
rect 9950 37312 9956 37324
rect 9911 37284 9956 37312
rect 9950 37272 9956 37284
rect 10008 37272 10014 37324
rect 12434 37272 12440 37324
rect 12492 37312 12498 37324
rect 12492 37284 12537 37312
rect 12492 37272 12498 37284
rect 13814 37272 13820 37324
rect 13872 37312 13878 37324
rect 15010 37312 15016 37324
rect 13872 37284 15016 37312
rect 13872 37272 13878 37284
rect 15010 37272 15016 37284
rect 15068 37272 15074 37324
rect 15562 37312 15568 37324
rect 15523 37284 15568 37312
rect 15562 37272 15568 37284
rect 15620 37272 15626 37324
rect 16945 37315 17003 37321
rect 16945 37281 16957 37315
rect 16991 37312 17003 37315
rect 17586 37312 17592 37324
rect 16991 37284 17592 37312
rect 16991 37281 17003 37284
rect 16945 37275 17003 37281
rect 17586 37272 17592 37284
rect 17644 37272 17650 37324
rect 18598 37312 18604 37324
rect 18559 37284 18604 37312
rect 18598 37272 18604 37284
rect 18656 37272 18662 37324
rect 26050 37272 26056 37324
rect 26108 37312 26114 37324
rect 26237 37315 26295 37321
rect 26237 37312 26249 37315
rect 26108 37284 26249 37312
rect 26108 37272 26114 37284
rect 26237 37281 26249 37284
rect 26283 37281 26295 37315
rect 26237 37275 26295 37281
rect 32401 37315 32459 37321
rect 32401 37281 32413 37315
rect 32447 37312 32459 37315
rect 33226 37312 33232 37324
rect 32447 37284 33232 37312
rect 32447 37281 32459 37284
rect 32401 37275 32459 37281
rect 33226 37272 33232 37284
rect 33284 37312 33290 37324
rect 33594 37312 33600 37324
rect 33284 37284 33600 37312
rect 33284 37272 33290 37284
rect 33594 37272 33600 37284
rect 33652 37272 33658 37324
rect 9692 37244 9720 37272
rect 10042 37244 10048 37256
rect 9692 37216 10048 37244
rect 10042 37204 10048 37216
rect 10100 37204 10106 37256
rect 12158 37244 12164 37256
rect 12119 37216 12164 37244
rect 12158 37204 12164 37216
rect 12216 37244 12222 37256
rect 12618 37244 12624 37256
rect 12216 37216 12624 37244
rect 12216 37204 12222 37216
rect 12618 37204 12624 37216
rect 12676 37204 12682 37256
rect 15286 37244 15292 37256
rect 15247 37216 15292 37244
rect 15286 37204 15292 37216
rect 15344 37204 15350 37256
rect 18138 37204 18144 37256
rect 18196 37244 18202 37256
rect 33796 37253 33824 37352
rect 33870 37272 33876 37324
rect 33928 37312 33934 37324
rect 34057 37315 34115 37321
rect 34057 37312 34069 37315
rect 33928 37284 34069 37312
rect 33928 37272 33934 37284
rect 34057 37281 34069 37284
rect 34103 37312 34115 37315
rect 34422 37312 34428 37324
rect 34103 37284 34428 37312
rect 34103 37281 34115 37284
rect 34057 37275 34115 37281
rect 34422 37272 34428 37284
rect 34480 37272 34486 37324
rect 34514 37272 34520 37324
rect 34572 37312 34578 37324
rect 35710 37312 35716 37324
rect 34572 37284 35716 37312
rect 34572 37272 34578 37284
rect 35710 37272 35716 37284
rect 35768 37312 35774 37324
rect 35805 37315 35863 37321
rect 35805 37312 35817 37315
rect 35768 37284 35817 37312
rect 35768 37272 35774 37284
rect 35805 37281 35817 37284
rect 35851 37281 35863 37315
rect 35805 37275 35863 37281
rect 18325 37247 18383 37253
rect 18325 37244 18337 37247
rect 18196 37216 18337 37244
rect 18196 37204 18202 37216
rect 18325 37213 18337 37216
rect 18371 37213 18383 37247
rect 18325 37207 18383 37213
rect 33781 37247 33839 37253
rect 33781 37213 33793 37247
rect 33827 37244 33839 37247
rect 34532 37244 34560 37272
rect 33827 37216 34560 37244
rect 33827 37213 33839 37216
rect 33781 37207 33839 37213
rect 7006 37108 7012 37120
rect 6967 37080 7012 37108
rect 7006 37068 7012 37080
rect 7064 37068 7070 37120
rect 11238 37108 11244 37120
rect 11199 37080 11244 37108
rect 11238 37068 11244 37080
rect 11296 37068 11302 37120
rect 13538 37108 13544 37120
rect 13499 37080 13544 37108
rect 13538 37068 13544 37080
rect 13596 37068 13602 37120
rect 19426 37068 19432 37120
rect 19484 37108 19490 37120
rect 19705 37111 19763 37117
rect 19705 37108 19717 37111
rect 19484 37080 19717 37108
rect 19484 37068 19490 37080
rect 19705 37077 19717 37080
rect 19751 37077 19763 37111
rect 19705 37071 19763 37077
rect 1104 37018 38548 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 38548 37018
rect 1104 36944 38548 36966
rect 1670 36904 1676 36916
rect 1631 36876 1676 36904
rect 1670 36864 1676 36876
rect 1728 36864 1734 36916
rect 2314 36904 2320 36916
rect 2275 36876 2320 36904
rect 2314 36864 2320 36876
rect 2372 36864 2378 36916
rect 5721 36907 5779 36913
rect 5721 36873 5733 36907
rect 5767 36904 5779 36907
rect 5994 36904 6000 36916
rect 5767 36876 6000 36904
rect 5767 36873 5779 36876
rect 5721 36867 5779 36873
rect 5994 36864 6000 36876
rect 6052 36864 6058 36916
rect 9769 36907 9827 36913
rect 9769 36873 9781 36907
rect 9815 36904 9827 36907
rect 9950 36904 9956 36916
rect 9815 36876 9956 36904
rect 9815 36873 9827 36876
rect 9769 36867 9827 36873
rect 9950 36864 9956 36876
rect 10008 36864 10014 36916
rect 10042 36864 10048 36916
rect 10100 36904 10106 36916
rect 10100 36876 10145 36904
rect 10100 36864 10106 36876
rect 11054 36864 11060 36916
rect 11112 36904 11118 36916
rect 12161 36907 12219 36913
rect 12161 36904 12173 36907
rect 11112 36876 12173 36904
rect 11112 36864 11118 36876
rect 12161 36873 12173 36876
rect 12207 36904 12219 36907
rect 12342 36904 12348 36916
rect 12207 36876 12348 36904
rect 12207 36873 12219 36876
rect 12161 36867 12219 36873
rect 12342 36864 12348 36876
rect 12400 36864 12406 36916
rect 12618 36904 12624 36916
rect 12579 36876 12624 36904
rect 12618 36864 12624 36876
rect 12676 36864 12682 36916
rect 15381 36907 15439 36913
rect 15381 36873 15393 36907
rect 15427 36904 15439 36907
rect 15562 36904 15568 36916
rect 15427 36876 15568 36904
rect 15427 36873 15439 36876
rect 15381 36867 15439 36873
rect 15562 36864 15568 36876
rect 15620 36864 15626 36916
rect 18417 36907 18475 36913
rect 18417 36873 18429 36907
rect 18463 36904 18475 36907
rect 18598 36904 18604 36916
rect 18463 36876 18604 36904
rect 18463 36873 18475 36876
rect 18417 36867 18475 36873
rect 18598 36864 18604 36876
rect 18656 36864 18662 36916
rect 26881 36907 26939 36913
rect 26881 36873 26893 36907
rect 26927 36904 26939 36907
rect 27522 36904 27528 36916
rect 26927 36876 27528 36904
rect 26927 36873 26939 36876
rect 26881 36867 26939 36873
rect 27522 36864 27528 36876
rect 27580 36864 27586 36916
rect 33870 36904 33876 36916
rect 33831 36876 33876 36904
rect 33870 36864 33876 36876
rect 33928 36864 33934 36916
rect 34241 36907 34299 36913
rect 34241 36873 34253 36907
rect 34287 36904 34299 36907
rect 34422 36904 34428 36916
rect 34287 36876 34428 36904
rect 34287 36873 34299 36876
rect 34241 36867 34299 36873
rect 34422 36864 34428 36876
rect 34480 36864 34486 36916
rect 35161 36907 35219 36913
rect 35161 36873 35173 36907
rect 35207 36904 35219 36907
rect 36538 36904 36544 36916
rect 35207 36876 36544 36904
rect 35207 36873 35219 36876
rect 35161 36867 35219 36873
rect 36538 36864 36544 36876
rect 36596 36864 36602 36916
rect 2332 36768 2360 36864
rect 1412 36740 2360 36768
rect 1412 36709 1440 36740
rect 5442 36728 5448 36780
rect 5500 36768 5506 36780
rect 5997 36771 6055 36777
rect 5997 36768 6009 36771
rect 5500 36740 6009 36768
rect 5500 36728 5506 36740
rect 5997 36737 6009 36740
rect 6043 36737 6055 36771
rect 5997 36731 6055 36737
rect 19061 36771 19119 36777
rect 19061 36737 19073 36771
rect 19107 36768 19119 36771
rect 19426 36768 19432 36780
rect 19107 36740 19432 36768
rect 19107 36737 19119 36740
rect 19061 36731 19119 36737
rect 19426 36728 19432 36740
rect 19484 36728 19490 36780
rect 25130 36768 25136 36780
rect 25091 36740 25136 36768
rect 25130 36728 25136 36740
rect 25188 36768 25194 36780
rect 25593 36771 25651 36777
rect 25593 36768 25605 36771
rect 25188 36740 25605 36768
rect 25188 36728 25194 36740
rect 25593 36737 25605 36740
rect 25639 36737 25651 36771
rect 35802 36768 35808 36780
rect 35763 36740 35808 36768
rect 25593 36731 25651 36737
rect 35802 36728 35808 36740
rect 35860 36728 35866 36780
rect 1397 36703 1455 36709
rect 1397 36669 1409 36703
rect 1443 36669 1455 36703
rect 1397 36663 1455 36669
rect 1581 36703 1639 36709
rect 1581 36669 1593 36703
rect 1627 36700 1639 36703
rect 1762 36700 1768 36712
rect 1627 36672 1768 36700
rect 1627 36669 1639 36672
rect 1581 36663 1639 36669
rect 1762 36660 1768 36672
rect 1820 36660 1826 36712
rect 18138 36660 18144 36712
rect 18196 36700 18202 36712
rect 19153 36703 19211 36709
rect 19153 36700 19165 36703
rect 18196 36672 19165 36700
rect 18196 36660 18202 36672
rect 19153 36669 19165 36672
rect 19199 36669 19211 36703
rect 19153 36663 19211 36669
rect 25317 36703 25375 36709
rect 25317 36669 25329 36703
rect 25363 36700 25375 36703
rect 26050 36700 26056 36712
rect 25363 36672 26056 36700
rect 25363 36669 25375 36672
rect 25317 36663 25375 36669
rect 20806 36632 20812 36644
rect 20767 36604 20812 36632
rect 20806 36592 20812 36604
rect 20864 36592 20870 36644
rect 25130 36592 25136 36644
rect 25188 36632 25194 36644
rect 25332 36632 25360 36663
rect 26050 36660 26056 36672
rect 26108 36660 26114 36712
rect 35713 36703 35771 36709
rect 35713 36700 35725 36703
rect 35452 36672 35725 36700
rect 25188 36604 25360 36632
rect 25188 36592 25194 36604
rect 35452 36576 35480 36672
rect 35713 36669 35725 36672
rect 35759 36669 35771 36703
rect 36403 36703 36461 36709
rect 36403 36700 36415 36703
rect 35713 36663 35771 36669
rect 35912 36672 36415 36700
rect 35526 36592 35532 36644
rect 35584 36632 35590 36644
rect 35912 36632 35940 36672
rect 36403 36669 36415 36672
rect 36449 36669 36461 36703
rect 36538 36700 36544 36712
rect 36499 36672 36544 36700
rect 36403 36663 36461 36669
rect 36538 36660 36544 36672
rect 36596 36660 36602 36712
rect 35584 36604 35940 36632
rect 35584 36592 35590 36604
rect 15286 36524 15292 36576
rect 15344 36564 15350 36576
rect 15749 36567 15807 36573
rect 15749 36564 15761 36567
rect 15344 36536 15761 36564
rect 15344 36524 15350 36536
rect 15749 36533 15761 36536
rect 15795 36564 15807 36567
rect 16482 36564 16488 36576
rect 15795 36536 16488 36564
rect 15795 36533 15807 36536
rect 15749 36527 15807 36533
rect 16482 36524 16488 36536
rect 16540 36524 16546 36576
rect 35434 36564 35440 36576
rect 35395 36536 35440 36564
rect 35434 36524 35440 36536
rect 35492 36524 35498 36576
rect 1104 36474 38548 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 38548 36474
rect 1104 36400 38548 36422
rect 10042 36320 10048 36372
rect 10100 36360 10106 36372
rect 10413 36363 10471 36369
rect 10413 36360 10425 36363
rect 10100 36332 10425 36360
rect 10100 36320 10106 36332
rect 10413 36329 10425 36332
rect 10459 36329 10471 36363
rect 10413 36323 10471 36329
rect 22830 36320 22836 36372
rect 22888 36360 22894 36372
rect 23014 36360 23020 36372
rect 22888 36332 23020 36360
rect 22888 36320 22894 36332
rect 23014 36320 23020 36332
rect 23072 36320 23078 36372
rect 37458 36320 37464 36372
rect 37516 36360 37522 36372
rect 38654 36360 38660 36372
rect 37516 36332 38660 36360
rect 37516 36320 37522 36332
rect 38654 36320 38660 36332
rect 38712 36320 38718 36372
rect 5166 36224 5172 36236
rect 5127 36196 5172 36224
rect 5166 36184 5172 36196
rect 5224 36184 5230 36236
rect 5442 36184 5448 36236
rect 5500 36184 5506 36236
rect 10594 36224 10600 36236
rect 10555 36196 10600 36224
rect 10594 36184 10600 36196
rect 10652 36184 10658 36236
rect 16393 36227 16451 36233
rect 16393 36193 16405 36227
rect 16439 36224 16451 36227
rect 16482 36224 16488 36236
rect 16439 36196 16488 36224
rect 16439 36193 16451 36196
rect 16393 36187 16451 36193
rect 16482 36184 16488 36196
rect 16540 36184 16546 36236
rect 4893 36159 4951 36165
rect 4893 36125 4905 36159
rect 4939 36156 4951 36159
rect 5460 36156 5488 36184
rect 16666 36156 16672 36168
rect 4939 36128 5488 36156
rect 16627 36128 16672 36156
rect 4939 36125 4951 36128
rect 4893 36119 4951 36125
rect 16666 36116 16672 36128
rect 16724 36116 16730 36168
rect 18046 36156 18052 36168
rect 18007 36128 18052 36156
rect 18046 36116 18052 36128
rect 18104 36116 18110 36168
rect 1673 36023 1731 36029
rect 1673 35989 1685 36023
rect 1719 36020 1731 36023
rect 1762 36020 1768 36032
rect 1719 35992 1768 36020
rect 1719 35989 1731 35992
rect 1673 35983 1731 35989
rect 1762 35980 1768 35992
rect 1820 35980 1826 36032
rect 6457 36023 6515 36029
rect 6457 35989 6469 36023
rect 6503 36020 6515 36023
rect 6914 36020 6920 36032
rect 6503 35992 6920 36020
rect 6503 35989 6515 35992
rect 6457 35983 6515 35989
rect 6914 35980 6920 35992
rect 6972 35980 6978 36032
rect 18138 35980 18144 36032
rect 18196 36020 18202 36032
rect 18325 36023 18383 36029
rect 18325 36020 18337 36023
rect 18196 35992 18337 36020
rect 18196 35980 18202 35992
rect 18325 35989 18337 35992
rect 18371 36020 18383 36023
rect 19153 36023 19211 36029
rect 19153 36020 19165 36023
rect 18371 35992 19165 36020
rect 18371 35989 18383 35992
rect 18325 35983 18383 35989
rect 19153 35989 19165 35992
rect 19199 35989 19211 36023
rect 19153 35983 19211 35989
rect 25130 35980 25136 36032
rect 25188 36020 25194 36032
rect 25317 36023 25375 36029
rect 25317 36020 25329 36023
rect 25188 35992 25329 36020
rect 25188 35980 25194 35992
rect 25317 35989 25329 35992
rect 25363 35989 25375 36023
rect 25317 35983 25375 35989
rect 35526 35980 35532 36032
rect 35584 36020 35590 36032
rect 35621 36023 35679 36029
rect 35621 36020 35633 36023
rect 35584 35992 35633 36020
rect 35584 35980 35590 35992
rect 35621 35989 35633 35992
rect 35667 35989 35679 36023
rect 35621 35983 35679 35989
rect 1104 35930 38548 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 38548 35930
rect 1104 35856 38548 35878
rect 4985 35819 5043 35825
rect 4985 35785 4997 35819
rect 5031 35816 5043 35819
rect 5166 35816 5172 35828
rect 5031 35788 5172 35816
rect 5031 35785 5043 35788
rect 4985 35779 5043 35785
rect 5166 35776 5172 35788
rect 5224 35776 5230 35828
rect 5353 35819 5411 35825
rect 5353 35785 5365 35819
rect 5399 35816 5411 35819
rect 5442 35816 5448 35828
rect 5399 35788 5448 35816
rect 5399 35785 5411 35788
rect 5353 35779 5411 35785
rect 5442 35776 5448 35788
rect 5500 35776 5506 35828
rect 10505 35819 10563 35825
rect 10505 35785 10517 35819
rect 10551 35816 10563 35819
rect 10594 35816 10600 35828
rect 10551 35788 10600 35816
rect 10551 35785 10563 35788
rect 10505 35779 10563 35785
rect 10594 35776 10600 35788
rect 10652 35776 10658 35828
rect 24946 35816 24952 35828
rect 24907 35788 24952 35816
rect 24946 35776 24952 35788
rect 25004 35776 25010 35828
rect 24964 35680 24992 35776
rect 25409 35683 25467 35689
rect 25409 35680 25421 35683
rect 24964 35652 25421 35680
rect 25409 35649 25421 35652
rect 25455 35649 25467 35683
rect 25409 35643 25467 35649
rect 35713 35683 35771 35689
rect 35713 35649 35725 35683
rect 35759 35680 35771 35683
rect 36078 35680 36084 35692
rect 35759 35652 36084 35680
rect 35759 35649 35771 35652
rect 35713 35643 35771 35649
rect 36078 35640 36084 35652
rect 36136 35640 36142 35692
rect 18046 35612 18052 35624
rect 18007 35584 18052 35612
rect 18046 35572 18052 35584
rect 18104 35572 18110 35624
rect 18325 35615 18383 35621
rect 18325 35612 18337 35615
rect 18156 35584 18337 35612
rect 16482 35504 16488 35556
rect 16540 35544 16546 35556
rect 17770 35544 17776 35556
rect 16540 35516 16896 35544
rect 17731 35516 17776 35544
rect 16540 35504 16546 35516
rect 15930 35436 15936 35488
rect 15988 35476 15994 35488
rect 16393 35479 16451 35485
rect 16393 35476 16405 35479
rect 15988 35448 16405 35476
rect 15988 35436 15994 35448
rect 16393 35445 16405 35448
rect 16439 35476 16451 35479
rect 16666 35476 16672 35488
rect 16439 35448 16672 35476
rect 16439 35445 16451 35448
rect 16393 35439 16451 35445
rect 16666 35436 16672 35448
rect 16724 35436 16730 35488
rect 16868 35485 16896 35516
rect 17770 35504 17776 35516
rect 17828 35544 17834 35556
rect 18156 35544 18184 35584
rect 18325 35581 18337 35584
rect 18371 35581 18383 35615
rect 25130 35612 25136 35624
rect 25091 35584 25136 35612
rect 18325 35575 18383 35581
rect 25130 35572 25136 35584
rect 25188 35572 25194 35624
rect 35805 35615 35863 35621
rect 35805 35581 35817 35615
rect 35851 35612 35863 35615
rect 35894 35612 35900 35624
rect 35851 35584 35900 35612
rect 35851 35581 35863 35584
rect 35805 35575 35863 35581
rect 35894 35572 35900 35584
rect 35952 35572 35958 35624
rect 17828 35516 18184 35544
rect 19705 35547 19763 35553
rect 17828 35504 17834 35516
rect 19705 35513 19717 35547
rect 19751 35544 19763 35547
rect 19886 35544 19892 35556
rect 19751 35516 19892 35544
rect 19751 35513 19763 35516
rect 19705 35507 19763 35513
rect 19886 35504 19892 35516
rect 19944 35504 19950 35556
rect 26786 35544 26792 35556
rect 26747 35516 26792 35544
rect 26786 35504 26792 35516
rect 26844 35504 26850 35556
rect 16853 35479 16911 35485
rect 16853 35445 16865 35479
rect 16899 35476 16911 35479
rect 18138 35476 18144 35488
rect 16899 35448 18144 35476
rect 16899 35445 16911 35448
rect 16853 35439 16911 35445
rect 18138 35436 18144 35448
rect 18196 35436 18202 35488
rect 36078 35436 36084 35488
rect 36136 35476 36142 35488
rect 37185 35479 37243 35485
rect 37185 35476 37197 35479
rect 36136 35448 37197 35476
rect 36136 35436 36142 35448
rect 37185 35445 37197 35448
rect 37231 35445 37243 35479
rect 37185 35439 37243 35445
rect 1104 35386 38548 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 38548 35386
rect 1104 35312 38548 35334
rect 10594 35232 10600 35284
rect 10652 35272 10658 35284
rect 11701 35275 11759 35281
rect 11701 35272 11713 35275
rect 10652 35244 11713 35272
rect 10652 35232 10658 35244
rect 11701 35241 11713 35244
rect 11747 35241 11759 35275
rect 11701 35235 11759 35241
rect 11716 35204 11744 35235
rect 29270 35232 29276 35284
rect 29328 35272 29334 35284
rect 29365 35275 29423 35281
rect 29365 35272 29377 35275
rect 29328 35244 29377 35272
rect 29328 35232 29334 35244
rect 29365 35241 29377 35244
rect 29411 35272 29423 35275
rect 30006 35272 30012 35284
rect 29411 35244 30012 35272
rect 29411 35241 29423 35244
rect 29365 35235 29423 35241
rect 30006 35232 30012 35244
rect 30064 35232 30070 35284
rect 13998 35204 14004 35216
rect 11716 35176 14004 35204
rect 13998 35164 14004 35176
rect 14056 35204 14062 35216
rect 14056 35176 14228 35204
rect 14056 35164 14062 35176
rect 6914 35096 6920 35148
rect 6972 35136 6978 35148
rect 7285 35139 7343 35145
rect 7285 35136 7297 35139
rect 6972 35108 7297 35136
rect 6972 35096 6978 35108
rect 7285 35105 7297 35108
rect 7331 35105 7343 35139
rect 11882 35136 11888 35148
rect 11843 35108 11888 35136
rect 7285 35099 7343 35105
rect 11882 35096 11888 35108
rect 11940 35096 11946 35148
rect 14200 35145 14228 35176
rect 14185 35139 14243 35145
rect 14185 35105 14197 35139
rect 14231 35105 14243 35139
rect 14185 35099 14243 35105
rect 7009 35071 7067 35077
rect 7009 35037 7021 35071
rect 7055 35068 7067 35071
rect 7374 35068 7380 35080
rect 7055 35040 7380 35068
rect 7055 35037 7067 35040
rect 7009 35031 7067 35037
rect 7374 35028 7380 35040
rect 7432 35028 7438 35080
rect 8573 34935 8631 34941
rect 8573 34901 8585 34935
rect 8619 34932 8631 34935
rect 9766 34932 9772 34944
rect 8619 34904 9772 34932
rect 8619 34901 8631 34904
rect 8573 34895 8631 34901
rect 9766 34892 9772 34904
rect 9824 34892 9830 34944
rect 14001 34935 14059 34941
rect 14001 34901 14013 34935
rect 14047 34932 14059 34935
rect 14734 34932 14740 34944
rect 14047 34904 14740 34932
rect 14047 34901 14059 34904
rect 14001 34895 14059 34901
rect 14734 34892 14740 34904
rect 14792 34892 14798 34944
rect 18138 34932 18144 34944
rect 18099 34904 18144 34932
rect 18138 34892 18144 34904
rect 18196 34892 18202 34944
rect 24029 34935 24087 34941
rect 24029 34901 24041 34935
rect 24075 34932 24087 34935
rect 24578 34932 24584 34944
rect 24075 34904 24584 34932
rect 24075 34901 24087 34904
rect 24029 34895 24087 34901
rect 24578 34892 24584 34904
rect 24636 34892 24642 34944
rect 25130 34932 25136 34944
rect 25091 34904 25136 34932
rect 25130 34892 25136 34904
rect 25188 34892 25194 34944
rect 35894 34932 35900 34944
rect 35855 34904 35900 34932
rect 35894 34892 35900 34904
rect 35952 34892 35958 34944
rect 1104 34842 38548 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 38548 34842
rect 1104 34768 38548 34790
rect 6914 34688 6920 34740
rect 6972 34728 6978 34740
rect 7009 34731 7067 34737
rect 7009 34728 7021 34731
rect 6972 34700 7021 34728
rect 6972 34688 6978 34700
rect 7009 34697 7021 34700
rect 7055 34697 7067 34731
rect 7374 34728 7380 34740
rect 7335 34700 7380 34728
rect 7009 34691 7067 34697
rect 7374 34688 7380 34700
rect 7432 34688 7438 34740
rect 11054 34688 11060 34740
rect 11112 34728 11118 34740
rect 11793 34731 11851 34737
rect 11793 34728 11805 34731
rect 11112 34700 11805 34728
rect 11112 34688 11118 34700
rect 11793 34697 11805 34700
rect 11839 34728 11851 34731
rect 11882 34728 11888 34740
rect 11839 34700 11888 34728
rect 11839 34697 11851 34700
rect 11793 34691 11851 34697
rect 11882 34688 11888 34700
rect 11940 34688 11946 34740
rect 13998 34728 14004 34740
rect 13959 34700 14004 34728
rect 13998 34688 14004 34700
rect 14056 34688 14062 34740
rect 25130 34688 25136 34740
rect 25188 34728 25194 34740
rect 25869 34731 25927 34737
rect 25869 34728 25881 34731
rect 25188 34700 25881 34728
rect 25188 34688 25194 34700
rect 25869 34697 25881 34700
rect 25915 34697 25927 34731
rect 37366 34728 37372 34740
rect 37327 34700 37372 34728
rect 25869 34691 25927 34697
rect 14734 34592 14740 34604
rect 14647 34564 14740 34592
rect 14734 34552 14740 34564
rect 14792 34592 14798 34604
rect 19705 34595 19763 34601
rect 14792 34564 15148 34592
rect 14792 34552 14798 34564
rect 15013 34527 15071 34533
rect 15013 34524 15025 34527
rect 14568 34496 15025 34524
rect 14568 34468 14596 34496
rect 15013 34493 15025 34496
rect 15059 34493 15071 34527
rect 15120 34524 15148 34564
rect 19705 34561 19717 34595
rect 19751 34592 19763 34595
rect 20070 34592 20076 34604
rect 19751 34564 20076 34592
rect 19751 34561 19763 34564
rect 19705 34555 19763 34561
rect 20070 34552 20076 34564
rect 20128 34552 20134 34604
rect 20898 34552 20904 34604
rect 20956 34592 20962 34604
rect 21177 34595 21235 34601
rect 21177 34592 21189 34595
rect 20956 34564 21189 34592
rect 20956 34552 20962 34564
rect 21177 34561 21189 34564
rect 21223 34561 21235 34595
rect 21177 34555 21235 34561
rect 15286 34524 15292 34536
rect 15120 34496 15292 34524
rect 15013 34487 15071 34493
rect 15286 34484 15292 34496
rect 15344 34484 15350 34536
rect 19426 34484 19432 34536
rect 19484 34524 19490 34536
rect 19797 34527 19855 34533
rect 19797 34524 19809 34527
rect 19484 34496 19809 34524
rect 19484 34484 19490 34496
rect 19797 34493 19809 34496
rect 19843 34493 19855 34527
rect 24578 34524 24584 34536
rect 24539 34496 24584 34524
rect 19797 34487 19855 34493
rect 24578 34484 24584 34496
rect 24636 34484 24642 34536
rect 25884 34524 25912 34691
rect 37366 34688 37372 34700
rect 37424 34688 37430 34740
rect 30650 34660 30656 34672
rect 30611 34632 30656 34660
rect 30650 34620 30656 34632
rect 30708 34620 30714 34672
rect 26329 34595 26387 34601
rect 26329 34561 26341 34595
rect 26375 34592 26387 34595
rect 26697 34595 26755 34601
rect 26697 34592 26709 34595
rect 26375 34564 26709 34592
rect 26375 34561 26387 34564
rect 26329 34555 26387 34561
rect 26697 34561 26709 34564
rect 26743 34592 26755 34595
rect 26878 34592 26884 34604
rect 26743 34564 26884 34592
rect 26743 34561 26755 34564
rect 26697 34555 26755 34561
rect 26878 34552 26884 34564
rect 26936 34552 26942 34604
rect 29089 34595 29147 34601
rect 29089 34561 29101 34595
rect 29135 34592 29147 34595
rect 29549 34595 29607 34601
rect 29549 34592 29561 34595
rect 29135 34564 29561 34592
rect 29135 34561 29147 34564
rect 29089 34555 29147 34561
rect 29549 34561 29561 34564
rect 29595 34592 29607 34595
rect 29914 34592 29920 34604
rect 29595 34564 29920 34592
rect 29595 34561 29607 34564
rect 29549 34555 29607 34561
rect 29914 34552 29920 34564
rect 29972 34552 29978 34604
rect 35713 34595 35771 34601
rect 35713 34561 35725 34595
rect 35759 34592 35771 34595
rect 36078 34592 36084 34604
rect 35759 34564 36084 34592
rect 35759 34561 35771 34564
rect 35713 34555 35771 34561
rect 36078 34552 36084 34564
rect 36136 34552 36142 34604
rect 26421 34527 26479 34533
rect 26421 34524 26433 34527
rect 25884 34496 26433 34524
rect 26421 34493 26433 34496
rect 26467 34524 26479 34527
rect 27154 34524 27160 34536
rect 26467 34496 27160 34524
rect 26467 34493 26479 34496
rect 26421 34487 26479 34493
rect 27154 34484 27160 34496
rect 27212 34484 27218 34536
rect 29270 34524 29276 34536
rect 29231 34496 29276 34524
rect 29270 34484 29276 34496
rect 29328 34484 29334 34536
rect 35805 34527 35863 34533
rect 35805 34493 35817 34527
rect 35851 34524 35863 34527
rect 35894 34524 35900 34536
rect 35851 34496 35900 34524
rect 35851 34493 35863 34496
rect 35805 34487 35863 34493
rect 35894 34484 35900 34496
rect 35952 34484 35958 34536
rect 14550 34456 14556 34468
rect 14511 34428 14556 34456
rect 14550 34416 14556 34428
rect 14608 34416 14614 34468
rect 15102 34348 15108 34400
rect 15160 34388 15166 34400
rect 16117 34391 16175 34397
rect 16117 34388 16129 34391
rect 15160 34360 16129 34388
rect 15160 34348 15166 34360
rect 16117 34357 16129 34360
rect 16163 34388 16175 34391
rect 16482 34388 16488 34400
rect 16163 34360 16488 34388
rect 16163 34357 16175 34360
rect 16117 34351 16175 34357
rect 16482 34348 16488 34360
rect 16540 34348 16546 34400
rect 24394 34388 24400 34400
rect 24355 34360 24400 34388
rect 24394 34348 24400 34360
rect 24452 34348 24458 34400
rect 26418 34348 26424 34400
rect 26476 34388 26482 34400
rect 27801 34391 27859 34397
rect 27801 34388 27813 34391
rect 26476 34360 27813 34388
rect 26476 34348 26482 34360
rect 27801 34357 27813 34360
rect 27847 34357 27859 34391
rect 27801 34351 27859 34357
rect 1104 34298 38548 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 38548 34298
rect 1104 34224 38548 34246
rect 15102 34184 15108 34196
rect 15063 34156 15108 34184
rect 15102 34144 15108 34156
rect 15160 34144 15166 34196
rect 15746 34184 15752 34196
rect 15707 34156 15752 34184
rect 15746 34144 15752 34156
rect 15804 34144 15810 34196
rect 27154 34144 27160 34196
rect 27212 34184 27218 34196
rect 27249 34187 27307 34193
rect 27249 34184 27261 34187
rect 27212 34156 27261 34184
rect 27212 34144 27218 34156
rect 27249 34153 27261 34156
rect 27295 34153 27307 34187
rect 27249 34147 27307 34153
rect 27801 34187 27859 34193
rect 27801 34153 27813 34187
rect 27847 34184 27859 34187
rect 27890 34184 27896 34196
rect 27847 34156 27896 34184
rect 27847 34153 27859 34156
rect 27801 34147 27859 34153
rect 27890 34144 27896 34156
rect 27948 34144 27954 34196
rect 9766 34008 9772 34060
rect 9824 34048 9830 34060
rect 9953 34051 10011 34057
rect 9953 34048 9965 34051
rect 9824 34020 9965 34048
rect 9824 34008 9830 34020
rect 9953 34017 9965 34020
rect 9999 34017 10011 34051
rect 9953 34011 10011 34017
rect 15654 34008 15660 34060
rect 15712 34048 15718 34060
rect 16117 34051 16175 34057
rect 16117 34048 16129 34051
rect 15712 34020 16129 34048
rect 15712 34008 15718 34020
rect 16117 34017 16129 34020
rect 16163 34017 16175 34051
rect 16482 34048 16488 34060
rect 16443 34020 16488 34048
rect 16117 34011 16175 34017
rect 16482 34008 16488 34020
rect 16540 34008 16546 34060
rect 16669 34051 16727 34057
rect 16669 34017 16681 34051
rect 16715 34048 16727 34051
rect 17126 34048 17132 34060
rect 16715 34020 17132 34048
rect 16715 34017 16727 34020
rect 16669 34011 16727 34017
rect 17126 34008 17132 34020
rect 17184 34008 17190 34060
rect 17954 34048 17960 34060
rect 17915 34020 17960 34048
rect 17954 34008 17960 34020
rect 18012 34008 18018 34060
rect 21818 34008 21824 34060
rect 21876 34048 21882 34060
rect 21913 34051 21971 34057
rect 21913 34048 21925 34051
rect 21876 34020 21925 34048
rect 21876 34008 21882 34020
rect 21913 34017 21925 34020
rect 21959 34017 21971 34051
rect 22462 34048 22468 34060
rect 22423 34020 22468 34048
rect 21913 34011 21971 34017
rect 22462 34008 22468 34020
rect 22520 34048 22526 34060
rect 23477 34051 23535 34057
rect 23477 34048 23489 34051
rect 22520 34020 23489 34048
rect 22520 34008 22526 34020
rect 23477 34017 23489 34020
rect 23523 34017 23535 34051
rect 23477 34011 23535 34017
rect 23658 34008 23664 34060
rect 23716 34048 23722 34060
rect 24305 34051 24363 34057
rect 24305 34048 24317 34051
rect 23716 34020 24317 34048
rect 23716 34008 23722 34020
rect 24305 34017 24317 34020
rect 24351 34017 24363 34051
rect 24305 34011 24363 34017
rect 24394 34008 24400 34060
rect 24452 34048 24458 34060
rect 24489 34051 24547 34057
rect 24489 34048 24501 34051
rect 24452 34020 24501 34048
rect 24452 34008 24458 34020
rect 24489 34017 24501 34020
rect 24535 34017 24547 34051
rect 24489 34011 24547 34017
rect 27433 34051 27491 34057
rect 27433 34017 27445 34051
rect 27479 34048 27491 34051
rect 27982 34048 27988 34060
rect 27479 34020 27988 34048
rect 27479 34017 27491 34020
rect 27433 34011 27491 34017
rect 27982 34008 27988 34020
rect 28040 34008 28046 34060
rect 30009 34051 30067 34057
rect 30009 34017 30021 34051
rect 30055 34017 30067 34051
rect 30282 34048 30288 34060
rect 30243 34020 30288 34048
rect 30009 34011 30067 34017
rect 9677 33983 9735 33989
rect 9677 33949 9689 33983
rect 9723 33980 9735 33983
rect 10042 33980 10048 33992
rect 9723 33952 10048 33980
rect 9723 33949 9735 33952
rect 9677 33943 9735 33949
rect 10042 33940 10048 33952
rect 10100 33940 10106 33992
rect 14550 33940 14556 33992
rect 14608 33980 14614 33992
rect 15102 33980 15108 33992
rect 14608 33952 15108 33980
rect 14608 33940 14614 33952
rect 15102 33940 15108 33952
rect 15160 33980 15166 33992
rect 15933 33983 15991 33989
rect 15933 33980 15945 33983
rect 15160 33952 15945 33980
rect 15160 33940 15166 33952
rect 15933 33949 15945 33952
rect 15979 33949 15991 33983
rect 15933 33943 15991 33949
rect 17681 33983 17739 33989
rect 17681 33949 17693 33983
rect 17727 33980 17739 33983
rect 18138 33980 18144 33992
rect 17727 33952 18144 33980
rect 17727 33949 17739 33952
rect 17681 33943 17739 33949
rect 18138 33940 18144 33952
rect 18196 33980 18202 33992
rect 19426 33980 19432 33992
rect 18196 33952 19432 33980
rect 18196 33940 18202 33952
rect 19426 33940 19432 33952
rect 19484 33980 19490 33992
rect 19797 33983 19855 33989
rect 19797 33980 19809 33983
rect 19484 33952 19809 33980
rect 19484 33940 19490 33952
rect 19797 33949 19809 33952
rect 19843 33949 19855 33983
rect 21726 33980 21732 33992
rect 21687 33952 21732 33980
rect 19797 33943 19855 33949
rect 21726 33940 21732 33952
rect 21784 33940 21790 33992
rect 23750 33940 23756 33992
rect 23808 33980 23814 33992
rect 24029 33983 24087 33989
rect 24029 33980 24041 33983
rect 23808 33952 24041 33980
rect 23808 33940 23814 33952
rect 24029 33949 24041 33952
rect 24075 33949 24087 33983
rect 29638 33980 29644 33992
rect 29599 33952 29644 33980
rect 24029 33943 24087 33949
rect 29638 33940 29644 33952
rect 29696 33940 29702 33992
rect 30024 33980 30052 34011
rect 30282 34008 30288 34020
rect 30340 34008 30346 34060
rect 30190 33980 30196 33992
rect 30024 33952 30196 33980
rect 30190 33940 30196 33952
rect 30248 33940 30254 33992
rect 30374 33980 30380 33992
rect 30335 33952 30380 33980
rect 30374 33940 30380 33952
rect 30432 33940 30438 33992
rect 22370 33912 22376 33924
rect 22331 33884 22376 33912
rect 22370 33872 22376 33884
rect 22428 33872 22434 33924
rect 11241 33847 11299 33853
rect 11241 33813 11253 33847
rect 11287 33844 11299 33847
rect 11974 33844 11980 33856
rect 11287 33816 11980 33844
rect 11287 33813 11299 33816
rect 11241 33807 11299 33813
rect 11974 33804 11980 33816
rect 12032 33804 12038 33856
rect 16666 33804 16672 33856
rect 16724 33844 16730 33856
rect 16945 33847 17003 33853
rect 16945 33844 16957 33847
rect 16724 33816 16957 33844
rect 16724 33804 16730 33816
rect 16945 33813 16957 33816
rect 16991 33813 17003 33847
rect 19058 33844 19064 33856
rect 19019 33816 19064 33844
rect 16945 33807 17003 33813
rect 19058 33804 19064 33816
rect 19116 33804 19122 33856
rect 20346 33844 20352 33856
rect 20307 33816 20352 33844
rect 20346 33804 20352 33816
rect 20404 33804 20410 33856
rect 25406 33844 25412 33856
rect 25367 33816 25412 33844
rect 25406 33804 25412 33816
rect 25464 33804 25470 33856
rect 27982 33804 27988 33856
rect 28040 33844 28046 33856
rect 28077 33847 28135 33853
rect 28077 33844 28089 33847
rect 28040 33816 28089 33844
rect 28040 33804 28046 33816
rect 28077 33813 28089 33816
rect 28123 33813 28135 33847
rect 28077 33807 28135 33813
rect 28994 33804 29000 33856
rect 29052 33844 29058 33856
rect 29365 33847 29423 33853
rect 29365 33844 29377 33847
rect 29052 33816 29377 33844
rect 29052 33804 29058 33816
rect 29365 33813 29377 33816
rect 29411 33844 29423 33847
rect 30098 33844 30104 33856
rect 29411 33816 30104 33844
rect 29411 33813 29423 33816
rect 29365 33807 29423 33813
rect 30098 33804 30104 33816
rect 30156 33804 30162 33856
rect 35894 33844 35900 33856
rect 35855 33816 35900 33844
rect 35894 33804 35900 33816
rect 35952 33804 35958 33856
rect 1104 33754 38548 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 38548 33754
rect 1104 33680 38548 33702
rect 9766 33640 9772 33652
rect 9727 33612 9772 33640
rect 9766 33600 9772 33612
rect 9824 33600 9830 33652
rect 10042 33640 10048 33652
rect 10003 33612 10048 33640
rect 10042 33600 10048 33612
rect 10100 33600 10106 33652
rect 14461 33643 14519 33649
rect 14461 33609 14473 33643
rect 14507 33640 14519 33643
rect 14550 33640 14556 33652
rect 14507 33612 14556 33640
rect 14507 33609 14519 33612
rect 14461 33603 14519 33609
rect 14550 33600 14556 33612
rect 14608 33600 14614 33652
rect 16206 33640 16212 33652
rect 16167 33612 16212 33640
rect 16206 33600 16212 33612
rect 16264 33600 16270 33652
rect 17773 33643 17831 33649
rect 17773 33609 17785 33643
rect 17819 33640 17831 33643
rect 17954 33640 17960 33652
rect 17819 33612 17960 33640
rect 17819 33609 17831 33612
rect 17773 33603 17831 33609
rect 17954 33600 17960 33612
rect 18012 33600 18018 33652
rect 21726 33600 21732 33652
rect 21784 33640 21790 33652
rect 22189 33643 22247 33649
rect 22189 33640 22201 33643
rect 21784 33612 22201 33640
rect 21784 33600 21790 33612
rect 22189 33609 22201 33612
rect 22235 33640 22247 33643
rect 24305 33643 24363 33649
rect 24305 33640 24317 33643
rect 22235 33612 24317 33640
rect 22235 33609 22247 33612
rect 22189 33603 22247 33609
rect 24305 33609 24317 33612
rect 24351 33640 24363 33643
rect 24394 33640 24400 33652
rect 24351 33612 24400 33640
rect 24351 33609 24363 33612
rect 24305 33603 24363 33609
rect 24394 33600 24400 33612
rect 24452 33600 24458 33652
rect 26234 33600 26240 33652
rect 26292 33640 26298 33652
rect 26697 33643 26755 33649
rect 26697 33640 26709 33643
rect 26292 33612 26709 33640
rect 26292 33600 26298 33612
rect 26697 33609 26709 33612
rect 26743 33609 26755 33643
rect 26697 33603 26755 33609
rect 22462 33572 22468 33584
rect 22423 33544 22468 33572
rect 22462 33532 22468 33544
rect 22520 33532 22526 33584
rect 16666 33504 16672 33516
rect 16627 33476 16672 33504
rect 16666 33464 16672 33476
rect 16724 33464 16730 33516
rect 20257 33507 20315 33513
rect 20257 33473 20269 33507
rect 20303 33504 20315 33507
rect 20438 33504 20444 33516
rect 20303 33476 20444 33504
rect 20303 33473 20315 33476
rect 20257 33467 20315 33473
rect 20438 33464 20444 33476
rect 20496 33464 20502 33516
rect 20530 33464 20536 33516
rect 20588 33504 20594 33516
rect 25498 33504 25504 33516
rect 20588 33476 20633 33504
rect 25459 33476 25504 33504
rect 20588 33464 20594 33476
rect 25498 33464 25504 33476
rect 25556 33464 25562 33516
rect 26418 33504 26424 33516
rect 26252 33476 26424 33504
rect 14829 33439 14887 33445
rect 14829 33405 14841 33439
rect 14875 33436 14887 33439
rect 16577 33439 16635 33445
rect 16577 33436 16589 33439
rect 14875 33408 16589 33436
rect 14875 33405 14887 33408
rect 14829 33399 14887 33405
rect 16577 33405 16589 33408
rect 16623 33405 16635 33439
rect 16942 33436 16948 33448
rect 16903 33408 16948 33436
rect 16577 33399 16635 33405
rect 16592 33368 16620 33399
rect 16942 33396 16948 33408
rect 17000 33396 17006 33448
rect 17126 33436 17132 33448
rect 17087 33408 17132 33436
rect 17126 33396 17132 33408
rect 17184 33396 17190 33448
rect 20346 33396 20352 33448
rect 20404 33436 20410 33448
rect 21269 33439 21327 33445
rect 21269 33436 21281 33439
rect 20404 33408 21281 33436
rect 20404 33396 20410 33408
rect 21269 33405 21281 33408
rect 21315 33405 21327 33439
rect 21269 33399 21327 33405
rect 21358 33396 21364 33448
rect 21416 33436 21422 33448
rect 22370 33436 22376 33448
rect 21416 33408 22376 33436
rect 21416 33396 21422 33408
rect 22370 33396 22376 33408
rect 22428 33396 22434 33448
rect 25406 33436 25412 33448
rect 25367 33408 25412 33436
rect 25406 33396 25412 33408
rect 25464 33396 25470 33448
rect 26252 33445 26280 33476
rect 26418 33464 26424 33476
rect 26476 33464 26482 33516
rect 26237 33439 26295 33445
rect 26237 33405 26249 33439
rect 26283 33405 26295 33439
rect 26237 33399 26295 33405
rect 26329 33439 26387 33445
rect 26329 33405 26341 33439
rect 26375 33405 26387 33439
rect 26712 33436 26740 33603
rect 27062 33464 27068 33516
rect 27120 33504 27126 33516
rect 27433 33507 27491 33513
rect 27433 33504 27445 33507
rect 27120 33476 27445 33504
rect 27120 33464 27126 33476
rect 27433 33473 27445 33476
rect 27479 33473 27491 33507
rect 27433 33467 27491 33473
rect 27246 33436 27252 33448
rect 26712 33408 27252 33436
rect 26329 33399 26387 33405
rect 17954 33368 17960 33380
rect 16592 33340 17960 33368
rect 17954 33328 17960 33340
rect 18012 33328 18018 33380
rect 23658 33328 23664 33380
rect 23716 33368 23722 33380
rect 23845 33371 23903 33377
rect 23845 33368 23857 33371
rect 23716 33340 23857 33368
rect 23716 33328 23722 33340
rect 23845 33337 23857 33340
rect 23891 33337 23903 33371
rect 23845 33331 23903 33337
rect 24857 33371 24915 33377
rect 24857 33337 24869 33371
rect 24903 33368 24915 33371
rect 26252 33368 26280 33399
rect 24903 33340 26280 33368
rect 26344 33368 26372 33399
rect 27246 33396 27252 33408
rect 27304 33436 27310 33448
rect 27341 33439 27399 33445
rect 27341 33436 27353 33439
rect 27304 33408 27353 33436
rect 27304 33396 27310 33408
rect 27341 33405 27353 33408
rect 27387 33405 27399 33439
rect 27341 33399 27399 33405
rect 27522 33396 27528 33448
rect 27580 33436 27586 33448
rect 27890 33436 27896 33448
rect 27580 33408 27896 33436
rect 27580 33396 27586 33408
rect 27890 33396 27896 33408
rect 27948 33436 27954 33448
rect 28169 33439 28227 33445
rect 28169 33436 28181 33439
rect 27948 33408 28181 33436
rect 27948 33396 27954 33408
rect 28169 33405 28181 33408
rect 28215 33405 28227 33439
rect 28169 33399 28227 33405
rect 28261 33439 28319 33445
rect 28261 33405 28273 33439
rect 28307 33405 28319 33439
rect 28261 33399 28319 33405
rect 29917 33439 29975 33445
rect 29917 33405 29929 33439
rect 29963 33436 29975 33439
rect 30098 33436 30104 33448
rect 29963 33408 30104 33436
rect 29963 33405 29975 33408
rect 29917 33399 29975 33405
rect 28276 33368 28304 33399
rect 30098 33396 30104 33408
rect 30156 33396 30162 33448
rect 30190 33396 30196 33448
rect 30248 33436 30254 33448
rect 30285 33439 30343 33445
rect 30285 33436 30297 33439
rect 30248 33408 30297 33436
rect 30248 33396 30254 33408
rect 30285 33405 30297 33408
rect 30331 33405 30343 33439
rect 30285 33399 30343 33405
rect 26344 33340 28304 33368
rect 29089 33371 29147 33377
rect 24903 33337 24915 33340
rect 24857 33331 24915 33337
rect 15197 33303 15255 33309
rect 15197 33269 15209 33303
rect 15243 33300 15255 33303
rect 15565 33303 15623 33309
rect 15565 33300 15577 33303
rect 15243 33272 15577 33300
rect 15243 33269 15255 33272
rect 15197 33263 15255 33269
rect 15565 33269 15577 33272
rect 15611 33300 15623 33303
rect 17126 33300 17132 33312
rect 15611 33272 17132 33300
rect 15611 33269 15623 33272
rect 15565 33263 15623 33269
rect 17126 33260 17132 33272
rect 17184 33260 17190 33312
rect 18138 33260 18144 33312
rect 18196 33300 18202 33312
rect 18233 33303 18291 33309
rect 18233 33300 18245 33303
rect 18196 33272 18245 33300
rect 18196 33260 18202 33272
rect 18233 33269 18245 33272
rect 18279 33269 18291 33303
rect 19058 33300 19064 33312
rect 19019 33272 19064 33300
rect 18233 33263 18291 33269
rect 19058 33260 19064 33272
rect 19116 33260 19122 33312
rect 21818 33300 21824 33312
rect 21779 33272 21824 33300
rect 21818 33260 21824 33272
rect 21876 33260 21882 33312
rect 23477 33303 23535 33309
rect 23477 33269 23489 33303
rect 23523 33300 23535 33303
rect 23750 33300 23756 33312
rect 23523 33272 23756 33300
rect 23523 33269 23535 33272
rect 23477 33263 23535 33269
rect 23750 33260 23756 33272
rect 23808 33260 23814 33312
rect 25225 33303 25283 33309
rect 25225 33269 25237 33303
rect 25271 33300 25283 33303
rect 26344 33300 26372 33340
rect 27172 33312 27200 33340
rect 29089 33337 29101 33371
rect 29135 33368 29147 33371
rect 29638 33368 29644 33380
rect 29135 33340 29644 33368
rect 29135 33337 29147 33340
rect 29089 33331 29147 33337
rect 29638 33328 29644 33340
rect 29696 33368 29702 33380
rect 30006 33368 30012 33380
rect 29696 33340 30012 33368
rect 29696 33328 29702 33340
rect 30006 33328 30012 33340
rect 30064 33328 30070 33380
rect 27154 33300 27160 33312
rect 25271 33272 26372 33300
rect 27115 33272 27160 33300
rect 25271 33269 25283 33272
rect 25225 33263 25283 33269
rect 27154 33260 27160 33272
rect 27212 33260 27218 33312
rect 28258 33260 28264 33312
rect 28316 33300 28322 33312
rect 28629 33303 28687 33309
rect 28629 33300 28641 33303
rect 28316 33272 28641 33300
rect 28316 33260 28322 33272
rect 28629 33269 28641 33272
rect 28675 33269 28687 33303
rect 30300 33300 30328 33399
rect 32030 33300 32036 33312
rect 30300 33272 32036 33300
rect 28629 33263 28687 33269
rect 32030 33260 32036 33272
rect 32088 33260 32094 33312
rect 1104 33210 38548 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 38548 33210
rect 1104 33136 38548 33158
rect 10873 33099 10931 33105
rect 10873 33065 10885 33099
rect 10919 33096 10931 33099
rect 10962 33096 10968 33108
rect 10919 33068 10968 33096
rect 10919 33065 10931 33068
rect 10873 33059 10931 33065
rect 10962 33056 10968 33068
rect 11020 33056 11026 33108
rect 15105 33099 15163 33105
rect 15105 33065 15117 33099
rect 15151 33096 15163 33099
rect 16942 33096 16948 33108
rect 15151 33068 16948 33096
rect 15151 33065 15163 33068
rect 15105 33059 15163 33065
rect 16942 33056 16948 33068
rect 17000 33096 17006 33108
rect 17129 33099 17187 33105
rect 17129 33096 17141 33099
rect 17000 33068 17141 33096
rect 17000 33056 17006 33068
rect 17129 33065 17141 33068
rect 17175 33065 17187 33099
rect 17129 33059 17187 33065
rect 20441 33099 20499 33105
rect 20441 33065 20453 33099
rect 20487 33096 20499 33099
rect 21358 33096 21364 33108
rect 20487 33068 21364 33096
rect 20487 33065 20499 33068
rect 20441 33059 20499 33065
rect 21358 33056 21364 33068
rect 21416 33056 21422 33108
rect 24578 33056 24584 33108
rect 24636 33096 24642 33108
rect 24949 33099 25007 33105
rect 24949 33096 24961 33099
rect 24636 33068 24961 33096
rect 24636 33056 24642 33068
rect 24949 33065 24961 33068
rect 24995 33096 25007 33099
rect 25406 33096 25412 33108
rect 24995 33068 25412 33096
rect 24995 33065 25007 33068
rect 24949 33059 25007 33065
rect 25406 33056 25412 33068
rect 25464 33056 25470 33108
rect 28166 33056 28172 33108
rect 28224 33096 28230 33108
rect 28261 33099 28319 33105
rect 28261 33096 28273 33099
rect 28224 33068 28273 33096
rect 28224 33056 28230 33068
rect 28261 33065 28273 33068
rect 28307 33096 28319 33099
rect 28902 33096 28908 33108
rect 28307 33068 28908 33096
rect 28307 33065 28319 33068
rect 28261 33059 28319 33065
rect 28902 33056 28908 33068
rect 28960 33056 28966 33108
rect 29270 33056 29276 33108
rect 29328 33096 29334 33108
rect 29917 33099 29975 33105
rect 29917 33096 29929 33099
rect 29328 33068 29929 33096
rect 29328 33056 29334 33068
rect 29917 33065 29929 33068
rect 29963 33065 29975 33099
rect 29917 33059 29975 33065
rect 15470 32988 15476 33040
rect 15528 33028 15534 33040
rect 15565 33031 15623 33037
rect 15565 33028 15577 33031
rect 15528 33000 15577 33028
rect 15528 32988 15534 33000
rect 15565 32997 15577 33000
rect 15611 33028 15623 33031
rect 15654 33028 15660 33040
rect 15611 33000 15660 33028
rect 15611 32997 15623 33000
rect 15565 32991 15623 32997
rect 15654 32988 15660 33000
rect 15712 32988 15718 33040
rect 19981 33031 20039 33037
rect 19981 32997 19993 33031
rect 20027 33028 20039 33031
rect 20346 33028 20352 33040
rect 20027 33000 20352 33028
rect 20027 32997 20039 33000
rect 19981 32991 20039 32997
rect 20346 32988 20352 33000
rect 20404 32988 20410 33040
rect 29549 33031 29607 33037
rect 29549 32997 29561 33031
rect 29595 33028 29607 33031
rect 30193 33031 30251 33037
rect 30193 33028 30205 33031
rect 29595 33000 30205 33028
rect 29595 32997 29607 33000
rect 29549 32991 29607 32997
rect 30193 32997 30205 33000
rect 30239 33028 30251 33031
rect 30282 33028 30288 33040
rect 30239 33000 30288 33028
rect 30239 32997 30251 33000
rect 30193 32991 30251 32997
rect 30282 32988 30288 33000
rect 30340 32988 30346 33040
rect 6086 32920 6092 32972
rect 6144 32960 6150 32972
rect 6273 32963 6331 32969
rect 6273 32960 6285 32963
rect 6144 32932 6285 32960
rect 6144 32920 6150 32932
rect 6273 32929 6285 32932
rect 6319 32929 6331 32963
rect 11054 32960 11060 32972
rect 11015 32932 11060 32960
rect 6273 32923 6331 32929
rect 11054 32920 11060 32932
rect 11112 32920 11118 32972
rect 15838 32920 15844 32972
rect 15896 32960 15902 32972
rect 16025 32963 16083 32969
rect 16025 32960 16037 32963
rect 15896 32932 16037 32960
rect 15896 32920 15902 32932
rect 16025 32929 16037 32932
rect 16071 32960 16083 32963
rect 16666 32960 16672 32972
rect 16071 32932 16672 32960
rect 16071 32929 16083 32932
rect 16025 32923 16083 32929
rect 16666 32920 16672 32932
rect 16724 32920 16730 32972
rect 24946 32960 24952 32972
rect 21652 32932 22048 32960
rect 24907 32932 24952 32960
rect 5997 32895 6055 32901
rect 5997 32861 6009 32895
rect 6043 32892 6055 32895
rect 6362 32892 6368 32904
rect 6043 32864 6368 32892
rect 6043 32861 6055 32864
rect 5997 32855 6055 32861
rect 6362 32852 6368 32864
rect 6420 32852 6426 32904
rect 12618 32892 12624 32904
rect 12579 32864 12624 32892
rect 12618 32852 12624 32864
rect 12676 32852 12682 32904
rect 12802 32852 12808 32904
rect 12860 32892 12866 32904
rect 12897 32895 12955 32901
rect 12897 32892 12909 32895
rect 12860 32864 12909 32892
rect 12860 32852 12866 32864
rect 12897 32861 12909 32864
rect 12943 32861 12955 32895
rect 12897 32855 12955 32861
rect 15654 32852 15660 32904
rect 15712 32892 15718 32904
rect 15749 32895 15807 32901
rect 15749 32892 15761 32895
rect 15712 32864 15761 32892
rect 15712 32852 15718 32864
rect 15749 32861 15761 32864
rect 15795 32892 15807 32895
rect 16482 32892 16488 32904
rect 15795 32864 16488 32892
rect 15795 32861 15807 32864
rect 15749 32855 15807 32861
rect 16482 32852 16488 32864
rect 16540 32852 16546 32904
rect 18138 32852 18144 32904
rect 18196 32892 18202 32904
rect 18325 32895 18383 32901
rect 18325 32892 18337 32895
rect 18196 32864 18337 32892
rect 18196 32852 18202 32864
rect 18325 32861 18337 32864
rect 18371 32861 18383 32895
rect 18598 32892 18604 32904
rect 18559 32864 18604 32892
rect 18325 32855 18383 32861
rect 18598 32852 18604 32864
rect 18656 32852 18662 32904
rect 21358 32852 21364 32904
rect 21416 32892 21422 32904
rect 21652 32901 21680 32932
rect 21637 32895 21695 32901
rect 21637 32892 21649 32895
rect 21416 32864 21649 32892
rect 21416 32852 21422 32864
rect 21637 32861 21649 32864
rect 21683 32861 21695 32895
rect 21910 32892 21916 32904
rect 21871 32864 21916 32892
rect 21637 32855 21695 32861
rect 21910 32852 21916 32864
rect 21968 32852 21974 32904
rect 22020 32892 22048 32932
rect 24946 32920 24952 32932
rect 25004 32920 25010 32972
rect 25314 32920 25320 32972
rect 25372 32960 25378 32972
rect 25409 32963 25467 32969
rect 25409 32960 25421 32963
rect 25372 32932 25421 32960
rect 25372 32920 25378 32932
rect 25409 32929 25421 32932
rect 25455 32960 25467 32963
rect 26513 32963 26571 32969
rect 26513 32960 26525 32963
rect 25455 32932 26525 32960
rect 25455 32929 25467 32932
rect 25409 32923 25467 32929
rect 26513 32929 26525 32932
rect 26559 32929 26571 32963
rect 26970 32960 26976 32972
rect 26931 32932 26976 32960
rect 26513 32923 26571 32929
rect 26970 32920 26976 32932
rect 27028 32920 27034 32972
rect 27338 32960 27344 32972
rect 27299 32932 27344 32960
rect 27338 32920 27344 32932
rect 27396 32920 27402 32972
rect 28350 32960 28356 32972
rect 28311 32932 28356 32960
rect 28350 32920 28356 32932
rect 28408 32920 28414 32972
rect 28905 32963 28963 32969
rect 28905 32929 28917 32963
rect 28951 32960 28963 32963
rect 28994 32960 29000 32972
rect 28951 32932 29000 32960
rect 28951 32929 28963 32932
rect 28905 32923 28963 32929
rect 28994 32920 29000 32932
rect 29052 32920 29058 32972
rect 30098 32960 30104 32972
rect 30059 32932 30104 32960
rect 30098 32920 30104 32932
rect 30156 32920 30162 32972
rect 31021 32963 31079 32969
rect 31021 32960 31033 32963
rect 30576 32932 31033 32960
rect 30576 32904 30604 32932
rect 31021 32929 31033 32932
rect 31067 32929 31079 32963
rect 31021 32923 31079 32929
rect 23290 32892 23296 32904
rect 22020 32864 23296 32892
rect 23290 32852 23296 32864
rect 23348 32852 23354 32904
rect 27430 32892 27436 32904
rect 27391 32864 27436 32892
rect 27430 32852 27436 32864
rect 27488 32852 27494 32904
rect 28813 32895 28871 32901
rect 28813 32861 28825 32895
rect 28859 32861 28871 32895
rect 28813 32855 28871 32861
rect 27246 32784 27252 32836
rect 27304 32824 27310 32836
rect 28828 32824 28856 32855
rect 29822 32852 29828 32904
rect 29880 32892 29886 32904
rect 30558 32892 30564 32904
rect 29880 32864 30564 32892
rect 29880 32852 29886 32864
rect 30558 32852 30564 32864
rect 30616 32852 30622 32904
rect 30742 32892 30748 32904
rect 30703 32864 30748 32892
rect 30742 32852 30748 32864
rect 30800 32852 30806 32904
rect 31202 32892 31208 32904
rect 31163 32864 31208 32892
rect 31202 32852 31208 32864
rect 31260 32852 31266 32904
rect 27304 32796 28856 32824
rect 27304 32784 27310 32796
rect 7561 32759 7619 32765
rect 7561 32725 7573 32759
rect 7607 32756 7619 32759
rect 7926 32756 7932 32768
rect 7607 32728 7932 32756
rect 7607 32725 7619 32728
rect 7561 32719 7619 32725
rect 7926 32716 7932 32728
rect 7984 32716 7990 32768
rect 13998 32756 14004 32768
rect 13959 32728 14004 32756
rect 13998 32716 14004 32728
rect 14056 32716 14062 32768
rect 23201 32759 23259 32765
rect 23201 32725 23213 32759
rect 23247 32756 23259 32759
rect 23290 32756 23296 32768
rect 23247 32728 23296 32756
rect 23247 32725 23259 32728
rect 23201 32719 23259 32725
rect 23290 32716 23296 32728
rect 23348 32716 23354 32768
rect 27798 32756 27804 32768
rect 27759 32728 27804 32756
rect 27798 32716 27804 32728
rect 27856 32716 27862 32768
rect 1104 32666 38548 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 38548 32666
rect 1104 32592 38548 32614
rect 5994 32552 6000 32564
rect 5955 32524 6000 32552
rect 5994 32512 6000 32524
rect 6052 32512 6058 32564
rect 6362 32552 6368 32564
rect 6323 32524 6368 32552
rect 6362 32512 6368 32524
rect 6420 32512 6426 32564
rect 12253 32555 12311 32561
rect 12253 32521 12265 32555
rect 12299 32552 12311 32555
rect 12618 32552 12624 32564
rect 12299 32524 12624 32552
rect 12299 32521 12311 32524
rect 12253 32515 12311 32521
rect 12618 32512 12624 32524
rect 12676 32512 12682 32564
rect 16482 32512 16488 32564
rect 16540 32552 16546 32564
rect 16669 32555 16727 32561
rect 16669 32552 16681 32555
rect 16540 32524 16681 32552
rect 16540 32512 16546 32524
rect 16669 32521 16681 32524
rect 16715 32521 16727 32555
rect 16669 32515 16727 32521
rect 15657 32487 15715 32493
rect 15657 32453 15669 32487
rect 15703 32484 15715 32487
rect 16298 32484 16304 32496
rect 15703 32456 16304 32484
rect 15703 32453 15715 32456
rect 15657 32447 15715 32453
rect 16298 32444 16304 32456
rect 16356 32444 16362 32496
rect 16684 32484 16712 32515
rect 17678 32512 17684 32564
rect 17736 32552 17742 32564
rect 17954 32552 17960 32564
rect 17736 32524 17960 32552
rect 17736 32512 17742 32524
rect 17954 32512 17960 32524
rect 18012 32552 18018 32564
rect 18233 32555 18291 32561
rect 18233 32552 18245 32555
rect 18012 32524 18245 32552
rect 18012 32512 18018 32524
rect 18233 32521 18245 32524
rect 18279 32521 18291 32555
rect 18966 32552 18972 32564
rect 18927 32524 18972 32552
rect 18233 32515 18291 32521
rect 18966 32512 18972 32524
rect 19024 32512 19030 32564
rect 21729 32555 21787 32561
rect 21729 32521 21741 32555
rect 21775 32552 21787 32555
rect 21910 32552 21916 32564
rect 21775 32524 21916 32552
rect 21775 32521 21787 32524
rect 21729 32515 21787 32521
rect 21910 32512 21916 32524
rect 21968 32512 21974 32564
rect 25314 32552 25320 32564
rect 25275 32524 25320 32552
rect 25314 32512 25320 32524
rect 25372 32512 25378 32564
rect 25869 32555 25927 32561
rect 25869 32521 25881 32555
rect 25915 32552 25927 32555
rect 27338 32552 27344 32564
rect 25915 32524 27344 32552
rect 25915 32521 25927 32524
rect 25869 32515 25927 32521
rect 27338 32512 27344 32524
rect 27396 32512 27402 32564
rect 28350 32512 28356 32564
rect 28408 32552 28414 32564
rect 28629 32555 28687 32561
rect 28629 32552 28641 32555
rect 28408 32524 28641 32552
rect 28408 32512 28414 32524
rect 28629 32521 28641 32524
rect 28675 32552 28687 32555
rect 29546 32552 29552 32564
rect 28675 32524 29552 32552
rect 28675 32521 28687 32524
rect 28629 32515 28687 32521
rect 29546 32512 29552 32524
rect 29604 32552 29610 32564
rect 29641 32555 29699 32561
rect 29641 32552 29653 32555
rect 29604 32524 29653 32552
rect 29604 32512 29610 32524
rect 29641 32521 29653 32524
rect 29687 32521 29699 32555
rect 29641 32515 29699 32521
rect 29822 32512 29828 32564
rect 29880 32552 29886 32564
rect 30009 32555 30067 32561
rect 30009 32552 30021 32555
rect 29880 32524 30021 32552
rect 29880 32512 29886 32524
rect 30009 32521 30021 32524
rect 30055 32521 30067 32555
rect 30009 32515 30067 32521
rect 30098 32512 30104 32564
rect 30156 32552 30162 32564
rect 31573 32555 31631 32561
rect 31573 32552 31585 32555
rect 30156 32524 31585 32552
rect 30156 32512 30162 32524
rect 31573 32521 31585 32524
rect 31619 32521 31631 32555
rect 31573 32515 31631 32521
rect 17773 32487 17831 32493
rect 17773 32484 17785 32487
rect 16684 32456 17785 32484
rect 17773 32453 17785 32456
rect 17819 32484 17831 32487
rect 18138 32484 18144 32496
rect 17819 32456 18144 32484
rect 17819 32453 17831 32456
rect 17773 32447 17831 32453
rect 18138 32444 18144 32456
rect 18196 32444 18202 32496
rect 25222 32484 25228 32496
rect 21928 32456 25228 32484
rect 13541 32419 13599 32425
rect 13541 32385 13553 32419
rect 13587 32416 13599 32419
rect 13722 32416 13728 32428
rect 13587 32388 13728 32416
rect 13587 32385 13599 32388
rect 13541 32379 13599 32385
rect 13722 32376 13728 32388
rect 13780 32376 13786 32428
rect 19334 32376 19340 32428
rect 19392 32416 19398 32428
rect 21928 32416 21956 32456
rect 25222 32444 25228 32456
rect 25280 32444 25286 32496
rect 27617 32487 27675 32493
rect 27617 32453 27629 32487
rect 27663 32484 27675 32487
rect 28994 32484 29000 32496
rect 27663 32456 29000 32484
rect 27663 32453 27675 32456
rect 27617 32447 27675 32453
rect 28994 32444 29000 32456
rect 29052 32444 29058 32496
rect 23750 32416 23756 32428
rect 19392 32388 21956 32416
rect 23711 32388 23756 32416
rect 19392 32376 19398 32388
rect 23750 32376 23756 32388
rect 23808 32376 23814 32428
rect 13630 32308 13636 32360
rect 13688 32348 13694 32360
rect 14001 32351 14059 32357
rect 14001 32348 14013 32351
rect 13688 32320 14013 32348
rect 13688 32308 13694 32320
rect 14001 32317 14013 32320
rect 14047 32317 14059 32351
rect 14001 32311 14059 32317
rect 14185 32351 14243 32357
rect 14185 32317 14197 32351
rect 14231 32317 14243 32351
rect 14185 32311 14243 32317
rect 14369 32351 14427 32357
rect 14369 32317 14381 32351
rect 14415 32317 14427 32351
rect 14369 32311 14427 32317
rect 14921 32351 14979 32357
rect 14921 32317 14933 32351
rect 14967 32348 14979 32351
rect 15286 32348 15292 32360
rect 14967 32320 15292 32348
rect 14967 32317 14979 32320
rect 14921 32311 14979 32317
rect 14200 32280 14228 32311
rect 13004 32252 14228 32280
rect 14384 32280 14412 32311
rect 15286 32308 15292 32320
rect 15344 32348 15350 32360
rect 15841 32351 15899 32357
rect 15841 32348 15853 32351
rect 15344 32320 15853 32348
rect 15344 32308 15350 32320
rect 15841 32317 15853 32320
rect 15887 32317 15899 32351
rect 16022 32348 16028 32360
rect 15983 32320 16028 32348
rect 15841 32311 15899 32317
rect 16022 32308 16028 32320
rect 16080 32308 16086 32360
rect 16209 32351 16267 32357
rect 16209 32317 16221 32351
rect 16255 32317 16267 32351
rect 16209 32311 16267 32317
rect 18049 32351 18107 32357
rect 18049 32317 18061 32351
rect 18095 32348 18107 32351
rect 18414 32348 18420 32360
rect 18095 32320 18420 32348
rect 18095 32317 18107 32320
rect 18049 32311 18107 32317
rect 15197 32283 15255 32289
rect 15197 32280 15209 32283
rect 14384 32252 15209 32280
rect 10965 32215 11023 32221
rect 10965 32181 10977 32215
rect 11011 32212 11023 32215
rect 11054 32212 11060 32224
rect 11011 32184 11060 32212
rect 11011 32181 11023 32184
rect 10965 32175 11023 32181
rect 11054 32172 11060 32184
rect 11112 32172 11118 32224
rect 12713 32215 12771 32221
rect 12713 32181 12725 32215
rect 12759 32212 12771 32215
rect 12802 32212 12808 32224
rect 12759 32184 12808 32212
rect 12759 32181 12771 32184
rect 12713 32175 12771 32181
rect 12802 32172 12808 32184
rect 12860 32212 12866 32224
rect 13004 32221 13032 32252
rect 12989 32215 13047 32221
rect 12989 32212 13001 32215
rect 12860 32184 13001 32212
rect 12860 32172 12866 32184
rect 12989 32181 13001 32184
rect 13035 32181 13047 32215
rect 13354 32212 13360 32224
rect 13315 32184 13360 32212
rect 12989 32175 13047 32181
rect 13354 32172 13360 32184
rect 13412 32212 13418 32224
rect 14384 32212 14412 32252
rect 15197 32249 15209 32252
rect 15243 32249 15255 32283
rect 15197 32243 15255 32249
rect 13412 32184 14412 32212
rect 15212 32212 15240 32243
rect 16224 32212 16252 32311
rect 18414 32308 18420 32320
rect 18472 32348 18478 32360
rect 18966 32348 18972 32360
rect 18472 32320 18972 32348
rect 18472 32308 18478 32320
rect 18966 32308 18972 32320
rect 19024 32308 19030 32360
rect 19058 32308 19064 32360
rect 19116 32348 19122 32360
rect 23477 32351 23535 32357
rect 19116 32320 19209 32348
rect 19116 32308 19122 32320
rect 23477 32317 23489 32351
rect 23523 32348 23535 32351
rect 24397 32351 24455 32357
rect 24397 32348 24409 32351
rect 23523 32320 24409 32348
rect 23523 32317 23535 32320
rect 23477 32311 23535 32317
rect 24397 32317 24409 32320
rect 24443 32348 24455 32351
rect 26237 32351 26295 32357
rect 24443 32320 24992 32348
rect 24443 32317 24455 32320
rect 24397 32311 24455 32317
rect 17954 32240 17960 32292
rect 18012 32280 18018 32292
rect 18509 32283 18567 32289
rect 18509 32280 18521 32283
rect 18012 32252 18521 32280
rect 18012 32240 18018 32252
rect 18509 32249 18521 32252
rect 18555 32280 18567 32283
rect 18598 32280 18604 32292
rect 18555 32252 18604 32280
rect 18555 32249 18567 32252
rect 18509 32243 18567 32249
rect 18598 32240 18604 32252
rect 18656 32240 18662 32292
rect 19076 32280 19104 32308
rect 18984 32252 19104 32280
rect 15212 32184 16252 32212
rect 13412 32172 13418 32184
rect 18138 32172 18144 32224
rect 18196 32212 18202 32224
rect 18984 32212 19012 32252
rect 24964 32224 24992 32320
rect 26237 32317 26249 32351
rect 26283 32348 26295 32351
rect 26970 32348 26976 32360
rect 26283 32320 26976 32348
rect 26283 32317 26295 32320
rect 26237 32311 26295 32317
rect 26970 32308 26976 32320
rect 27028 32308 27034 32360
rect 27798 32348 27804 32360
rect 27759 32320 27804 32348
rect 27798 32308 27804 32320
rect 27856 32308 27862 32360
rect 28166 32348 28172 32360
rect 28127 32320 28172 32348
rect 28166 32308 28172 32320
rect 28224 32308 28230 32360
rect 28261 32351 28319 32357
rect 28261 32317 28273 32351
rect 28307 32348 28319 32351
rect 28718 32348 28724 32360
rect 28307 32320 28724 32348
rect 28307 32317 28319 32320
rect 28261 32311 28319 32317
rect 26605 32283 26663 32289
rect 26605 32249 26617 32283
rect 26651 32280 26663 32283
rect 27249 32283 27307 32289
rect 27249 32280 27261 32283
rect 26651 32252 27261 32280
rect 26651 32249 26663 32252
rect 26605 32243 26663 32249
rect 27249 32249 27261 32252
rect 27295 32280 27307 32283
rect 27430 32280 27436 32292
rect 27295 32252 27436 32280
rect 27295 32249 27307 32252
rect 27249 32243 27307 32249
rect 27430 32240 27436 32252
rect 27488 32280 27494 32292
rect 28276 32280 28304 32311
rect 28718 32308 28724 32320
rect 28776 32308 28782 32360
rect 29546 32308 29552 32360
rect 29604 32348 29610 32360
rect 30285 32351 30343 32357
rect 30285 32348 30297 32351
rect 29604 32320 30297 32348
rect 29604 32308 29610 32320
rect 30285 32317 30297 32320
rect 30331 32317 30343 32351
rect 30285 32311 30343 32317
rect 27488 32252 28304 32280
rect 27488 32240 27494 32252
rect 30742 32240 30748 32292
rect 30800 32280 30806 32292
rect 30929 32283 30987 32289
rect 30929 32280 30941 32283
rect 30800 32252 30941 32280
rect 30800 32240 30806 32252
rect 30929 32249 30941 32252
rect 30975 32249 30987 32283
rect 30929 32243 30987 32249
rect 18196 32184 19012 32212
rect 18196 32172 18202 32184
rect 20070 32172 20076 32224
rect 20128 32212 20134 32224
rect 20441 32215 20499 32221
rect 20441 32212 20453 32215
rect 20128 32184 20453 32212
rect 20128 32172 20134 32184
rect 20441 32181 20453 32184
rect 20487 32181 20499 32215
rect 20441 32175 20499 32181
rect 21358 32172 21364 32224
rect 21416 32212 21422 32224
rect 22005 32215 22063 32221
rect 22005 32212 22017 32215
rect 21416 32184 22017 32212
rect 21416 32172 21422 32184
rect 22005 32181 22017 32184
rect 22051 32181 22063 32215
rect 24946 32212 24952 32224
rect 24907 32184 24952 32212
rect 22005 32175 22063 32181
rect 24946 32172 24952 32184
rect 25004 32172 25010 32224
rect 30944 32212 30972 32243
rect 31297 32215 31355 32221
rect 31297 32212 31309 32215
rect 30944 32184 31309 32212
rect 31297 32181 31309 32184
rect 31343 32212 31355 32215
rect 31386 32212 31392 32224
rect 31343 32184 31392 32212
rect 31343 32181 31355 32184
rect 31297 32175 31355 32181
rect 31386 32172 31392 32184
rect 31444 32172 31450 32224
rect 1104 32122 38548 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 38548 32122
rect 1104 32048 38548 32070
rect 13630 32008 13636 32020
rect 13591 31980 13636 32008
rect 13630 31968 13636 31980
rect 13688 32008 13694 32020
rect 13688 31980 14412 32008
rect 13688 31968 13694 31980
rect 14384 31949 14412 31980
rect 15378 31968 15384 32020
rect 15436 32008 15442 32020
rect 16022 32008 16028 32020
rect 15436 31980 16028 32008
rect 15436 31968 15442 31980
rect 16022 31968 16028 31980
rect 16080 32008 16086 32020
rect 16117 32011 16175 32017
rect 16117 32008 16129 32011
rect 16080 31980 16129 32008
rect 16080 31968 16086 31980
rect 16117 31977 16129 31980
rect 16163 31977 16175 32011
rect 16117 31971 16175 31977
rect 18506 31968 18512 32020
rect 18564 32008 18570 32020
rect 18601 32011 18659 32017
rect 18601 32008 18613 32011
rect 18564 31980 18613 32008
rect 18564 31968 18570 31980
rect 18601 31977 18613 31980
rect 18647 31977 18659 32011
rect 18601 31971 18659 31977
rect 19153 32011 19211 32017
rect 19153 31977 19165 32011
rect 19199 32008 19211 32011
rect 19334 32008 19340 32020
rect 19199 31980 19340 32008
rect 19199 31977 19211 31980
rect 19153 31971 19211 31977
rect 19334 31968 19340 31980
rect 19392 31968 19398 32020
rect 19426 31968 19432 32020
rect 19484 32008 19490 32020
rect 19613 32011 19671 32017
rect 19613 32008 19625 32011
rect 19484 31980 19625 32008
rect 19484 31968 19490 31980
rect 19613 31977 19625 31980
rect 19659 31977 19671 32011
rect 19613 31971 19671 31977
rect 26329 32011 26387 32017
rect 26329 31977 26341 32011
rect 26375 32008 26387 32011
rect 26418 32008 26424 32020
rect 26375 31980 26424 32008
rect 26375 31977 26387 31980
rect 26329 31971 26387 31977
rect 26418 31968 26424 31980
rect 26476 32008 26482 32020
rect 26476 31980 26924 32008
rect 26476 31968 26482 31980
rect 14369 31943 14427 31949
rect 14369 31909 14381 31943
rect 14415 31909 14427 31943
rect 15746 31940 15752 31952
rect 15707 31912 15752 31940
rect 14369 31903 14427 31909
rect 15746 31900 15752 31912
rect 15804 31900 15810 31952
rect 16574 31940 16580 31952
rect 16535 31912 16580 31940
rect 16574 31900 16580 31912
rect 16632 31900 16638 31952
rect 17494 31900 17500 31952
rect 17552 31940 17558 31952
rect 18138 31940 18144 31952
rect 17552 31912 18144 31940
rect 17552 31900 17558 31912
rect 18138 31900 18144 31912
rect 18196 31900 18202 31952
rect 24394 31940 24400 31952
rect 24307 31912 24400 31940
rect 24394 31900 24400 31912
rect 24452 31940 24458 31952
rect 26896 31949 26924 31980
rect 27982 31968 27988 32020
rect 28040 32008 28046 32020
rect 28077 32011 28135 32017
rect 28077 32008 28089 32011
rect 28040 31980 28089 32008
rect 28040 31968 28046 31980
rect 28077 31977 28089 31980
rect 28123 32008 28135 32011
rect 28123 31980 29132 32008
rect 28123 31977 28135 31980
rect 28077 31971 28135 31977
rect 26881 31943 26939 31949
rect 24452 31912 25544 31940
rect 24452 31900 24458 31912
rect 25516 31884 25544 31912
rect 26881 31909 26893 31943
rect 26927 31909 26939 31943
rect 26881 31903 26939 31909
rect 26970 31900 26976 31952
rect 27028 31940 27034 31952
rect 27249 31943 27307 31949
rect 27249 31940 27261 31943
rect 27028 31912 27261 31940
rect 27028 31900 27034 31912
rect 27249 31909 27261 31912
rect 27295 31909 27307 31943
rect 27249 31903 27307 31909
rect 28718 31900 28724 31952
rect 28776 31940 28782 31952
rect 29104 31940 29132 31980
rect 30006 31968 30012 32020
rect 30064 32008 30070 32020
rect 30285 32011 30343 32017
rect 30285 32008 30297 32011
rect 30064 31980 30297 32008
rect 30064 31968 30070 31980
rect 30285 31977 30297 31980
rect 30331 32008 30343 32011
rect 31202 32008 31208 32020
rect 30331 31980 31208 32008
rect 30331 31977 30343 31980
rect 30285 31971 30343 31977
rect 31202 31968 31208 31980
rect 31260 31968 31266 32020
rect 30098 31940 30104 31952
rect 28776 31912 29040 31940
rect 29104 31912 30104 31940
rect 28776 31900 28782 31912
rect 13909 31875 13967 31881
rect 13909 31841 13921 31875
rect 13955 31872 13967 31875
rect 13998 31872 14004 31884
rect 13955 31844 14004 31872
rect 13955 31841 13967 31844
rect 13909 31835 13967 31841
rect 13998 31832 14004 31844
rect 14056 31832 14062 31884
rect 17034 31872 17040 31884
rect 16995 31844 17040 31872
rect 17034 31832 17040 31844
rect 17092 31832 17098 31884
rect 17218 31872 17224 31884
rect 17179 31844 17224 31872
rect 17218 31832 17224 31844
rect 17276 31832 17282 31884
rect 17405 31875 17463 31881
rect 17405 31841 17417 31875
rect 17451 31841 17463 31875
rect 18414 31872 18420 31884
rect 18375 31844 18420 31872
rect 17405 31835 17463 31841
rect 13814 31804 13820 31816
rect 13775 31776 13820 31804
rect 13814 31764 13820 31776
rect 13872 31764 13878 31816
rect 16390 31764 16396 31816
rect 16448 31804 16454 31816
rect 17420 31804 17448 31835
rect 18414 31832 18420 31844
rect 18472 31832 18478 31884
rect 19334 31832 19340 31884
rect 19392 31872 19398 31884
rect 19429 31875 19487 31881
rect 19429 31872 19441 31875
rect 19392 31844 19441 31872
rect 19392 31832 19398 31844
rect 19429 31841 19441 31844
rect 19475 31841 19487 31875
rect 24670 31872 24676 31884
rect 24631 31844 24676 31872
rect 19429 31835 19487 31841
rect 24670 31832 24676 31844
rect 24728 31832 24734 31884
rect 25406 31872 25412 31884
rect 25367 31844 25412 31872
rect 25406 31832 25412 31844
rect 25464 31832 25470 31884
rect 25498 31832 25504 31884
rect 25556 31872 25562 31884
rect 26694 31872 26700 31884
rect 25556 31844 25601 31872
rect 26655 31844 26700 31872
rect 25556 31832 25562 31844
rect 26694 31832 26700 31844
rect 26752 31832 26758 31884
rect 26789 31875 26847 31881
rect 26789 31841 26801 31875
rect 26835 31872 26847 31875
rect 27430 31872 27436 31884
rect 26835 31844 27436 31872
rect 26835 31841 26847 31844
rect 26789 31835 26847 31841
rect 27430 31832 27436 31844
rect 27488 31872 27494 31884
rect 27893 31875 27951 31881
rect 27893 31872 27905 31875
rect 27488 31844 27905 31872
rect 27488 31832 27494 31844
rect 27893 31841 27905 31844
rect 27939 31841 27951 31875
rect 28258 31872 28264 31884
rect 28219 31844 28264 31872
rect 27893 31835 27951 31841
rect 28258 31832 28264 31844
rect 28316 31832 28322 31884
rect 28810 31872 28816 31884
rect 28771 31844 28816 31872
rect 28810 31832 28816 31844
rect 28868 31832 28874 31884
rect 29012 31881 29040 31912
rect 30098 31900 30104 31912
rect 30156 31900 30162 31952
rect 28997 31875 29055 31881
rect 28997 31841 29009 31875
rect 29043 31841 29055 31875
rect 29178 31872 29184 31884
rect 29139 31844 29184 31872
rect 28997 31835 29055 31841
rect 29178 31832 29184 31844
rect 29236 31872 29242 31884
rect 29825 31875 29883 31881
rect 29825 31872 29837 31875
rect 29236 31844 29837 31872
rect 29236 31832 29242 31844
rect 29825 31841 29837 31844
rect 29871 31872 29883 31875
rect 30561 31875 30619 31881
rect 30561 31872 30573 31875
rect 29871 31844 30573 31872
rect 29871 31841 29883 31844
rect 29825 31835 29883 31841
rect 30561 31841 30573 31844
rect 30607 31841 30619 31875
rect 30561 31835 30619 31841
rect 19981 31807 20039 31813
rect 19981 31804 19993 31807
rect 16448 31776 17448 31804
rect 19352 31776 19993 31804
rect 16448 31764 16454 31776
rect 12526 31696 12532 31748
rect 12584 31736 12590 31748
rect 16114 31736 16120 31748
rect 12584 31708 16120 31736
rect 12584 31696 12590 31708
rect 16114 31696 16120 31708
rect 16172 31696 16178 31748
rect 19242 31696 19248 31748
rect 19300 31736 19306 31748
rect 19352 31736 19380 31776
rect 19981 31773 19993 31776
rect 20027 31804 20039 31807
rect 20438 31804 20444 31816
rect 20027 31776 20444 31804
rect 20027 31773 20039 31776
rect 19981 31767 20039 31773
rect 20438 31764 20444 31776
rect 20496 31764 20502 31816
rect 24578 31804 24584 31816
rect 24539 31776 24584 31804
rect 24578 31764 24584 31776
rect 24636 31764 24642 31816
rect 26510 31804 26516 31816
rect 26471 31776 26516 31804
rect 26510 31764 26516 31776
rect 26568 31764 26574 31816
rect 28353 31807 28411 31813
rect 28353 31773 28365 31807
rect 28399 31804 28411 31807
rect 28399 31776 28948 31804
rect 28399 31773 28411 31776
rect 28353 31767 28411 31773
rect 19300 31708 19380 31736
rect 28920 31736 28948 31776
rect 29730 31736 29736 31748
rect 28920 31708 29736 31736
rect 19300 31696 19306 31708
rect 29730 31696 29736 31708
rect 29788 31696 29794 31748
rect 3237 31671 3295 31677
rect 3237 31637 3249 31671
rect 3283 31668 3295 31671
rect 3786 31668 3792 31680
rect 3283 31640 3792 31668
rect 3283 31637 3295 31640
rect 3237 31631 3295 31637
rect 3786 31628 3792 31640
rect 3844 31628 3850 31680
rect 12894 31668 12900 31680
rect 12855 31640 12900 31668
rect 12894 31628 12900 31640
rect 12952 31628 12958 31680
rect 23658 31668 23664 31680
rect 23619 31640 23664 31668
rect 23658 31628 23664 31640
rect 23716 31668 23722 31680
rect 25869 31671 25927 31677
rect 25869 31668 25881 31671
rect 23716 31640 25881 31668
rect 23716 31628 23722 31640
rect 25869 31637 25881 31640
rect 25915 31668 25927 31671
rect 25958 31668 25964 31680
rect 25915 31640 25964 31668
rect 25915 31637 25927 31640
rect 25869 31631 25927 31637
rect 25958 31628 25964 31640
rect 26016 31628 26022 31680
rect 27246 31628 27252 31680
rect 27304 31668 27310 31680
rect 27525 31671 27583 31677
rect 27525 31668 27537 31671
rect 27304 31640 27537 31668
rect 27304 31628 27310 31640
rect 27525 31637 27537 31640
rect 27571 31637 27583 31671
rect 30926 31668 30932 31680
rect 30887 31640 30932 31668
rect 27525 31631 27583 31637
rect 30926 31628 30932 31640
rect 30984 31628 30990 31680
rect 1104 31578 38548 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 38548 31578
rect 1104 31504 38548 31526
rect 10873 31467 10931 31473
rect 10873 31433 10885 31467
rect 10919 31464 10931 31467
rect 10962 31464 10968 31476
rect 10919 31436 10968 31464
rect 10919 31433 10931 31436
rect 10873 31427 10931 31433
rect 3050 31396 3056 31408
rect 2963 31368 3056 31396
rect 3050 31356 3056 31368
rect 3108 31396 3114 31408
rect 7742 31396 7748 31408
rect 3108 31368 7748 31396
rect 3108 31356 3114 31368
rect 2774 31288 2780 31340
rect 2832 31328 2838 31340
rect 3896 31337 3924 31368
rect 7742 31356 7748 31368
rect 7800 31356 7806 31408
rect 3145 31331 3203 31337
rect 3145 31328 3157 31331
rect 2832 31300 3157 31328
rect 2832 31288 2838 31300
rect 3145 31297 3157 31300
rect 3191 31297 3203 31331
rect 3145 31291 3203 31297
rect 3881 31331 3939 31337
rect 3881 31297 3893 31331
rect 3927 31297 3939 31331
rect 4062 31328 4068 31340
rect 4023 31300 4068 31328
rect 3881 31291 3939 31297
rect 4062 31288 4068 31300
rect 4120 31288 4126 31340
rect 3786 31260 3792 31272
rect 3747 31232 3792 31260
rect 3786 31220 3792 31232
rect 3844 31220 3850 31272
rect 4157 31263 4215 31269
rect 4157 31229 4169 31263
rect 4203 31229 4215 31263
rect 4157 31223 4215 31229
rect 10505 31263 10563 31269
rect 10505 31229 10517 31263
rect 10551 31260 10563 31263
rect 10888 31260 10916 31427
rect 10962 31424 10968 31436
rect 11020 31424 11026 31476
rect 16117 31467 16175 31473
rect 16117 31433 16129 31467
rect 16163 31464 16175 31467
rect 16853 31467 16911 31473
rect 16853 31464 16865 31467
rect 16163 31436 16865 31464
rect 16163 31433 16175 31436
rect 16117 31427 16175 31433
rect 16853 31433 16865 31436
rect 16899 31464 16911 31467
rect 17034 31464 17040 31476
rect 16899 31436 17040 31464
rect 16899 31433 16911 31436
rect 16853 31427 16911 31433
rect 17034 31424 17040 31436
rect 17092 31424 17098 31476
rect 23109 31467 23167 31473
rect 23109 31433 23121 31467
rect 23155 31464 23167 31467
rect 25406 31464 25412 31476
rect 23155 31436 25412 31464
rect 23155 31433 23167 31436
rect 23109 31427 23167 31433
rect 25406 31424 25412 31436
rect 25464 31424 25470 31476
rect 28629 31467 28687 31473
rect 28629 31433 28641 31467
rect 28675 31464 28687 31467
rect 28718 31464 28724 31476
rect 28675 31436 28724 31464
rect 28675 31433 28687 31436
rect 28629 31427 28687 31433
rect 28718 31424 28724 31436
rect 28776 31424 28782 31476
rect 30653 31467 30711 31473
rect 30653 31433 30665 31467
rect 30699 31464 30711 31467
rect 30926 31464 30932 31476
rect 30699 31436 30932 31464
rect 30699 31433 30711 31436
rect 30653 31427 30711 31433
rect 30926 31424 30932 31436
rect 30984 31464 30990 31476
rect 35618 31464 35624 31476
rect 30984 31436 32076 31464
rect 35579 31436 35624 31464
rect 30984 31424 30990 31436
rect 16390 31396 16396 31408
rect 16351 31368 16396 31396
rect 16390 31356 16396 31368
rect 16448 31396 16454 31408
rect 17586 31396 17592 31408
rect 16448 31368 17592 31396
rect 16448 31356 16454 31368
rect 17586 31356 17592 31368
rect 17644 31396 17650 31408
rect 18233 31399 18291 31405
rect 18233 31396 18245 31399
rect 17644 31368 18245 31396
rect 17644 31356 17650 31368
rect 18233 31365 18245 31368
rect 18279 31365 18291 31399
rect 18233 31359 18291 31365
rect 18874 31356 18880 31408
rect 18932 31396 18938 31408
rect 19150 31396 19156 31408
rect 18932 31368 19156 31396
rect 18932 31356 18938 31368
rect 19150 31356 19156 31368
rect 19208 31356 19214 31408
rect 23658 31356 23664 31408
rect 23716 31396 23722 31408
rect 23716 31368 24624 31396
rect 23716 31356 23722 31368
rect 12894 31328 12900 31340
rect 12855 31300 12900 31328
rect 12894 31288 12900 31300
rect 12952 31288 12958 31340
rect 15749 31331 15807 31337
rect 15749 31297 15761 31331
rect 15795 31328 15807 31331
rect 19889 31331 19947 31337
rect 15795 31300 16712 31328
rect 15795 31297 15807 31300
rect 15749 31291 15807 31297
rect 16684 31272 16712 31300
rect 19889 31297 19901 31331
rect 19935 31328 19947 31331
rect 20070 31328 20076 31340
rect 19935 31300 20076 31328
rect 19935 31297 19947 31300
rect 19889 31291 19947 31297
rect 20070 31288 20076 31300
rect 20128 31288 20134 31340
rect 23842 31328 23848 31340
rect 23803 31300 23848 31328
rect 23842 31288 23848 31300
rect 23900 31288 23906 31340
rect 13173 31263 13231 31269
rect 13173 31260 13185 31263
rect 10551 31232 10916 31260
rect 13004 31232 13185 31260
rect 10551 31229 10563 31232
rect 10505 31223 10563 31229
rect 4172 31192 4200 31223
rect 4614 31192 4620 31204
rect 4172 31164 4620 31192
rect 4614 31152 4620 31164
rect 4672 31152 4678 31204
rect 13004 31136 13032 31232
rect 13173 31229 13185 31232
rect 13219 31229 13231 31263
rect 13173 31223 13231 31229
rect 16390 31220 16396 31272
rect 16448 31260 16454 31272
rect 16577 31263 16635 31269
rect 16577 31260 16589 31263
rect 16448 31232 16589 31260
rect 16448 31220 16454 31232
rect 16577 31229 16589 31232
rect 16623 31229 16635 31263
rect 16577 31223 16635 31229
rect 14550 31192 14556 31204
rect 14511 31164 14556 31192
rect 14550 31152 14556 31164
rect 14608 31152 14614 31204
rect 16592 31192 16620 31223
rect 16666 31220 16672 31272
rect 16724 31260 16730 31272
rect 16724 31232 16817 31260
rect 16724 31220 16730 31232
rect 16942 31220 16948 31272
rect 17000 31260 17006 31272
rect 17862 31260 17868 31272
rect 17000 31232 17868 31260
rect 17000 31220 17006 31232
rect 17862 31220 17868 31232
rect 17920 31220 17926 31272
rect 18049 31263 18107 31269
rect 18049 31229 18061 31263
rect 18095 31260 18107 31263
rect 18138 31260 18144 31272
rect 18095 31232 18144 31260
rect 18095 31229 18107 31232
rect 18049 31223 18107 31229
rect 18138 31220 18144 31232
rect 18196 31260 18202 31272
rect 18874 31260 18880 31272
rect 18196 31232 18880 31260
rect 18196 31220 18202 31232
rect 18874 31220 18880 31232
rect 18932 31220 18938 31272
rect 19242 31260 19248 31272
rect 19203 31232 19248 31260
rect 19242 31220 19248 31232
rect 19300 31220 19306 31272
rect 19613 31263 19671 31269
rect 19613 31229 19625 31263
rect 19659 31260 19671 31263
rect 20254 31260 20260 31272
rect 19659 31232 20260 31260
rect 19659 31229 19671 31232
rect 19613 31223 19671 31229
rect 20254 31220 20260 31232
rect 20312 31220 20318 31272
rect 23750 31260 23756 31272
rect 23711 31232 23756 31260
rect 23750 31220 23756 31232
rect 23808 31220 23814 31272
rect 24596 31269 24624 31368
rect 25501 31331 25559 31337
rect 25501 31297 25513 31331
rect 25547 31328 25559 31331
rect 25593 31331 25651 31337
rect 25593 31328 25605 31331
rect 25547 31300 25605 31328
rect 25547 31297 25559 31300
rect 25501 31291 25559 31297
rect 25593 31297 25605 31300
rect 25639 31328 25651 31331
rect 26510 31328 26516 31340
rect 25639 31300 26516 31328
rect 25639 31297 25651 31300
rect 25593 31291 25651 31297
rect 26510 31288 26516 31300
rect 26568 31288 26574 31340
rect 27798 31288 27804 31340
rect 27856 31328 27862 31340
rect 27893 31331 27951 31337
rect 27893 31328 27905 31331
rect 27856 31300 27905 31328
rect 27856 31288 27862 31300
rect 27893 31297 27905 31300
rect 27939 31297 27951 31331
rect 30006 31328 30012 31340
rect 29967 31300 30012 31328
rect 27893 31291 27951 31297
rect 30006 31288 30012 31300
rect 30064 31288 30070 31340
rect 30558 31288 30564 31340
rect 30616 31328 30622 31340
rect 30926 31328 30932 31340
rect 30616 31300 30932 31328
rect 30616 31288 30622 31300
rect 30926 31288 30932 31300
rect 30984 31328 30990 31340
rect 32048 31328 32076 31436
rect 35618 31424 35624 31436
rect 35676 31424 35682 31476
rect 32122 31328 32128 31340
rect 30984 31300 31984 31328
rect 32035 31300 32128 31328
rect 30984 31288 30990 31300
rect 24581 31263 24639 31269
rect 24581 31229 24593 31263
rect 24627 31229 24639 31263
rect 24581 31223 24639 31229
rect 24673 31263 24731 31269
rect 24673 31229 24685 31263
rect 24719 31229 24731 31263
rect 25777 31263 25835 31269
rect 25777 31260 25789 31263
rect 24673 31223 24731 31229
rect 25056 31232 25789 31260
rect 17405 31195 17463 31201
rect 17405 31192 17417 31195
rect 16592 31164 17417 31192
rect 17405 31161 17417 31164
rect 17451 31161 17463 31195
rect 18506 31192 18512 31204
rect 17405 31155 17463 31161
rect 18064 31164 18512 31192
rect 2682 31124 2688 31136
rect 2643 31096 2688 31124
rect 2682 31084 2688 31096
rect 2740 31084 2746 31136
rect 10318 31124 10324 31136
rect 10279 31096 10324 31124
rect 10318 31084 10324 31096
rect 10376 31084 10382 31136
rect 12805 31127 12863 31133
rect 12805 31093 12817 31127
rect 12851 31124 12863 31127
rect 12986 31124 12992 31136
rect 12851 31096 12992 31124
rect 12851 31093 12863 31096
rect 12805 31087 12863 31093
rect 12986 31084 12992 31096
rect 13044 31084 13050 31136
rect 17420 31124 17448 31155
rect 18064 31136 18092 31164
rect 18506 31152 18512 31164
rect 18564 31152 18570 31204
rect 24688 31192 24716 31223
rect 23676 31164 24716 31192
rect 23676 31136 23704 31164
rect 25056 31136 25084 31232
rect 25777 31229 25789 31232
rect 25823 31229 25835 31263
rect 25777 31223 25835 31229
rect 26329 31263 26387 31269
rect 26329 31229 26341 31263
rect 26375 31260 26387 31263
rect 28810 31260 28816 31272
rect 26375 31232 28816 31260
rect 26375 31229 26387 31232
rect 26329 31223 26387 31229
rect 28810 31220 28816 31232
rect 28868 31220 28874 31272
rect 29549 31263 29607 31269
rect 29549 31229 29561 31263
rect 29595 31229 29607 31263
rect 29730 31260 29736 31272
rect 29691 31232 29736 31260
rect 29549 31223 29607 31229
rect 25958 31192 25964 31204
rect 25919 31164 25964 31192
rect 25958 31152 25964 31164
rect 26016 31152 26022 31204
rect 27157 31195 27215 31201
rect 27157 31161 27169 31195
rect 27203 31161 27215 31195
rect 27522 31192 27528 31204
rect 27483 31164 27528 31192
rect 27157 31155 27215 31161
rect 18046 31124 18052 31136
rect 17420 31096 18052 31124
rect 18046 31084 18052 31096
rect 18104 31084 18110 31136
rect 18414 31084 18420 31136
rect 18472 31124 18478 31136
rect 18601 31127 18659 31133
rect 18601 31124 18613 31127
rect 18472 31096 18613 31124
rect 18472 31084 18478 31096
rect 18601 31093 18613 31096
rect 18647 31124 18659 31127
rect 18690 31124 18696 31136
rect 18647 31096 18696 31124
rect 18647 31093 18659 31096
rect 18601 31087 18659 31093
rect 18690 31084 18696 31096
rect 18748 31084 18754 31136
rect 19058 31124 19064 31136
rect 19019 31096 19064 31124
rect 19058 31084 19064 31096
rect 19116 31084 19122 31136
rect 20990 31124 20996 31136
rect 20951 31096 20996 31124
rect 20990 31084 20996 31096
rect 21048 31084 21054 31136
rect 23477 31127 23535 31133
rect 23477 31093 23489 31127
rect 23523 31124 23535 31127
rect 23658 31124 23664 31136
rect 23523 31096 23664 31124
rect 23523 31093 23535 31096
rect 23477 31087 23535 31093
rect 23658 31084 23664 31096
rect 23716 31084 23722 31136
rect 25038 31124 25044 31136
rect 24999 31096 25044 31124
rect 25038 31084 25044 31096
rect 25096 31084 25102 31136
rect 25869 31127 25927 31133
rect 25869 31093 25881 31127
rect 25915 31124 25927 31127
rect 26050 31124 26056 31136
rect 25915 31096 26056 31124
rect 25915 31093 25927 31096
rect 25869 31087 25927 31093
rect 26050 31084 26056 31096
rect 26108 31084 26114 31136
rect 26510 31084 26516 31136
rect 26568 31124 26574 31136
rect 26605 31127 26663 31133
rect 26605 31124 26617 31127
rect 26568 31096 26617 31124
rect 26568 31084 26574 31096
rect 26605 31093 26617 31096
rect 26651 31093 26663 31127
rect 26970 31124 26976 31136
rect 26931 31096 26976 31124
rect 26605 31087 26663 31093
rect 26970 31084 26976 31096
rect 27028 31124 27034 31136
rect 27172 31124 27200 31155
rect 27522 31152 27528 31164
rect 27580 31152 27586 31204
rect 29089 31195 29147 31201
rect 29089 31161 29101 31195
rect 29135 31192 29147 31195
rect 29564 31192 29592 31223
rect 29730 31220 29736 31232
rect 29788 31220 29794 31272
rect 31478 31220 31484 31272
rect 31536 31260 31542 31272
rect 31956 31269 31984 31300
rect 32122 31288 32128 31300
rect 32180 31288 32186 31340
rect 35636 31328 35664 31424
rect 36081 31331 36139 31337
rect 36081 31328 36093 31331
rect 35636 31300 36093 31328
rect 36081 31297 36093 31300
rect 36127 31297 36139 31331
rect 36081 31291 36139 31297
rect 31665 31263 31723 31269
rect 31665 31260 31677 31263
rect 31536 31232 31677 31260
rect 31536 31220 31542 31232
rect 31665 31229 31677 31232
rect 31711 31229 31723 31263
rect 31665 31223 31723 31229
rect 31941 31263 31999 31269
rect 31941 31229 31953 31263
rect 31987 31229 31999 31263
rect 31941 31223 31999 31229
rect 35805 31263 35863 31269
rect 35805 31229 35817 31263
rect 35851 31260 35863 31263
rect 35894 31260 35900 31272
rect 35851 31232 35900 31260
rect 35851 31229 35863 31232
rect 35805 31223 35863 31229
rect 35894 31220 35900 31232
rect 35952 31220 35958 31272
rect 30742 31192 30748 31204
rect 29135 31164 30748 31192
rect 29135 31161 29147 31164
rect 29089 31155 29147 31161
rect 30742 31152 30748 31164
rect 30800 31152 30806 31204
rect 31113 31195 31171 31201
rect 31113 31161 31125 31195
rect 31159 31161 31171 31195
rect 31113 31155 31171 31161
rect 27028 31096 27200 31124
rect 27028 31084 27034 31096
rect 27246 31084 27252 31136
rect 27304 31124 27310 31136
rect 27341 31127 27399 31133
rect 27341 31124 27353 31127
rect 27304 31096 27353 31124
rect 27304 31084 27310 31096
rect 27341 31093 27353 31096
rect 27387 31093 27399 31127
rect 27341 31087 27399 31093
rect 27430 31084 27436 31136
rect 27488 31124 27494 31136
rect 28166 31124 28172 31136
rect 27488 31096 28172 31124
rect 27488 31084 27494 31096
rect 28166 31084 28172 31096
rect 28224 31084 28230 31136
rect 31128 31124 31156 31155
rect 31662 31124 31668 31136
rect 31128 31096 31668 31124
rect 31662 31084 31668 31096
rect 31720 31084 31726 31136
rect 37274 31084 37280 31136
rect 37332 31124 37338 31136
rect 37369 31127 37427 31133
rect 37369 31124 37381 31127
rect 37332 31096 37381 31124
rect 37332 31084 37338 31096
rect 37369 31093 37381 31096
rect 37415 31093 37427 31127
rect 37369 31087 37427 31093
rect 1104 31034 38548 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 38548 31034
rect 1104 30960 38548 30982
rect 3237 30923 3295 30929
rect 3237 30889 3249 30923
rect 3283 30920 3295 30923
rect 4062 30920 4068 30932
rect 3283 30892 4068 30920
rect 3283 30889 3295 30892
rect 3237 30883 3295 30889
rect 4062 30880 4068 30892
rect 4120 30880 4126 30932
rect 13814 30880 13820 30932
rect 13872 30920 13878 30932
rect 13909 30923 13967 30929
rect 13909 30920 13921 30923
rect 13872 30892 13921 30920
rect 13872 30880 13878 30892
rect 13909 30889 13921 30892
rect 13955 30889 13967 30923
rect 13909 30883 13967 30889
rect 13081 30855 13139 30861
rect 13081 30821 13093 30855
rect 13127 30852 13139 30855
rect 13722 30852 13728 30864
rect 13127 30824 13728 30852
rect 13127 30821 13139 30824
rect 13081 30815 13139 30821
rect 11977 30787 12035 30793
rect 11977 30753 11989 30787
rect 12023 30784 12035 30787
rect 13096 30784 13124 30815
rect 13722 30812 13728 30824
rect 13780 30812 13786 30864
rect 13924 30852 13952 30883
rect 13998 30880 14004 30932
rect 14056 30920 14062 30932
rect 14277 30923 14335 30929
rect 14277 30920 14289 30923
rect 14056 30892 14289 30920
rect 14056 30880 14062 30892
rect 14277 30889 14289 30892
rect 14323 30889 14335 30923
rect 16666 30920 16672 30932
rect 16627 30892 16672 30920
rect 14277 30883 14335 30889
rect 16666 30880 16672 30892
rect 16724 30880 16730 30932
rect 17218 30920 17224 30932
rect 17179 30892 17224 30920
rect 17218 30880 17224 30892
rect 17276 30880 17282 30932
rect 18874 30880 18880 30932
rect 18932 30920 18938 30932
rect 19334 30920 19340 30932
rect 18932 30892 19340 30920
rect 18932 30880 18938 30892
rect 19334 30880 19340 30892
rect 19392 30920 19398 30932
rect 19429 30923 19487 30929
rect 19429 30920 19441 30923
rect 19392 30892 19441 30920
rect 19392 30880 19398 30892
rect 19429 30889 19441 30892
rect 19475 30889 19487 30923
rect 19429 30883 19487 30889
rect 19889 30923 19947 30929
rect 19889 30889 19901 30923
rect 19935 30920 19947 30923
rect 20070 30920 20076 30932
rect 19935 30892 20076 30920
rect 19935 30889 19947 30892
rect 19889 30883 19947 30889
rect 20070 30880 20076 30892
rect 20128 30880 20134 30932
rect 23750 30920 23756 30932
rect 23711 30892 23756 30920
rect 23750 30880 23756 30892
rect 23808 30880 23814 30932
rect 24578 30920 24584 30932
rect 24539 30892 24584 30920
rect 24578 30880 24584 30892
rect 24636 30880 24642 30932
rect 26329 30923 26387 30929
rect 26329 30889 26341 30923
rect 26375 30920 26387 30923
rect 27522 30920 27528 30932
rect 26375 30892 27528 30920
rect 26375 30889 26387 30892
rect 26329 30883 26387 30889
rect 27522 30880 27528 30892
rect 27580 30880 27586 30932
rect 28534 30880 28540 30932
rect 28592 30920 28598 30932
rect 28721 30923 28779 30929
rect 28721 30920 28733 30923
rect 28592 30892 28733 30920
rect 28592 30880 28598 30892
rect 28721 30889 28733 30892
rect 28767 30889 28779 30923
rect 29730 30920 29736 30932
rect 29691 30892 29736 30920
rect 28721 30883 28779 30889
rect 29730 30880 29736 30892
rect 29788 30880 29794 30932
rect 35894 30920 35900 30932
rect 35855 30892 35900 30920
rect 35894 30880 35900 30892
rect 35952 30880 35958 30932
rect 14734 30852 14740 30864
rect 13924 30824 14740 30852
rect 14734 30812 14740 30824
rect 14792 30812 14798 30864
rect 17586 30812 17592 30864
rect 17644 30852 17650 30864
rect 25225 30855 25283 30861
rect 25225 30852 25237 30855
rect 17644 30824 18920 30852
rect 17644 30812 17650 30824
rect 12023 30756 13124 30784
rect 12023 30753 12035 30756
rect 11977 30747 12035 30753
rect 13170 30744 13176 30796
rect 13228 30784 13234 30796
rect 13228 30756 13273 30784
rect 13228 30744 13234 30756
rect 18414 30744 18420 30796
rect 18472 30784 18478 30796
rect 18509 30787 18567 30793
rect 18509 30784 18521 30787
rect 18472 30756 18521 30784
rect 18472 30744 18478 30756
rect 18509 30753 18521 30756
rect 18555 30753 18567 30787
rect 18509 30747 18567 30753
rect 18598 30744 18604 30796
rect 18656 30784 18662 30796
rect 18892 30793 18920 30824
rect 24136 30824 25237 30852
rect 18693 30787 18751 30793
rect 18693 30784 18705 30787
rect 18656 30756 18705 30784
rect 18656 30744 18662 30756
rect 18693 30753 18705 30756
rect 18739 30753 18751 30787
rect 18693 30747 18751 30753
rect 18877 30787 18935 30793
rect 18877 30753 18889 30787
rect 18923 30753 18935 30787
rect 20254 30784 20260 30796
rect 20167 30756 20260 30784
rect 18877 30747 18935 30753
rect 20254 30744 20260 30756
rect 20312 30784 20318 30796
rect 21358 30784 21364 30796
rect 20312 30756 21364 30784
rect 20312 30744 20318 30756
rect 21358 30744 21364 30756
rect 21416 30744 21422 30796
rect 23014 30784 23020 30796
rect 22975 30756 23020 30784
rect 23014 30744 23020 30756
rect 23072 30744 23078 30796
rect 12066 30716 12072 30728
rect 12027 30688 12072 30716
rect 12066 30676 12072 30688
rect 12124 30676 12130 30728
rect 15289 30719 15347 30725
rect 15289 30685 15301 30719
rect 15335 30716 15347 30719
rect 15470 30716 15476 30728
rect 15335 30688 15476 30716
rect 15335 30685 15347 30688
rect 15289 30679 15347 30685
rect 15470 30676 15476 30688
rect 15528 30676 15534 30728
rect 15562 30676 15568 30728
rect 15620 30716 15626 30728
rect 15620 30688 15665 30716
rect 15620 30676 15626 30688
rect 21266 30676 21272 30728
rect 21324 30716 21330 30728
rect 21637 30719 21695 30725
rect 21637 30716 21649 30719
rect 21324 30688 21649 30716
rect 21324 30676 21330 30688
rect 21637 30685 21649 30688
rect 21683 30685 21695 30719
rect 21637 30679 21695 30685
rect 4062 30608 4068 30660
rect 4120 30648 4126 30660
rect 9582 30648 9588 30660
rect 4120 30620 9588 30648
rect 4120 30608 4126 30620
rect 9582 30608 9588 30620
rect 9640 30608 9646 30660
rect 18322 30648 18328 30660
rect 18283 30620 18328 30648
rect 18322 30608 18328 30620
rect 18380 30608 18386 30660
rect 6914 30580 6920 30592
rect 6875 30552 6920 30580
rect 6914 30540 6920 30552
rect 6972 30540 6978 30592
rect 10410 30580 10416 30592
rect 10371 30552 10416 30580
rect 10410 30540 10416 30552
rect 10468 30540 10474 30592
rect 12529 30583 12587 30589
rect 12529 30549 12541 30583
rect 12575 30580 12587 30583
rect 12710 30580 12716 30592
rect 12575 30552 12716 30580
rect 12575 30549 12587 30552
rect 12529 30543 12587 30549
rect 12710 30540 12716 30552
rect 12768 30580 12774 30592
rect 12897 30583 12955 30589
rect 12897 30580 12909 30583
rect 12768 30552 12909 30580
rect 12768 30540 12774 30552
rect 12897 30549 12909 30552
rect 12943 30549 12955 30583
rect 13354 30580 13360 30592
rect 13315 30552 13360 30580
rect 12897 30543 12955 30549
rect 13354 30540 13360 30552
rect 13412 30540 13418 30592
rect 23198 30540 23204 30592
rect 23256 30580 23262 30592
rect 24136 30589 24164 30824
rect 25225 30821 25237 30824
rect 25271 30821 25283 30855
rect 27338 30852 27344 30864
rect 27299 30824 27344 30852
rect 25225 30815 25283 30821
rect 27338 30812 27344 30824
rect 27396 30812 27402 30864
rect 27433 30855 27491 30861
rect 27433 30821 27445 30855
rect 27479 30821 27491 30855
rect 27433 30815 27491 30821
rect 28445 30855 28503 30861
rect 28445 30821 28457 30855
rect 28491 30852 28503 30855
rect 28810 30852 28816 30864
rect 28491 30824 28816 30852
rect 28491 30821 28503 30824
rect 28445 30815 28503 30821
rect 25038 30784 25044 30796
rect 24999 30756 25044 30784
rect 25038 30744 25044 30756
rect 25096 30744 25102 30796
rect 25133 30787 25191 30793
rect 25133 30753 25145 30787
rect 25179 30753 25191 30787
rect 27246 30784 27252 30796
rect 27207 30756 27252 30784
rect 25133 30747 25191 30753
rect 24854 30716 24860 30728
rect 24815 30688 24860 30716
rect 24854 30676 24860 30688
rect 24912 30676 24918 30728
rect 24121 30583 24179 30589
rect 24121 30580 24133 30583
rect 23256 30552 24133 30580
rect 23256 30540 23262 30552
rect 24121 30549 24133 30552
rect 24167 30549 24179 30583
rect 25148 30580 25176 30747
rect 27246 30744 27252 30756
rect 27304 30744 27310 30796
rect 27448 30784 27476 30815
rect 28810 30812 28816 30824
rect 28868 30812 28874 30864
rect 27522 30784 27528 30796
rect 27448 30756 27528 30784
rect 25590 30716 25596 30728
rect 25551 30688 25596 30716
rect 25590 30676 25596 30688
rect 25648 30676 25654 30728
rect 26970 30676 26976 30728
rect 27028 30716 27034 30728
rect 27065 30719 27123 30725
rect 27065 30716 27077 30719
rect 27028 30688 27077 30716
rect 27028 30676 27034 30688
rect 27065 30685 27077 30688
rect 27111 30685 27123 30719
rect 27065 30679 27123 30685
rect 26786 30608 26792 30660
rect 26844 30648 26850 30660
rect 27448 30648 27476 30756
rect 27522 30744 27528 30756
rect 27580 30744 27586 30796
rect 30006 30784 30012 30796
rect 29967 30756 30012 30784
rect 30006 30744 30012 30756
rect 30064 30744 30070 30796
rect 30742 30784 30748 30796
rect 30703 30756 30748 30784
rect 30742 30744 30748 30756
rect 30800 30744 30806 30796
rect 31205 30787 31263 30793
rect 31205 30753 31217 30787
rect 31251 30784 31263 30787
rect 31478 30784 31484 30796
rect 31251 30756 31484 30784
rect 31251 30753 31263 30756
rect 31205 30747 31263 30753
rect 31478 30744 31484 30756
rect 31536 30744 31542 30796
rect 27798 30716 27804 30728
rect 27759 30688 27804 30716
rect 27798 30676 27804 30688
rect 27856 30676 27862 30728
rect 26844 30620 27476 30648
rect 26844 30608 26850 30620
rect 25961 30583 26019 30589
rect 25961 30580 25973 30583
rect 25148 30552 25973 30580
rect 24121 30543 24179 30549
rect 25961 30549 25973 30552
rect 26007 30580 26019 30583
rect 26050 30580 26056 30592
rect 26007 30552 26056 30580
rect 26007 30549 26019 30552
rect 25961 30543 26019 30549
rect 26050 30540 26056 30552
rect 26108 30540 26114 30592
rect 26694 30580 26700 30592
rect 26655 30552 26700 30580
rect 26694 30540 26700 30552
rect 26752 30540 26758 30592
rect 29270 30580 29276 30592
rect 29231 30552 29276 30580
rect 29270 30540 29276 30552
rect 29328 30540 29334 30592
rect 1104 30490 38548 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 38548 30490
rect 1104 30416 38548 30438
rect 3786 30336 3792 30388
rect 3844 30376 3850 30388
rect 10318 30376 10324 30388
rect 3844 30348 4108 30376
rect 3844 30336 3850 30348
rect 4080 30308 4108 30348
rect 9600 30348 10324 30376
rect 4525 30311 4583 30317
rect 4525 30308 4537 30311
rect 4080 30280 4537 30308
rect 4525 30277 4537 30280
rect 4571 30277 4583 30311
rect 4525 30271 4583 30277
rect 9217 30311 9275 30317
rect 9217 30277 9229 30311
rect 9263 30308 9275 30311
rect 9600 30308 9628 30348
rect 10318 30336 10324 30348
rect 10376 30336 10382 30388
rect 12894 30336 12900 30388
rect 12952 30376 12958 30388
rect 13446 30376 13452 30388
rect 12952 30348 13452 30376
rect 12952 30336 12958 30348
rect 13446 30336 13452 30348
rect 13504 30376 13510 30388
rect 14001 30379 14059 30385
rect 14001 30376 14013 30379
rect 13504 30348 14013 30376
rect 13504 30336 13510 30348
rect 14001 30345 14013 30348
rect 14047 30345 14059 30379
rect 14550 30376 14556 30388
rect 14511 30348 14556 30376
rect 14001 30339 14059 30345
rect 14550 30336 14556 30348
rect 14608 30336 14614 30388
rect 15562 30336 15568 30388
rect 15620 30376 15626 30388
rect 16025 30379 16083 30385
rect 16025 30376 16037 30379
rect 15620 30348 16037 30376
rect 15620 30336 15626 30348
rect 16025 30345 16037 30348
rect 16071 30376 16083 30379
rect 17218 30376 17224 30388
rect 16071 30348 17224 30376
rect 16071 30345 16083 30348
rect 16025 30339 16083 30345
rect 17218 30336 17224 30348
rect 17276 30336 17282 30388
rect 17586 30336 17592 30388
rect 17644 30376 17650 30388
rect 17773 30379 17831 30385
rect 17773 30376 17785 30379
rect 17644 30348 17785 30376
rect 17644 30336 17650 30348
rect 17773 30345 17785 30348
rect 17819 30345 17831 30379
rect 18322 30376 18328 30388
rect 18283 30348 18328 30376
rect 17773 30339 17831 30345
rect 9263 30280 9628 30308
rect 9263 30277 9275 30280
rect 9217 30271 9275 30277
rect 2774 30200 2780 30252
rect 2832 30240 2838 30252
rect 3053 30243 3111 30249
rect 3053 30240 3065 30243
rect 2832 30212 3065 30240
rect 2832 30200 2838 30212
rect 3053 30209 3065 30212
rect 3099 30240 3111 30243
rect 3099 30212 3464 30240
rect 3099 30209 3111 30212
rect 3053 30203 3111 30209
rect 2685 30175 2743 30181
rect 2685 30141 2697 30175
rect 2731 30172 2743 30175
rect 3145 30175 3203 30181
rect 3145 30172 3157 30175
rect 2731 30144 3157 30172
rect 2731 30141 2743 30144
rect 2685 30135 2743 30141
rect 3145 30141 3157 30144
rect 3191 30172 3203 30175
rect 3234 30172 3240 30184
rect 3191 30144 3240 30172
rect 3191 30141 3203 30144
rect 3145 30135 3203 30141
rect 3234 30132 3240 30144
rect 3292 30132 3298 30184
rect 3436 30181 3464 30212
rect 6914 30200 6920 30252
rect 6972 30240 6978 30252
rect 7837 30243 7895 30249
rect 7837 30240 7849 30243
rect 6972 30212 7849 30240
rect 6972 30200 6978 30212
rect 7837 30209 7849 30212
rect 7883 30209 7895 30243
rect 7837 30203 7895 30209
rect 3421 30175 3479 30181
rect 3421 30141 3433 30175
rect 3467 30172 3479 30175
rect 4614 30172 4620 30184
rect 3467 30144 4620 30172
rect 3467 30141 3479 30144
rect 3421 30135 3479 30141
rect 4614 30132 4620 30144
rect 4672 30132 4678 30184
rect 7374 30172 7380 30184
rect 7335 30144 7380 30172
rect 7374 30132 7380 30144
rect 7432 30132 7438 30184
rect 7653 30175 7711 30181
rect 7653 30141 7665 30175
rect 7699 30172 7711 30175
rect 8018 30172 8024 30184
rect 7699 30144 8024 30172
rect 7699 30141 7711 30144
rect 7653 30135 7711 30141
rect 6825 30107 6883 30113
rect 6825 30073 6837 30107
rect 6871 30104 6883 30107
rect 7098 30104 7104 30116
rect 6871 30076 7104 30104
rect 6871 30073 6883 30076
rect 6825 30067 6883 30073
rect 7098 30064 7104 30076
rect 7156 30064 7162 30116
rect 6641 30039 6699 30045
rect 6641 30005 6653 30039
rect 6687 30036 6699 30039
rect 7668 30036 7696 30135
rect 8018 30132 8024 30144
rect 8076 30132 8082 30184
rect 8849 30175 8907 30181
rect 8849 30141 8861 30175
rect 8895 30172 8907 30175
rect 9232 30172 9260 30271
rect 9674 30268 9680 30320
rect 9732 30308 9738 30320
rect 10413 30311 10471 30317
rect 10413 30308 10425 30311
rect 9732 30280 10425 30308
rect 9732 30268 9738 30280
rect 10413 30277 10425 30280
rect 10459 30308 10471 30311
rect 10502 30308 10508 30320
rect 10459 30280 10508 30308
rect 10459 30277 10471 30280
rect 10413 30271 10471 30277
rect 10502 30268 10508 30280
rect 10560 30268 10566 30320
rect 11885 30311 11943 30317
rect 11885 30277 11897 30311
rect 11931 30308 11943 30311
rect 12526 30308 12532 30320
rect 11931 30280 12532 30308
rect 11931 30277 11943 30280
rect 11885 30271 11943 30277
rect 12526 30268 12532 30280
rect 12584 30308 12590 30320
rect 13906 30308 13912 30320
rect 12584 30280 13912 30308
rect 12584 30268 12590 30280
rect 13906 30268 13912 30280
rect 13964 30268 13970 30320
rect 10229 30243 10287 30249
rect 10229 30209 10241 30243
rect 10275 30240 10287 30243
rect 12066 30240 12072 30252
rect 10275 30212 12072 30240
rect 10275 30209 10287 30212
rect 10229 30203 10287 30209
rect 10410 30172 10416 30184
rect 8895 30144 9260 30172
rect 10371 30144 10416 30172
rect 8895 30141 8907 30144
rect 8849 30135 8907 30141
rect 10410 30132 10416 30144
rect 10468 30132 10474 30184
rect 10980 30181 11008 30212
rect 12066 30200 12072 30212
rect 12124 30200 12130 30252
rect 13170 30200 13176 30252
rect 13228 30240 13234 30252
rect 13449 30243 13507 30249
rect 13449 30240 13461 30243
rect 13228 30212 13461 30240
rect 13228 30200 13234 30212
rect 13449 30209 13461 30212
rect 13495 30209 13507 30243
rect 14568 30240 14596 30336
rect 17788 30308 17816 30339
rect 18322 30336 18328 30348
rect 18380 30336 18386 30388
rect 21266 30336 21272 30388
rect 21324 30376 21330 30388
rect 21361 30379 21419 30385
rect 21361 30376 21373 30379
rect 21324 30348 21373 30376
rect 21324 30336 21330 30348
rect 21361 30345 21373 30348
rect 21407 30345 21419 30379
rect 21361 30339 21419 30345
rect 28166 30336 28172 30388
rect 28224 30376 28230 30388
rect 28261 30379 28319 30385
rect 28261 30376 28273 30379
rect 28224 30348 28273 30376
rect 28224 30336 28230 30348
rect 28261 30345 28273 30348
rect 28307 30345 28319 30379
rect 28261 30339 28319 30345
rect 31757 30379 31815 30385
rect 31757 30345 31769 30379
rect 31803 30376 31815 30379
rect 32122 30376 32128 30388
rect 31803 30348 32128 30376
rect 31803 30345 31815 30348
rect 31757 30339 31815 30345
rect 32122 30336 32128 30348
rect 32180 30336 32186 30388
rect 18414 30308 18420 30320
rect 17788 30280 18420 30308
rect 18414 30268 18420 30280
rect 18472 30268 18478 30320
rect 26789 30311 26847 30317
rect 26789 30277 26801 30311
rect 26835 30308 26847 30311
rect 27154 30308 27160 30320
rect 26835 30280 27160 30308
rect 26835 30277 26847 30280
rect 26789 30271 26847 30277
rect 27154 30268 27160 30280
rect 27212 30308 27218 30320
rect 27890 30308 27896 30320
rect 27212 30280 27896 30308
rect 27212 30268 27218 30280
rect 27890 30268 27896 30280
rect 27948 30268 27954 30320
rect 28350 30268 28356 30320
rect 28408 30308 28414 30320
rect 28810 30308 28816 30320
rect 28408 30280 28816 30308
rect 28408 30268 28414 30280
rect 28810 30268 28816 30280
rect 28868 30268 28874 30320
rect 15286 30240 15292 30252
rect 14568 30212 14872 30240
rect 15247 30212 15292 30240
rect 13449 30203 13507 30209
rect 10965 30175 11023 30181
rect 10965 30141 10977 30175
rect 11011 30141 11023 30175
rect 10965 30135 11023 30141
rect 11057 30175 11115 30181
rect 11057 30141 11069 30175
rect 11103 30172 11115 30175
rect 11698 30172 11704 30184
rect 11103 30144 11704 30172
rect 11103 30141 11115 30144
rect 11057 30135 11115 30141
rect 9861 30107 9919 30113
rect 9861 30073 9873 30107
rect 9907 30104 9919 30107
rect 11072 30104 11100 30135
rect 11698 30132 11704 30144
rect 11756 30132 11762 30184
rect 12437 30175 12495 30181
rect 12437 30172 12449 30175
rect 12176 30144 12449 30172
rect 9907 30076 11100 30104
rect 9907 30073 9919 30076
rect 9861 30067 9919 30073
rect 12176 30048 12204 30144
rect 12437 30141 12449 30144
rect 12483 30141 12495 30175
rect 12710 30172 12716 30184
rect 12671 30144 12716 30172
rect 12437 30135 12495 30141
rect 12710 30132 12716 30144
rect 12768 30132 12774 30184
rect 14182 30172 14188 30184
rect 14143 30144 14188 30172
rect 14182 30132 14188 30144
rect 14240 30132 14246 30184
rect 14734 30172 14740 30184
rect 14695 30144 14740 30172
rect 14734 30132 14740 30144
rect 14792 30132 14798 30184
rect 14844 30181 14872 30212
rect 15286 30200 15292 30212
rect 15344 30200 15350 30252
rect 18046 30240 18052 30252
rect 18007 30212 18052 30240
rect 18046 30200 18052 30212
rect 18104 30240 18110 30252
rect 18598 30240 18604 30252
rect 18104 30212 18604 30240
rect 18104 30200 18110 30212
rect 18598 30200 18604 30212
rect 18656 30240 18662 30252
rect 18877 30243 18935 30249
rect 18877 30240 18889 30243
rect 18656 30212 18889 30240
rect 18656 30200 18662 30212
rect 18877 30209 18889 30212
rect 18923 30209 18935 30243
rect 18877 30203 18935 30209
rect 19150 30200 19156 30252
rect 19208 30240 19214 30252
rect 19429 30243 19487 30249
rect 19429 30240 19441 30243
rect 19208 30212 19441 30240
rect 19208 30200 19214 30212
rect 19429 30209 19441 30212
rect 19475 30240 19487 30243
rect 20162 30240 20168 30252
rect 19475 30212 20168 30240
rect 19475 30209 19487 30212
rect 19429 30203 19487 30209
rect 20162 30200 20168 30212
rect 20220 30200 20226 30252
rect 21082 30240 21088 30252
rect 21043 30212 21088 30240
rect 21082 30200 21088 30212
rect 21140 30200 21146 30252
rect 24581 30243 24639 30249
rect 24581 30209 24593 30243
rect 24627 30240 24639 30243
rect 24854 30240 24860 30252
rect 24627 30212 24860 30240
rect 24627 30209 24639 30212
rect 24581 30203 24639 30209
rect 24854 30200 24860 30212
rect 24912 30200 24918 30252
rect 24949 30243 25007 30249
rect 24949 30209 24961 30243
rect 24995 30240 25007 30243
rect 25961 30243 26019 30249
rect 25961 30240 25973 30243
rect 24995 30212 25973 30240
rect 24995 30209 25007 30212
rect 24949 30203 25007 30209
rect 25961 30209 25973 30212
rect 26007 30240 26019 30243
rect 26602 30240 26608 30252
rect 26007 30212 26608 30240
rect 26007 30209 26019 30212
rect 25961 30203 26019 30209
rect 26602 30200 26608 30212
rect 26660 30200 26666 30252
rect 26973 30243 27031 30249
rect 26973 30209 26985 30243
rect 27019 30240 27031 30243
rect 28258 30240 28264 30252
rect 27019 30212 28264 30240
rect 27019 30209 27031 30212
rect 26973 30203 27031 30209
rect 28258 30200 28264 30212
rect 28316 30240 28322 30252
rect 28629 30243 28687 30249
rect 28629 30240 28641 30243
rect 28316 30212 28641 30240
rect 28316 30200 28322 30212
rect 28629 30209 28641 30212
rect 28675 30240 28687 30243
rect 29270 30240 29276 30252
rect 28675 30212 29276 30240
rect 28675 30209 28687 30212
rect 28629 30203 28687 30209
rect 29270 30200 29276 30212
rect 29328 30240 29334 30252
rect 29365 30243 29423 30249
rect 29365 30240 29377 30243
rect 29328 30212 29377 30240
rect 29328 30200 29334 30212
rect 29365 30209 29377 30212
rect 29411 30209 29423 30243
rect 29365 30203 29423 30209
rect 29730 30200 29736 30252
rect 29788 30240 29794 30252
rect 30285 30243 30343 30249
rect 30285 30240 30297 30243
rect 29788 30212 30297 30240
rect 29788 30200 29794 30212
rect 30285 30209 30297 30212
rect 30331 30209 30343 30243
rect 32140 30240 32168 30336
rect 35713 30311 35771 30317
rect 35713 30277 35725 30311
rect 35759 30308 35771 30311
rect 35802 30308 35808 30320
rect 35759 30280 35808 30308
rect 35759 30277 35771 30280
rect 35713 30271 35771 30277
rect 35802 30268 35808 30280
rect 35860 30268 35866 30320
rect 32309 30243 32367 30249
rect 32309 30240 32321 30243
rect 32140 30212 32321 30240
rect 30285 30203 30343 30209
rect 32309 30209 32321 30212
rect 32355 30209 32367 30243
rect 35820 30240 35848 30268
rect 36081 30243 36139 30249
rect 36081 30240 36093 30243
rect 35820 30212 36093 30240
rect 32309 30203 32367 30209
rect 36081 30209 36093 30212
rect 36127 30209 36139 30243
rect 36081 30203 36139 30209
rect 14829 30175 14887 30181
rect 14829 30141 14841 30175
rect 14875 30141 14887 30175
rect 14829 30135 14887 30141
rect 18141 30175 18199 30181
rect 18141 30141 18153 30175
rect 18187 30141 18199 30175
rect 19705 30175 19763 30181
rect 19705 30172 19717 30175
rect 18141 30135 18199 30141
rect 19352 30144 19717 30172
rect 13173 30107 13231 30113
rect 13173 30073 13185 30107
rect 13219 30104 13231 30107
rect 13262 30104 13268 30116
rect 13219 30076 13268 30104
rect 13219 30073 13231 30076
rect 13173 30067 13231 30073
rect 13262 30064 13268 30076
rect 13320 30064 13326 30116
rect 14752 30104 14780 30132
rect 15565 30107 15623 30113
rect 15565 30104 15577 30107
rect 14752 30076 15577 30104
rect 15565 30073 15577 30076
rect 15611 30104 15623 30107
rect 16390 30104 16396 30116
rect 15611 30076 16396 30104
rect 15611 30073 15623 30076
rect 15565 30067 15623 30073
rect 16390 30064 16396 30076
rect 16448 30064 16454 30116
rect 18156 30104 18184 30135
rect 17604 30076 18184 30104
rect 17604 30048 17632 30076
rect 19352 30048 19380 30144
rect 19705 30141 19717 30144
rect 19751 30141 19763 30175
rect 19705 30135 19763 30141
rect 21913 30175 21971 30181
rect 21913 30141 21925 30175
rect 21959 30172 21971 30175
rect 22278 30172 22284 30184
rect 21959 30144 22284 30172
rect 21959 30141 21971 30144
rect 21913 30135 21971 30141
rect 22278 30132 22284 30144
rect 22336 30132 22342 30184
rect 22557 30175 22615 30181
rect 22557 30141 22569 30175
rect 22603 30141 22615 30175
rect 22557 30135 22615 30141
rect 22186 30064 22192 30116
rect 22244 30104 22250 30116
rect 22572 30104 22600 30135
rect 24210 30132 24216 30184
rect 24268 30172 24274 30184
rect 25501 30175 25559 30181
rect 25501 30172 25513 30175
rect 24268 30144 25513 30172
rect 24268 30132 24274 30144
rect 25501 30141 25513 30144
rect 25547 30172 25559 30175
rect 25590 30172 25596 30184
rect 25547 30144 25596 30172
rect 25547 30141 25559 30144
rect 25501 30135 25559 30141
rect 25590 30132 25596 30144
rect 25648 30132 25654 30184
rect 25869 30175 25927 30181
rect 25869 30141 25881 30175
rect 25915 30172 25927 30175
rect 26142 30172 26148 30184
rect 25915 30144 26148 30172
rect 25915 30141 25927 30144
rect 25869 30135 25927 30141
rect 26142 30132 26148 30144
rect 26200 30132 26206 30184
rect 27706 30132 27712 30184
rect 27764 30172 27770 30184
rect 27801 30175 27859 30181
rect 27801 30172 27813 30175
rect 27764 30144 27813 30172
rect 27764 30132 27770 30144
rect 27801 30141 27813 30144
rect 27847 30141 27859 30175
rect 27801 30135 27859 30141
rect 27890 30132 27896 30184
rect 27948 30181 27954 30184
rect 27948 30175 27997 30181
rect 27948 30141 27951 30175
rect 27985 30141 27997 30175
rect 28994 30172 29000 30184
rect 28955 30144 29000 30172
rect 27948 30135 27997 30141
rect 27948 30132 27954 30135
rect 28994 30132 29000 30144
rect 29052 30172 29058 30184
rect 29052 30144 29592 30172
rect 29052 30132 29058 30144
rect 25041 30107 25099 30113
rect 25041 30104 25053 30107
rect 22244 30076 25053 30104
rect 22244 30064 22250 30076
rect 25041 30073 25053 30076
rect 25087 30073 25099 30107
rect 25041 30067 25099 30073
rect 27065 30107 27123 30113
rect 27065 30073 27077 30107
rect 27111 30104 27123 30107
rect 27522 30104 27528 30116
rect 27111 30076 27528 30104
rect 27111 30073 27123 30076
rect 27065 30067 27123 30073
rect 27522 30064 27528 30076
rect 27580 30064 27586 30116
rect 29362 30064 29368 30116
rect 29420 30104 29426 30116
rect 29457 30107 29515 30113
rect 29457 30104 29469 30107
rect 29420 30076 29469 30104
rect 29420 30064 29426 30076
rect 29457 30073 29469 30076
rect 29503 30073 29515 30107
rect 29564 30104 29592 30144
rect 30006 30132 30012 30184
rect 30064 30172 30070 30184
rect 30193 30175 30251 30181
rect 30193 30172 30205 30175
rect 30064 30144 30205 30172
rect 30064 30132 30070 30144
rect 30193 30141 30205 30144
rect 30239 30141 30251 30175
rect 30193 30135 30251 30141
rect 32030 30132 32036 30184
rect 32088 30172 32094 30184
rect 32125 30175 32183 30181
rect 32125 30172 32137 30175
rect 32088 30144 32137 30172
rect 32088 30132 32094 30144
rect 32125 30141 32137 30144
rect 32171 30172 32183 30175
rect 32769 30175 32827 30181
rect 32769 30172 32781 30175
rect 32171 30144 32781 30172
rect 32171 30141 32183 30144
rect 32125 30135 32183 30141
rect 32769 30141 32781 30144
rect 32815 30172 32827 30175
rect 32858 30172 32864 30184
rect 32815 30144 32864 30172
rect 32815 30141 32827 30144
rect 32769 30135 32827 30141
rect 32858 30132 32864 30144
rect 32916 30132 32922 30184
rect 32950 30132 32956 30184
rect 33008 30172 33014 30184
rect 33045 30175 33103 30181
rect 33045 30172 33057 30175
rect 33008 30144 33057 30172
rect 33008 30132 33014 30144
rect 33045 30141 33057 30144
rect 33091 30141 33103 30175
rect 33045 30135 33103 30141
rect 35805 30175 35863 30181
rect 35805 30141 35817 30175
rect 35851 30172 35863 30175
rect 35894 30172 35900 30184
rect 35851 30144 35900 30172
rect 35851 30141 35863 30144
rect 35805 30135 35863 30141
rect 35894 30132 35900 30144
rect 35952 30132 35958 30184
rect 31021 30107 31079 30113
rect 31021 30104 31033 30107
rect 29564 30076 31033 30104
rect 29457 30067 29515 30073
rect 31021 30073 31033 30076
rect 31067 30073 31079 30107
rect 31021 30067 31079 30073
rect 33321 30107 33379 30113
rect 33321 30073 33333 30107
rect 33367 30104 33379 30107
rect 33410 30104 33416 30116
rect 33367 30076 33416 30104
rect 33367 30073 33379 30076
rect 33321 30067 33379 30073
rect 33410 30064 33416 30076
rect 33468 30064 33474 30116
rect 6687 30008 7696 30036
rect 6687 30005 6699 30008
rect 6641 29999 6699 30005
rect 8570 29996 8576 30048
rect 8628 30036 8634 30048
rect 8665 30039 8723 30045
rect 8665 30036 8677 30039
rect 8628 30008 8677 30036
rect 8628 29996 8634 30008
rect 8665 30005 8677 30008
rect 8711 30005 8723 30039
rect 8665 29999 8723 30005
rect 11422 29996 11428 30048
rect 11480 30036 11486 30048
rect 12158 30036 12164 30048
rect 11480 30008 12164 30036
rect 11480 29996 11486 30008
rect 12158 29996 12164 30008
rect 12216 29996 12222 30048
rect 17497 30039 17555 30045
rect 17497 30005 17509 30039
rect 17543 30036 17555 30039
rect 17586 30036 17592 30048
rect 17543 30008 17592 30036
rect 17543 30005 17555 30008
rect 17497 29999 17555 30005
rect 17586 29996 17592 30008
rect 17644 29996 17650 30048
rect 19334 30036 19340 30048
rect 19295 30008 19340 30036
rect 19334 29996 19340 30008
rect 19392 29996 19398 30048
rect 22278 30036 22284 30048
rect 22239 30008 22284 30036
rect 22278 29996 22284 30008
rect 22336 29996 22342 30048
rect 23474 30036 23480 30048
rect 23435 30008 23480 30036
rect 23474 29996 23480 30008
rect 23532 29996 23538 30048
rect 24118 30036 24124 30048
rect 24079 30008 24124 30036
rect 24118 29996 24124 30008
rect 24176 29996 24182 30048
rect 26418 30036 26424 30048
rect 26379 30008 26424 30036
rect 26418 29996 26424 30008
rect 26476 30036 26482 30048
rect 27246 30036 27252 30048
rect 26476 30008 27252 30036
rect 26476 29996 26482 30008
rect 27246 29996 27252 30008
rect 27304 29996 27310 30048
rect 30742 30036 30748 30048
rect 30703 30008 30748 30036
rect 30742 29996 30748 30008
rect 30800 29996 30806 30048
rect 37366 30036 37372 30048
rect 37327 30008 37372 30036
rect 37366 29996 37372 30008
rect 37424 29996 37430 30048
rect 1104 29946 38548 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 38548 29946
rect 1104 29872 38548 29894
rect 3418 29832 3424 29844
rect 3379 29804 3424 29832
rect 3418 29792 3424 29804
rect 3476 29792 3482 29844
rect 6917 29835 6975 29841
rect 6917 29801 6929 29835
rect 6963 29832 6975 29835
rect 7374 29832 7380 29844
rect 6963 29804 7380 29832
rect 6963 29801 6975 29804
rect 6917 29795 6975 29801
rect 7374 29792 7380 29804
rect 7432 29792 7438 29844
rect 12526 29832 12532 29844
rect 12487 29804 12532 29832
rect 12526 29792 12532 29804
rect 12584 29792 12590 29844
rect 12710 29792 12716 29844
rect 12768 29832 12774 29844
rect 12805 29835 12863 29841
rect 12805 29832 12817 29835
rect 12768 29804 12817 29832
rect 12768 29792 12774 29804
rect 12805 29801 12817 29804
rect 12851 29801 12863 29835
rect 12805 29795 12863 29801
rect 14093 29835 14151 29841
rect 14093 29801 14105 29835
rect 14139 29832 14151 29835
rect 14182 29832 14188 29844
rect 14139 29804 14188 29832
rect 14139 29801 14151 29804
rect 14093 29795 14151 29801
rect 14182 29792 14188 29804
rect 14240 29792 14246 29844
rect 15470 29832 15476 29844
rect 15431 29804 15476 29832
rect 15470 29792 15476 29804
rect 15528 29792 15534 29844
rect 17586 29832 17592 29844
rect 17547 29804 17592 29832
rect 17586 29792 17592 29804
rect 17644 29792 17650 29844
rect 18233 29835 18291 29841
rect 18233 29801 18245 29835
rect 18279 29832 18291 29835
rect 18322 29832 18328 29844
rect 18279 29804 18328 29832
rect 18279 29801 18291 29804
rect 18233 29795 18291 29801
rect 18322 29792 18328 29804
rect 18380 29792 18386 29844
rect 18506 29832 18512 29844
rect 18467 29804 18512 29832
rect 18506 29792 18512 29804
rect 18564 29792 18570 29844
rect 19150 29832 19156 29844
rect 19111 29804 19156 29832
rect 19150 29792 19156 29804
rect 19208 29792 19214 29844
rect 21358 29832 21364 29844
rect 21319 29804 21364 29832
rect 21358 29792 21364 29804
rect 21416 29792 21422 29844
rect 22097 29835 22155 29841
rect 22097 29801 22109 29835
rect 22143 29832 22155 29835
rect 22186 29832 22192 29844
rect 22143 29804 22192 29832
rect 22143 29801 22155 29804
rect 22097 29795 22155 29801
rect 22186 29792 22192 29804
rect 22244 29792 22250 29844
rect 23290 29792 23296 29844
rect 23348 29832 23354 29844
rect 23753 29835 23811 29841
rect 23753 29832 23765 29835
rect 23348 29804 23765 29832
rect 23348 29792 23354 29804
rect 23753 29801 23765 29804
rect 23799 29801 23811 29835
rect 24210 29832 24216 29844
rect 24171 29804 24216 29832
rect 23753 29795 23811 29801
rect 12158 29724 12164 29776
rect 12216 29764 12222 29776
rect 12989 29767 13047 29773
rect 12989 29764 13001 29767
rect 12216 29736 13001 29764
rect 12216 29724 12222 29736
rect 12989 29733 13001 29736
rect 13035 29764 13047 29767
rect 13170 29764 13176 29776
rect 13035 29736 13176 29764
rect 13035 29733 13047 29736
rect 12989 29727 13047 29733
rect 13170 29724 13176 29736
rect 13228 29724 13234 29776
rect 1670 29696 1676 29708
rect 1631 29668 1676 29696
rect 1670 29656 1676 29668
rect 1728 29656 1734 29708
rect 7558 29696 7564 29708
rect 7519 29668 7564 29696
rect 7558 29656 7564 29668
rect 7616 29656 7622 29708
rect 7929 29699 7987 29705
rect 7929 29665 7941 29699
rect 7975 29696 7987 29699
rect 8018 29696 8024 29708
rect 7975 29668 8024 29696
rect 7975 29665 7987 29668
rect 7929 29659 7987 29665
rect 8018 29656 8024 29668
rect 8076 29656 8082 29708
rect 10137 29699 10195 29705
rect 10137 29665 10149 29699
rect 10183 29696 10195 29699
rect 10318 29696 10324 29708
rect 10183 29668 10324 29696
rect 10183 29665 10195 29668
rect 10137 29659 10195 29665
rect 10318 29656 10324 29668
rect 10376 29656 10382 29708
rect 10410 29656 10416 29708
rect 10468 29696 10474 29708
rect 11422 29696 11428 29708
rect 10468 29668 11428 29696
rect 10468 29656 10474 29668
rect 11422 29656 11428 29668
rect 11480 29656 11486 29708
rect 11698 29656 11704 29708
rect 11756 29696 11762 29708
rect 13630 29696 13636 29708
rect 11756 29668 11801 29696
rect 13591 29668 13636 29696
rect 11756 29656 11762 29668
rect 13630 29656 13636 29668
rect 13688 29656 13694 29708
rect 16298 29656 16304 29708
rect 16356 29696 16362 29708
rect 16485 29699 16543 29705
rect 16485 29696 16497 29699
rect 16356 29668 16497 29696
rect 16356 29656 16362 29668
rect 16485 29665 16497 29668
rect 16531 29696 16543 29699
rect 18524 29696 18552 29792
rect 19886 29696 19892 29708
rect 16531 29668 18552 29696
rect 19847 29668 19892 29696
rect 16531 29665 16543 29668
rect 16485 29659 16543 29665
rect 19886 29656 19892 29668
rect 19944 29656 19950 29708
rect 22554 29696 22560 29708
rect 22515 29668 22560 29696
rect 22554 29656 22560 29668
rect 22612 29656 22618 29708
rect 22738 29656 22744 29708
rect 22796 29696 22802 29708
rect 23198 29696 23204 29708
rect 22796 29668 23204 29696
rect 22796 29656 22802 29668
rect 23198 29656 23204 29668
rect 23256 29696 23262 29708
rect 23293 29699 23351 29705
rect 23293 29696 23305 29699
rect 23256 29668 23305 29696
rect 23256 29656 23262 29668
rect 23293 29665 23305 29668
rect 23339 29665 23351 29699
rect 23658 29696 23664 29708
rect 23293 29659 23351 29665
rect 23400 29668 23664 29696
rect 1397 29631 1455 29637
rect 1397 29597 1409 29631
rect 1443 29628 1455 29631
rect 2038 29628 2044 29640
rect 1443 29600 2044 29628
rect 1443 29597 1455 29600
rect 1397 29591 1455 29597
rect 2038 29588 2044 29600
rect 2096 29588 2102 29640
rect 7190 29628 7196 29640
rect 7151 29600 7196 29628
rect 7190 29588 7196 29600
rect 7248 29588 7254 29640
rect 10045 29631 10103 29637
rect 10045 29597 10057 29631
rect 10091 29597 10103 29631
rect 10594 29628 10600 29640
rect 10555 29600 10600 29628
rect 10045 29591 10103 29597
rect 7834 29560 7840 29572
rect 7795 29532 7840 29560
rect 7834 29520 7840 29532
rect 7892 29520 7898 29572
rect 10060 29560 10088 29591
rect 10594 29588 10600 29600
rect 10652 29588 10658 29640
rect 11238 29588 11244 29640
rect 11296 29628 11302 29640
rect 11885 29631 11943 29637
rect 11885 29628 11897 29631
rect 11296 29600 11897 29628
rect 11296 29588 11302 29600
rect 11885 29597 11897 29600
rect 11931 29597 11943 29631
rect 11885 29591 11943 29597
rect 15470 29588 15476 29640
rect 15528 29628 15534 29640
rect 16209 29631 16267 29637
rect 16209 29628 16221 29631
rect 15528 29600 16221 29628
rect 15528 29588 15534 29600
rect 16209 29597 16221 29600
rect 16255 29597 16267 29631
rect 16209 29591 16267 29597
rect 19981 29631 20039 29637
rect 19981 29597 19993 29631
rect 20027 29628 20039 29631
rect 20346 29628 20352 29640
rect 20027 29600 20352 29628
rect 20027 29597 20039 29600
rect 19981 29591 20039 29597
rect 20346 29588 20352 29600
rect 20404 29588 20410 29640
rect 22278 29588 22284 29640
rect 22336 29628 22342 29640
rect 22465 29631 22523 29637
rect 22465 29628 22477 29631
rect 22336 29600 22477 29628
rect 22336 29588 22342 29600
rect 22465 29597 22477 29600
rect 22511 29597 22523 29631
rect 22465 29591 22523 29597
rect 10134 29560 10140 29572
rect 10047 29532 10140 29560
rect 10134 29520 10140 29532
rect 10192 29560 10198 29572
rect 10873 29563 10931 29569
rect 10873 29560 10885 29563
rect 10192 29532 10885 29560
rect 10192 29520 10198 29532
rect 10873 29529 10885 29532
rect 10919 29529 10931 29563
rect 10873 29523 10931 29529
rect 11517 29563 11575 29569
rect 11517 29529 11529 29563
rect 11563 29560 11575 29563
rect 12066 29560 12072 29572
rect 11563 29532 12072 29560
rect 11563 29529 11575 29532
rect 11517 29523 11575 29529
rect 12066 29520 12072 29532
rect 12124 29520 12130 29572
rect 22480 29560 22508 29591
rect 22830 29588 22836 29640
rect 22888 29628 22894 29640
rect 23400 29637 23428 29668
rect 23658 29656 23664 29668
rect 23716 29656 23722 29708
rect 23768 29696 23796 29795
rect 24210 29792 24216 29804
rect 24268 29792 24274 29844
rect 27798 29832 27804 29844
rect 27759 29804 27804 29832
rect 27798 29792 27804 29804
rect 27856 29792 27862 29844
rect 28258 29832 28264 29844
rect 28219 29804 28264 29832
rect 28258 29792 28264 29804
rect 28316 29792 28322 29844
rect 29730 29832 29736 29844
rect 29691 29804 29736 29832
rect 29730 29792 29736 29804
rect 29788 29792 29794 29844
rect 31754 29792 31760 29844
rect 31812 29832 31818 29844
rect 32309 29835 32367 29841
rect 32309 29832 32321 29835
rect 31812 29804 32321 29832
rect 31812 29792 31818 29804
rect 32309 29801 32321 29804
rect 32355 29832 32367 29835
rect 32950 29832 32956 29844
rect 32355 29804 32956 29832
rect 32355 29801 32367 29804
rect 32309 29795 32367 29801
rect 32950 29792 32956 29804
rect 33008 29792 33014 29844
rect 27816 29764 27844 29792
rect 27816 29736 28488 29764
rect 25225 29699 25283 29705
rect 25225 29696 25237 29699
rect 23768 29668 25237 29696
rect 25225 29665 25237 29668
rect 25271 29665 25283 29699
rect 26510 29696 26516 29708
rect 26471 29668 26516 29696
rect 25225 29659 25283 29665
rect 26510 29656 26516 29668
rect 26568 29656 26574 29708
rect 28258 29696 28264 29708
rect 28219 29668 28264 29696
rect 28258 29656 28264 29668
rect 28316 29656 28322 29708
rect 28460 29705 28488 29736
rect 28445 29699 28503 29705
rect 28445 29665 28457 29699
rect 28491 29665 28503 29699
rect 28445 29659 28503 29665
rect 28813 29699 28871 29705
rect 28813 29665 28825 29699
rect 28859 29665 28871 29699
rect 28813 29659 28871 29665
rect 23385 29631 23443 29637
rect 23385 29628 23397 29631
rect 22888 29600 23397 29628
rect 22888 29588 22894 29600
rect 23385 29597 23397 29600
rect 23431 29597 23443 29631
rect 23385 29591 23443 29597
rect 23474 29588 23480 29640
rect 23532 29628 23538 29640
rect 24397 29631 24455 29637
rect 24397 29628 24409 29631
rect 23532 29600 24409 29628
rect 23532 29588 23538 29600
rect 24397 29597 24409 29600
rect 24443 29597 24455 29631
rect 24397 29591 24455 29597
rect 24489 29631 24547 29637
rect 24489 29597 24501 29631
rect 24535 29628 24547 29631
rect 24578 29628 24584 29640
rect 24535 29600 24584 29628
rect 24535 29597 24547 29600
rect 24489 29591 24547 29597
rect 24578 29588 24584 29600
rect 24636 29588 24642 29640
rect 24762 29588 24768 29640
rect 24820 29628 24826 29640
rect 25317 29631 25375 29637
rect 25317 29628 25329 29631
rect 24820 29600 25329 29628
rect 24820 29588 24826 29600
rect 25317 29597 25329 29600
rect 25363 29597 25375 29631
rect 25317 29591 25375 29597
rect 27982 29588 27988 29640
rect 28040 29628 28046 29640
rect 28828 29628 28856 29659
rect 29730 29656 29736 29708
rect 29788 29696 29794 29708
rect 30009 29699 30067 29705
rect 30009 29696 30021 29699
rect 29788 29668 30021 29696
rect 29788 29656 29794 29668
rect 30009 29665 30021 29668
rect 30055 29665 30067 29699
rect 30466 29696 30472 29708
rect 30427 29668 30472 29696
rect 30009 29659 30067 29665
rect 29270 29628 29276 29640
rect 28040 29600 29276 29628
rect 28040 29588 28046 29600
rect 29270 29588 29276 29600
rect 29328 29588 29334 29640
rect 29914 29628 29920 29640
rect 29875 29600 29920 29628
rect 29914 29588 29920 29600
rect 29972 29588 29978 29640
rect 30024 29628 30052 29659
rect 30466 29656 30472 29668
rect 30524 29656 30530 29708
rect 33686 29656 33692 29708
rect 33744 29696 33750 29708
rect 34885 29699 34943 29705
rect 34885 29696 34897 29699
rect 33744 29668 34897 29696
rect 33744 29656 33750 29668
rect 34885 29665 34897 29668
rect 34931 29696 34943 29699
rect 36538 29696 36544 29708
rect 34931 29668 36544 29696
rect 34931 29665 34943 29668
rect 34885 29659 34943 29665
rect 36538 29656 36544 29668
rect 36596 29656 36602 29708
rect 30745 29631 30803 29637
rect 30745 29628 30757 29631
rect 30024 29600 30757 29628
rect 30745 29597 30757 29600
rect 30791 29597 30803 29631
rect 30745 29591 30803 29597
rect 32950 29588 32956 29640
rect 33008 29628 33014 29640
rect 33962 29628 33968 29640
rect 33008 29600 33968 29628
rect 33008 29588 33014 29600
rect 33962 29588 33968 29600
rect 34020 29628 34026 29640
rect 34057 29631 34115 29637
rect 34057 29628 34069 29631
rect 34020 29600 34069 29628
rect 34020 29588 34026 29600
rect 34057 29597 34069 29600
rect 34103 29597 34115 29631
rect 34057 29591 34115 29597
rect 34146 29588 34152 29640
rect 34204 29628 34210 29640
rect 34204 29600 34249 29628
rect 34204 29588 34210 29600
rect 34330 29588 34336 29640
rect 34388 29628 34394 29640
rect 34977 29631 35035 29637
rect 34977 29628 34989 29631
rect 34388 29600 34989 29628
rect 34388 29588 34394 29600
rect 34977 29597 34989 29600
rect 35023 29597 35035 29631
rect 34977 29591 35035 29597
rect 23492 29560 23520 29588
rect 22480 29532 23520 29560
rect 25130 29520 25136 29572
rect 25188 29560 25194 29572
rect 25777 29563 25835 29569
rect 25777 29560 25789 29563
rect 25188 29532 25789 29560
rect 25188 29520 25194 29532
rect 25777 29529 25789 29532
rect 25823 29560 25835 29563
rect 26050 29560 26056 29572
rect 25823 29532 26056 29560
rect 25823 29529 25835 29532
rect 25777 29523 25835 29529
rect 26050 29520 26056 29532
rect 26108 29560 26114 29572
rect 27430 29560 27436 29572
rect 26108 29532 27436 29560
rect 26108 29520 26114 29532
rect 27430 29520 27436 29532
rect 27488 29520 27494 29572
rect 2774 29452 2780 29504
rect 2832 29492 2838 29504
rect 8570 29492 8576 29504
rect 2832 29464 2877 29492
rect 8531 29464 8576 29492
rect 2832 29452 2838 29464
rect 8570 29452 8576 29464
rect 8628 29452 8634 29504
rect 11698 29452 11704 29504
rect 11756 29492 11762 29504
rect 12710 29492 12716 29504
rect 11756 29464 12716 29492
rect 11756 29452 11762 29464
rect 12710 29452 12716 29464
rect 12768 29452 12774 29504
rect 20441 29495 20499 29501
rect 20441 29461 20453 29495
rect 20487 29492 20499 29495
rect 21266 29492 21272 29504
rect 20487 29464 21272 29492
rect 20487 29461 20499 29464
rect 20441 29455 20499 29461
rect 21266 29452 21272 29464
rect 21324 29452 21330 29504
rect 22922 29452 22928 29504
rect 22980 29492 22986 29504
rect 23290 29492 23296 29504
rect 22980 29464 23296 29492
rect 22980 29452 22986 29464
rect 23290 29452 23296 29464
rect 23348 29452 23354 29504
rect 26142 29492 26148 29504
rect 26103 29464 26148 29492
rect 26142 29452 26148 29464
rect 26200 29452 26206 29504
rect 26326 29452 26332 29504
rect 26384 29492 26390 29504
rect 26697 29495 26755 29501
rect 26697 29492 26709 29495
rect 26384 29464 26709 29492
rect 26384 29452 26390 29464
rect 26697 29461 26709 29464
rect 26743 29492 26755 29495
rect 26970 29492 26976 29504
rect 26743 29464 26976 29492
rect 26743 29461 26755 29464
rect 26697 29455 26755 29461
rect 26970 29452 26976 29464
rect 27028 29492 27034 29504
rect 27065 29495 27123 29501
rect 27065 29492 27077 29495
rect 27028 29464 27077 29492
rect 27028 29452 27034 29464
rect 27065 29461 27077 29464
rect 27111 29461 27123 29495
rect 29454 29492 29460 29504
rect 29415 29464 29460 29492
rect 27065 29455 27123 29461
rect 29454 29452 29460 29464
rect 29512 29452 29518 29504
rect 31202 29492 31208 29504
rect 31163 29464 31208 29492
rect 31202 29452 31208 29464
rect 31260 29452 31266 29504
rect 35437 29495 35495 29501
rect 35437 29461 35449 29495
rect 35483 29492 35495 29495
rect 35894 29492 35900 29504
rect 35483 29464 35900 29492
rect 35483 29461 35495 29464
rect 35437 29455 35495 29461
rect 35894 29452 35900 29464
rect 35952 29452 35958 29504
rect 1104 29402 38548 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 38548 29402
rect 1104 29328 38548 29350
rect 1670 29288 1676 29300
rect 1631 29260 1676 29288
rect 1670 29248 1676 29260
rect 1728 29248 1734 29300
rect 4890 29288 4896 29300
rect 4851 29260 4896 29288
rect 4890 29248 4896 29260
rect 4948 29248 4954 29300
rect 7837 29291 7895 29297
rect 7837 29257 7849 29291
rect 7883 29288 7895 29291
rect 8018 29288 8024 29300
rect 7883 29260 8024 29288
rect 7883 29257 7895 29260
rect 7837 29251 7895 29257
rect 8018 29248 8024 29260
rect 8076 29248 8082 29300
rect 10134 29288 10140 29300
rect 10095 29260 10140 29288
rect 10134 29248 10140 29260
rect 10192 29248 10198 29300
rect 11238 29288 11244 29300
rect 11199 29260 11244 29288
rect 11238 29248 11244 29260
rect 11296 29248 11302 29300
rect 12158 29288 12164 29300
rect 12119 29260 12164 29288
rect 12158 29248 12164 29260
rect 12216 29248 12222 29300
rect 13262 29288 13268 29300
rect 13223 29260 13268 29288
rect 13262 29248 13268 29260
rect 13320 29248 13326 29300
rect 15194 29288 15200 29300
rect 15155 29260 15200 29288
rect 15194 29248 15200 29260
rect 15252 29248 15258 29300
rect 16298 29288 16304 29300
rect 16259 29260 16304 29288
rect 16298 29248 16304 29260
rect 16356 29248 16362 29300
rect 22097 29291 22155 29297
rect 22097 29257 22109 29291
rect 22143 29288 22155 29291
rect 22738 29288 22744 29300
rect 22143 29260 22744 29288
rect 22143 29257 22155 29260
rect 22097 29251 22155 29257
rect 22738 29248 22744 29260
rect 22796 29248 22802 29300
rect 22833 29291 22891 29297
rect 22833 29257 22845 29291
rect 22879 29288 22891 29291
rect 23474 29288 23480 29300
rect 22879 29260 23480 29288
rect 22879 29257 22891 29260
rect 22833 29251 22891 29257
rect 23474 29248 23480 29260
rect 23532 29248 23538 29300
rect 27982 29288 27988 29300
rect 27943 29260 27988 29288
rect 27982 29248 27988 29260
rect 28040 29248 28046 29300
rect 28902 29288 28908 29300
rect 28863 29260 28908 29288
rect 28902 29248 28908 29260
rect 28960 29248 28966 29300
rect 33686 29288 33692 29300
rect 33647 29260 33692 29288
rect 33686 29248 33692 29260
rect 33744 29248 33750 29300
rect 33962 29288 33968 29300
rect 33923 29260 33968 29288
rect 33962 29248 33968 29260
rect 34020 29248 34026 29300
rect 34330 29288 34336 29300
rect 34291 29260 34336 29288
rect 34330 29248 34336 29260
rect 34388 29248 34394 29300
rect 36538 29288 36544 29300
rect 36499 29260 36544 29288
rect 36538 29248 36544 29260
rect 36596 29248 36602 29300
rect 2038 29152 2044 29164
rect 1951 29124 2044 29152
rect 2038 29112 2044 29124
rect 2096 29152 2102 29164
rect 3326 29152 3332 29164
rect 2096 29124 3332 29152
rect 2096 29112 2102 29124
rect 3326 29112 3332 29124
rect 3384 29112 3390 29164
rect 8481 29155 8539 29161
rect 8481 29121 8493 29155
rect 8527 29152 8539 29155
rect 8527 29124 8892 29152
rect 8527 29121 8539 29124
rect 8481 29115 8539 29121
rect 3605 29087 3663 29093
rect 3605 29084 3617 29087
rect 3436 29056 3617 29084
rect 3142 29016 3148 29028
rect 3103 28988 3148 29016
rect 3142 28976 3148 28988
rect 3200 29016 3206 29028
rect 3436 29016 3464 29056
rect 3605 29053 3617 29056
rect 3651 29053 3663 29087
rect 8570 29084 8576 29096
rect 8531 29056 8576 29084
rect 3605 29047 3663 29053
rect 8570 29044 8576 29056
rect 8628 29044 8634 29096
rect 8864 29093 8892 29124
rect 8849 29087 8907 29093
rect 8849 29053 8861 29087
rect 8895 29084 8907 29087
rect 8938 29084 8944 29096
rect 8895 29056 8944 29084
rect 8895 29053 8907 29056
rect 8849 29047 8907 29053
rect 8938 29044 8944 29056
rect 8996 29044 9002 29096
rect 11256 29084 11284 29248
rect 11514 29220 11520 29232
rect 11475 29192 11520 29220
rect 11514 29180 11520 29192
rect 11572 29180 11578 29232
rect 11333 29087 11391 29093
rect 11333 29084 11345 29087
rect 11256 29056 11345 29084
rect 11333 29053 11345 29056
rect 11379 29053 11391 29087
rect 11333 29047 11391 29053
rect 12805 29087 12863 29093
rect 12805 29053 12817 29087
rect 12851 29084 12863 29087
rect 13280 29084 13308 29248
rect 21174 29220 21180 29232
rect 21135 29192 21180 29220
rect 21174 29180 21180 29192
rect 21232 29180 21238 29232
rect 24765 29223 24823 29229
rect 24765 29189 24777 29223
rect 24811 29220 24823 29223
rect 24854 29220 24860 29232
rect 24811 29192 24860 29220
rect 24811 29189 24823 29192
rect 24765 29183 24823 29189
rect 24854 29180 24860 29192
rect 24912 29220 24918 29232
rect 27617 29223 27675 29229
rect 24912 29192 26556 29220
rect 24912 29180 24918 29192
rect 26528 29164 26556 29192
rect 27617 29189 27629 29223
rect 27663 29220 27675 29223
rect 28166 29220 28172 29232
rect 27663 29192 28172 29220
rect 27663 29189 27675 29192
rect 27617 29183 27675 29189
rect 28166 29180 28172 29192
rect 28224 29180 28230 29232
rect 29914 29220 29920 29232
rect 29380 29192 29920 29220
rect 13725 29155 13783 29161
rect 13725 29121 13737 29155
rect 13771 29152 13783 29155
rect 13771 29124 14136 29152
rect 13771 29121 13783 29124
rect 13725 29115 13783 29121
rect 14108 29096 14136 29124
rect 18598 29112 18604 29164
rect 18656 29152 18662 29164
rect 18785 29155 18843 29161
rect 18785 29152 18797 29155
rect 18656 29124 18797 29152
rect 18656 29112 18662 29124
rect 18785 29121 18797 29124
rect 18831 29152 18843 29155
rect 19613 29155 19671 29161
rect 19613 29152 19625 29155
rect 18831 29124 19625 29152
rect 18831 29121 18843 29124
rect 18785 29115 18843 29121
rect 19613 29121 19625 29124
rect 19659 29121 19671 29155
rect 19613 29115 19671 29121
rect 20257 29155 20315 29161
rect 20257 29121 20269 29155
rect 20303 29152 20315 29155
rect 21450 29152 21456 29164
rect 20303 29124 21456 29152
rect 20303 29121 20315 29124
rect 20257 29115 20315 29121
rect 12851 29056 13308 29084
rect 12851 29053 12863 29056
rect 12805 29047 12863 29053
rect 13446 29044 13452 29096
rect 13504 29084 13510 29096
rect 13817 29087 13875 29093
rect 13817 29084 13829 29087
rect 13504 29056 13829 29084
rect 13504 29044 13510 29056
rect 13817 29053 13829 29056
rect 13863 29084 13875 29087
rect 13906 29084 13912 29096
rect 13863 29056 13912 29084
rect 13863 29053 13875 29056
rect 13817 29047 13875 29053
rect 13906 29044 13912 29056
rect 13964 29044 13970 29096
rect 14090 29084 14096 29096
rect 14051 29056 14096 29084
rect 14090 29044 14096 29056
rect 14148 29044 14154 29096
rect 14458 29044 14464 29096
rect 14516 29084 14522 29096
rect 15746 29084 15752 29096
rect 14516 29056 15752 29084
rect 14516 29044 14522 29056
rect 15746 29044 15752 29056
rect 15804 29044 15810 29096
rect 18877 29087 18935 29093
rect 18877 29053 18889 29087
rect 18923 29084 18935 29087
rect 19242 29084 19248 29096
rect 18923 29056 19248 29084
rect 18923 29053 18935 29056
rect 18877 29047 18935 29053
rect 3200 28988 3464 29016
rect 7101 29019 7159 29025
rect 3200 28976 3206 28988
rect 7101 28985 7113 29019
rect 7147 29016 7159 29019
rect 7190 29016 7196 29028
rect 7147 28988 7196 29016
rect 7147 28985 7159 28988
rect 7101 28979 7159 28985
rect 7190 28976 7196 28988
rect 7248 28976 7254 29028
rect 7469 29019 7527 29025
rect 7469 28985 7481 29019
rect 7515 29016 7527 29019
rect 7558 29016 7564 29028
rect 7515 28988 7564 29016
rect 7515 28985 7527 28988
rect 7469 28979 7527 28985
rect 7558 28976 7564 28988
rect 7616 28976 7622 29028
rect 10410 28976 10416 29028
rect 10468 29016 10474 29028
rect 10505 29019 10563 29025
rect 10505 29016 10517 29019
rect 10468 28988 10517 29016
rect 10468 28976 10474 28988
rect 10505 28985 10517 28988
rect 10551 28985 10563 29019
rect 10505 28979 10563 28985
rect 11885 29019 11943 29025
rect 11885 28985 11897 29019
rect 11931 29016 11943 29019
rect 12066 29016 12072 29028
rect 11931 28988 12072 29016
rect 11931 28985 11943 28988
rect 11885 28979 11943 28985
rect 12066 28976 12072 28988
rect 12124 28976 12130 29028
rect 12342 28976 12348 29028
rect 12400 29016 12406 29028
rect 12713 29019 12771 29025
rect 12713 29016 12725 29019
rect 12400 28988 12725 29016
rect 12400 28976 12406 28988
rect 12713 28985 12725 28988
rect 12759 29016 12771 29019
rect 13630 29016 13636 29028
rect 12759 28988 13636 29016
rect 12759 28985 12771 28988
rect 12713 28979 12771 28985
rect 13630 28976 13636 28988
rect 13688 28976 13694 29028
rect 15102 28976 15108 29028
rect 15160 29016 15166 29028
rect 15838 29016 15844 29028
rect 15160 28988 15844 29016
rect 15160 28976 15166 28988
rect 15838 28976 15844 28988
rect 15896 28976 15902 29028
rect 16022 28976 16028 29028
rect 16080 29016 16086 29028
rect 16298 29016 16304 29028
rect 16080 28988 16304 29016
rect 16080 28976 16086 28988
rect 16298 28976 16304 28988
rect 16356 28976 16362 29028
rect 18693 29019 18751 29025
rect 18693 28985 18705 29019
rect 18739 29016 18751 29019
rect 18892 29016 18920 29047
rect 19242 29044 19248 29056
rect 19300 29044 19306 29096
rect 20346 29084 20352 29096
rect 20307 29056 20352 29084
rect 20346 29044 20352 29056
rect 20404 29044 20410 29096
rect 20916 29093 20944 29124
rect 21450 29112 21456 29124
rect 21508 29152 21514 29164
rect 21818 29152 21824 29164
rect 21508 29124 21824 29152
rect 21508 29112 21514 29124
rect 21818 29112 21824 29124
rect 21876 29112 21882 29164
rect 24029 29155 24087 29161
rect 24029 29121 24041 29155
rect 24075 29152 24087 29155
rect 24118 29152 24124 29164
rect 24075 29124 24124 29152
rect 24075 29121 24087 29124
rect 24029 29115 24087 29121
rect 24118 29112 24124 29124
rect 24176 29152 24182 29164
rect 25038 29152 25044 29164
rect 24176 29124 25044 29152
rect 24176 29112 24182 29124
rect 25038 29112 25044 29124
rect 25096 29152 25102 29164
rect 25096 29124 26464 29152
rect 25096 29112 25102 29124
rect 20901 29087 20959 29093
rect 20901 29053 20913 29087
rect 20947 29053 20959 29087
rect 21266 29084 21272 29096
rect 21227 29056 21272 29084
rect 20901 29047 20959 29053
rect 21266 29044 21272 29056
rect 21324 29044 21330 29096
rect 24854 29084 24860 29096
rect 24815 29056 24860 29084
rect 24854 29044 24860 29056
rect 24912 29044 24918 29096
rect 24946 29044 24952 29096
rect 25004 29084 25010 29096
rect 25593 29087 25651 29093
rect 25593 29084 25605 29087
rect 25004 29056 25605 29084
rect 25004 29044 25010 29056
rect 25593 29053 25605 29056
rect 25639 29053 25651 29087
rect 25593 29047 25651 29053
rect 25961 29087 26019 29093
rect 25961 29053 25973 29087
rect 26007 29084 26019 29087
rect 26050 29084 26056 29096
rect 26007 29056 26056 29084
rect 26007 29053 26019 29056
rect 25961 29047 26019 29053
rect 26050 29044 26056 29056
rect 26108 29044 26114 29096
rect 26436 29093 26464 29124
rect 26510 29112 26516 29164
rect 26568 29152 26574 29164
rect 26973 29155 27031 29161
rect 26973 29152 26985 29155
rect 26568 29124 26985 29152
rect 26568 29112 26574 29124
rect 26973 29121 26985 29124
rect 27019 29152 27031 29155
rect 27798 29152 27804 29164
rect 27019 29124 27804 29152
rect 27019 29121 27031 29124
rect 26973 29115 27031 29121
rect 27798 29112 27804 29124
rect 27856 29112 27862 29164
rect 29270 29152 29276 29164
rect 29231 29124 29276 29152
rect 29270 29112 29276 29124
rect 29328 29112 29334 29164
rect 26421 29087 26479 29093
rect 26421 29053 26433 29087
rect 26467 29053 26479 29087
rect 27430 29084 27436 29096
rect 27391 29056 27436 29084
rect 26421 29047 26479 29053
rect 18739 28988 18920 29016
rect 19337 29019 19395 29025
rect 18739 28985 18751 28988
rect 18693 28979 18751 28985
rect 19337 28985 19349 29019
rect 19383 28985 19395 29019
rect 19337 28979 19395 28985
rect 7742 28908 7748 28960
rect 7800 28948 7806 28960
rect 9582 28948 9588 28960
rect 7800 28920 9588 28948
rect 7800 28908 7806 28920
rect 9582 28908 9588 28920
rect 9640 28908 9646 28960
rect 12894 28908 12900 28960
rect 12952 28948 12958 28960
rect 12989 28951 13047 28957
rect 12989 28948 13001 28951
rect 12952 28920 13001 28948
rect 12952 28908 12958 28920
rect 12989 28917 13001 28920
rect 13035 28917 13047 28951
rect 12989 28911 13047 28917
rect 16669 28951 16727 28957
rect 16669 28917 16681 28951
rect 16715 28948 16727 28951
rect 17494 28948 17500 28960
rect 16715 28920 17500 28948
rect 16715 28917 16727 28920
rect 16669 28911 16727 28917
rect 17494 28908 17500 28920
rect 17552 28908 17558 28960
rect 19242 28908 19248 28960
rect 19300 28948 19306 28960
rect 19352 28948 19380 28979
rect 23106 28976 23112 29028
rect 23164 29016 23170 29028
rect 24026 29016 24032 29028
rect 23164 28988 24032 29016
rect 23164 28976 23170 28988
rect 24026 28976 24032 28988
rect 24084 28976 24090 29028
rect 24397 29019 24455 29025
rect 24397 28985 24409 29019
rect 24443 29016 24455 29019
rect 24762 29016 24768 29028
rect 24443 28988 24768 29016
rect 24443 28985 24455 28988
rect 24397 28979 24455 28985
rect 24762 28976 24768 28988
rect 24820 28976 24826 29028
rect 25038 29016 25044 29028
rect 24999 28988 25044 29016
rect 25038 28976 25044 28988
rect 25096 28976 25102 29028
rect 25222 29016 25228 29028
rect 25183 28988 25228 29016
rect 25222 28976 25228 28988
rect 25280 29016 25286 29028
rect 26237 29019 26295 29025
rect 26237 29016 26249 29019
rect 25280 28988 26249 29016
rect 25280 28976 25286 28988
rect 26237 28985 26249 28988
rect 26283 28985 26295 29019
rect 26436 29016 26464 29047
rect 27430 29044 27436 29056
rect 27488 29044 27494 29096
rect 29089 29087 29147 29093
rect 29089 29053 29101 29087
rect 29135 29084 29147 29087
rect 29178 29084 29184 29096
rect 29135 29056 29184 29084
rect 29135 29053 29147 29056
rect 29089 29047 29147 29053
rect 29178 29044 29184 29056
rect 29236 29084 29242 29096
rect 29380 29084 29408 29192
rect 29914 29180 29920 29192
rect 29972 29220 29978 29232
rect 30561 29223 30619 29229
rect 30561 29220 30573 29223
rect 29972 29192 30573 29220
rect 29972 29180 29978 29192
rect 30561 29189 30573 29192
rect 30607 29220 30619 29223
rect 30929 29223 30987 29229
rect 30929 29220 30941 29223
rect 30607 29192 30941 29220
rect 30607 29189 30619 29192
rect 30561 29183 30619 29189
rect 30929 29189 30941 29192
rect 30975 29189 30987 29223
rect 30929 29183 30987 29189
rect 29454 29112 29460 29164
rect 29512 29152 29518 29164
rect 30285 29155 30343 29161
rect 30285 29152 30297 29155
rect 29512 29124 30297 29152
rect 29512 29112 29518 29124
rect 30285 29121 30297 29124
rect 30331 29152 30343 29155
rect 30374 29152 30380 29164
rect 30331 29124 30380 29152
rect 30331 29121 30343 29124
rect 30285 29115 30343 29121
rect 30374 29112 30380 29124
rect 30432 29112 30438 29164
rect 29825 29087 29883 29093
rect 29825 29084 29837 29087
rect 29236 29056 29837 29084
rect 29236 29044 29242 29056
rect 29825 29053 29837 29056
rect 29871 29053 29883 29087
rect 30098 29084 30104 29096
rect 30059 29056 30104 29084
rect 29825 29047 29883 29053
rect 30098 29044 30104 29056
rect 30156 29044 30162 29096
rect 26694 29016 26700 29028
rect 26436 28988 26700 29016
rect 26237 28979 26295 28985
rect 26694 28976 26700 28988
rect 26752 29016 26758 29028
rect 27154 29016 27160 29028
rect 26752 28988 27160 29016
rect 26752 28976 26758 28988
rect 27154 28976 27160 28988
rect 27212 29016 27218 29028
rect 27249 29019 27307 29025
rect 27249 29016 27261 29019
rect 27212 28988 27261 29016
rect 27212 28976 27218 28988
rect 27249 28985 27261 28988
rect 27295 28985 27307 29019
rect 27249 28979 27307 28985
rect 28721 29019 28779 29025
rect 28721 28985 28733 29019
rect 28767 29016 28779 29019
rect 30116 29016 30144 29044
rect 28767 28988 30144 29016
rect 30944 29016 30972 29183
rect 31294 29152 31300 29164
rect 31255 29124 31300 29152
rect 31294 29112 31300 29124
rect 31352 29112 31358 29164
rect 35434 29152 35440 29164
rect 35395 29124 35440 29152
rect 35434 29112 35440 29124
rect 35492 29112 35498 29164
rect 31202 29084 31208 29096
rect 31163 29056 31208 29084
rect 31202 29044 31208 29056
rect 31260 29084 31266 29096
rect 31754 29084 31760 29096
rect 31260 29056 31760 29084
rect 31260 29044 31266 29056
rect 31754 29044 31760 29056
rect 31812 29044 31818 29096
rect 32033 29087 32091 29093
rect 32033 29053 32045 29087
rect 32079 29053 32091 29087
rect 32033 29047 32091 29053
rect 32125 29087 32183 29093
rect 32125 29053 32137 29087
rect 32171 29084 32183 29087
rect 32214 29084 32220 29096
rect 32171 29056 32220 29084
rect 32171 29053 32183 29056
rect 32125 29047 32183 29053
rect 32048 29016 32076 29047
rect 32214 29044 32220 29056
rect 32272 29044 32278 29096
rect 35161 29087 35219 29093
rect 35161 29053 35173 29087
rect 35207 29084 35219 29087
rect 35894 29084 35900 29096
rect 35207 29056 35900 29084
rect 35207 29053 35219 29056
rect 35161 29047 35219 29053
rect 35894 29044 35900 29056
rect 35952 29044 35958 29096
rect 30944 28988 32076 29016
rect 28767 28985 28779 28988
rect 28721 28979 28779 28985
rect 19300 28920 19380 28948
rect 22465 28951 22523 28957
rect 19300 28908 19306 28920
rect 22465 28917 22477 28951
rect 22511 28948 22523 28951
rect 22738 28948 22744 28960
rect 22511 28920 22744 28948
rect 22511 28917 22523 28920
rect 22465 28911 22523 28917
rect 22738 28908 22744 28920
rect 22796 28908 22802 28960
rect 25130 28948 25136 28960
rect 25091 28920 25136 28948
rect 25130 28908 25136 28920
rect 25188 28908 25194 28960
rect 26418 28908 26424 28960
rect 26476 28948 26482 28960
rect 26605 28951 26663 28957
rect 26605 28948 26617 28951
rect 26476 28920 26617 28948
rect 26476 28908 26482 28920
rect 26605 28917 26617 28920
rect 26651 28917 26663 28951
rect 28902 28948 28908 28960
rect 28863 28920 28908 28948
rect 26605 28911 26663 28917
rect 28902 28908 28908 28920
rect 28960 28908 28966 28960
rect 1104 28858 38548 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 38548 28858
rect 1104 28784 38548 28806
rect 3970 28704 3976 28756
rect 4028 28744 4034 28756
rect 4893 28747 4951 28753
rect 4893 28744 4905 28747
rect 4028 28716 4905 28744
rect 4028 28704 4034 28716
rect 4893 28713 4905 28716
rect 4939 28744 4951 28747
rect 4982 28744 4988 28756
rect 4939 28716 4988 28744
rect 4939 28713 4951 28716
rect 4893 28707 4951 28713
rect 4982 28704 4988 28716
rect 5040 28704 5046 28756
rect 11517 28747 11575 28753
rect 11517 28713 11529 28747
rect 11563 28744 11575 28747
rect 11698 28744 11704 28756
rect 11563 28716 11704 28744
rect 11563 28713 11575 28716
rect 11517 28707 11575 28713
rect 11698 28704 11704 28716
rect 11756 28704 11762 28756
rect 13449 28747 13507 28753
rect 13449 28713 13461 28747
rect 13495 28744 13507 28747
rect 14366 28744 14372 28756
rect 13495 28716 14372 28744
rect 13495 28713 13507 28716
rect 13449 28707 13507 28713
rect 14366 28704 14372 28716
rect 14424 28704 14430 28756
rect 16666 28744 16672 28756
rect 16627 28716 16672 28744
rect 16666 28704 16672 28716
rect 16724 28704 16730 28756
rect 19334 28744 19340 28756
rect 19295 28716 19340 28744
rect 19334 28704 19340 28716
rect 19392 28704 19398 28756
rect 20346 28744 20352 28756
rect 20307 28716 20352 28744
rect 20346 28704 20352 28716
rect 20404 28704 20410 28756
rect 26234 28744 26240 28756
rect 26195 28716 26240 28744
rect 26234 28704 26240 28716
rect 26292 28704 26298 28756
rect 28077 28747 28135 28753
rect 28077 28713 28089 28747
rect 28123 28744 28135 28747
rect 28258 28744 28264 28756
rect 28123 28716 28264 28744
rect 28123 28713 28135 28716
rect 28077 28707 28135 28713
rect 28258 28704 28264 28716
rect 28316 28704 28322 28756
rect 30374 28704 30380 28756
rect 30432 28744 30438 28756
rect 31202 28744 31208 28756
rect 30432 28716 31208 28744
rect 30432 28704 30438 28716
rect 31202 28704 31208 28716
rect 31260 28704 31266 28756
rect 35253 28747 35311 28753
rect 35253 28713 35265 28747
rect 35299 28744 35311 28747
rect 35434 28744 35440 28756
rect 35299 28716 35440 28744
rect 35299 28713 35311 28716
rect 35253 28707 35311 28713
rect 35434 28704 35440 28716
rect 35492 28704 35498 28756
rect 26602 28676 26608 28688
rect 25424 28648 26608 28676
rect 25424 28620 25452 28648
rect 26602 28636 26608 28648
rect 26660 28636 26666 28688
rect 26878 28676 26884 28688
rect 26839 28648 26884 28676
rect 26878 28636 26884 28648
rect 26936 28636 26942 28688
rect 30558 28636 30564 28688
rect 30616 28676 30622 28688
rect 30745 28679 30803 28685
rect 30745 28676 30757 28679
rect 30616 28648 30757 28676
rect 30616 28636 30622 28648
rect 30745 28645 30757 28648
rect 30791 28676 30803 28679
rect 31846 28676 31852 28688
rect 30791 28648 31852 28676
rect 30791 28645 30803 28648
rect 30745 28639 30803 28645
rect 31846 28636 31852 28648
rect 31904 28636 31910 28688
rect 1394 28568 1400 28620
rect 1452 28608 1458 28620
rect 1765 28611 1823 28617
rect 1765 28608 1777 28611
rect 1452 28580 1777 28608
rect 1452 28568 1458 28580
rect 1765 28577 1777 28580
rect 1811 28577 1823 28611
rect 1765 28571 1823 28577
rect 2038 28568 2044 28620
rect 2096 28568 2102 28620
rect 4706 28608 4712 28620
rect 4667 28580 4712 28608
rect 4706 28568 4712 28580
rect 4764 28568 4770 28620
rect 5350 28568 5356 28620
rect 5408 28608 5414 28620
rect 6641 28611 6699 28617
rect 6641 28608 6653 28611
rect 5408 28580 6653 28608
rect 5408 28568 5414 28580
rect 6641 28577 6653 28580
rect 6687 28577 6699 28611
rect 7006 28608 7012 28620
rect 6919 28580 7012 28608
rect 6641 28571 6699 28577
rect 7006 28568 7012 28580
rect 7064 28608 7070 28620
rect 7834 28608 7840 28620
rect 7064 28580 7840 28608
rect 7064 28568 7070 28580
rect 7834 28568 7840 28580
rect 7892 28568 7898 28620
rect 8662 28608 8668 28620
rect 8623 28580 8668 28608
rect 8662 28568 8668 28580
rect 8720 28568 8726 28620
rect 10594 28608 10600 28620
rect 10555 28580 10600 28608
rect 10594 28568 10600 28580
rect 10652 28568 10658 28620
rect 10870 28568 10876 28620
rect 10928 28608 10934 28620
rect 10965 28611 11023 28617
rect 10965 28608 10977 28611
rect 10928 28580 10977 28608
rect 10928 28568 10934 28580
rect 10965 28577 10977 28580
rect 11011 28577 11023 28611
rect 12894 28608 12900 28620
rect 12855 28580 12900 28608
rect 10965 28571 11023 28577
rect 12894 28568 12900 28580
rect 12952 28568 12958 28620
rect 13814 28608 13820 28620
rect 13775 28580 13820 28608
rect 13814 28568 13820 28580
rect 13872 28568 13878 28620
rect 15378 28568 15384 28620
rect 15436 28608 15442 28620
rect 15565 28611 15623 28617
rect 15565 28608 15577 28611
rect 15436 28580 15577 28608
rect 15436 28568 15442 28580
rect 15565 28577 15577 28580
rect 15611 28577 15623 28611
rect 22186 28608 22192 28620
rect 22147 28580 22192 28608
rect 15565 28571 15623 28577
rect 22186 28568 22192 28580
rect 22244 28568 22250 28620
rect 22922 28608 22928 28620
rect 22883 28580 22928 28608
rect 22922 28568 22928 28580
rect 22980 28568 22986 28620
rect 24397 28611 24455 28617
rect 24397 28577 24409 28611
rect 24443 28608 24455 28611
rect 24946 28608 24952 28620
rect 24443 28580 24952 28608
rect 24443 28577 24455 28580
rect 24397 28571 24455 28577
rect 24946 28568 24952 28580
rect 25004 28568 25010 28620
rect 25314 28608 25320 28620
rect 25275 28580 25320 28608
rect 25314 28568 25320 28580
rect 25372 28568 25378 28620
rect 25406 28568 25412 28620
rect 25464 28608 25470 28620
rect 25464 28580 25557 28608
rect 25464 28568 25470 28580
rect 26418 28568 26424 28620
rect 26476 28608 26482 28620
rect 26697 28611 26755 28617
rect 26697 28608 26709 28611
rect 26476 28580 26709 28608
rect 26476 28568 26482 28580
rect 26697 28577 26709 28580
rect 26743 28577 26755 28611
rect 26697 28571 26755 28577
rect 26789 28611 26847 28617
rect 26789 28577 26801 28611
rect 26835 28608 26847 28611
rect 28166 28608 28172 28620
rect 26835 28580 28172 28608
rect 26835 28577 26847 28580
rect 26789 28571 26847 28577
rect 28166 28568 28172 28580
rect 28224 28568 28230 28620
rect 28626 28608 28632 28620
rect 28587 28580 28632 28608
rect 28626 28568 28632 28580
rect 28684 28568 28690 28620
rect 28718 28568 28724 28620
rect 28776 28608 28782 28620
rect 28813 28611 28871 28617
rect 28813 28608 28825 28611
rect 28776 28580 28825 28608
rect 28776 28568 28782 28580
rect 28813 28577 28825 28580
rect 28859 28577 28871 28611
rect 28813 28571 28871 28577
rect 28997 28611 29055 28617
rect 28997 28577 29009 28611
rect 29043 28608 29055 28611
rect 29273 28611 29331 28617
rect 29273 28608 29285 28611
rect 29043 28580 29285 28608
rect 29043 28577 29055 28580
rect 28997 28571 29055 28577
rect 29273 28577 29285 28580
rect 29319 28577 29331 28611
rect 30282 28608 30288 28620
rect 30243 28580 30288 28608
rect 29273 28571 29331 28577
rect 30282 28568 30288 28580
rect 30340 28568 30346 28620
rect 30469 28611 30527 28617
rect 30469 28577 30481 28611
rect 30515 28577 30527 28611
rect 33778 28608 33784 28620
rect 33739 28580 33784 28608
rect 30469 28571 30527 28577
rect 1489 28543 1547 28549
rect 1489 28509 1501 28543
rect 1535 28540 1547 28543
rect 2056 28540 2084 28568
rect 1535 28512 2084 28540
rect 6733 28543 6791 28549
rect 1535 28509 1547 28512
rect 1489 28503 1547 28509
rect 6733 28509 6745 28543
rect 6779 28509 6791 28543
rect 7098 28540 7104 28552
rect 7059 28512 7104 28540
rect 6733 28503 6791 28509
rect 6748 28472 6776 28503
rect 7098 28500 7104 28512
rect 7156 28500 7162 28552
rect 8018 28540 8024 28552
rect 7979 28512 8024 28540
rect 8018 28500 8024 28512
rect 8076 28500 8082 28552
rect 11057 28543 11115 28549
rect 11057 28509 11069 28543
rect 11103 28540 11115 28543
rect 11238 28540 11244 28552
rect 11103 28512 11244 28540
rect 11103 28509 11115 28512
rect 11057 28503 11115 28509
rect 11238 28500 11244 28512
rect 11296 28500 11302 28552
rect 12989 28543 13047 28549
rect 12989 28509 13001 28543
rect 13035 28540 13047 28543
rect 13262 28540 13268 28552
rect 13035 28512 13268 28540
rect 13035 28509 13047 28512
rect 12989 28503 13047 28509
rect 13262 28500 13268 28512
rect 13320 28500 13326 28552
rect 13906 28500 13912 28552
rect 13964 28540 13970 28552
rect 14369 28543 14427 28549
rect 14369 28540 14381 28543
rect 13964 28512 14381 28540
rect 13964 28500 13970 28512
rect 14369 28509 14381 28512
rect 14415 28540 14427 28543
rect 15289 28543 15347 28549
rect 15289 28540 15301 28543
rect 14415 28512 15301 28540
rect 14415 28509 14427 28512
rect 14369 28503 14427 28509
rect 15289 28509 15301 28512
rect 15335 28540 15347 28543
rect 15470 28540 15476 28552
rect 15335 28512 15476 28540
rect 15335 28509 15347 28512
rect 15289 28503 15347 28509
rect 15470 28500 15476 28512
rect 15528 28500 15534 28552
rect 17494 28500 17500 28552
rect 17552 28540 17558 28552
rect 17773 28543 17831 28549
rect 17773 28540 17785 28543
rect 17552 28512 17785 28540
rect 17552 28500 17558 28512
rect 17773 28509 17785 28512
rect 17819 28509 17831 28543
rect 18046 28540 18052 28552
rect 18007 28512 18052 28540
rect 17773 28503 17831 28509
rect 18046 28500 18052 28512
rect 18104 28500 18110 28552
rect 22094 28500 22100 28552
rect 22152 28540 22158 28552
rect 22152 28512 22197 28540
rect 22152 28500 22158 28512
rect 22738 28500 22744 28552
rect 22796 28540 22802 28552
rect 23014 28540 23020 28552
rect 22796 28512 23020 28540
rect 22796 28500 22802 28512
rect 23014 28500 23020 28512
rect 23072 28500 23078 28552
rect 23753 28543 23811 28549
rect 23753 28509 23765 28543
rect 23799 28540 23811 28543
rect 24210 28540 24216 28552
rect 23799 28512 24216 28540
rect 23799 28509 23811 28512
rect 23753 28503 23811 28509
rect 24210 28500 24216 28512
rect 24268 28540 24274 28552
rect 24489 28543 24547 28549
rect 24489 28540 24501 28543
rect 24268 28512 24501 28540
rect 24268 28500 24274 28512
rect 24489 28509 24501 28512
rect 24535 28509 24547 28543
rect 24489 28503 24547 28509
rect 26326 28500 26332 28552
rect 26384 28540 26390 28552
rect 26513 28543 26571 28549
rect 26513 28540 26525 28543
rect 26384 28512 26525 28540
rect 26384 28500 26390 28512
rect 26513 28509 26525 28512
rect 26559 28509 26571 28543
rect 26513 28503 26571 28509
rect 26878 28500 26884 28552
rect 26936 28540 26942 28552
rect 27249 28543 27307 28549
rect 27249 28540 27261 28543
rect 26936 28512 27261 28540
rect 26936 28500 26942 28512
rect 27249 28509 27261 28512
rect 27295 28509 27307 28543
rect 27249 28503 27307 28509
rect 8036 28472 8064 28500
rect 10410 28472 10416 28484
rect 6748 28444 8064 28472
rect 10371 28444 10416 28472
rect 10410 28432 10416 28444
rect 10468 28432 10474 28484
rect 28445 28475 28503 28481
rect 28445 28441 28457 28475
rect 28491 28472 28503 28475
rect 30484 28472 30512 28571
rect 33778 28568 33784 28580
rect 33836 28568 33842 28620
rect 34149 28611 34207 28617
rect 34149 28577 34161 28611
rect 34195 28608 34207 28611
rect 34790 28608 34796 28620
rect 34195 28580 34796 28608
rect 34195 28577 34207 28580
rect 34149 28571 34207 28577
rect 34790 28568 34796 28580
rect 34848 28568 34854 28620
rect 33686 28540 33692 28552
rect 33647 28512 33692 28540
rect 33686 28500 33692 28512
rect 33744 28500 33750 28552
rect 34241 28543 34299 28549
rect 34241 28509 34253 28543
rect 34287 28509 34299 28543
rect 34241 28503 34299 28509
rect 31662 28472 31668 28484
rect 28491 28444 31668 28472
rect 28491 28441 28503 28444
rect 28445 28435 28503 28441
rect 31662 28432 31668 28444
rect 31720 28432 31726 28484
rect 32769 28475 32827 28481
rect 32769 28441 32781 28475
rect 32815 28472 32827 28475
rect 33134 28472 33140 28484
rect 32815 28444 33140 28472
rect 32815 28441 32827 28444
rect 32769 28435 32827 28441
rect 33134 28432 33140 28444
rect 33192 28472 33198 28484
rect 34256 28472 34284 28503
rect 33192 28444 34284 28472
rect 33192 28432 33198 28444
rect 3050 28404 3056 28416
rect 3011 28376 3056 28404
rect 3050 28364 3056 28376
rect 3108 28364 3114 28416
rect 6086 28404 6092 28416
rect 6047 28376 6092 28404
rect 6086 28364 6092 28376
rect 6144 28364 6150 28416
rect 9030 28364 9036 28416
rect 9088 28404 9094 28416
rect 9125 28407 9183 28413
rect 9125 28404 9137 28407
rect 9088 28376 9137 28404
rect 9088 28364 9094 28376
rect 9125 28373 9137 28376
rect 9171 28404 9183 28407
rect 9398 28404 9404 28416
rect 9171 28376 9404 28404
rect 9171 28373 9183 28376
rect 9125 28367 9183 28373
rect 9398 28364 9404 28376
rect 9456 28364 9462 28416
rect 13998 28404 14004 28416
rect 13959 28376 14004 28404
rect 13998 28364 14004 28376
rect 14056 28364 14062 28416
rect 19794 28404 19800 28416
rect 19755 28376 19800 28404
rect 19794 28364 19800 28376
rect 19852 28364 19858 28416
rect 27338 28364 27344 28416
rect 27396 28404 27402 28416
rect 27525 28407 27583 28413
rect 27525 28404 27537 28407
rect 27396 28376 27537 28404
rect 27396 28364 27402 28376
rect 27525 28373 27537 28376
rect 27571 28373 27583 28407
rect 27525 28367 27583 28373
rect 29273 28407 29331 28413
rect 29273 28373 29285 28407
rect 29319 28404 29331 28407
rect 29549 28407 29607 28413
rect 29549 28404 29561 28407
rect 29319 28376 29561 28404
rect 29319 28373 29331 28376
rect 29273 28367 29331 28373
rect 29549 28373 29561 28376
rect 29595 28404 29607 28407
rect 29917 28407 29975 28413
rect 29917 28404 29929 28407
rect 29595 28376 29929 28404
rect 29595 28373 29607 28376
rect 29549 28367 29607 28373
rect 29917 28373 29929 28376
rect 29963 28404 29975 28407
rect 30834 28404 30840 28416
rect 29963 28376 30840 28404
rect 29963 28373 29975 28376
rect 29917 28367 29975 28373
rect 30834 28364 30840 28376
rect 30892 28364 30898 28416
rect 31202 28404 31208 28416
rect 31115 28376 31208 28404
rect 31202 28364 31208 28376
rect 31260 28404 31266 28416
rect 32214 28404 32220 28416
rect 31260 28376 32220 28404
rect 31260 28364 31266 28376
rect 32214 28364 32220 28376
rect 32272 28364 32278 28416
rect 33226 28404 33232 28416
rect 33187 28376 33232 28404
rect 33226 28364 33232 28376
rect 33284 28364 33290 28416
rect 35802 28404 35808 28416
rect 35763 28376 35808 28404
rect 35802 28364 35808 28376
rect 35860 28364 35866 28416
rect 1104 28314 38548 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 38548 28314
rect 1104 28240 38548 28262
rect 1394 28160 1400 28212
rect 1452 28200 1458 28212
rect 1581 28203 1639 28209
rect 1581 28200 1593 28203
rect 1452 28172 1593 28200
rect 1452 28160 1458 28172
rect 1581 28169 1593 28172
rect 1627 28169 1639 28203
rect 2038 28200 2044 28212
rect 1999 28172 2044 28200
rect 1581 28163 1639 28169
rect 2038 28160 2044 28172
rect 2096 28160 2102 28212
rect 3694 28160 3700 28212
rect 3752 28200 3758 28212
rect 4706 28200 4712 28212
rect 3752 28172 4712 28200
rect 3752 28160 3758 28172
rect 4706 28160 4712 28172
rect 4764 28160 4770 28212
rect 6457 28203 6515 28209
rect 6457 28169 6469 28203
rect 6503 28200 6515 28203
rect 7006 28200 7012 28212
rect 6503 28172 7012 28200
rect 6503 28169 6515 28172
rect 6457 28163 6515 28169
rect 7006 28160 7012 28172
rect 7064 28160 7070 28212
rect 7377 28203 7435 28209
rect 7377 28169 7389 28203
rect 7423 28200 7435 28203
rect 8662 28200 8668 28212
rect 7423 28172 8668 28200
rect 7423 28169 7435 28172
rect 7377 28163 7435 28169
rect 8662 28160 8668 28172
rect 8720 28160 8726 28212
rect 10594 28200 10600 28212
rect 10555 28172 10600 28200
rect 10594 28160 10600 28172
rect 10652 28160 10658 28212
rect 11238 28200 11244 28212
rect 11199 28172 11244 28200
rect 11238 28160 11244 28172
rect 11296 28160 11302 28212
rect 11698 28160 11704 28212
rect 11756 28200 11762 28212
rect 11793 28203 11851 28209
rect 11793 28200 11805 28203
rect 11756 28172 11805 28200
rect 11756 28160 11762 28172
rect 11793 28169 11805 28172
rect 11839 28169 11851 28203
rect 11793 28163 11851 28169
rect 23109 28203 23167 28209
rect 23109 28169 23121 28203
rect 23155 28200 23167 28203
rect 23198 28200 23204 28212
rect 23155 28172 23204 28200
rect 23155 28169 23167 28172
rect 23109 28163 23167 28169
rect 23198 28160 23204 28172
rect 23256 28160 23262 28212
rect 24765 28203 24823 28209
rect 24765 28169 24777 28203
rect 24811 28200 24823 28203
rect 25406 28200 25412 28212
rect 24811 28172 25412 28200
rect 24811 28169 24823 28172
rect 24765 28163 24823 28169
rect 25406 28160 25412 28172
rect 25464 28160 25470 28212
rect 28166 28200 28172 28212
rect 28127 28172 28172 28200
rect 28166 28160 28172 28172
rect 28224 28160 28230 28212
rect 28258 28160 28264 28212
rect 28316 28200 28322 28212
rect 28629 28203 28687 28209
rect 28629 28200 28641 28203
rect 28316 28172 28641 28200
rect 28316 28160 28322 28172
rect 28629 28169 28641 28172
rect 28675 28200 28687 28203
rect 28718 28200 28724 28212
rect 28675 28172 28724 28200
rect 28675 28169 28687 28172
rect 28629 28163 28687 28169
rect 28718 28160 28724 28172
rect 28776 28160 28782 28212
rect 31662 28200 31668 28212
rect 31623 28172 31668 28200
rect 31662 28160 31668 28172
rect 31720 28160 31726 28212
rect 31754 28160 31760 28212
rect 31812 28200 31818 28212
rect 32493 28203 32551 28209
rect 32493 28200 32505 28203
rect 31812 28172 32505 28200
rect 31812 28160 31818 28172
rect 32493 28169 32505 28172
rect 32539 28169 32551 28203
rect 32493 28163 32551 28169
rect 34517 28203 34575 28209
rect 34517 28169 34529 28203
rect 34563 28200 34575 28203
rect 34790 28200 34796 28212
rect 34563 28172 34796 28200
rect 34563 28169 34575 28172
rect 34517 28163 34575 28169
rect 5721 28135 5779 28141
rect 5721 28101 5733 28135
rect 5767 28132 5779 28135
rect 7098 28132 7104 28144
rect 5767 28104 7104 28132
rect 5767 28101 5779 28104
rect 5721 28095 5779 28101
rect 7098 28092 7104 28104
rect 7156 28092 7162 28144
rect 8297 28135 8355 28141
rect 8297 28101 8309 28135
rect 8343 28132 8355 28135
rect 9766 28132 9772 28144
rect 8343 28104 9772 28132
rect 8343 28101 8355 28104
rect 8297 28095 8355 28101
rect 9766 28092 9772 28104
rect 9824 28092 9830 28144
rect 10229 28135 10287 28141
rect 10229 28101 10241 28135
rect 10275 28132 10287 28135
rect 10870 28132 10876 28144
rect 10275 28104 10876 28132
rect 10275 28101 10287 28104
rect 10229 28095 10287 28101
rect 10870 28092 10876 28104
rect 10928 28132 10934 28144
rect 18601 28135 18659 28141
rect 18601 28132 18613 28135
rect 10928 28104 18613 28132
rect 10928 28092 10934 28104
rect 18601 28101 18613 28104
rect 18647 28101 18659 28135
rect 19058 28132 19064 28144
rect 19019 28104 19064 28132
rect 18601 28095 18659 28101
rect 8938 28064 8944 28076
rect 8851 28036 8944 28064
rect 8938 28024 8944 28036
rect 8996 28064 9002 28076
rect 11238 28064 11244 28076
rect 8996 28036 11244 28064
rect 8996 28024 9002 28036
rect 11238 28024 11244 28036
rect 11296 28024 11302 28076
rect 13541 28067 13599 28073
rect 13541 28064 13553 28067
rect 11348 28036 13553 28064
rect 6089 27999 6147 28005
rect 6089 27965 6101 27999
rect 6135 27996 6147 27999
rect 7466 27996 7472 28008
rect 6135 27968 7472 27996
rect 6135 27965 6147 27968
rect 6089 27959 6147 27965
rect 7466 27956 7472 27968
rect 7524 27996 7530 28008
rect 8018 27996 8024 28008
rect 7524 27968 8024 27996
rect 7524 27956 7530 27968
rect 8018 27956 8024 27968
rect 8076 27956 8082 28008
rect 8846 27996 8852 28008
rect 8807 27968 8852 27996
rect 8846 27956 8852 27968
rect 8904 27956 8910 28008
rect 9677 27999 9735 28005
rect 9677 27965 9689 27999
rect 9723 27965 9735 27999
rect 9677 27959 9735 27965
rect 9692 27928 9720 27959
rect 9766 27956 9772 28008
rect 9824 27996 9830 28008
rect 9824 27968 9869 27996
rect 9824 27956 9830 27968
rect 10226 27956 10232 28008
rect 10284 27996 10290 28008
rect 11348 27996 11376 28036
rect 13541 28033 13553 28036
rect 13587 28033 13599 28067
rect 14366 28064 14372 28076
rect 14327 28036 14372 28064
rect 13541 28027 13599 28033
rect 14366 28024 14372 28036
rect 14424 28024 14430 28076
rect 18616 28064 18644 28095
rect 19058 28092 19064 28104
rect 19116 28092 19122 28144
rect 19426 28092 19432 28144
rect 19484 28092 19490 28144
rect 22002 28092 22008 28144
rect 22060 28092 22066 28144
rect 27614 28092 27620 28144
rect 27672 28132 27678 28144
rect 28905 28135 28963 28141
rect 28905 28132 28917 28135
rect 27672 28104 28917 28132
rect 27672 28092 27678 28104
rect 28905 28101 28917 28104
rect 28951 28101 28963 28135
rect 30282 28132 30288 28144
rect 30195 28104 30288 28132
rect 28905 28095 28963 28101
rect 30282 28092 30288 28104
rect 30340 28132 30346 28144
rect 30742 28132 30748 28144
rect 30340 28104 30748 28132
rect 30340 28092 30346 28104
rect 30742 28092 30748 28104
rect 30800 28132 30806 28144
rect 31297 28135 31355 28141
rect 31297 28132 31309 28135
rect 30800 28104 31309 28132
rect 30800 28092 30806 28104
rect 31297 28101 31309 28104
rect 31343 28101 31355 28135
rect 31297 28095 31355 28101
rect 19444 28064 19472 28092
rect 20901 28067 20959 28073
rect 18616 28036 19656 28064
rect 10284 27968 11376 27996
rect 13265 27999 13323 28005
rect 10284 27956 10290 27968
rect 13265 27965 13277 27999
rect 13311 27996 13323 27999
rect 13446 27996 13452 28008
rect 13311 27968 13452 27996
rect 13311 27965 13323 27968
rect 13265 27959 13323 27965
rect 13446 27956 13452 27968
rect 13504 27956 13510 28008
rect 13630 27956 13636 28008
rect 13688 27996 13694 28008
rect 14182 27996 14188 28008
rect 13688 27968 14188 27996
rect 13688 27956 13694 27968
rect 14182 27956 14188 27968
rect 14240 27996 14246 28008
rect 14277 27999 14335 28005
rect 14277 27996 14289 27999
rect 14240 27968 14289 27996
rect 14240 27956 14246 27968
rect 14277 27965 14289 27968
rect 14323 27965 14335 27999
rect 14277 27959 14335 27965
rect 18325 27999 18383 28005
rect 18325 27965 18337 27999
rect 18371 27996 18383 27999
rect 19242 27996 19248 28008
rect 18371 27968 19248 27996
rect 18371 27965 18383 27968
rect 18325 27959 18383 27965
rect 19242 27956 19248 27968
rect 19300 27956 19306 28008
rect 19628 28005 19656 28036
rect 20901 28033 20913 28067
rect 20947 28064 20959 28067
rect 22020 28064 22048 28092
rect 20947 28036 22048 28064
rect 22741 28067 22799 28073
rect 20947 28033 20959 28036
rect 20901 28027 20959 28033
rect 19429 27999 19487 28005
rect 19429 27965 19441 27999
rect 19475 27965 19487 27999
rect 19429 27959 19487 27965
rect 19613 27999 19671 28005
rect 19613 27965 19625 27999
rect 19659 27996 19671 27999
rect 19886 27996 19892 28008
rect 19659 27968 19892 27996
rect 19659 27965 19671 27968
rect 19613 27959 19671 27965
rect 8588 27900 9720 27928
rect 12713 27931 12771 27937
rect 5350 27860 5356 27872
rect 5311 27832 5356 27860
rect 5350 27820 5356 27832
rect 5408 27820 5414 27872
rect 7650 27860 7656 27872
rect 7611 27832 7656 27860
rect 7650 27820 7656 27832
rect 7708 27820 7714 27872
rect 8386 27820 8392 27872
rect 8444 27860 8450 27872
rect 8588 27869 8616 27900
rect 12713 27897 12725 27931
rect 12759 27928 12771 27931
rect 12894 27928 12900 27940
rect 12759 27900 12900 27928
rect 12759 27897 12771 27900
rect 12713 27891 12771 27897
rect 12894 27888 12900 27900
rect 12952 27928 12958 27940
rect 13354 27928 13360 27940
rect 12952 27900 13360 27928
rect 12952 27888 12958 27900
rect 13354 27888 13360 27900
rect 13412 27888 13418 27940
rect 16850 27888 16856 27940
rect 16908 27928 16914 27940
rect 17773 27931 17831 27937
rect 17773 27928 17785 27931
rect 16908 27900 17785 27928
rect 16908 27888 16914 27900
rect 17773 27897 17785 27900
rect 17819 27928 17831 27931
rect 18046 27928 18052 27940
rect 17819 27900 18052 27928
rect 17819 27897 17831 27900
rect 17773 27891 17831 27897
rect 18046 27888 18052 27900
rect 18104 27928 18110 27940
rect 19444 27928 19472 27959
rect 19886 27956 19892 27968
rect 19944 27956 19950 28008
rect 20533 27999 20591 28005
rect 20533 27965 20545 27999
rect 20579 27996 20591 27999
rect 21082 27996 21088 28008
rect 20579 27968 21088 27996
rect 20579 27965 20591 27968
rect 20533 27959 20591 27965
rect 21082 27956 21088 27968
rect 21140 27996 21146 28008
rect 21836 28005 21864 28036
rect 22741 28033 22753 28067
rect 22787 28064 22799 28067
rect 23014 28064 23020 28076
rect 22787 28036 23020 28064
rect 22787 28033 22799 28036
rect 22741 28027 22799 28033
rect 23014 28024 23020 28036
rect 23072 28064 23078 28076
rect 24854 28064 24860 28076
rect 23072 28036 24860 28064
rect 23072 28024 23078 28036
rect 24854 28024 24860 28036
rect 24912 28024 24918 28076
rect 21545 27999 21603 28005
rect 21545 27996 21557 27999
rect 21140 27968 21557 27996
rect 21140 27956 21146 27968
rect 21545 27965 21557 27968
rect 21591 27965 21603 27999
rect 21545 27959 21603 27965
rect 21821 27999 21879 28005
rect 21821 27965 21833 27999
rect 21867 27965 21879 27999
rect 21821 27959 21879 27965
rect 22005 27999 22063 28005
rect 22005 27965 22017 27999
rect 22051 27965 22063 27999
rect 22005 27959 22063 27965
rect 23937 27999 23995 28005
rect 23937 27965 23949 27999
rect 23983 27965 23995 27999
rect 24210 27996 24216 28008
rect 24171 27968 24216 27996
rect 23937 27959 23995 27965
rect 20073 27931 20131 27937
rect 20073 27928 20085 27931
rect 18104 27900 20085 27928
rect 18104 27888 18110 27900
rect 20073 27897 20085 27900
rect 20119 27897 20131 27931
rect 20073 27891 20131 27897
rect 20993 27931 21051 27937
rect 20993 27897 21005 27931
rect 21039 27928 21051 27931
rect 21266 27928 21272 27940
rect 21039 27900 21272 27928
rect 21039 27897 21051 27900
rect 20993 27891 21051 27897
rect 21266 27888 21272 27900
rect 21324 27888 21330 27940
rect 21358 27888 21364 27940
rect 21416 27928 21422 27940
rect 22020 27928 22048 27959
rect 23474 27928 23480 27940
rect 21416 27900 22048 27928
rect 23387 27900 23480 27928
rect 21416 27888 21422 27900
rect 23474 27888 23480 27900
rect 23532 27928 23538 27940
rect 23952 27928 23980 27959
rect 24210 27956 24216 27968
rect 24268 27956 24274 28008
rect 25317 27999 25375 28005
rect 25317 27965 25329 27999
rect 25363 27965 25375 27999
rect 25317 27959 25375 27965
rect 25225 27931 25283 27937
rect 25225 27928 25237 27931
rect 23532 27900 25237 27928
rect 23532 27888 23538 27900
rect 25225 27897 25237 27900
rect 25271 27928 25283 27931
rect 25332 27928 25360 27959
rect 25406 27956 25412 28008
rect 25464 27996 25470 28008
rect 25777 27999 25835 28005
rect 25777 27996 25789 27999
rect 25464 27968 25789 27996
rect 25464 27956 25470 27968
rect 25777 27965 25789 27968
rect 25823 27965 25835 27999
rect 25777 27959 25835 27965
rect 26418 27956 26424 28008
rect 26476 27996 26482 28008
rect 27338 27996 27344 28008
rect 26476 27968 27344 27996
rect 26476 27956 26482 27968
rect 27338 27956 27344 27968
rect 27396 27956 27402 28008
rect 27433 27999 27491 28005
rect 27433 27965 27445 27999
rect 27479 27996 27491 27999
rect 27706 27996 27712 28008
rect 27479 27968 27712 27996
rect 27479 27965 27491 27968
rect 27433 27959 27491 27965
rect 27706 27956 27712 27968
rect 27764 27996 27770 28008
rect 28166 27996 28172 28008
rect 27764 27968 28172 27996
rect 27764 27956 27770 27968
rect 28166 27956 28172 27968
rect 28224 27956 28230 28008
rect 28810 27956 28816 28008
rect 28868 27996 28874 28008
rect 29089 27999 29147 28005
rect 29089 27996 29101 27999
rect 28868 27968 29101 27996
rect 28868 27956 28874 27968
rect 29089 27965 29101 27968
rect 29135 27996 29147 27999
rect 29638 27996 29644 28008
rect 29135 27968 29644 27996
rect 29135 27965 29147 27968
rect 29089 27959 29147 27965
rect 29638 27956 29644 27968
rect 29696 27956 29702 28008
rect 29917 27999 29975 28005
rect 29917 27965 29929 27999
rect 29963 27996 29975 27999
rect 30466 27996 30472 28008
rect 29963 27968 30472 27996
rect 29963 27965 29975 27968
rect 29917 27959 29975 27965
rect 30466 27956 30472 27968
rect 30524 27956 30530 28008
rect 30558 27956 30564 28008
rect 30616 27996 30622 28008
rect 30653 27999 30711 28005
rect 30653 27996 30665 27999
rect 30616 27968 30665 27996
rect 30616 27956 30622 27968
rect 30653 27965 30665 27968
rect 30699 27965 30711 27999
rect 30834 27996 30840 28008
rect 30747 27968 30840 27996
rect 30653 27959 30711 27965
rect 30834 27956 30840 27968
rect 30892 27996 30898 28008
rect 31110 27996 31116 28008
rect 30892 27968 31116 27996
rect 30892 27956 30898 27968
rect 31110 27956 31116 27968
rect 31168 27956 31174 28008
rect 32508 27996 32536 28163
rect 34790 28160 34796 28172
rect 34848 28160 34854 28212
rect 33413 28067 33471 28073
rect 33413 28033 33425 28067
rect 33459 28064 33471 28067
rect 33778 28064 33784 28076
rect 33459 28036 33784 28064
rect 33459 28033 33471 28036
rect 33413 28027 33471 28033
rect 33778 28024 33784 28036
rect 33836 28064 33842 28076
rect 34057 28067 34115 28073
rect 34057 28064 34069 28067
rect 33836 28036 34069 28064
rect 33836 28024 33842 28036
rect 34057 28033 34069 28036
rect 34103 28033 34115 28067
rect 34057 28027 34115 28033
rect 35713 28067 35771 28073
rect 35713 28033 35725 28067
rect 35759 28064 35771 28067
rect 36078 28064 36084 28076
rect 35759 28036 36084 28064
rect 35759 28033 35771 28036
rect 35713 28027 35771 28033
rect 36078 28024 36084 28036
rect 36136 28024 36142 28076
rect 32674 27996 32680 28008
rect 32508 27968 32680 27996
rect 32674 27956 32680 27968
rect 32732 27956 32738 28008
rect 33134 27996 33140 28008
rect 33095 27968 33140 27996
rect 33134 27956 33140 27968
rect 33192 27956 33198 28008
rect 35802 27996 35808 28008
rect 35763 27968 35808 27996
rect 35802 27956 35808 27968
rect 35860 27956 35866 28008
rect 25498 27928 25504 27940
rect 25271 27900 25504 27928
rect 25271 27897 25283 27900
rect 25225 27891 25283 27897
rect 25498 27888 25504 27900
rect 25556 27888 25562 27940
rect 27157 27931 27215 27937
rect 27157 27897 27169 27931
rect 27203 27897 27215 27931
rect 27157 27891 27215 27897
rect 8573 27863 8631 27869
rect 8573 27860 8585 27863
rect 8444 27832 8585 27860
rect 8444 27820 8450 27832
rect 8573 27829 8585 27832
rect 8619 27829 8631 27863
rect 10962 27860 10968 27872
rect 10923 27832 10968 27860
rect 8573 27823 8631 27829
rect 10962 27820 10968 27832
rect 11020 27820 11026 27872
rect 15378 27860 15384 27872
rect 15339 27832 15384 27860
rect 15378 27820 15384 27832
rect 15436 27820 15442 27872
rect 15470 27820 15476 27872
rect 15528 27860 15534 27872
rect 15749 27863 15807 27869
rect 15749 27860 15761 27863
rect 15528 27832 15761 27860
rect 15528 27820 15534 27832
rect 15749 27829 15761 27832
rect 15795 27860 15807 27863
rect 16298 27860 16304 27872
rect 15795 27832 16304 27860
rect 15795 27829 15807 27832
rect 15749 27823 15807 27829
rect 16298 27820 16304 27832
rect 16356 27820 16362 27872
rect 17494 27860 17500 27872
rect 17455 27832 17500 27860
rect 17494 27820 17500 27832
rect 17552 27820 17558 27872
rect 22094 27820 22100 27872
rect 22152 27860 22158 27872
rect 22281 27863 22339 27869
rect 22281 27860 22293 27863
rect 22152 27832 22293 27860
rect 22152 27820 22158 27832
rect 22281 27829 22293 27832
rect 22327 27829 22339 27863
rect 23750 27860 23756 27872
rect 23711 27832 23756 27860
rect 22281 27823 22339 27829
rect 23750 27820 23756 27832
rect 23808 27820 23814 27872
rect 25314 27820 25320 27872
rect 25372 27860 25378 27872
rect 25409 27863 25467 27869
rect 25409 27860 25421 27863
rect 25372 27832 25421 27860
rect 25372 27820 25378 27832
rect 25409 27829 25421 27832
rect 25455 27829 25467 27863
rect 25409 27823 25467 27829
rect 26326 27820 26332 27872
rect 26384 27860 26390 27872
rect 26513 27863 26571 27869
rect 26513 27860 26525 27863
rect 26384 27832 26525 27860
rect 26384 27820 26390 27832
rect 26513 27829 26525 27832
rect 26559 27860 26571 27863
rect 26973 27863 27031 27869
rect 26973 27860 26985 27863
rect 26559 27832 26985 27860
rect 26559 27829 26571 27832
rect 26513 27823 26571 27829
rect 26973 27829 26985 27832
rect 27019 27860 27031 27863
rect 27172 27860 27200 27891
rect 27246 27888 27252 27940
rect 27304 27928 27310 27940
rect 27525 27931 27583 27937
rect 27525 27928 27537 27931
rect 27304 27900 27537 27928
rect 27304 27888 27310 27900
rect 27525 27897 27537 27900
rect 27571 27897 27583 27931
rect 27525 27891 27583 27897
rect 27893 27931 27951 27937
rect 27893 27897 27905 27931
rect 27939 27928 27951 27931
rect 28626 27928 28632 27940
rect 27939 27900 28632 27928
rect 27939 27897 27951 27900
rect 27893 27891 27951 27897
rect 28626 27888 28632 27900
rect 28684 27888 28690 27940
rect 29549 27931 29607 27937
rect 29549 27897 29561 27931
rect 29595 27928 29607 27931
rect 30098 27928 30104 27940
rect 29595 27900 30104 27928
rect 29595 27897 29607 27900
rect 29549 27891 29607 27897
rect 30098 27888 30104 27900
rect 30156 27928 30162 27940
rect 30576 27928 30604 27956
rect 30156 27900 30604 27928
rect 30156 27888 30162 27900
rect 33686 27860 33692 27872
rect 27019 27832 27200 27860
rect 33647 27832 33692 27860
rect 27019 27829 27031 27832
rect 26973 27823 27031 27829
rect 33686 27820 33692 27832
rect 33744 27820 33750 27872
rect 37366 27860 37372 27872
rect 37327 27832 37372 27860
rect 37366 27820 37372 27832
rect 37424 27820 37430 27872
rect 1104 27770 38548 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 38548 27770
rect 1104 27696 38548 27718
rect 7466 27656 7472 27668
rect 7427 27628 7472 27656
rect 7466 27616 7472 27628
rect 7524 27616 7530 27668
rect 8846 27656 8852 27668
rect 8588 27628 8852 27656
rect 6086 27548 6092 27600
rect 6144 27588 6150 27600
rect 8588 27597 8616 27628
rect 8846 27616 8852 27628
rect 8904 27616 8910 27668
rect 14182 27656 14188 27668
rect 14143 27628 14188 27656
rect 14182 27616 14188 27628
rect 14240 27616 14246 27668
rect 20346 27616 20352 27668
rect 20404 27656 20410 27668
rect 21085 27659 21143 27665
rect 21085 27656 21097 27659
rect 20404 27628 21097 27656
rect 20404 27616 20410 27628
rect 21085 27625 21097 27628
rect 21131 27656 21143 27659
rect 21358 27656 21364 27668
rect 21131 27628 21364 27656
rect 21131 27625 21143 27628
rect 21085 27619 21143 27625
rect 21358 27616 21364 27628
rect 21416 27616 21422 27668
rect 21545 27659 21603 27665
rect 21545 27625 21557 27659
rect 21591 27656 21603 27659
rect 21726 27656 21732 27668
rect 21591 27628 21732 27656
rect 21591 27625 21603 27628
rect 21545 27619 21603 27625
rect 21726 27616 21732 27628
rect 21784 27656 21790 27668
rect 22002 27656 22008 27668
rect 21784 27628 22008 27656
rect 21784 27616 21790 27628
rect 22002 27616 22008 27628
rect 22060 27616 22066 27668
rect 22097 27659 22155 27665
rect 22097 27625 22109 27659
rect 22143 27656 22155 27659
rect 22922 27656 22928 27668
rect 22143 27628 22928 27656
rect 22143 27625 22155 27628
rect 22097 27619 22155 27625
rect 22922 27616 22928 27628
rect 22980 27616 22986 27668
rect 23474 27656 23480 27668
rect 23400 27628 23480 27656
rect 8573 27591 8631 27597
rect 6144 27560 6868 27588
rect 6144 27548 6150 27560
rect 1486 27480 1492 27532
rect 1544 27520 1550 27532
rect 1673 27523 1731 27529
rect 1673 27520 1685 27523
rect 1544 27492 1685 27520
rect 1544 27480 1550 27492
rect 1673 27489 1685 27492
rect 1719 27489 1731 27523
rect 5718 27520 5724 27532
rect 5679 27492 5724 27520
rect 1673 27483 1731 27489
rect 5718 27480 5724 27492
rect 5776 27480 5782 27532
rect 5810 27480 5816 27532
rect 5868 27520 5874 27532
rect 5997 27523 6055 27529
rect 5997 27520 6009 27523
rect 5868 27492 6009 27520
rect 5868 27480 5874 27492
rect 5997 27489 6009 27492
rect 6043 27489 6055 27523
rect 6638 27520 6644 27532
rect 6599 27492 6644 27520
rect 5997 27483 6055 27489
rect 6638 27480 6644 27492
rect 6696 27480 6702 27532
rect 6840 27529 6868 27560
rect 8573 27557 8585 27591
rect 8619 27557 8631 27591
rect 8573 27551 8631 27557
rect 11701 27591 11759 27597
rect 11701 27557 11713 27591
rect 11747 27588 11759 27591
rect 11793 27591 11851 27597
rect 11793 27588 11805 27591
rect 11747 27560 11805 27588
rect 11747 27557 11759 27560
rect 11701 27551 11759 27557
rect 11793 27557 11805 27560
rect 11839 27588 11851 27591
rect 12342 27588 12348 27600
rect 11839 27560 12348 27588
rect 11839 27557 11851 27560
rect 11793 27551 11851 27557
rect 12342 27548 12348 27560
rect 12400 27548 12406 27600
rect 12529 27591 12587 27597
rect 12529 27557 12541 27591
rect 12575 27588 12587 27591
rect 13814 27588 13820 27600
rect 12575 27560 13820 27588
rect 12575 27557 12587 27560
rect 12529 27551 12587 27557
rect 13814 27548 13820 27560
rect 13872 27548 13878 27600
rect 6825 27523 6883 27529
rect 6825 27489 6837 27523
rect 6871 27489 6883 27523
rect 8018 27520 8024 27532
rect 6825 27483 6883 27489
rect 7116 27492 8024 27520
rect 1397 27455 1455 27461
rect 1397 27421 1409 27455
rect 1443 27452 1455 27455
rect 2038 27452 2044 27464
rect 1443 27424 2044 27452
rect 1443 27421 1455 27424
rect 1397 27415 1455 27421
rect 2038 27412 2044 27424
rect 2096 27412 2102 27464
rect 3050 27452 3056 27464
rect 3011 27424 3056 27452
rect 3050 27412 3056 27424
rect 3108 27412 3114 27464
rect 5537 27455 5595 27461
rect 5537 27421 5549 27455
rect 5583 27452 5595 27455
rect 7116 27452 7144 27492
rect 8018 27480 8024 27492
rect 8076 27480 8082 27532
rect 8110 27480 8116 27532
rect 8168 27520 8174 27532
rect 8205 27523 8263 27529
rect 8205 27520 8217 27523
rect 8168 27492 8217 27520
rect 8168 27480 8174 27492
rect 8205 27489 8217 27492
rect 8251 27489 8263 27523
rect 11054 27520 11060 27532
rect 11015 27492 11060 27520
rect 8205 27483 8263 27489
rect 11054 27480 11060 27492
rect 11112 27520 11118 27532
rect 11514 27520 11520 27532
rect 11112 27492 11520 27520
rect 11112 27480 11118 27492
rect 11514 27480 11520 27492
rect 11572 27480 11578 27532
rect 13354 27520 13360 27532
rect 13315 27492 13360 27520
rect 13354 27480 13360 27492
rect 13412 27480 13418 27532
rect 15286 27520 15292 27532
rect 15247 27492 15292 27520
rect 15286 27480 15292 27492
rect 15344 27480 15350 27532
rect 16390 27480 16396 27532
rect 16448 27520 16454 27532
rect 16577 27523 16635 27529
rect 16577 27520 16589 27523
rect 16448 27492 16589 27520
rect 16448 27480 16454 27492
rect 16577 27489 16589 27492
rect 16623 27489 16635 27523
rect 16577 27483 16635 27489
rect 17034 27480 17040 27532
rect 17092 27520 17098 27532
rect 17678 27520 17684 27532
rect 17092 27492 17684 27520
rect 17092 27480 17098 27492
rect 17678 27480 17684 27492
rect 17736 27480 17742 27532
rect 18690 27480 18696 27532
rect 18748 27520 18754 27532
rect 18785 27523 18843 27529
rect 18785 27520 18797 27523
rect 18748 27492 18797 27520
rect 18748 27480 18754 27492
rect 18785 27489 18797 27492
rect 18831 27489 18843 27523
rect 22830 27520 22836 27532
rect 22743 27492 22836 27520
rect 18785 27483 18843 27489
rect 22830 27480 22836 27492
rect 22888 27520 22894 27532
rect 23400 27520 23428 27628
rect 23474 27616 23480 27628
rect 23532 27616 23538 27668
rect 27246 27656 27252 27668
rect 26160 27628 27252 27656
rect 23934 27588 23940 27600
rect 23895 27560 23940 27588
rect 23934 27548 23940 27560
rect 23992 27548 23998 27600
rect 25961 27591 26019 27597
rect 25961 27557 25973 27591
rect 26007 27588 26019 27591
rect 26160 27588 26188 27628
rect 27246 27616 27252 27628
rect 27304 27616 27310 27668
rect 27706 27656 27712 27668
rect 27667 27628 27712 27656
rect 27706 27616 27712 27628
rect 27764 27616 27770 27668
rect 28258 27656 28264 27668
rect 27816 27628 28264 27656
rect 27816 27588 27844 27628
rect 28258 27616 28264 27628
rect 28316 27616 28322 27668
rect 28626 27616 28632 27668
rect 28684 27656 28690 27668
rect 28684 27628 28948 27656
rect 28684 27616 28690 27628
rect 26007 27560 26188 27588
rect 27540 27560 27844 27588
rect 28920 27588 28948 27628
rect 28994 27616 29000 27668
rect 29052 27656 29058 27668
rect 29362 27656 29368 27668
rect 29052 27628 29368 27656
rect 29052 27616 29058 27628
rect 29362 27616 29368 27628
rect 29420 27616 29426 27668
rect 29638 27656 29644 27668
rect 29599 27628 29644 27656
rect 29638 27616 29644 27628
rect 29696 27616 29702 27668
rect 29273 27591 29331 27597
rect 29273 27588 29285 27591
rect 28920 27560 29285 27588
rect 26007 27557 26019 27560
rect 25961 27551 26019 27557
rect 22888 27492 23428 27520
rect 22888 27480 22894 27492
rect 23750 27480 23756 27532
rect 23808 27520 23814 27532
rect 23845 27523 23903 27529
rect 23845 27520 23857 27523
rect 23808 27492 23857 27520
rect 23808 27480 23814 27492
rect 23845 27489 23857 27492
rect 23891 27489 23903 27523
rect 24670 27520 24676 27532
rect 24631 27492 24676 27520
rect 23845 27483 23903 27489
rect 24670 27480 24676 27492
rect 24728 27480 24734 27532
rect 26602 27480 26608 27532
rect 26660 27520 26666 27532
rect 26881 27523 26939 27529
rect 26881 27520 26893 27523
rect 26660 27492 26893 27520
rect 26660 27480 26666 27492
rect 26881 27489 26893 27492
rect 26927 27489 26939 27523
rect 26881 27483 26939 27489
rect 5583 27424 7144 27452
rect 5583 27421 5595 27424
rect 5537 27415 5595 27421
rect 11698 27412 11704 27464
rect 11756 27452 11762 27464
rect 12161 27455 12219 27461
rect 12161 27452 12173 27455
rect 11756 27424 12173 27452
rect 11756 27412 11762 27424
rect 12161 27421 12173 27424
rect 12207 27421 12219 27455
rect 16298 27452 16304 27464
rect 16211 27424 16304 27452
rect 12161 27415 12219 27421
rect 16298 27412 16304 27424
rect 16356 27452 16362 27464
rect 17494 27452 17500 27464
rect 16356 27424 17500 27452
rect 16356 27412 16362 27424
rect 17494 27412 17500 27424
rect 17552 27412 17558 27464
rect 22186 27452 22192 27464
rect 22147 27424 22192 27452
rect 22186 27412 22192 27424
rect 22244 27412 22250 27464
rect 23661 27455 23719 27461
rect 23661 27421 23673 27455
rect 23707 27452 23719 27455
rect 24688 27452 24716 27480
rect 23707 27424 24716 27452
rect 23707 27421 23719 27424
rect 23661 27415 23719 27421
rect 24762 27412 24768 27464
rect 24820 27452 24826 27464
rect 24820 27424 24865 27452
rect 24820 27412 24826 27424
rect 5169 27387 5227 27393
rect 5169 27353 5181 27387
rect 5215 27353 5227 27387
rect 5169 27347 5227 27353
rect 9953 27387 10011 27393
rect 9953 27353 9965 27387
rect 9999 27384 10011 27387
rect 10502 27384 10508 27396
rect 9999 27356 10508 27384
rect 9999 27353 10011 27356
rect 9953 27347 10011 27353
rect 3418 27316 3424 27328
rect 3379 27288 3424 27316
rect 3418 27276 3424 27288
rect 3476 27276 3482 27328
rect 4890 27276 4896 27328
rect 4948 27316 4954 27328
rect 4985 27319 5043 27325
rect 4985 27316 4997 27319
rect 4948 27288 4997 27316
rect 4948 27276 4954 27288
rect 4985 27285 4997 27288
rect 5031 27316 5043 27319
rect 5184 27316 5212 27347
rect 10502 27344 10508 27356
rect 10560 27344 10566 27396
rect 18598 27344 18604 27396
rect 18656 27384 18662 27396
rect 18874 27384 18880 27396
rect 18656 27356 18880 27384
rect 18656 27344 18662 27356
rect 18874 27344 18880 27356
rect 18932 27384 18938 27396
rect 18969 27387 19027 27393
rect 18969 27384 18981 27387
rect 18932 27356 18981 27384
rect 18932 27344 18938 27356
rect 18969 27353 18981 27356
rect 19015 27353 19027 27387
rect 18969 27347 19027 27353
rect 26329 27387 26387 27393
rect 26329 27353 26341 27387
rect 26375 27384 26387 27387
rect 26786 27384 26792 27396
rect 26375 27356 26792 27384
rect 26375 27353 26387 27356
rect 26329 27347 26387 27353
rect 26786 27344 26792 27356
rect 26844 27344 26850 27396
rect 5031 27288 5212 27316
rect 7929 27319 7987 27325
rect 5031 27285 5043 27288
rect 4985 27279 5043 27285
rect 7929 27285 7941 27319
rect 7975 27316 7987 27319
rect 8202 27316 8208 27328
rect 7975 27288 8208 27316
rect 7975 27285 7987 27288
rect 7929 27279 7987 27285
rect 8202 27276 8208 27288
rect 8260 27276 8266 27328
rect 9306 27316 9312 27328
rect 9267 27288 9312 27316
rect 9306 27276 9312 27288
rect 9364 27276 9370 27328
rect 10318 27316 10324 27328
rect 10279 27288 10324 27316
rect 10318 27276 10324 27288
rect 10376 27276 10382 27328
rect 10778 27316 10784 27328
rect 10739 27288 10784 27316
rect 10778 27276 10784 27288
rect 10836 27276 10842 27328
rect 11698 27276 11704 27328
rect 11756 27316 11762 27328
rect 11931 27319 11989 27325
rect 11931 27316 11943 27319
rect 11756 27288 11943 27316
rect 11756 27276 11762 27288
rect 11931 27285 11943 27288
rect 11977 27285 11989 27319
rect 12066 27316 12072 27328
rect 12027 27288 12072 27316
rect 11931 27279 11989 27285
rect 12066 27276 12072 27288
rect 12124 27276 12130 27328
rect 13538 27316 13544 27328
rect 13499 27288 13544 27316
rect 13538 27276 13544 27288
rect 13596 27276 13602 27328
rect 15470 27316 15476 27328
rect 15431 27288 15476 27316
rect 15470 27276 15476 27288
rect 15528 27276 15534 27328
rect 17678 27316 17684 27328
rect 17639 27288 17684 27316
rect 17678 27276 17684 27288
rect 17736 27276 17742 27328
rect 19334 27316 19340 27328
rect 19295 27288 19340 27316
rect 19334 27276 19340 27288
rect 19392 27276 19398 27328
rect 25406 27316 25412 27328
rect 25367 27288 25412 27316
rect 25406 27276 25412 27288
rect 25464 27276 25470 27328
rect 26418 27276 26424 27328
rect 26476 27316 26482 27328
rect 26697 27319 26755 27325
rect 26697 27316 26709 27319
rect 26476 27288 26709 27316
rect 26476 27276 26482 27288
rect 26697 27285 26709 27288
rect 26743 27285 26755 27319
rect 26896 27316 26924 27483
rect 26970 27344 26976 27396
rect 27028 27384 27034 27396
rect 27065 27387 27123 27393
rect 27065 27384 27077 27387
rect 27028 27356 27077 27384
rect 27028 27344 27034 27356
rect 27065 27353 27077 27356
rect 27111 27384 27123 27387
rect 27540 27384 27568 27560
rect 29273 27557 29285 27560
rect 29319 27557 29331 27591
rect 32674 27588 32680 27600
rect 32635 27560 32680 27588
rect 29273 27551 29331 27557
rect 32674 27548 32680 27560
rect 32732 27548 32738 27600
rect 33594 27548 33600 27600
rect 33652 27588 33658 27600
rect 36078 27588 36084 27600
rect 33652 27560 36084 27588
rect 33652 27548 33658 27560
rect 36078 27548 36084 27560
rect 36136 27588 36142 27600
rect 36136 27560 36584 27588
rect 36136 27548 36142 27560
rect 27982 27520 27988 27532
rect 27943 27492 27988 27520
rect 27982 27480 27988 27492
rect 28040 27480 28046 27532
rect 28810 27520 28816 27532
rect 28771 27492 28816 27520
rect 28810 27480 28816 27492
rect 28868 27480 28874 27532
rect 28994 27480 29000 27532
rect 29052 27520 29058 27532
rect 29362 27520 29368 27532
rect 29052 27492 29368 27520
rect 29052 27480 29058 27492
rect 29362 27480 29368 27492
rect 29420 27480 29426 27532
rect 31110 27520 31116 27532
rect 31071 27492 31116 27520
rect 31110 27480 31116 27492
rect 31168 27480 31174 27532
rect 32125 27523 32183 27529
rect 32125 27489 32137 27523
rect 32171 27520 32183 27523
rect 32214 27520 32220 27532
rect 32171 27492 32220 27520
rect 32171 27489 32183 27492
rect 32125 27483 32183 27489
rect 32214 27480 32220 27492
rect 32272 27480 32278 27532
rect 32309 27523 32367 27529
rect 32309 27489 32321 27523
rect 32355 27489 32367 27523
rect 32309 27483 32367 27489
rect 33505 27523 33563 27529
rect 33505 27489 33517 27523
rect 33551 27520 33563 27523
rect 34514 27520 34520 27532
rect 33551 27492 34520 27520
rect 33551 27489 33563 27492
rect 33505 27483 33563 27489
rect 28074 27452 28080 27464
rect 28035 27424 28080 27452
rect 28074 27412 28080 27424
rect 28132 27412 28138 27464
rect 28905 27455 28963 27461
rect 28905 27421 28917 27455
rect 28951 27421 28963 27455
rect 28905 27415 28963 27421
rect 31205 27455 31263 27461
rect 31205 27421 31217 27455
rect 31251 27452 31263 27455
rect 31846 27452 31852 27464
rect 31251 27424 31852 27452
rect 31251 27421 31263 27424
rect 31205 27415 31263 27421
rect 27111 27356 27568 27384
rect 27111 27353 27123 27356
rect 27065 27347 27123 27353
rect 27890 27344 27896 27396
rect 27948 27384 27954 27396
rect 28920 27384 28948 27415
rect 31846 27412 31852 27424
rect 31904 27452 31910 27464
rect 32324 27452 32352 27483
rect 34514 27480 34520 27492
rect 34572 27480 34578 27532
rect 35618 27480 35624 27532
rect 35676 27520 35682 27532
rect 35805 27523 35863 27529
rect 35805 27520 35817 27523
rect 35676 27492 35817 27520
rect 35676 27480 35682 27492
rect 35805 27489 35817 27492
rect 35851 27489 35863 27523
rect 35805 27483 35863 27489
rect 31904 27424 32352 27452
rect 35897 27455 35955 27461
rect 31904 27412 31910 27424
rect 35897 27421 35909 27455
rect 35943 27452 35955 27455
rect 35986 27452 35992 27464
rect 35943 27424 35992 27452
rect 35943 27421 35955 27424
rect 35897 27415 35955 27421
rect 35986 27412 35992 27424
rect 36044 27412 36050 27464
rect 36556 27452 36584 27560
rect 36633 27523 36691 27529
rect 36633 27489 36645 27523
rect 36679 27520 36691 27523
rect 37182 27520 37188 27532
rect 36679 27492 37188 27520
rect 36679 27489 36691 27492
rect 36633 27483 36691 27489
rect 37182 27480 37188 27492
rect 37240 27480 37246 27532
rect 36725 27455 36783 27461
rect 36725 27452 36737 27455
rect 36556 27424 36737 27452
rect 36725 27421 36737 27424
rect 36771 27421 36783 27455
rect 36725 27415 36783 27421
rect 34701 27387 34759 27393
rect 34701 27384 34713 27387
rect 27948 27356 28948 27384
rect 33152 27356 34713 27384
rect 27948 27344 27954 27356
rect 33152 27328 33180 27356
rect 34701 27353 34713 27356
rect 34747 27353 34759 27387
rect 34701 27347 34759 27353
rect 27433 27319 27491 27325
rect 27433 27316 27445 27319
rect 26896 27288 27445 27316
rect 26697 27279 26755 27285
rect 27433 27285 27445 27288
rect 27479 27316 27491 27319
rect 29730 27316 29736 27328
rect 27479 27288 29736 27316
rect 27479 27285 27491 27288
rect 27433 27279 27491 27285
rect 29730 27276 29736 27288
rect 29788 27276 29794 27328
rect 29822 27276 29828 27328
rect 29880 27316 29886 27328
rect 30193 27319 30251 27325
rect 30193 27316 30205 27319
rect 29880 27288 30205 27316
rect 29880 27276 29886 27288
rect 30193 27285 30205 27288
rect 30239 27316 30251 27319
rect 30466 27316 30472 27328
rect 30239 27288 30472 27316
rect 30239 27285 30251 27288
rect 30193 27279 30251 27285
rect 30466 27276 30472 27288
rect 30524 27316 30530 27328
rect 30834 27316 30840 27328
rect 30524 27288 30840 27316
rect 30524 27276 30530 27288
rect 30834 27276 30840 27288
rect 30892 27276 30898 27328
rect 31202 27276 31208 27328
rect 31260 27316 31266 27328
rect 31481 27319 31539 27325
rect 31481 27316 31493 27319
rect 31260 27288 31493 27316
rect 31260 27276 31266 27288
rect 31481 27285 31493 27288
rect 31527 27285 31539 27319
rect 33134 27316 33140 27328
rect 33095 27288 33140 27316
rect 31481 27279 31539 27285
rect 33134 27276 33140 27288
rect 33192 27276 33198 27328
rect 33594 27276 33600 27328
rect 33652 27316 33658 27328
rect 33689 27319 33747 27325
rect 33689 27316 33701 27319
rect 33652 27288 33701 27316
rect 33652 27276 33658 27288
rect 33689 27285 33701 27288
rect 33735 27285 33747 27319
rect 33689 27279 33747 27285
rect 34790 27276 34796 27328
rect 34848 27316 34854 27328
rect 34977 27319 35035 27325
rect 34977 27316 34989 27319
rect 34848 27288 34989 27316
rect 34848 27276 34854 27288
rect 34977 27285 34989 27288
rect 35023 27285 35035 27319
rect 34977 27279 35035 27285
rect 1104 27226 38548 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 38548 27226
rect 1104 27152 38548 27174
rect 2038 27112 2044 27124
rect 1999 27084 2044 27112
rect 2038 27072 2044 27084
rect 2096 27072 2102 27124
rect 4525 27115 4583 27121
rect 4525 27081 4537 27115
rect 4571 27112 4583 27115
rect 4614 27112 4620 27124
rect 4571 27084 4620 27112
rect 4571 27081 4583 27084
rect 4525 27075 4583 27081
rect 4614 27072 4620 27084
rect 4672 27072 4678 27124
rect 5261 27115 5319 27121
rect 5261 27081 5273 27115
rect 5307 27112 5319 27115
rect 5810 27112 5816 27124
rect 5307 27084 5816 27112
rect 5307 27081 5319 27084
rect 5261 27075 5319 27081
rect 5810 27072 5816 27084
rect 5868 27072 5874 27124
rect 5997 27115 6055 27121
rect 5997 27081 6009 27115
rect 6043 27112 6055 27115
rect 6086 27112 6092 27124
rect 6043 27084 6092 27112
rect 6043 27081 6055 27084
rect 5997 27075 6055 27081
rect 6086 27072 6092 27084
rect 6144 27072 6150 27124
rect 7098 27112 7104 27124
rect 7059 27084 7104 27112
rect 7098 27072 7104 27084
rect 7156 27072 7162 27124
rect 11885 27115 11943 27121
rect 11885 27081 11897 27115
rect 11931 27112 11943 27115
rect 12066 27112 12072 27124
rect 11931 27084 12072 27112
rect 11931 27081 11943 27084
rect 11885 27075 11943 27081
rect 12066 27072 12072 27084
rect 12124 27072 12130 27124
rect 13354 27112 13360 27124
rect 13315 27084 13360 27112
rect 13354 27072 13360 27084
rect 13412 27072 13418 27124
rect 20993 27115 21051 27121
rect 20993 27081 21005 27115
rect 21039 27112 21051 27115
rect 21082 27112 21088 27124
rect 21039 27084 21088 27112
rect 21039 27081 21051 27084
rect 20993 27075 21051 27081
rect 21082 27072 21088 27084
rect 21140 27072 21146 27124
rect 22830 27112 22836 27124
rect 22791 27084 22836 27112
rect 22830 27072 22836 27084
rect 22888 27072 22894 27124
rect 23477 27115 23535 27121
rect 23477 27081 23489 27115
rect 23523 27112 23535 27115
rect 24762 27112 24768 27124
rect 23523 27084 24768 27112
rect 23523 27081 23535 27084
rect 23477 27075 23535 27081
rect 24762 27072 24768 27084
rect 24820 27072 24826 27124
rect 25961 27115 26019 27121
rect 25961 27081 25973 27115
rect 26007 27112 26019 27115
rect 26970 27112 26976 27124
rect 26007 27084 26976 27112
rect 26007 27081 26019 27084
rect 25961 27075 26019 27081
rect 26970 27072 26976 27084
rect 27028 27072 27034 27124
rect 27890 27112 27896 27124
rect 27851 27084 27896 27112
rect 27890 27072 27896 27084
rect 27948 27112 27954 27124
rect 28353 27115 28411 27121
rect 28353 27112 28365 27115
rect 27948 27084 28365 27112
rect 27948 27072 27954 27084
rect 28353 27081 28365 27084
rect 28399 27081 28411 27115
rect 28353 27075 28411 27081
rect 29546 27072 29552 27124
rect 29604 27112 29610 27124
rect 30193 27115 30251 27121
rect 30193 27112 30205 27115
rect 29604 27084 30205 27112
rect 29604 27072 29610 27084
rect 30193 27081 30205 27084
rect 30239 27081 30251 27115
rect 31846 27112 31852 27124
rect 31807 27084 31852 27112
rect 30193 27075 30251 27081
rect 31846 27072 31852 27084
rect 31904 27072 31910 27124
rect 32490 27072 32496 27124
rect 32548 27112 32554 27124
rect 33965 27115 34023 27121
rect 33965 27112 33977 27115
rect 32548 27084 33977 27112
rect 32548 27072 32554 27084
rect 33965 27081 33977 27084
rect 34011 27112 34023 27115
rect 34330 27112 34336 27124
rect 34011 27084 34336 27112
rect 34011 27081 34023 27084
rect 33965 27075 34023 27081
rect 34330 27072 34336 27084
rect 34388 27072 34394 27124
rect 36262 27112 36268 27124
rect 36223 27084 36268 27112
rect 36262 27072 36268 27084
rect 36320 27072 36326 27124
rect 5718 27004 5724 27056
rect 5776 27044 5782 27056
rect 6270 27044 6276 27056
rect 5776 27016 6276 27044
rect 5776 27004 5782 27016
rect 6270 27004 6276 27016
rect 6328 27004 6334 27056
rect 8110 27044 8116 27056
rect 8071 27016 8116 27044
rect 8110 27004 8116 27016
rect 8168 27004 8174 27056
rect 8573 27047 8631 27053
rect 8573 27013 8585 27047
rect 8619 27044 8631 27047
rect 10318 27044 10324 27056
rect 8619 27016 10324 27044
rect 8619 27013 8631 27016
rect 8573 27007 8631 27013
rect 10318 27004 10324 27016
rect 10376 27004 10382 27056
rect 12621 27047 12679 27053
rect 12621 27044 12633 27047
rect 11164 27016 12633 27044
rect 3418 26976 3424 26988
rect 3379 26948 3424 26976
rect 3418 26936 3424 26948
rect 3476 26936 3482 26988
rect 10336 26976 10364 27004
rect 10336 26948 10732 26976
rect 3237 26911 3295 26917
rect 3237 26877 3249 26911
rect 3283 26908 3295 26911
rect 3326 26908 3332 26920
rect 3283 26880 3332 26908
rect 3283 26877 3295 26880
rect 3237 26871 3295 26877
rect 3326 26868 3332 26880
rect 3384 26908 3390 26920
rect 3513 26911 3571 26917
rect 3513 26908 3525 26911
rect 3384 26880 3525 26908
rect 3384 26868 3390 26880
rect 3513 26877 3525 26880
rect 3559 26908 3571 26911
rect 3878 26908 3884 26920
rect 3559 26880 3884 26908
rect 3559 26877 3571 26880
rect 3513 26871 3571 26877
rect 3878 26868 3884 26880
rect 3936 26908 3942 26920
rect 4065 26911 4123 26917
rect 4065 26908 4077 26911
rect 3936 26880 4077 26908
rect 3936 26868 3942 26880
rect 4065 26877 4077 26880
rect 4111 26877 4123 26911
rect 4065 26871 4123 26877
rect 4249 26911 4307 26917
rect 4249 26877 4261 26911
rect 4295 26877 4307 26911
rect 4249 26871 4307 26877
rect 2869 26843 2927 26849
rect 2869 26809 2881 26843
rect 2915 26840 2927 26843
rect 4264 26840 4292 26871
rect 6454 26868 6460 26920
rect 6512 26908 6518 26920
rect 6825 26911 6883 26917
rect 6825 26908 6837 26911
rect 6512 26880 6837 26908
rect 6512 26868 6518 26880
rect 6825 26877 6837 26880
rect 6871 26877 6883 26911
rect 6825 26871 6883 26877
rect 6917 26911 6975 26917
rect 6917 26877 6929 26911
rect 6963 26877 6975 26911
rect 6917 26871 6975 26877
rect 8481 26911 8539 26917
rect 8481 26877 8493 26911
rect 8527 26877 8539 26911
rect 8846 26908 8852 26920
rect 8807 26880 8852 26908
rect 8481 26871 8539 26877
rect 4522 26840 4528 26852
rect 2915 26812 4528 26840
rect 2915 26809 2927 26812
rect 2869 26803 2927 26809
rect 4522 26800 4528 26812
rect 4580 26800 4586 26852
rect 5629 26843 5687 26849
rect 5629 26809 5641 26843
rect 5675 26840 5687 26843
rect 6638 26840 6644 26852
rect 5675 26812 6644 26840
rect 5675 26809 5687 26812
rect 5629 26803 5687 26809
rect 6638 26800 6644 26812
rect 6696 26800 6702 26852
rect 1486 26732 1492 26784
rect 1544 26772 1550 26784
rect 1581 26775 1639 26781
rect 1581 26772 1593 26775
rect 1544 26744 1593 26772
rect 1544 26732 1550 26744
rect 1581 26741 1593 26744
rect 1627 26741 1639 26775
rect 6932 26772 6960 26871
rect 8496 26840 8524 26871
rect 8846 26868 8852 26880
rect 8904 26868 8910 26920
rect 9122 26908 9128 26920
rect 9083 26880 9128 26908
rect 9122 26868 9128 26880
rect 9180 26868 9186 26920
rect 10704 26917 10732 26948
rect 10321 26911 10379 26917
rect 10321 26908 10333 26911
rect 10152 26880 10333 26908
rect 9674 26840 9680 26852
rect 8496 26812 9680 26840
rect 9674 26800 9680 26812
rect 9732 26800 9738 26852
rect 10152 26784 10180 26880
rect 10321 26877 10333 26880
rect 10367 26877 10379 26911
rect 10321 26871 10379 26877
rect 10689 26911 10747 26917
rect 10689 26877 10701 26911
rect 10735 26877 10747 26911
rect 10689 26871 10747 26877
rect 10778 26868 10784 26920
rect 10836 26908 10842 26920
rect 11164 26917 11192 27016
rect 12621 27013 12633 27016
rect 12667 27044 12679 27047
rect 15010 27044 15016 27056
rect 12667 27016 15016 27044
rect 12667 27013 12679 27016
rect 12621 27007 12679 27013
rect 15010 27004 15016 27016
rect 15068 27004 15074 27056
rect 15746 27004 15752 27056
rect 15804 27044 15810 27056
rect 18874 27044 18880 27056
rect 15804 27016 18880 27044
rect 15804 27004 15810 27016
rect 18874 27004 18880 27016
rect 18932 27004 18938 27056
rect 15470 26936 15476 26988
rect 15528 26976 15534 26988
rect 15528 26948 16160 26976
rect 15528 26936 15534 26948
rect 11149 26911 11207 26917
rect 11149 26908 11161 26911
rect 10836 26880 11161 26908
rect 10836 26868 10842 26880
rect 11149 26877 11161 26880
rect 11195 26877 11207 26911
rect 11149 26871 11207 26877
rect 12437 26911 12495 26917
rect 12437 26877 12449 26911
rect 12483 26908 12495 26911
rect 13998 26908 14004 26920
rect 12483 26880 12572 26908
rect 13911 26880 14004 26908
rect 12483 26877 12495 26880
rect 12437 26871 12495 26877
rect 11422 26840 11428 26852
rect 11383 26812 11428 26840
rect 11422 26800 11428 26812
rect 11480 26800 11486 26852
rect 12544 26784 12572 26880
rect 13998 26868 14004 26880
rect 14056 26908 14062 26920
rect 14458 26908 14464 26920
rect 14056 26880 14464 26908
rect 14056 26868 14062 26880
rect 14458 26868 14464 26880
rect 14516 26868 14522 26920
rect 15838 26908 15844 26920
rect 15751 26880 15844 26908
rect 15838 26868 15844 26880
rect 15896 26908 15902 26920
rect 16132 26917 16160 26948
rect 19334 26936 19340 26988
rect 19392 26976 19398 26988
rect 19392 26948 19748 26976
rect 19392 26936 19398 26948
rect 16025 26911 16083 26917
rect 16025 26908 16037 26911
rect 15896 26880 16037 26908
rect 15896 26868 15902 26880
rect 16025 26877 16037 26880
rect 16071 26877 16083 26911
rect 16025 26871 16083 26877
rect 16117 26911 16175 26917
rect 16117 26877 16129 26911
rect 16163 26908 16175 26911
rect 16853 26911 16911 26917
rect 16853 26908 16865 26911
rect 16163 26880 16865 26908
rect 16163 26877 16175 26880
rect 16117 26871 16175 26877
rect 16853 26877 16865 26880
rect 16899 26877 16911 26911
rect 16853 26871 16911 26877
rect 18509 26911 18567 26917
rect 18509 26877 18521 26911
rect 18555 26908 18567 26911
rect 19426 26908 19432 26920
rect 18555 26880 19432 26908
rect 18555 26877 18567 26880
rect 18509 26871 18567 26877
rect 19426 26868 19432 26880
rect 19484 26908 19490 26920
rect 19720 26917 19748 26948
rect 19521 26911 19579 26917
rect 19521 26908 19533 26911
rect 19484 26880 19533 26908
rect 19484 26868 19490 26880
rect 19521 26877 19533 26880
rect 19567 26877 19579 26911
rect 19521 26871 19579 26877
rect 19705 26911 19763 26917
rect 19705 26877 19717 26911
rect 19751 26877 19763 26911
rect 19886 26908 19892 26920
rect 19847 26880 19892 26908
rect 19705 26871 19763 26877
rect 19886 26868 19892 26880
rect 19944 26868 19950 26920
rect 21100 26908 21128 27072
rect 22002 27044 22008 27056
rect 21468 27016 22008 27044
rect 21468 26985 21496 27016
rect 22002 27004 22008 27016
rect 22060 27004 22066 27056
rect 28718 27044 28724 27056
rect 28679 27016 28724 27044
rect 28718 27004 28724 27016
rect 28776 27004 28782 27056
rect 30009 27047 30067 27053
rect 30009 27013 30021 27047
rect 30055 27044 30067 27047
rect 30466 27044 30472 27056
rect 30055 27016 30472 27044
rect 30055 27013 30067 27016
rect 30009 27007 30067 27013
rect 30466 27004 30472 27016
rect 30524 27044 30530 27056
rect 30524 27016 31248 27044
rect 30524 27004 30530 27016
rect 21453 26979 21511 26985
rect 21453 26945 21465 26979
rect 21499 26945 21511 26979
rect 21453 26939 21511 26945
rect 21726 26936 21732 26988
rect 21784 26976 21790 26988
rect 23750 26976 23756 26988
rect 21784 26948 22324 26976
rect 23711 26948 23756 26976
rect 21784 26936 21790 26948
rect 22005 26911 22063 26917
rect 22005 26908 22017 26911
rect 21100 26880 22017 26908
rect 22005 26877 22017 26880
rect 22051 26908 22063 26911
rect 22186 26908 22192 26920
rect 22051 26880 22192 26908
rect 22051 26877 22063 26880
rect 22005 26871 22063 26877
rect 22186 26868 22192 26880
rect 22244 26868 22250 26920
rect 22296 26917 22324 26948
rect 23750 26936 23756 26948
rect 23808 26936 23814 26988
rect 25041 26979 25099 26985
rect 25041 26976 25053 26979
rect 24596 26948 25053 26976
rect 22281 26911 22339 26917
rect 22281 26877 22293 26911
rect 22327 26877 22339 26911
rect 22462 26908 22468 26920
rect 22423 26880 22468 26908
rect 22281 26871 22339 26877
rect 22462 26868 22468 26880
rect 22520 26868 22526 26920
rect 24486 26868 24492 26920
rect 24544 26908 24550 26920
rect 24596 26917 24624 26948
rect 25041 26945 25053 26948
rect 25087 26976 25099 26979
rect 25222 26976 25228 26988
rect 25087 26948 25228 26976
rect 25087 26945 25099 26948
rect 25041 26939 25099 26945
rect 25222 26936 25228 26948
rect 25280 26936 25286 26988
rect 25406 26936 25412 26988
rect 25464 26976 25470 26988
rect 26329 26979 26387 26985
rect 26329 26976 26341 26979
rect 25464 26948 26341 26976
rect 25464 26936 25470 26948
rect 26329 26945 26341 26948
rect 26375 26945 26387 26979
rect 27614 26976 27620 26988
rect 26329 26939 26387 26945
rect 26712 26948 27620 26976
rect 24581 26911 24639 26917
rect 24581 26908 24593 26911
rect 24544 26880 24593 26908
rect 24544 26868 24550 26880
rect 24581 26877 24593 26880
rect 24627 26877 24639 26911
rect 24581 26871 24639 26877
rect 24673 26911 24731 26917
rect 24673 26877 24685 26911
rect 24719 26908 24731 26911
rect 24854 26908 24860 26920
rect 24719 26880 24860 26908
rect 24719 26877 24731 26880
rect 24673 26871 24731 26877
rect 24854 26868 24860 26880
rect 24912 26868 24918 26920
rect 25958 26868 25964 26920
rect 26016 26908 26022 26920
rect 26237 26911 26295 26917
rect 26237 26908 26249 26911
rect 26016 26880 26249 26908
rect 26016 26868 26022 26880
rect 26237 26877 26249 26880
rect 26283 26908 26295 26911
rect 26712 26908 26740 26948
rect 27614 26936 27620 26948
rect 27672 26936 27678 26988
rect 26283 26880 26740 26908
rect 26789 26911 26847 26917
rect 26283 26877 26295 26880
rect 26237 26871 26295 26877
rect 26789 26877 26801 26911
rect 26835 26908 26847 26911
rect 26878 26908 26884 26920
rect 26835 26880 26884 26908
rect 26835 26877 26847 26880
rect 26789 26871 26847 26877
rect 14829 26843 14887 26849
rect 14829 26809 14841 26843
rect 14875 26840 14887 26843
rect 15286 26840 15292 26852
rect 14875 26812 15292 26840
rect 14875 26809 14887 26812
rect 14829 26803 14887 26809
rect 15286 26800 15292 26812
rect 15344 26800 15350 26852
rect 7374 26772 7380 26784
rect 6932 26744 7380 26772
rect 1581 26735 1639 26741
rect 7374 26732 7380 26744
rect 7432 26772 7438 26784
rect 7653 26775 7711 26781
rect 7653 26772 7665 26775
rect 7432 26744 7665 26772
rect 7432 26732 7438 26744
rect 7653 26741 7665 26744
rect 7699 26741 7711 26775
rect 10134 26772 10140 26784
rect 10095 26744 10140 26772
rect 7653 26735 7711 26741
rect 10134 26732 10140 26744
rect 10192 26732 10198 26784
rect 11698 26732 11704 26784
rect 11756 26772 11762 26784
rect 12161 26775 12219 26781
rect 12161 26772 12173 26775
rect 11756 26744 12173 26772
rect 11756 26732 11762 26744
rect 12161 26741 12173 26744
rect 12207 26741 12219 26775
rect 12161 26735 12219 26741
rect 12526 26732 12532 26784
rect 12584 26772 12590 26784
rect 12897 26775 12955 26781
rect 12897 26772 12909 26775
rect 12584 26744 12909 26772
rect 12584 26732 12590 26744
rect 12897 26741 12909 26744
rect 12943 26772 12955 26775
rect 13538 26772 13544 26784
rect 12943 26744 13544 26772
rect 12943 26741 12955 26744
rect 12897 26735 12955 26741
rect 13538 26732 13544 26744
rect 13596 26732 13602 26784
rect 15562 26732 15568 26784
rect 15620 26772 15626 26784
rect 15856 26781 15884 26868
rect 16574 26840 16580 26852
rect 16535 26812 16580 26840
rect 16574 26800 16580 26812
rect 16632 26800 16638 26852
rect 17313 26843 17371 26849
rect 17313 26809 17325 26843
rect 17359 26840 17371 26843
rect 17494 26840 17500 26852
rect 17359 26812 17500 26840
rect 17359 26809 17371 26812
rect 17313 26803 17371 26809
rect 17494 26800 17500 26812
rect 17552 26840 17558 26852
rect 18322 26840 18328 26852
rect 17552 26812 18328 26840
rect 17552 26800 17558 26812
rect 18322 26800 18328 26812
rect 18380 26800 18386 26852
rect 19061 26843 19119 26849
rect 19061 26809 19073 26843
rect 19107 26840 19119 26843
rect 19242 26840 19248 26852
rect 19107 26812 19248 26840
rect 19107 26809 19119 26812
rect 19061 26803 19119 26809
rect 19242 26800 19248 26812
rect 19300 26800 19306 26852
rect 21082 26800 21088 26852
rect 21140 26840 21146 26852
rect 21361 26843 21419 26849
rect 21361 26840 21373 26843
rect 21140 26812 21373 26840
rect 21140 26800 21146 26812
rect 21361 26809 21373 26812
rect 21407 26840 21419 26843
rect 22480 26840 22508 26868
rect 23845 26843 23903 26849
rect 23845 26840 23857 26843
rect 21407 26812 22508 26840
rect 23768 26812 23857 26840
rect 21407 26809 21419 26812
rect 21361 26803 21419 26809
rect 23768 26784 23796 26812
rect 23845 26809 23857 26812
rect 23891 26809 23903 26843
rect 23845 26803 23903 26809
rect 25593 26843 25651 26849
rect 25593 26809 25605 26843
rect 25639 26840 25651 26843
rect 26804 26840 26832 26871
rect 26878 26868 26884 26880
rect 26936 26868 26942 26920
rect 26970 26868 26976 26920
rect 27028 26908 27034 26920
rect 27157 26911 27215 26917
rect 27028 26880 27073 26908
rect 27028 26868 27034 26880
rect 27157 26877 27169 26911
rect 27203 26877 27215 26911
rect 27157 26871 27215 26877
rect 28169 26911 28227 26917
rect 28169 26877 28181 26911
rect 28215 26908 28227 26911
rect 28736 26908 28764 27004
rect 30834 26976 30840 26988
rect 30795 26948 30840 26976
rect 30834 26936 30840 26948
rect 30892 26936 30898 26988
rect 31220 26985 31248 27016
rect 31205 26979 31263 26985
rect 31205 26945 31217 26979
rect 31251 26945 31263 26979
rect 31205 26939 31263 26945
rect 34701 26979 34759 26985
rect 34701 26945 34713 26979
rect 34747 26976 34759 26979
rect 34747 26948 35204 26976
rect 34747 26945 34759 26948
rect 34701 26939 34759 26945
rect 28215 26880 28764 26908
rect 29641 26911 29699 26917
rect 28215 26877 28227 26880
rect 28169 26871 28227 26877
rect 29641 26877 29653 26911
rect 29687 26908 29699 26911
rect 30742 26908 30748 26920
rect 29687 26880 30748 26908
rect 29687 26877 29699 26880
rect 29641 26871 29699 26877
rect 25639 26812 26832 26840
rect 25639 26809 25651 26812
rect 25593 26803 25651 26809
rect 15841 26775 15899 26781
rect 15841 26772 15853 26775
rect 15620 26744 15853 26772
rect 15620 26732 15626 26744
rect 15841 26741 15853 26744
rect 15887 26741 15899 26775
rect 15841 26735 15899 26741
rect 18046 26732 18052 26784
rect 18104 26772 18110 26784
rect 18690 26772 18696 26784
rect 18104 26744 18696 26772
rect 18104 26732 18110 26744
rect 18690 26732 18696 26744
rect 18748 26772 18754 26784
rect 18785 26775 18843 26781
rect 18785 26772 18797 26775
rect 18748 26744 18797 26772
rect 18748 26732 18754 26744
rect 18785 26741 18797 26744
rect 18831 26741 18843 26775
rect 18785 26735 18843 26741
rect 23750 26732 23756 26784
rect 23808 26732 23814 26784
rect 26053 26775 26111 26781
rect 26053 26741 26065 26775
rect 26099 26772 26111 26775
rect 26142 26772 26148 26784
rect 26099 26744 26148 26772
rect 26099 26741 26111 26744
rect 26053 26735 26111 26741
rect 26142 26732 26148 26744
rect 26200 26732 26206 26784
rect 26234 26732 26240 26784
rect 26292 26772 26298 26784
rect 27172 26772 27200 26871
rect 30742 26868 30748 26880
rect 30800 26868 30806 26920
rect 31110 26908 31116 26920
rect 30852 26880 31116 26908
rect 30852 26852 30880 26880
rect 31110 26868 31116 26880
rect 31168 26868 31174 26920
rect 32398 26908 32404 26920
rect 32359 26880 32404 26908
rect 32398 26868 32404 26880
rect 32456 26868 32462 26920
rect 32493 26911 32551 26917
rect 32493 26877 32505 26911
rect 32539 26908 32551 26911
rect 33781 26911 33839 26917
rect 33781 26908 33793 26911
rect 32539 26880 33793 26908
rect 32539 26877 32551 26880
rect 32493 26871 32551 26877
rect 33781 26877 33793 26880
rect 33827 26908 33839 26911
rect 34882 26908 34888 26920
rect 33827 26880 33861 26908
rect 34843 26880 34888 26908
rect 33827 26877 33839 26880
rect 33781 26871 33839 26877
rect 30834 26800 30840 26852
rect 30892 26800 30898 26852
rect 32950 26840 32956 26852
rect 32911 26812 32956 26840
rect 32950 26800 32956 26812
rect 33008 26800 33014 26852
rect 33597 26843 33655 26849
rect 33597 26809 33609 26843
rect 33643 26840 33655 26843
rect 33796 26840 33824 26871
rect 34882 26868 34888 26880
rect 34940 26868 34946 26920
rect 35176 26917 35204 26948
rect 35161 26911 35219 26917
rect 35161 26877 35173 26911
rect 35207 26908 35219 26911
rect 36170 26908 36176 26920
rect 35207 26880 36176 26908
rect 35207 26877 35219 26880
rect 35161 26871 35219 26877
rect 36170 26868 36176 26880
rect 36228 26868 36234 26920
rect 33643 26812 34376 26840
rect 33643 26809 33655 26812
rect 33597 26803 33655 26809
rect 26292 26744 27200 26772
rect 26292 26732 26298 26744
rect 27430 26732 27436 26784
rect 27488 26772 27494 26784
rect 32214 26772 32220 26784
rect 27488 26744 32220 26772
rect 27488 26732 27494 26744
rect 32214 26732 32220 26744
rect 32272 26732 32278 26784
rect 34348 26781 34376 26812
rect 34333 26775 34391 26781
rect 34333 26741 34345 26775
rect 34379 26772 34391 26775
rect 34514 26772 34520 26784
rect 34379 26744 34520 26772
rect 34379 26741 34391 26744
rect 34333 26735 34391 26741
rect 34514 26732 34520 26744
rect 34572 26732 34578 26784
rect 36909 26775 36967 26781
rect 36909 26741 36921 26775
rect 36955 26772 36967 26775
rect 37182 26772 37188 26784
rect 36955 26744 37188 26772
rect 36955 26741 36967 26744
rect 36909 26735 36967 26741
rect 37182 26732 37188 26744
rect 37240 26732 37246 26784
rect 1104 26682 38548 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 38548 26682
rect 1104 26608 38548 26630
rect 1394 26528 1400 26580
rect 1452 26568 1458 26580
rect 1673 26571 1731 26577
rect 1673 26568 1685 26571
rect 1452 26540 1685 26568
rect 1452 26528 1458 26540
rect 1673 26537 1685 26540
rect 1719 26568 1731 26571
rect 2038 26568 2044 26580
rect 1719 26540 2044 26568
rect 1719 26537 1731 26540
rect 1673 26531 1731 26537
rect 2038 26528 2044 26540
rect 2096 26528 2102 26580
rect 3326 26568 3332 26580
rect 3287 26540 3332 26568
rect 3326 26528 3332 26540
rect 3384 26528 3390 26580
rect 4522 26568 4528 26580
rect 4483 26540 4528 26568
rect 4522 26528 4528 26540
rect 4580 26528 4586 26580
rect 6181 26571 6239 26577
rect 6181 26537 6193 26571
rect 6227 26568 6239 26571
rect 7098 26568 7104 26580
rect 6227 26540 7104 26568
rect 6227 26537 6239 26540
rect 6181 26531 6239 26537
rect 7098 26528 7104 26540
rect 7156 26528 7162 26580
rect 8018 26568 8024 26580
rect 7979 26540 8024 26568
rect 8018 26528 8024 26540
rect 8076 26528 8082 26580
rect 14274 26568 14280 26580
rect 14235 26540 14280 26568
rect 14274 26528 14280 26540
rect 14332 26528 14338 26580
rect 16390 26568 16396 26580
rect 16351 26540 16396 26568
rect 16390 26528 16396 26540
rect 16448 26568 16454 26580
rect 16666 26568 16672 26580
rect 16448 26540 16672 26568
rect 16448 26528 16454 26540
rect 16666 26528 16672 26540
rect 16724 26568 16730 26580
rect 16853 26571 16911 26577
rect 16853 26568 16865 26571
rect 16724 26540 16865 26568
rect 16724 26528 16730 26540
rect 16853 26537 16865 26540
rect 16899 26568 16911 26571
rect 16899 26540 18000 26568
rect 16899 26537 16911 26540
rect 16853 26531 16911 26537
rect 4540 26500 4568 26528
rect 9674 26500 9680 26512
rect 4540 26472 5304 26500
rect 9635 26472 9680 26500
rect 4893 26435 4951 26441
rect 4893 26401 4905 26435
rect 4939 26432 4951 26435
rect 5074 26432 5080 26444
rect 4939 26404 5080 26432
rect 4939 26401 4951 26404
rect 4893 26395 4951 26401
rect 5074 26392 5080 26404
rect 5132 26392 5138 26444
rect 5276 26441 5304 26472
rect 9674 26460 9680 26472
rect 9732 26460 9738 26512
rect 16758 26460 16764 26512
rect 16816 26500 16822 26512
rect 16945 26503 17003 26509
rect 16945 26500 16957 26503
rect 16816 26472 16957 26500
rect 16816 26460 16822 26472
rect 16945 26469 16957 26472
rect 16991 26469 17003 26503
rect 16945 26463 17003 26469
rect 5261 26435 5319 26441
rect 5261 26401 5273 26435
rect 5307 26432 5319 26435
rect 6454 26432 6460 26444
rect 5307 26404 6460 26432
rect 5307 26401 5319 26404
rect 5261 26395 5319 26401
rect 6454 26392 6460 26404
rect 6512 26392 6518 26444
rect 6546 26392 6552 26444
rect 6604 26432 6610 26444
rect 6641 26435 6699 26441
rect 6641 26432 6653 26435
rect 6604 26404 6653 26432
rect 6604 26392 6610 26404
rect 6641 26401 6653 26404
rect 6687 26401 6699 26435
rect 6641 26395 6699 26401
rect 7009 26435 7067 26441
rect 7009 26401 7021 26435
rect 7055 26401 7067 26435
rect 7466 26432 7472 26444
rect 7427 26404 7472 26432
rect 7009 26395 7067 26401
rect 5537 26367 5595 26373
rect 5537 26333 5549 26367
rect 5583 26333 5595 26367
rect 5537 26327 5595 26333
rect 4982 26296 4988 26308
rect 4943 26268 4988 26296
rect 4982 26256 4988 26268
rect 5040 26256 5046 26308
rect 5258 26256 5264 26308
rect 5316 26296 5322 26308
rect 5552 26296 5580 26327
rect 5994 26324 6000 26376
rect 6052 26364 6058 26376
rect 7024 26364 7052 26395
rect 7466 26392 7472 26404
rect 7524 26432 7530 26444
rect 7650 26432 7656 26444
rect 7524 26404 7656 26432
rect 7524 26392 7530 26404
rect 7650 26392 7656 26404
rect 7708 26392 7714 26444
rect 10042 26392 10048 26444
rect 10100 26432 10106 26444
rect 10137 26435 10195 26441
rect 10137 26432 10149 26435
rect 10100 26404 10149 26432
rect 10100 26392 10106 26404
rect 10137 26401 10149 26404
rect 10183 26401 10195 26435
rect 10502 26432 10508 26444
rect 10463 26404 10508 26432
rect 10137 26395 10195 26401
rect 10502 26392 10508 26404
rect 10560 26392 10566 26444
rect 10594 26392 10600 26444
rect 10652 26432 10658 26444
rect 10652 26404 10697 26432
rect 10652 26392 10658 26404
rect 11422 26392 11428 26444
rect 11480 26432 11486 26444
rect 12066 26432 12072 26444
rect 11480 26404 12072 26432
rect 11480 26392 11486 26404
rect 12066 26392 12072 26404
rect 12124 26432 12130 26444
rect 12253 26435 12311 26441
rect 12253 26432 12265 26435
rect 12124 26404 12265 26432
rect 12124 26392 12130 26404
rect 12253 26401 12265 26404
rect 12299 26401 12311 26435
rect 12253 26395 12311 26401
rect 12434 26392 12440 26444
rect 12492 26432 12498 26444
rect 12710 26432 12716 26444
rect 12492 26404 12537 26432
rect 12671 26404 12716 26432
rect 12492 26392 12498 26404
rect 12710 26392 12716 26404
rect 12768 26392 12774 26444
rect 14090 26432 14096 26444
rect 14051 26404 14096 26432
rect 14090 26392 14096 26404
rect 14148 26392 14154 26444
rect 15286 26432 15292 26444
rect 15247 26404 15292 26432
rect 15286 26392 15292 26404
rect 15344 26392 15350 26444
rect 17589 26435 17647 26441
rect 17589 26401 17601 26435
rect 17635 26432 17647 26435
rect 17678 26432 17684 26444
rect 17635 26404 17684 26432
rect 17635 26401 17647 26404
rect 17589 26395 17647 26401
rect 17678 26392 17684 26404
rect 17736 26392 17742 26444
rect 17972 26441 18000 26540
rect 23842 26528 23848 26580
rect 23900 26568 23906 26580
rect 24029 26571 24087 26577
rect 24029 26568 24041 26571
rect 23900 26540 24041 26568
rect 23900 26528 23906 26540
rect 24029 26537 24041 26540
rect 24075 26568 24087 26571
rect 24397 26571 24455 26577
rect 24397 26568 24409 26571
rect 24075 26540 24409 26568
rect 24075 26537 24087 26540
rect 24029 26531 24087 26537
rect 24397 26537 24409 26540
rect 24443 26537 24455 26571
rect 25958 26568 25964 26580
rect 25919 26540 25964 26568
rect 24397 26531 24455 26537
rect 25958 26528 25964 26540
rect 26016 26528 26022 26580
rect 27982 26568 27988 26580
rect 27943 26540 27988 26568
rect 27982 26528 27988 26540
rect 28040 26528 28046 26580
rect 31018 26528 31024 26580
rect 31076 26568 31082 26580
rect 31941 26571 31999 26577
rect 31941 26568 31953 26571
rect 31076 26540 31953 26568
rect 31076 26528 31082 26540
rect 31941 26537 31953 26540
rect 31987 26568 31999 26571
rect 32398 26568 32404 26580
rect 31987 26540 32404 26568
rect 31987 26537 31999 26540
rect 31941 26531 31999 26537
rect 32398 26528 32404 26540
rect 32456 26528 32462 26580
rect 34698 26568 34704 26580
rect 34659 26540 34704 26568
rect 34698 26528 34704 26540
rect 34756 26528 34762 26580
rect 35618 26528 35624 26580
rect 35676 26568 35682 26580
rect 35713 26571 35771 26577
rect 35713 26568 35725 26571
rect 35676 26540 35725 26568
rect 35676 26528 35682 26540
rect 35713 26537 35725 26540
rect 35759 26537 35771 26571
rect 36078 26568 36084 26580
rect 36039 26540 36084 26568
rect 35713 26531 35771 26537
rect 36078 26528 36084 26540
rect 36136 26528 36142 26580
rect 19426 26460 19432 26512
rect 19484 26500 19490 26512
rect 19981 26503 20039 26509
rect 19981 26500 19993 26503
rect 19484 26472 19993 26500
rect 19484 26460 19490 26472
rect 19981 26469 19993 26472
rect 20027 26469 20039 26503
rect 19981 26463 20039 26469
rect 23753 26503 23811 26509
rect 23753 26469 23765 26503
rect 23799 26500 23811 26503
rect 24854 26500 24860 26512
rect 23799 26472 24860 26500
rect 23799 26469 23811 26472
rect 23753 26463 23811 26469
rect 24854 26460 24860 26472
rect 24912 26460 24918 26512
rect 26234 26500 26240 26512
rect 26195 26472 26240 26500
rect 26234 26460 26240 26472
rect 26292 26460 26298 26512
rect 26602 26460 26608 26512
rect 26660 26500 26666 26512
rect 27246 26500 27252 26512
rect 26660 26472 27252 26500
rect 26660 26460 26666 26472
rect 27246 26460 27252 26472
rect 27304 26500 27310 26512
rect 28261 26503 28319 26509
rect 28261 26500 28273 26503
rect 27304 26472 28273 26500
rect 27304 26460 27310 26472
rect 28261 26469 28273 26472
rect 28307 26500 28319 26503
rect 28810 26500 28816 26512
rect 28307 26472 28816 26500
rect 28307 26469 28319 26472
rect 28261 26463 28319 26469
rect 28810 26460 28816 26472
rect 28868 26460 28874 26512
rect 29086 26500 29092 26512
rect 29047 26472 29092 26500
rect 29086 26460 29092 26472
rect 29144 26460 29150 26512
rect 32861 26503 32919 26509
rect 32861 26469 32873 26503
rect 32907 26500 32919 26503
rect 32907 26472 33732 26500
rect 32907 26469 32919 26472
rect 32861 26463 32919 26469
rect 17957 26435 18015 26441
rect 17957 26401 17969 26435
rect 18003 26401 18015 26435
rect 17957 26395 18015 26401
rect 18141 26435 18199 26441
rect 18141 26401 18153 26435
rect 18187 26432 18199 26435
rect 19518 26432 19524 26444
rect 18187 26404 19380 26432
rect 19479 26404 19524 26432
rect 18187 26401 18199 26404
rect 18141 26395 18199 26401
rect 9122 26364 9128 26376
rect 6052 26336 7052 26364
rect 9083 26336 9128 26364
rect 6052 26324 6058 26336
rect 9122 26324 9128 26336
rect 9180 26324 9186 26376
rect 11790 26364 11796 26376
rect 11751 26336 11796 26364
rect 11790 26324 11796 26336
rect 11848 26324 11854 26376
rect 12986 26364 12992 26376
rect 12947 26336 12992 26364
rect 12986 26324 12992 26336
rect 13044 26324 13050 26376
rect 13170 26364 13176 26376
rect 13131 26336 13176 26364
rect 13170 26324 13176 26336
rect 13228 26324 13234 26376
rect 17402 26364 17408 26376
rect 17363 26336 17408 26364
rect 17402 26324 17408 26336
rect 17460 26324 17466 26376
rect 17494 26324 17500 26376
rect 17552 26364 17558 26376
rect 18156 26364 18184 26395
rect 17552 26336 18184 26364
rect 19352 26364 19380 26404
rect 19518 26392 19524 26404
rect 19576 26392 19582 26444
rect 21082 26432 21088 26444
rect 21043 26404 21088 26432
rect 21082 26392 21088 26404
rect 21140 26392 21146 26444
rect 21450 26432 21456 26444
rect 21411 26404 21456 26432
rect 21450 26392 21456 26404
rect 21508 26392 21514 26444
rect 21821 26435 21879 26441
rect 21821 26401 21833 26435
rect 21867 26432 21879 26435
rect 22002 26432 22008 26444
rect 21867 26404 22008 26432
rect 21867 26401 21879 26404
rect 21821 26395 21879 26401
rect 22002 26392 22008 26404
rect 22060 26392 22066 26444
rect 26786 26392 26792 26444
rect 26844 26432 26850 26444
rect 27433 26435 27491 26441
rect 27433 26432 27445 26435
rect 26844 26404 27445 26432
rect 26844 26392 26850 26404
rect 27433 26401 27445 26404
rect 27479 26401 27491 26435
rect 27433 26395 27491 26401
rect 27525 26435 27583 26441
rect 27525 26401 27537 26435
rect 27571 26432 27583 26435
rect 27890 26432 27896 26444
rect 27571 26404 27896 26432
rect 27571 26401 27583 26404
rect 27525 26395 27583 26401
rect 19429 26367 19487 26373
rect 19429 26364 19441 26367
rect 19352 26336 19441 26364
rect 17552 26324 17558 26336
rect 19429 26333 19441 26336
rect 19475 26364 19487 26367
rect 20346 26364 20352 26376
rect 19475 26336 20352 26364
rect 19475 26333 19487 26336
rect 19429 26327 19487 26333
rect 20346 26324 20352 26336
rect 20404 26324 20410 26376
rect 26234 26324 26240 26376
rect 26292 26364 26298 26376
rect 26605 26367 26663 26373
rect 26605 26364 26617 26367
rect 26292 26336 26617 26364
rect 26292 26324 26298 26336
rect 26605 26333 26617 26336
rect 26651 26333 26663 26367
rect 26605 26327 26663 26333
rect 26697 26367 26755 26373
rect 26697 26333 26709 26367
rect 26743 26333 26755 26367
rect 26697 26327 26755 26333
rect 5316 26268 5580 26296
rect 5316 26256 5322 26268
rect 6638 26256 6644 26308
rect 6696 26296 6702 26308
rect 7469 26299 7527 26305
rect 7469 26296 7481 26299
rect 6696 26268 7481 26296
rect 6696 26256 6702 26268
rect 7469 26265 7481 26268
rect 7515 26265 7527 26299
rect 8389 26299 8447 26305
rect 8389 26296 8401 26299
rect 7469 26259 7527 26265
rect 7944 26268 8401 26296
rect 7742 26188 7748 26240
rect 7800 26228 7806 26240
rect 7944 26228 7972 26268
rect 8389 26265 8401 26268
rect 8435 26265 8447 26299
rect 8389 26259 8447 26265
rect 8478 26256 8484 26308
rect 8536 26296 8542 26308
rect 8757 26299 8815 26305
rect 8757 26296 8769 26299
rect 8536 26268 8769 26296
rect 8536 26256 8542 26268
rect 8757 26265 8769 26268
rect 8803 26296 8815 26299
rect 8846 26296 8852 26308
rect 8803 26268 8852 26296
rect 8803 26265 8815 26268
rect 8757 26259 8815 26265
rect 8846 26256 8852 26268
rect 8904 26256 8910 26308
rect 11330 26296 11336 26308
rect 11291 26268 11336 26296
rect 11330 26256 11336 26268
rect 11388 26256 11394 26308
rect 13446 26256 13452 26308
rect 13504 26296 13510 26308
rect 13541 26299 13599 26305
rect 13541 26296 13553 26299
rect 13504 26268 13553 26296
rect 13504 26256 13510 26268
rect 13541 26265 13553 26268
rect 13587 26265 13599 26299
rect 13541 26259 13599 26265
rect 15102 26256 15108 26308
rect 15160 26296 15166 26308
rect 15473 26299 15531 26305
rect 15473 26296 15485 26299
rect 15160 26268 15485 26296
rect 15160 26256 15166 26268
rect 15473 26265 15485 26268
rect 15519 26265 15531 26299
rect 15473 26259 15531 26265
rect 19153 26299 19211 26305
rect 19153 26265 19165 26299
rect 19199 26296 19211 26299
rect 19886 26296 19892 26308
rect 19199 26268 19892 26296
rect 19199 26265 19211 26268
rect 19153 26259 19211 26265
rect 19886 26256 19892 26268
rect 19944 26256 19950 26308
rect 21174 26256 21180 26308
rect 21232 26296 21238 26308
rect 21729 26299 21787 26305
rect 21729 26296 21741 26299
rect 21232 26268 21741 26296
rect 21232 26256 21238 26268
rect 21729 26265 21741 26268
rect 21775 26265 21787 26299
rect 26712 26296 26740 26327
rect 26878 26324 26884 26376
rect 26936 26364 26942 26376
rect 27540 26364 27568 26395
rect 27890 26392 27896 26404
rect 27948 26392 27954 26444
rect 29546 26392 29552 26444
rect 29604 26432 29610 26444
rect 29733 26435 29791 26441
rect 29733 26432 29745 26435
rect 29604 26404 29745 26432
rect 29604 26392 29610 26404
rect 29733 26401 29745 26404
rect 29779 26401 29791 26435
rect 29733 26395 29791 26401
rect 29822 26392 29828 26444
rect 29880 26432 29886 26444
rect 29880 26404 29925 26432
rect 29880 26392 29886 26404
rect 30006 26392 30012 26444
rect 30064 26432 30070 26444
rect 30101 26435 30159 26441
rect 30101 26432 30113 26435
rect 30064 26404 30113 26432
rect 30064 26392 30070 26404
rect 30101 26401 30113 26404
rect 30147 26401 30159 26435
rect 30101 26395 30159 26401
rect 30285 26435 30343 26441
rect 30285 26401 30297 26435
rect 30331 26432 30343 26435
rect 30466 26432 30472 26444
rect 30331 26404 30472 26432
rect 30331 26401 30343 26404
rect 30285 26395 30343 26401
rect 30466 26392 30472 26404
rect 30524 26392 30530 26444
rect 31202 26392 31208 26444
rect 31260 26432 31266 26444
rect 33704 26441 33732 26472
rect 31297 26435 31355 26441
rect 31297 26432 31309 26435
rect 31260 26404 31309 26432
rect 31260 26392 31266 26404
rect 31297 26401 31309 26404
rect 31343 26401 31355 26435
rect 31297 26395 31355 26401
rect 33045 26435 33103 26441
rect 33045 26401 33057 26435
rect 33091 26401 33103 26435
rect 33045 26395 33103 26401
rect 33689 26435 33747 26441
rect 33689 26401 33701 26435
rect 33735 26432 33747 26435
rect 34514 26432 34520 26444
rect 33735 26404 34520 26432
rect 33735 26401 33747 26404
rect 33689 26395 33747 26401
rect 26936 26336 27568 26364
rect 26936 26324 26942 26336
rect 28997 26299 29055 26305
rect 26712 26268 28028 26296
rect 21729 26259 21787 26265
rect 28000 26240 28028 26268
rect 28997 26265 29009 26299
rect 29043 26296 29055 26299
rect 29086 26296 29092 26308
rect 29043 26268 29092 26296
rect 29043 26265 29055 26268
rect 28997 26259 29055 26265
rect 29086 26256 29092 26268
rect 29144 26256 29150 26308
rect 32493 26299 32551 26305
rect 32493 26265 32505 26299
rect 32539 26296 32551 26299
rect 33060 26296 33088 26395
rect 34514 26392 34520 26404
rect 34572 26432 34578 26444
rect 34977 26435 35035 26441
rect 34977 26432 34989 26435
rect 34572 26404 34989 26432
rect 34572 26392 34578 26404
rect 34977 26401 34989 26404
rect 35023 26401 35035 26435
rect 34977 26395 35035 26401
rect 33502 26296 33508 26308
rect 32539 26268 33508 26296
rect 32539 26265 32551 26268
rect 32493 26259 32551 26265
rect 33502 26256 33508 26268
rect 33560 26256 33566 26308
rect 10962 26228 10968 26240
rect 7800 26200 7972 26228
rect 10923 26200 10968 26228
rect 7800 26188 7806 26200
rect 10962 26188 10968 26200
rect 11020 26188 11026 26240
rect 11606 26188 11612 26240
rect 11664 26228 11670 26240
rect 15746 26228 15752 26240
rect 11664 26200 15752 26228
rect 11664 26188 11670 26200
rect 15746 26188 15752 26200
rect 15804 26188 15810 26240
rect 18322 26188 18328 26240
rect 18380 26228 18386 26240
rect 18417 26231 18475 26237
rect 18417 26228 18429 26231
rect 18380 26200 18429 26228
rect 18380 26188 18386 26200
rect 18417 26197 18429 26200
rect 18463 26197 18475 26231
rect 18417 26191 18475 26197
rect 22373 26231 22431 26237
rect 22373 26197 22385 26231
rect 22419 26228 22431 26231
rect 22830 26228 22836 26240
rect 22419 26200 22836 26228
rect 22419 26197 22431 26200
rect 22373 26191 22431 26197
rect 22830 26188 22836 26200
rect 22888 26188 22894 26240
rect 27982 26188 27988 26240
rect 28040 26188 28046 26240
rect 30653 26231 30711 26237
rect 30653 26197 30665 26231
rect 30699 26228 30711 26231
rect 30834 26228 30840 26240
rect 30699 26200 30840 26228
rect 30699 26197 30711 26200
rect 30653 26191 30711 26197
rect 30834 26188 30840 26200
rect 30892 26228 30898 26240
rect 30929 26231 30987 26237
rect 30929 26228 30941 26231
rect 30892 26200 30941 26228
rect 30892 26188 30898 26200
rect 30929 26197 30941 26200
rect 30975 26197 30987 26231
rect 30929 26191 30987 26197
rect 31113 26231 31171 26237
rect 31113 26197 31125 26231
rect 31159 26228 31171 26231
rect 35802 26228 35808 26240
rect 31159 26200 35808 26228
rect 31159 26197 31171 26200
rect 31113 26191 31171 26197
rect 35802 26188 35808 26200
rect 35860 26188 35866 26240
rect 1104 26138 38548 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 38548 26138
rect 1104 26064 38548 26086
rect 2774 25984 2780 26036
rect 2832 26024 2838 26036
rect 4985 26027 5043 26033
rect 2832 25996 2877 26024
rect 2832 25984 2838 25996
rect 4985 25993 4997 26027
rect 5031 26024 5043 26027
rect 5074 26024 5080 26036
rect 5031 25996 5080 26024
rect 5031 25993 5043 25996
rect 4985 25987 5043 25993
rect 5074 25984 5080 25996
rect 5132 25984 5138 26036
rect 8938 26024 8944 26036
rect 8899 25996 8944 26024
rect 8938 25984 8944 25996
rect 8996 25984 9002 26036
rect 11790 26024 11796 26036
rect 11751 25996 11796 26024
rect 11790 25984 11796 25996
rect 11848 25984 11854 26036
rect 13814 26024 13820 26036
rect 13727 25996 13820 26024
rect 13814 25984 13820 25996
rect 13872 26024 13878 26036
rect 14642 26024 14648 26036
rect 13872 25996 14648 26024
rect 13872 25984 13878 25996
rect 14642 25984 14648 25996
rect 14700 25984 14706 26036
rect 15286 26024 15292 26036
rect 15247 25996 15292 26024
rect 15286 25984 15292 25996
rect 15344 25984 15350 26036
rect 15930 25984 15936 26036
rect 15988 26024 15994 26036
rect 16390 26024 16396 26036
rect 15988 25996 16396 26024
rect 15988 25984 15994 25996
rect 16390 25984 16396 25996
rect 16448 25984 16454 26036
rect 17037 26027 17095 26033
rect 17037 25993 17049 26027
rect 17083 26024 17095 26027
rect 17494 26024 17500 26036
rect 17083 25996 17500 26024
rect 17083 25993 17095 25996
rect 17037 25987 17095 25993
rect 17494 25984 17500 25996
rect 17552 25984 17558 26036
rect 17678 26024 17684 26036
rect 17639 25996 17684 26024
rect 17678 25984 17684 25996
rect 17736 25984 17742 26036
rect 19518 25984 19524 26036
rect 19576 26024 19582 26036
rect 19613 26027 19671 26033
rect 19613 26024 19625 26027
rect 19576 25996 19625 26024
rect 19576 25984 19582 25996
rect 19613 25993 19625 25996
rect 19659 25993 19671 26027
rect 19613 25987 19671 25993
rect 20993 26027 21051 26033
rect 20993 25993 21005 26027
rect 21039 26024 21051 26027
rect 21082 26024 21088 26036
rect 21039 25996 21088 26024
rect 21039 25993 21051 25996
rect 20993 25987 21051 25993
rect 21082 25984 21088 25996
rect 21140 25984 21146 26036
rect 21361 26027 21419 26033
rect 21361 25993 21373 26027
rect 21407 26024 21419 26027
rect 21450 26024 21456 26036
rect 21407 25996 21456 26024
rect 21407 25993 21419 25996
rect 21361 25987 21419 25993
rect 21450 25984 21456 25996
rect 21508 25984 21514 26036
rect 21729 26027 21787 26033
rect 21729 25993 21741 26027
rect 21775 26024 21787 26027
rect 22002 26024 22008 26036
rect 21775 25996 22008 26024
rect 21775 25993 21787 25996
rect 21729 25987 21787 25993
rect 22002 25984 22008 25996
rect 22060 25984 22066 26036
rect 22462 26024 22468 26036
rect 22423 25996 22468 26024
rect 22462 25984 22468 25996
rect 22520 25984 22526 26036
rect 25314 25984 25320 26036
rect 25372 26024 25378 26036
rect 26053 26027 26111 26033
rect 26053 26024 26065 26027
rect 25372 25996 26065 26024
rect 25372 25984 25378 25996
rect 26053 25993 26065 25996
rect 26099 26024 26111 26027
rect 26142 26024 26148 26036
rect 26099 25996 26148 26024
rect 26099 25993 26111 25996
rect 26053 25987 26111 25993
rect 26142 25984 26148 25996
rect 26200 25984 26206 26036
rect 26513 26027 26571 26033
rect 26513 25993 26525 26027
rect 26559 26024 26571 26027
rect 26878 26024 26884 26036
rect 26559 25996 26884 26024
rect 26559 25993 26571 25996
rect 26513 25987 26571 25993
rect 26878 25984 26884 25996
rect 26936 25984 26942 26036
rect 27798 26024 27804 26036
rect 27759 25996 27804 26024
rect 27798 25984 27804 25996
rect 27856 25984 27862 26036
rect 29546 26024 29552 26036
rect 29507 25996 29552 26024
rect 29546 25984 29552 25996
rect 29604 25984 29610 26036
rect 29822 25984 29828 26036
rect 29880 26024 29886 26036
rect 30101 26027 30159 26033
rect 30101 26024 30113 26027
rect 29880 25996 30113 26024
rect 29880 25984 29886 25996
rect 30101 25993 30113 25996
rect 30147 25993 30159 26027
rect 30101 25987 30159 25993
rect 30742 25984 30748 26036
rect 30800 26024 30806 26036
rect 30929 26027 30987 26033
rect 30929 26024 30941 26027
rect 30800 25996 30941 26024
rect 30800 25984 30806 25996
rect 30929 25993 30941 25996
rect 30975 25993 30987 26027
rect 34514 26024 34520 26036
rect 34475 25996 34520 26024
rect 30929 25987 30987 25993
rect 34514 25984 34520 25996
rect 34572 25984 34578 26036
rect 37274 25984 37280 26036
rect 37332 26024 37338 26036
rect 37369 26027 37427 26033
rect 37369 26024 37381 26027
rect 37332 25996 37381 26024
rect 37332 25984 37338 25996
rect 37369 25993 37381 25996
rect 37415 25993 37427 26027
rect 37369 25987 37427 25993
rect 10413 25959 10471 25965
rect 10413 25925 10425 25959
rect 10459 25956 10471 25959
rect 12434 25956 12440 25968
rect 10459 25928 12440 25956
rect 10459 25925 10471 25928
rect 10413 25919 10471 25925
rect 12434 25916 12440 25928
rect 12492 25956 12498 25968
rect 12621 25959 12679 25965
rect 12621 25956 12633 25959
rect 12492 25928 12633 25956
rect 12492 25916 12498 25928
rect 12621 25925 12633 25928
rect 12667 25925 12679 25959
rect 12621 25919 12679 25925
rect 12710 25916 12716 25968
rect 12768 25916 12774 25968
rect 17402 25956 17408 25968
rect 17363 25928 17408 25956
rect 17402 25916 17408 25928
rect 17460 25916 17466 25968
rect 26789 25959 26847 25965
rect 26789 25925 26801 25959
rect 26835 25956 26847 25959
rect 27154 25956 27160 25968
rect 26835 25928 27160 25956
rect 26835 25925 26847 25928
rect 26789 25919 26847 25925
rect 27154 25916 27160 25928
rect 27212 25916 27218 25968
rect 29089 25959 29147 25965
rect 29089 25925 29101 25959
rect 29135 25956 29147 25959
rect 29178 25956 29184 25968
rect 29135 25928 29184 25956
rect 29135 25925 29147 25928
rect 29089 25919 29147 25925
rect 29178 25916 29184 25928
rect 29236 25956 29242 25968
rect 30006 25956 30012 25968
rect 29236 25928 30012 25956
rect 29236 25916 29242 25928
rect 30006 25916 30012 25928
rect 30064 25956 30070 25968
rect 32306 25956 32312 25968
rect 30064 25928 32312 25956
rect 30064 25916 30070 25928
rect 32306 25916 32312 25928
rect 32364 25916 32370 25968
rect 1394 25888 1400 25900
rect 1355 25860 1400 25888
rect 1394 25848 1400 25860
rect 1452 25848 1458 25900
rect 4614 25888 4620 25900
rect 4575 25860 4620 25888
rect 4614 25848 4620 25860
rect 4672 25848 4678 25900
rect 6825 25891 6883 25897
rect 6825 25857 6837 25891
rect 6871 25888 6883 25891
rect 7006 25888 7012 25900
rect 6871 25860 7012 25888
rect 6871 25857 6883 25860
rect 6825 25851 6883 25857
rect 7006 25848 7012 25860
rect 7064 25848 7070 25900
rect 7098 25848 7104 25900
rect 7156 25888 7162 25900
rect 7837 25891 7895 25897
rect 7837 25888 7849 25891
rect 7156 25860 7849 25888
rect 7156 25848 7162 25860
rect 7837 25857 7849 25860
rect 7883 25857 7895 25891
rect 7837 25851 7895 25857
rect 8202 25848 8208 25900
rect 8260 25888 8266 25900
rect 8665 25891 8723 25897
rect 8665 25888 8677 25891
rect 8260 25860 8677 25888
rect 8260 25848 8266 25860
rect 8665 25857 8677 25860
rect 8711 25888 8723 25891
rect 9122 25888 9128 25900
rect 8711 25860 9128 25888
rect 8711 25857 8723 25860
rect 8665 25851 8723 25857
rect 9122 25848 9128 25860
rect 9180 25848 9186 25900
rect 10226 25888 10232 25900
rect 10139 25860 10232 25888
rect 10226 25848 10232 25860
rect 10284 25888 10290 25900
rect 10870 25888 10876 25900
rect 10284 25860 10876 25888
rect 10284 25848 10290 25860
rect 10870 25848 10876 25860
rect 10928 25848 10934 25900
rect 11256 25860 11560 25888
rect 1670 25820 1676 25832
rect 1631 25792 1676 25820
rect 1670 25780 1676 25792
rect 1728 25780 1734 25832
rect 3789 25823 3847 25829
rect 3789 25789 3801 25823
rect 3835 25820 3847 25823
rect 4522 25820 4528 25832
rect 3835 25792 4528 25820
rect 3835 25789 3847 25792
rect 3789 25783 3847 25789
rect 4522 25780 4528 25792
rect 4580 25780 4586 25832
rect 5905 25823 5963 25829
rect 5905 25789 5917 25823
rect 5951 25820 5963 25823
rect 7377 25823 7435 25829
rect 7377 25820 7389 25823
rect 5951 25792 7389 25820
rect 5951 25789 5963 25792
rect 5905 25783 5963 25789
rect 7377 25789 7389 25792
rect 7423 25820 7435 25823
rect 7466 25820 7472 25832
rect 7423 25792 7472 25820
rect 7423 25789 7435 25792
rect 7377 25783 7435 25789
rect 5258 25684 5264 25696
rect 5219 25656 5264 25684
rect 5258 25644 5264 25656
rect 5316 25644 5322 25696
rect 5994 25644 6000 25696
rect 6052 25684 6058 25696
rect 6181 25687 6239 25693
rect 6181 25684 6193 25687
rect 6052 25656 6193 25684
rect 6052 25644 6058 25656
rect 6181 25653 6193 25656
rect 6227 25653 6239 25687
rect 6546 25684 6552 25696
rect 6507 25656 6552 25684
rect 6181 25647 6239 25653
rect 6546 25644 6552 25656
rect 6604 25644 6610 25696
rect 7392 25684 7420 25783
rect 7466 25780 7472 25792
rect 7524 25780 7530 25832
rect 7653 25823 7711 25829
rect 7653 25789 7665 25823
rect 7699 25820 7711 25823
rect 7742 25820 7748 25832
rect 7699 25792 7748 25820
rect 7699 25789 7711 25792
rect 7653 25783 7711 25789
rect 7742 25780 7748 25792
rect 7800 25780 7806 25832
rect 8757 25823 8815 25829
rect 8757 25789 8769 25823
rect 8803 25789 8815 25823
rect 10962 25820 10968 25832
rect 10923 25792 10968 25820
rect 8757 25783 8815 25789
rect 8202 25684 8208 25696
rect 7392 25656 8208 25684
rect 8202 25644 8208 25656
rect 8260 25644 8266 25696
rect 8573 25687 8631 25693
rect 8573 25653 8585 25687
rect 8619 25684 8631 25687
rect 8772 25684 8800 25783
rect 10962 25780 10968 25792
rect 11020 25780 11026 25832
rect 11054 25780 11060 25832
rect 11112 25820 11118 25832
rect 11256 25820 11284 25860
rect 11532 25829 11560 25860
rect 11112 25792 11284 25820
rect 11333 25823 11391 25829
rect 11112 25780 11118 25792
rect 11333 25789 11345 25823
rect 11379 25789 11391 25823
rect 11333 25783 11391 25789
rect 11517 25823 11575 25829
rect 11517 25789 11529 25823
rect 11563 25820 11575 25823
rect 12158 25820 12164 25832
rect 11563 25792 12164 25820
rect 11563 25789 11575 25792
rect 11517 25783 11575 25789
rect 11348 25752 11376 25783
rect 12158 25780 12164 25792
rect 12216 25780 12222 25832
rect 12253 25823 12311 25829
rect 12253 25789 12265 25823
rect 12299 25820 12311 25823
rect 12728 25820 12756 25916
rect 14090 25848 14096 25900
rect 14148 25888 14154 25900
rect 14185 25891 14243 25897
rect 14185 25888 14197 25891
rect 14148 25860 14197 25888
rect 14148 25848 14154 25860
rect 14185 25857 14197 25860
rect 14231 25888 14243 25891
rect 15102 25888 15108 25900
rect 14231 25860 15108 25888
rect 14231 25857 14243 25860
rect 14185 25851 14243 25857
rect 15102 25848 15108 25860
rect 15160 25848 15166 25900
rect 15746 25848 15752 25900
rect 15804 25888 15810 25900
rect 16393 25891 16451 25897
rect 16393 25888 16405 25891
rect 15804 25860 16405 25888
rect 15804 25848 15810 25860
rect 16393 25857 16405 25860
rect 16439 25857 16451 25891
rect 18506 25888 18512 25900
rect 18467 25860 18512 25888
rect 16393 25851 16451 25857
rect 18506 25848 18512 25860
rect 18564 25848 18570 25900
rect 23477 25891 23535 25897
rect 23477 25857 23489 25891
rect 23523 25888 23535 25891
rect 23523 25860 23980 25888
rect 23523 25857 23535 25860
rect 23477 25851 23535 25857
rect 23952 25832 23980 25860
rect 29638 25848 29644 25900
rect 29696 25888 29702 25900
rect 30190 25888 30196 25900
rect 29696 25860 30196 25888
rect 29696 25848 29702 25860
rect 30190 25848 30196 25860
rect 30248 25888 30254 25900
rect 30653 25891 30711 25897
rect 30653 25888 30665 25891
rect 30248 25860 30665 25888
rect 30248 25848 30254 25860
rect 30653 25857 30665 25860
rect 30699 25888 30711 25891
rect 31846 25888 31852 25900
rect 30699 25860 31852 25888
rect 30699 25857 30711 25860
rect 30653 25851 30711 25857
rect 31846 25848 31852 25860
rect 31904 25848 31910 25900
rect 35713 25891 35771 25897
rect 35713 25857 35725 25891
rect 35759 25888 35771 25891
rect 35759 25860 36124 25888
rect 35759 25857 35771 25860
rect 35713 25851 35771 25857
rect 36096 25832 36124 25860
rect 13538 25820 13544 25832
rect 12299 25792 13544 25820
rect 12299 25789 12311 25792
rect 12253 25783 12311 25789
rect 13538 25780 13544 25792
rect 13596 25780 13602 25832
rect 14366 25820 14372 25832
rect 14327 25792 14372 25820
rect 14366 25780 14372 25792
rect 14424 25820 14430 25832
rect 14829 25823 14887 25829
rect 14829 25820 14841 25823
rect 14424 25792 14841 25820
rect 14424 25780 14430 25792
rect 14829 25789 14841 25792
rect 14875 25820 14887 25823
rect 15194 25820 15200 25832
rect 14875 25792 15200 25820
rect 14875 25789 14887 25792
rect 14829 25783 14887 25789
rect 15194 25780 15200 25792
rect 15252 25820 15258 25832
rect 15252 25792 15884 25820
rect 15252 25780 15258 25792
rect 11606 25752 11612 25764
rect 11348 25724 11612 25752
rect 11606 25712 11612 25724
rect 11664 25712 11670 25764
rect 12989 25755 13047 25761
rect 12989 25721 13001 25755
rect 13035 25752 13047 25755
rect 13170 25752 13176 25764
rect 13035 25724 13176 25752
rect 13035 25721 13047 25724
rect 12989 25715 13047 25721
rect 13170 25712 13176 25724
rect 13228 25752 13234 25764
rect 15378 25752 15384 25764
rect 13228 25724 14320 25752
rect 15339 25724 15384 25752
rect 13228 25712 13234 25724
rect 14292 25696 14320 25724
rect 15378 25712 15384 25724
rect 15436 25712 15442 25764
rect 15856 25752 15884 25792
rect 15930 25780 15936 25832
rect 15988 25820 15994 25832
rect 16209 25823 16267 25829
rect 15988 25792 16033 25820
rect 15988 25780 15994 25792
rect 16209 25789 16221 25823
rect 16255 25789 16267 25823
rect 18230 25820 18236 25832
rect 18191 25792 18236 25820
rect 16209 25783 16267 25789
rect 16224 25752 16252 25783
rect 18230 25780 18236 25792
rect 18288 25780 18294 25832
rect 22649 25823 22707 25829
rect 22649 25789 22661 25823
rect 22695 25820 22707 25823
rect 22830 25820 22836 25832
rect 22695 25792 22836 25820
rect 22695 25789 22707 25792
rect 22649 25783 22707 25789
rect 22830 25780 22836 25792
rect 22888 25780 22894 25832
rect 23658 25820 23664 25832
rect 23619 25792 23664 25820
rect 23658 25780 23664 25792
rect 23716 25780 23722 25832
rect 23934 25820 23940 25832
rect 23895 25792 23940 25820
rect 23934 25780 23940 25792
rect 23992 25780 23998 25832
rect 26605 25823 26663 25829
rect 26605 25789 26617 25823
rect 26651 25820 26663 25823
rect 26878 25820 26884 25832
rect 26651 25792 26884 25820
rect 26651 25789 26663 25792
rect 26605 25783 26663 25789
rect 26878 25780 26884 25792
rect 26936 25820 26942 25832
rect 27065 25823 27123 25829
rect 27065 25820 27077 25823
rect 26936 25792 27077 25820
rect 26936 25780 26942 25792
rect 27065 25789 27077 25792
rect 27111 25789 27123 25823
rect 27065 25783 27123 25789
rect 27617 25823 27675 25829
rect 27617 25789 27629 25823
rect 27663 25820 27675 25823
rect 27663 25792 28212 25820
rect 27663 25789 27675 25792
rect 27617 25783 27675 25789
rect 15856 25724 16252 25752
rect 8846 25684 8852 25696
rect 8619 25656 8852 25684
rect 8619 25653 8631 25656
rect 8573 25647 8631 25653
rect 8846 25644 8852 25656
rect 8904 25644 8910 25696
rect 9769 25687 9827 25693
rect 9769 25653 9781 25687
rect 9815 25684 9827 25687
rect 10042 25684 10048 25696
rect 9815 25656 10048 25684
rect 9815 25653 9827 25656
rect 9769 25647 9827 25653
rect 10042 25644 10048 25656
rect 10100 25684 10106 25696
rect 10778 25684 10784 25696
rect 10100 25656 10784 25684
rect 10100 25644 10106 25656
rect 10778 25644 10784 25656
rect 10836 25644 10842 25696
rect 13078 25644 13084 25696
rect 13136 25684 13142 25696
rect 13357 25687 13415 25693
rect 13357 25684 13369 25687
rect 13136 25656 13369 25684
rect 13136 25644 13142 25656
rect 13357 25653 13369 25656
rect 13403 25653 13415 25687
rect 13357 25647 13415 25653
rect 14274 25644 14280 25696
rect 14332 25684 14338 25696
rect 14553 25687 14611 25693
rect 14553 25684 14565 25687
rect 14332 25656 14565 25684
rect 14332 25644 14338 25656
rect 14553 25653 14565 25656
rect 14599 25653 14611 25687
rect 14553 25647 14611 25653
rect 20257 25687 20315 25693
rect 20257 25653 20269 25687
rect 20303 25684 20315 25687
rect 20346 25684 20352 25696
rect 20303 25656 20352 25684
rect 20303 25653 20315 25656
rect 20257 25647 20315 25653
rect 20346 25644 20352 25656
rect 20404 25644 20410 25696
rect 25038 25684 25044 25696
rect 24999 25656 25044 25684
rect 25038 25644 25044 25656
rect 25096 25644 25102 25696
rect 28184 25693 28212 25792
rect 29086 25780 29092 25832
rect 29144 25820 29150 25832
rect 29273 25823 29331 25829
rect 29273 25820 29285 25823
rect 29144 25792 29285 25820
rect 29144 25780 29150 25792
rect 29273 25789 29285 25792
rect 29319 25789 29331 25823
rect 29273 25783 29331 25789
rect 29362 25780 29368 25832
rect 29420 25820 29426 25832
rect 30745 25823 30803 25829
rect 29420 25792 30236 25820
rect 29420 25780 29426 25792
rect 30208 25764 30236 25792
rect 30745 25789 30757 25823
rect 30791 25820 30803 25823
rect 31481 25823 31539 25829
rect 31481 25820 31493 25823
rect 30791 25792 31493 25820
rect 30791 25789 30803 25792
rect 30745 25783 30803 25789
rect 31481 25789 31493 25792
rect 31527 25789 31539 25823
rect 31481 25783 31539 25789
rect 31941 25823 31999 25829
rect 31941 25789 31953 25823
rect 31987 25820 31999 25823
rect 32861 25823 32919 25829
rect 32861 25820 32873 25823
rect 31987 25792 32873 25820
rect 31987 25789 31999 25792
rect 31941 25783 31999 25789
rect 32861 25789 32873 25792
rect 32907 25820 32919 25823
rect 32950 25820 32956 25832
rect 32907 25792 32956 25820
rect 32907 25789 32919 25792
rect 32861 25783 32919 25789
rect 30190 25712 30196 25764
rect 30248 25752 30254 25764
rect 30561 25755 30619 25761
rect 30561 25752 30573 25755
rect 30248 25724 30573 25752
rect 30248 25712 30254 25724
rect 30561 25721 30573 25724
rect 30607 25752 30619 25755
rect 30760 25752 30788 25783
rect 32950 25780 32956 25792
rect 33008 25780 33014 25832
rect 33229 25823 33287 25829
rect 33229 25789 33241 25823
rect 33275 25789 33287 25823
rect 33229 25783 33287 25789
rect 33321 25823 33379 25829
rect 33321 25789 33333 25823
rect 33367 25820 33379 25823
rect 33502 25820 33508 25832
rect 33367 25792 33508 25820
rect 33367 25789 33379 25792
rect 33321 25783 33379 25789
rect 32398 25752 32404 25764
rect 30607 25724 30788 25752
rect 32359 25724 32404 25752
rect 30607 25721 30619 25724
rect 30561 25715 30619 25721
rect 32398 25712 32404 25724
rect 32456 25712 32462 25764
rect 28169 25687 28227 25693
rect 28169 25653 28181 25687
rect 28215 25684 28227 25687
rect 28258 25684 28264 25696
rect 28215 25656 28264 25684
rect 28215 25653 28227 25656
rect 28169 25647 28227 25653
rect 28258 25644 28264 25656
rect 28316 25644 28322 25696
rect 28718 25684 28724 25696
rect 28679 25656 28724 25684
rect 28718 25644 28724 25656
rect 28776 25644 28782 25696
rect 32306 25684 32312 25696
rect 32267 25656 32312 25684
rect 32306 25644 32312 25656
rect 32364 25684 32370 25696
rect 33244 25684 33272 25783
rect 33502 25780 33508 25792
rect 33560 25820 33566 25832
rect 33689 25823 33747 25829
rect 33689 25820 33701 25823
rect 33560 25792 33701 25820
rect 33560 25780 33566 25792
rect 33689 25789 33701 25792
rect 33735 25789 33747 25823
rect 35802 25820 35808 25832
rect 35763 25792 35808 25820
rect 33689 25783 33747 25789
rect 35802 25780 35808 25792
rect 35860 25780 35866 25832
rect 36078 25820 36084 25832
rect 36039 25792 36084 25820
rect 36078 25780 36084 25792
rect 36136 25780 36142 25832
rect 32364 25656 33272 25684
rect 32364 25644 32370 25656
rect 1104 25594 38548 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 38548 25594
rect 1104 25520 38548 25542
rect 6181 25483 6239 25489
rect 6181 25449 6193 25483
rect 6227 25480 6239 25483
rect 7098 25480 7104 25492
rect 6227 25452 7104 25480
rect 6227 25449 6239 25452
rect 6181 25443 6239 25449
rect 7098 25440 7104 25452
rect 7156 25480 7162 25492
rect 9953 25483 10011 25489
rect 7156 25452 7788 25480
rect 7156 25440 7162 25452
rect 7190 25412 7196 25424
rect 7151 25384 7196 25412
rect 7190 25372 7196 25384
rect 7248 25372 7254 25424
rect 7760 25412 7788 25452
rect 9953 25449 9965 25483
rect 9999 25480 10011 25483
rect 10594 25480 10600 25492
rect 9999 25452 10600 25480
rect 9999 25449 10011 25452
rect 9953 25443 10011 25449
rect 10594 25440 10600 25452
rect 10652 25440 10658 25492
rect 12066 25480 12072 25492
rect 12027 25452 12072 25480
rect 12066 25440 12072 25452
rect 12124 25440 12130 25492
rect 12529 25483 12587 25489
rect 12529 25449 12541 25483
rect 12575 25480 12587 25483
rect 12618 25480 12624 25492
rect 12575 25452 12624 25480
rect 12575 25449 12587 25452
rect 12529 25443 12587 25449
rect 12618 25440 12624 25452
rect 12676 25440 12682 25492
rect 14366 25480 14372 25492
rect 14327 25452 14372 25480
rect 14366 25440 14372 25452
rect 14424 25440 14430 25492
rect 15010 25440 15016 25492
rect 15068 25480 15074 25492
rect 15473 25483 15531 25489
rect 15473 25480 15485 25483
rect 15068 25452 15485 25480
rect 15068 25440 15074 25452
rect 15473 25449 15485 25452
rect 15519 25480 15531 25483
rect 15930 25480 15936 25492
rect 15519 25452 15936 25480
rect 15519 25449 15531 25452
rect 15473 25443 15531 25449
rect 15930 25440 15936 25452
rect 15988 25480 15994 25492
rect 16758 25480 16764 25492
rect 15988 25452 16764 25480
rect 15988 25440 15994 25452
rect 16758 25440 16764 25452
rect 16816 25440 16822 25492
rect 18325 25483 18383 25489
rect 18325 25449 18337 25483
rect 18371 25480 18383 25483
rect 18506 25480 18512 25492
rect 18371 25452 18512 25480
rect 18371 25449 18383 25452
rect 18325 25443 18383 25449
rect 18506 25440 18512 25452
rect 18564 25440 18570 25492
rect 19426 25480 19432 25492
rect 19387 25452 19432 25480
rect 19426 25440 19432 25452
rect 19484 25440 19490 25492
rect 21177 25483 21235 25489
rect 21177 25449 21189 25483
rect 21223 25480 21235 25483
rect 21542 25480 21548 25492
rect 21223 25452 21548 25480
rect 21223 25449 21235 25452
rect 21177 25443 21235 25449
rect 21542 25440 21548 25452
rect 21600 25440 21606 25492
rect 23198 25440 23204 25492
rect 23256 25480 23262 25492
rect 23658 25480 23664 25492
rect 23256 25452 23664 25480
rect 23256 25440 23262 25452
rect 23658 25440 23664 25452
rect 23716 25440 23722 25492
rect 28997 25483 29055 25489
rect 28997 25449 29009 25483
rect 29043 25480 29055 25483
rect 29546 25480 29552 25492
rect 29043 25452 29552 25480
rect 29043 25449 29055 25452
rect 28997 25443 29055 25449
rect 29546 25440 29552 25452
rect 29604 25440 29610 25492
rect 30190 25480 30196 25492
rect 29840 25452 30196 25480
rect 8941 25415 8999 25421
rect 8941 25412 8953 25415
rect 7760 25384 8953 25412
rect 4341 25347 4399 25353
rect 4341 25313 4353 25347
rect 4387 25344 4399 25347
rect 4617 25347 4675 25353
rect 4617 25344 4629 25347
rect 4387 25316 4629 25344
rect 4387 25313 4399 25316
rect 4341 25307 4399 25313
rect 4617 25313 4629 25316
rect 4663 25344 4675 25347
rect 5074 25344 5080 25356
rect 4663 25316 5080 25344
rect 4663 25313 4675 25316
rect 4617 25307 4675 25313
rect 5074 25304 5080 25316
rect 5132 25304 5138 25356
rect 5169 25347 5227 25353
rect 5169 25313 5181 25347
rect 5215 25344 5227 25347
rect 5442 25344 5448 25356
rect 5215 25316 5448 25344
rect 5215 25313 5227 25316
rect 5169 25307 5227 25313
rect 5442 25304 5448 25316
rect 5500 25304 5506 25356
rect 7653 25347 7711 25353
rect 7653 25344 7665 25347
rect 7208 25316 7665 25344
rect 7208 25288 7236 25316
rect 7653 25313 7665 25316
rect 7699 25313 7711 25347
rect 7760 25344 7788 25384
rect 8941 25381 8953 25384
rect 8987 25412 8999 25415
rect 9490 25412 9496 25424
rect 8987 25384 9496 25412
rect 8987 25381 8999 25384
rect 8941 25375 8999 25381
rect 9490 25372 9496 25384
rect 9548 25372 9554 25424
rect 10413 25415 10471 25421
rect 10413 25381 10425 25415
rect 10459 25412 10471 25415
rect 16666 25412 16672 25424
rect 10459 25384 11652 25412
rect 16627 25384 16672 25412
rect 10459 25381 10471 25384
rect 10413 25375 10471 25381
rect 11624 25356 11652 25384
rect 16666 25372 16672 25384
rect 16724 25372 16730 25424
rect 27249 25415 27307 25421
rect 27249 25381 27261 25415
rect 27295 25412 27307 25415
rect 27430 25412 27436 25424
rect 27295 25384 27436 25412
rect 27295 25381 27307 25384
rect 27249 25375 27307 25381
rect 27430 25372 27436 25384
rect 27488 25372 27494 25424
rect 29840 25421 29868 25452
rect 30190 25440 30196 25452
rect 30248 25440 30254 25492
rect 30558 25440 30564 25492
rect 30616 25480 30622 25492
rect 30929 25483 30987 25489
rect 30929 25480 30941 25483
rect 30616 25452 30941 25480
rect 30616 25440 30622 25452
rect 30929 25449 30941 25452
rect 30975 25449 30987 25483
rect 31846 25480 31852 25492
rect 31807 25452 31852 25480
rect 30929 25443 30987 25449
rect 31846 25440 31852 25452
rect 31904 25440 31910 25492
rect 32858 25440 32864 25492
rect 32916 25480 32922 25492
rect 33689 25483 33747 25489
rect 33689 25480 33701 25483
rect 32916 25452 33701 25480
rect 32916 25440 32922 25452
rect 33689 25449 33701 25452
rect 33735 25449 33747 25483
rect 35802 25480 35808 25492
rect 35763 25452 35808 25480
rect 33689 25443 33747 25449
rect 35802 25440 35808 25452
rect 35860 25440 35866 25492
rect 29825 25415 29883 25421
rect 29825 25381 29837 25415
rect 29871 25381 29883 25415
rect 32674 25412 32680 25424
rect 32635 25384 32680 25412
rect 29825 25375 29883 25381
rect 32674 25372 32680 25384
rect 32732 25372 32738 25424
rect 7837 25347 7895 25353
rect 7837 25344 7849 25347
rect 7760 25316 7849 25344
rect 7653 25307 7711 25313
rect 7837 25313 7849 25316
rect 7883 25313 7895 25347
rect 8110 25344 8116 25356
rect 8071 25316 8116 25344
rect 7837 25307 7895 25313
rect 8110 25304 8116 25316
rect 8168 25304 8174 25356
rect 8665 25347 8723 25353
rect 8665 25313 8677 25347
rect 8711 25344 8723 25347
rect 8846 25344 8852 25356
rect 8711 25316 8852 25344
rect 8711 25313 8723 25316
rect 8665 25307 8723 25313
rect 8846 25304 8852 25316
rect 8904 25304 8910 25356
rect 11238 25344 11244 25356
rect 11199 25316 11244 25344
rect 11238 25304 11244 25316
rect 11296 25304 11302 25356
rect 11606 25344 11612 25356
rect 11567 25316 11612 25344
rect 11606 25304 11612 25316
rect 11664 25304 11670 25356
rect 12621 25347 12679 25353
rect 12621 25313 12633 25347
rect 12667 25344 12679 25347
rect 12894 25344 12900 25356
rect 12667 25316 12900 25344
rect 12667 25313 12679 25316
rect 12621 25307 12679 25313
rect 12894 25304 12900 25316
rect 12952 25304 12958 25356
rect 13170 25344 13176 25356
rect 13131 25316 13176 25344
rect 13170 25304 13176 25316
rect 13228 25304 13234 25356
rect 13354 25344 13360 25356
rect 13315 25316 13360 25344
rect 13354 25304 13360 25316
rect 13412 25304 13418 25356
rect 13538 25344 13544 25356
rect 13499 25316 13544 25344
rect 13538 25304 13544 25316
rect 13596 25304 13602 25356
rect 14090 25344 14096 25356
rect 14051 25316 14096 25344
rect 14090 25304 14096 25316
rect 14148 25304 14154 25356
rect 16574 25304 16580 25356
rect 16632 25344 16638 25356
rect 17129 25347 17187 25353
rect 17129 25344 17141 25347
rect 16632 25316 17141 25344
rect 16632 25304 16638 25316
rect 17129 25313 17141 25316
rect 17175 25344 17187 25347
rect 17402 25344 17408 25356
rect 17175 25316 17408 25344
rect 17175 25313 17187 25316
rect 17129 25307 17187 25313
rect 17402 25304 17408 25316
rect 17460 25304 17466 25356
rect 17494 25304 17500 25356
rect 17552 25344 17558 25356
rect 17862 25344 17868 25356
rect 17552 25316 17868 25344
rect 17552 25304 17558 25316
rect 17862 25304 17868 25316
rect 17920 25304 17926 25356
rect 21082 25304 21088 25356
rect 21140 25344 21146 25356
rect 21545 25347 21603 25353
rect 21545 25344 21557 25347
rect 21140 25316 21557 25344
rect 21140 25304 21146 25316
rect 21545 25313 21557 25316
rect 21591 25313 21603 25347
rect 21910 25344 21916 25356
rect 21871 25316 21916 25344
rect 21545 25307 21603 25313
rect 21910 25304 21916 25316
rect 21968 25304 21974 25356
rect 25409 25347 25467 25353
rect 25409 25313 25421 25347
rect 25455 25344 25467 25347
rect 25590 25344 25596 25356
rect 25455 25316 25596 25344
rect 25455 25313 25467 25316
rect 25409 25307 25467 25313
rect 25590 25304 25596 25316
rect 25648 25344 25654 25356
rect 25958 25344 25964 25356
rect 25648 25316 25964 25344
rect 25648 25304 25654 25316
rect 25958 25304 25964 25316
rect 26016 25304 26022 25356
rect 28077 25347 28135 25353
rect 28077 25313 28089 25347
rect 28123 25344 28135 25347
rect 29270 25344 29276 25356
rect 28123 25316 29276 25344
rect 28123 25313 28135 25316
rect 28077 25307 28135 25313
rect 29270 25304 29276 25316
rect 29328 25304 29334 25356
rect 29365 25347 29423 25353
rect 29365 25313 29377 25347
rect 29411 25344 29423 25347
rect 29454 25344 29460 25356
rect 29411 25316 29460 25344
rect 29411 25313 29423 25316
rect 29365 25307 29423 25313
rect 29454 25304 29460 25316
rect 29512 25304 29518 25356
rect 30558 25304 30564 25356
rect 30616 25344 30622 25356
rect 30653 25347 30711 25353
rect 30653 25344 30665 25347
rect 30616 25316 30665 25344
rect 30616 25304 30622 25316
rect 30653 25313 30665 25316
rect 30699 25313 30711 25347
rect 30653 25307 30711 25313
rect 30837 25347 30895 25353
rect 30837 25313 30849 25347
rect 30883 25313 30895 25347
rect 32214 25344 32220 25356
rect 32127 25316 32220 25344
rect 30837 25307 30895 25313
rect 4798 25236 4804 25288
rect 4856 25276 4862 25288
rect 5258 25276 5264 25288
rect 4856 25248 5264 25276
rect 4856 25236 4862 25248
rect 5258 25236 5264 25248
rect 5316 25236 5322 25288
rect 7190 25236 7196 25288
rect 7248 25236 7254 25288
rect 8297 25279 8355 25285
rect 8297 25245 8309 25279
rect 8343 25276 8355 25279
rect 8386 25276 8392 25288
rect 8343 25248 8392 25276
rect 8343 25245 8355 25248
rect 8297 25239 8355 25245
rect 4709 25211 4767 25217
rect 4709 25177 4721 25211
rect 4755 25208 4767 25211
rect 4982 25208 4988 25220
rect 4755 25180 4988 25208
rect 4755 25177 4767 25180
rect 4709 25171 4767 25177
rect 4982 25168 4988 25180
rect 5040 25168 5046 25220
rect 7006 25208 7012 25220
rect 6472 25180 7012 25208
rect 6472 25152 6500 25180
rect 7006 25168 7012 25180
rect 7064 25168 7070 25220
rect 7834 25168 7840 25220
rect 7892 25208 7898 25220
rect 8312 25208 8340 25239
rect 8386 25236 8392 25248
rect 8444 25236 8450 25288
rect 10870 25236 10876 25288
rect 10928 25276 10934 25288
rect 11333 25279 11391 25285
rect 11333 25276 11345 25279
rect 10928 25248 11345 25276
rect 10928 25236 10934 25248
rect 11333 25245 11345 25248
rect 11379 25276 11391 25279
rect 11422 25276 11428 25288
rect 11379 25248 11428 25276
rect 11379 25245 11391 25248
rect 11333 25239 11391 25245
rect 11422 25236 11428 25248
rect 11480 25236 11486 25288
rect 11514 25236 11520 25288
rect 11572 25276 11578 25288
rect 11701 25279 11759 25285
rect 11701 25276 11713 25279
rect 11572 25248 11713 25276
rect 11572 25236 11578 25248
rect 11701 25245 11713 25248
rect 11747 25276 11759 25279
rect 11882 25276 11888 25288
rect 11747 25248 11888 25276
rect 11747 25245 11759 25248
rect 11701 25239 11759 25245
rect 11882 25236 11888 25248
rect 11940 25236 11946 25288
rect 13722 25276 13728 25288
rect 13683 25248 13728 25276
rect 13722 25236 13728 25248
rect 13780 25236 13786 25288
rect 15930 25276 15936 25288
rect 15843 25248 15936 25276
rect 15930 25236 15936 25248
rect 15988 25276 15994 25288
rect 17218 25276 17224 25288
rect 15988 25248 17224 25276
rect 15988 25236 15994 25248
rect 17218 25236 17224 25248
rect 17276 25276 17282 25288
rect 17589 25279 17647 25285
rect 17589 25276 17601 25279
rect 17276 25248 17601 25276
rect 17276 25236 17282 25248
rect 17589 25245 17601 25248
rect 17635 25245 17647 25279
rect 21358 25276 21364 25288
rect 21319 25248 21364 25276
rect 17589 25239 17647 25245
rect 21358 25236 21364 25248
rect 21416 25236 21422 25288
rect 21726 25236 21732 25288
rect 21784 25276 21790 25288
rect 21821 25279 21879 25285
rect 21821 25276 21833 25279
rect 21784 25248 21833 25276
rect 21784 25236 21790 25248
rect 21821 25245 21833 25248
rect 21867 25245 21879 25279
rect 21821 25239 21879 25245
rect 27614 25236 27620 25288
rect 27672 25276 27678 25288
rect 27801 25279 27859 25285
rect 27801 25276 27813 25279
rect 27672 25248 27813 25276
rect 27672 25236 27678 25248
rect 27801 25245 27813 25248
rect 27847 25245 27859 25279
rect 28258 25276 28264 25288
rect 28219 25248 28264 25276
rect 27801 25239 27859 25245
rect 28258 25236 28264 25248
rect 28316 25276 28322 25288
rect 29089 25279 29147 25285
rect 29089 25276 29101 25279
rect 28316 25248 29101 25276
rect 28316 25236 28322 25248
rect 29089 25245 29101 25248
rect 29135 25245 29147 25279
rect 30852 25276 30880 25307
rect 32214 25304 32220 25316
rect 32272 25344 32278 25356
rect 32582 25344 32588 25356
rect 32272 25316 32588 25344
rect 32272 25304 32278 25316
rect 32582 25304 32588 25316
rect 32640 25304 32646 25356
rect 33502 25344 33508 25356
rect 33463 25316 33508 25344
rect 33502 25304 33508 25316
rect 33560 25304 33566 25356
rect 31481 25279 31539 25285
rect 31481 25276 31493 25279
rect 29089 25239 29147 25245
rect 30484 25248 31493 25276
rect 30484 25220 30512 25248
rect 31481 25245 31493 25248
rect 31527 25245 31539 25279
rect 31481 25239 31539 25245
rect 32125 25279 32183 25285
rect 32125 25245 32137 25279
rect 32171 25276 32183 25279
rect 32171 25248 32260 25276
rect 32171 25245 32183 25248
rect 32125 25239 32183 25245
rect 32232 25220 32260 25248
rect 7892 25180 8340 25208
rect 10689 25211 10747 25217
rect 7892 25168 7898 25180
rect 10689 25177 10701 25211
rect 10735 25208 10747 25211
rect 13354 25208 13360 25220
rect 10735 25180 13360 25208
rect 10735 25177 10747 25180
rect 10689 25171 10747 25177
rect 13354 25168 13360 25180
rect 13412 25168 13418 25220
rect 15105 25211 15163 25217
rect 15105 25177 15117 25211
rect 15151 25208 15163 25211
rect 15378 25208 15384 25220
rect 15151 25180 15384 25208
rect 15151 25177 15163 25180
rect 15105 25171 15163 25177
rect 15378 25168 15384 25180
rect 15436 25208 15442 25220
rect 16298 25208 16304 25220
rect 15436 25180 16304 25208
rect 15436 25168 15442 25180
rect 16298 25168 16304 25180
rect 16356 25168 16362 25220
rect 16666 25168 16672 25220
rect 16724 25208 16730 25220
rect 17770 25208 17776 25220
rect 16724 25180 17776 25208
rect 16724 25168 16730 25180
rect 17770 25168 17776 25180
rect 17828 25168 17834 25220
rect 25041 25211 25099 25217
rect 25041 25177 25053 25211
rect 25087 25208 25099 25211
rect 25682 25208 25688 25220
rect 25087 25180 25688 25208
rect 25087 25177 25099 25180
rect 25041 25171 25099 25177
rect 25682 25168 25688 25180
rect 25740 25208 25746 25220
rect 26418 25208 26424 25220
rect 25740 25180 26424 25208
rect 25740 25168 25746 25180
rect 26418 25168 26424 25180
rect 26476 25168 26482 25220
rect 30466 25168 30472 25220
rect 30524 25168 30530 25220
rect 32214 25168 32220 25220
rect 32272 25168 32278 25220
rect 1670 25140 1676 25152
rect 1583 25112 1676 25140
rect 1670 25100 1676 25112
rect 1728 25140 1734 25152
rect 2958 25140 2964 25152
rect 1728 25112 2964 25140
rect 1728 25100 1734 25112
rect 2958 25100 2964 25112
rect 3016 25100 3022 25152
rect 6454 25140 6460 25152
rect 6415 25112 6460 25140
rect 6454 25100 6460 25112
rect 6512 25100 6518 25152
rect 6914 25140 6920 25152
rect 6875 25112 6920 25140
rect 6914 25100 6920 25112
rect 6972 25100 6978 25152
rect 9493 25143 9551 25149
rect 9493 25109 9505 25143
rect 9539 25140 9551 25143
rect 9582 25140 9588 25152
rect 9539 25112 9588 25140
rect 9539 25109 9551 25112
rect 9493 25103 9551 25109
rect 9582 25100 9588 25112
rect 9640 25100 9646 25152
rect 11422 25100 11428 25152
rect 11480 25140 11486 25152
rect 12618 25140 12624 25152
rect 11480 25112 12624 25140
rect 11480 25100 11486 25112
rect 12618 25100 12624 25112
rect 12676 25100 12682 25152
rect 16206 25140 16212 25152
rect 16167 25112 16212 25140
rect 16206 25100 16212 25112
rect 16264 25100 16270 25152
rect 25593 25143 25651 25149
rect 25593 25109 25605 25143
rect 25639 25140 25651 25143
rect 25866 25140 25872 25152
rect 25639 25112 25872 25140
rect 25639 25109 25651 25112
rect 25593 25103 25651 25109
rect 25866 25100 25872 25112
rect 25924 25100 25930 25152
rect 26786 25140 26792 25152
rect 26747 25112 26792 25140
rect 26786 25100 26792 25112
rect 26844 25100 26850 25152
rect 27062 25140 27068 25152
rect 27023 25112 27068 25140
rect 27062 25100 27068 25112
rect 27120 25100 27126 25152
rect 30561 25143 30619 25149
rect 30561 25109 30573 25143
rect 30607 25140 30619 25143
rect 31110 25140 31116 25152
rect 30607 25112 31116 25140
rect 30607 25109 30619 25112
rect 30561 25103 30619 25109
rect 31110 25100 31116 25112
rect 31168 25140 31174 25152
rect 31570 25140 31576 25152
rect 31168 25112 31576 25140
rect 31168 25100 31174 25112
rect 31570 25100 31576 25112
rect 31628 25100 31634 25152
rect 1104 25050 38548 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 38548 25050
rect 1104 24976 38548 24998
rect 6914 24896 6920 24948
rect 6972 24896 6978 24948
rect 10781 24939 10839 24945
rect 10781 24905 10793 24939
rect 10827 24936 10839 24939
rect 10962 24936 10968 24948
rect 10827 24908 10968 24936
rect 10827 24905 10839 24908
rect 10781 24899 10839 24905
rect 10962 24896 10968 24908
rect 11020 24896 11026 24948
rect 13722 24936 13728 24948
rect 12452 24908 13728 24936
rect 3326 24828 3332 24880
rect 3384 24868 3390 24880
rect 3510 24868 3516 24880
rect 3384 24840 3516 24868
rect 3384 24828 3390 24840
rect 3510 24828 3516 24840
rect 3568 24828 3574 24880
rect 6932 24868 6960 24896
rect 8110 24868 8116 24880
rect 6840 24840 8116 24868
rect 4249 24803 4307 24809
rect 4249 24769 4261 24803
rect 4295 24800 4307 24803
rect 4617 24803 4675 24809
rect 4617 24800 4629 24803
rect 4295 24772 4629 24800
rect 4295 24769 4307 24772
rect 4249 24763 4307 24769
rect 4617 24769 4629 24772
rect 4663 24800 4675 24803
rect 5261 24803 5319 24809
rect 5261 24800 5273 24803
rect 4663 24772 5273 24800
rect 4663 24769 4675 24772
rect 4617 24763 4675 24769
rect 5261 24769 5273 24772
rect 5307 24800 5319 24803
rect 5442 24800 5448 24812
rect 5307 24772 5448 24800
rect 5307 24769 5319 24772
rect 5261 24763 5319 24769
rect 5442 24760 5448 24772
rect 5500 24760 5506 24812
rect 5813 24803 5871 24809
rect 5813 24769 5825 24803
rect 5859 24800 5871 24803
rect 6546 24800 6552 24812
rect 5859 24772 6552 24800
rect 5859 24769 5871 24772
rect 5813 24763 5871 24769
rect 6546 24760 6552 24772
rect 6604 24760 6610 24812
rect 3421 24735 3479 24741
rect 3421 24701 3433 24735
rect 3467 24732 3479 24735
rect 3510 24732 3516 24744
rect 3467 24704 3516 24732
rect 3467 24701 3479 24704
rect 3421 24695 3479 24701
rect 3510 24692 3516 24704
rect 3568 24732 3574 24744
rect 4157 24735 4215 24741
rect 4157 24732 4169 24735
rect 3568 24704 4169 24732
rect 3568 24692 3574 24704
rect 4157 24701 4169 24704
rect 4203 24732 4215 24735
rect 5166 24732 5172 24744
rect 4203 24704 5172 24732
rect 4203 24701 4215 24704
rect 4157 24695 4215 24701
rect 5166 24692 5172 24704
rect 5224 24692 5230 24744
rect 5353 24735 5411 24741
rect 5353 24701 5365 24735
rect 5399 24701 5411 24735
rect 5460 24732 5488 24760
rect 6089 24735 6147 24741
rect 6089 24732 6101 24735
rect 5460 24704 6101 24732
rect 5353 24695 5411 24701
rect 6089 24701 6101 24704
rect 6135 24701 6147 24735
rect 6089 24695 6147 24701
rect 5368 24664 5396 24695
rect 5092 24636 5396 24664
rect 5092 24608 5120 24636
rect 5626 24624 5632 24676
rect 5684 24664 5690 24676
rect 6840 24673 6868 24840
rect 8110 24828 8116 24840
rect 8168 24868 8174 24880
rect 8205 24871 8263 24877
rect 8205 24868 8217 24871
rect 8168 24840 8217 24868
rect 8168 24828 8174 24840
rect 8205 24837 8217 24840
rect 8251 24837 8263 24871
rect 8205 24831 8263 24837
rect 8220 24800 8248 24831
rect 9490 24828 9496 24880
rect 9548 24868 9554 24880
rect 9548 24840 9628 24868
rect 9548 24828 9554 24840
rect 8757 24803 8815 24809
rect 8757 24800 8769 24803
rect 8220 24772 8769 24800
rect 8757 24769 8769 24772
rect 8803 24800 8815 24803
rect 9600 24800 9628 24840
rect 10870 24828 10876 24880
rect 10928 24868 10934 24880
rect 12452 24868 12480 24908
rect 13722 24896 13728 24908
rect 13780 24936 13786 24948
rect 13909 24939 13967 24945
rect 13909 24936 13921 24939
rect 13780 24908 13921 24936
rect 13780 24896 13786 24908
rect 13909 24905 13921 24908
rect 13955 24905 13967 24939
rect 17218 24936 17224 24948
rect 17179 24908 17224 24936
rect 13909 24899 13967 24905
rect 17218 24896 17224 24908
rect 17276 24896 17282 24948
rect 17402 24896 17408 24948
rect 17460 24936 17466 24948
rect 17497 24939 17555 24945
rect 17497 24936 17509 24939
rect 17460 24908 17509 24936
rect 17460 24896 17466 24908
rect 17497 24905 17509 24908
rect 17543 24905 17555 24939
rect 17497 24899 17555 24905
rect 26973 24939 27031 24945
rect 26973 24905 26985 24939
rect 27019 24936 27031 24939
rect 27246 24936 27252 24948
rect 27019 24908 27252 24936
rect 27019 24905 27031 24908
rect 26973 24899 27031 24905
rect 27246 24896 27252 24908
rect 27304 24936 27310 24948
rect 29089 24939 29147 24945
rect 29089 24936 29101 24939
rect 27304 24908 29101 24936
rect 27304 24896 27310 24908
rect 29089 24905 29101 24908
rect 29135 24936 29147 24939
rect 29270 24936 29276 24948
rect 29135 24908 29276 24936
rect 29135 24905 29147 24908
rect 29089 24899 29147 24905
rect 29270 24896 29276 24908
rect 29328 24896 29334 24948
rect 10928 24840 12480 24868
rect 12529 24871 12587 24877
rect 10928 24828 10934 24840
rect 12529 24837 12541 24871
rect 12575 24868 12587 24871
rect 13170 24868 13176 24880
rect 12575 24840 13176 24868
rect 12575 24837 12587 24840
rect 12529 24831 12587 24837
rect 13170 24828 13176 24840
rect 13228 24828 13234 24880
rect 13354 24828 13360 24880
rect 13412 24868 13418 24880
rect 13412 24840 13768 24868
rect 13412 24828 13418 24840
rect 9858 24800 9864 24812
rect 8803 24772 9536 24800
rect 9600 24772 9864 24800
rect 8803 24769 8815 24772
rect 8757 24763 8815 24769
rect 7006 24692 7012 24744
rect 7064 24732 7070 24744
rect 7101 24735 7159 24741
rect 7101 24732 7113 24735
rect 7064 24704 7113 24732
rect 7064 24692 7070 24704
rect 7101 24701 7113 24704
rect 7147 24701 7159 24735
rect 7101 24695 7159 24701
rect 7282 24692 7288 24744
rect 7340 24732 7346 24744
rect 7561 24735 7619 24741
rect 7561 24732 7573 24735
rect 7340 24704 7573 24732
rect 7340 24692 7346 24704
rect 7561 24701 7573 24704
rect 7607 24732 7619 24735
rect 8202 24732 8208 24744
rect 7607 24704 8208 24732
rect 7607 24701 7619 24704
rect 7561 24695 7619 24701
rect 8202 24692 8208 24704
rect 8260 24692 8266 24744
rect 9398 24732 9404 24744
rect 9359 24704 9404 24732
rect 9398 24692 9404 24704
rect 9456 24692 9462 24744
rect 6825 24667 6883 24673
rect 6825 24664 6837 24667
rect 5684 24636 6837 24664
rect 5684 24624 5690 24636
rect 6825 24633 6837 24636
rect 6871 24633 6883 24667
rect 7190 24664 7196 24676
rect 7151 24636 7196 24664
rect 6825 24627 6883 24633
rect 7190 24624 7196 24636
rect 7248 24624 7254 24676
rect 8938 24664 8944 24676
rect 8899 24636 8944 24664
rect 8938 24624 8944 24636
rect 8996 24624 9002 24676
rect 9508 24664 9536 24772
rect 9692 24741 9720 24772
rect 9858 24760 9864 24772
rect 9916 24760 9922 24812
rect 11790 24800 11796 24812
rect 11751 24772 11796 24800
rect 11790 24760 11796 24772
rect 11848 24760 11854 24812
rect 12710 24760 12716 24812
rect 12768 24800 12774 24812
rect 13541 24803 13599 24809
rect 13541 24800 13553 24803
rect 12768 24772 13553 24800
rect 12768 24760 12774 24772
rect 13541 24769 13553 24772
rect 13587 24769 13599 24803
rect 13740 24800 13768 24840
rect 14277 24803 14335 24809
rect 14277 24800 14289 24803
rect 13740 24772 14289 24800
rect 13541 24763 13599 24769
rect 14277 24769 14289 24772
rect 14323 24769 14335 24803
rect 15286 24800 15292 24812
rect 15247 24772 15292 24800
rect 14277 24763 14335 24769
rect 15286 24760 15292 24772
rect 15344 24760 15350 24812
rect 16206 24800 16212 24812
rect 16167 24772 16212 24800
rect 16206 24760 16212 24772
rect 16264 24760 16270 24812
rect 17236 24800 17264 24896
rect 27062 24828 27068 24880
rect 27120 24868 27126 24880
rect 27706 24868 27712 24880
rect 27120 24840 27712 24868
rect 27120 24828 27126 24840
rect 27706 24828 27712 24840
rect 27764 24828 27770 24880
rect 31570 24868 31576 24880
rect 31483 24840 31576 24868
rect 31570 24828 31576 24840
rect 31628 24868 31634 24880
rect 32769 24871 32827 24877
rect 32769 24868 32781 24871
rect 31628 24840 32781 24868
rect 31628 24828 31634 24840
rect 32769 24837 32781 24840
rect 32815 24837 32827 24871
rect 32769 24831 32827 24837
rect 16684 24772 17264 24800
rect 19797 24803 19855 24809
rect 9677 24735 9735 24741
rect 9677 24701 9689 24735
rect 9723 24701 9735 24735
rect 9766 24732 9772 24744
rect 9677 24695 9735 24701
rect 9765 24692 9772 24732
rect 9824 24732 9830 24744
rect 10042 24732 10048 24744
rect 9824 24704 9869 24732
rect 10003 24704 10048 24732
rect 9824 24692 9830 24704
rect 10042 24692 10048 24704
rect 10100 24692 10106 24744
rect 10413 24735 10471 24741
rect 10413 24701 10425 24735
rect 10459 24732 10471 24735
rect 10502 24732 10508 24744
rect 10459 24704 10508 24732
rect 10459 24701 10471 24704
rect 10413 24695 10471 24701
rect 10502 24692 10508 24704
rect 10560 24692 10566 24744
rect 11333 24735 11391 24741
rect 11333 24732 11345 24735
rect 11164 24704 11345 24732
rect 9765 24664 9793 24692
rect 9508 24636 9793 24664
rect 10060 24664 10088 24692
rect 11164 24673 11192 24704
rect 11333 24701 11345 24704
rect 11379 24732 11391 24735
rect 11422 24732 11428 24744
rect 11379 24704 11428 24732
rect 11379 24701 11391 24704
rect 11333 24695 11391 24701
rect 11422 24692 11428 24704
rect 11480 24692 11486 24744
rect 11514 24692 11520 24744
rect 11572 24732 11578 24744
rect 13078 24732 13084 24744
rect 11572 24704 13084 24732
rect 11572 24692 11578 24704
rect 13078 24692 13084 24704
rect 13136 24692 13142 24744
rect 13173 24735 13231 24741
rect 13173 24701 13185 24735
rect 13219 24732 13231 24735
rect 13262 24732 13268 24744
rect 13219 24704 13268 24732
rect 13219 24701 13231 24704
rect 13173 24695 13231 24701
rect 11149 24667 11207 24673
rect 11149 24664 11161 24667
rect 10060 24636 11161 24664
rect 11149 24633 11161 24636
rect 11195 24633 11207 24667
rect 11149 24627 11207 24633
rect 11790 24624 11796 24676
rect 11848 24664 11854 24676
rect 13188 24664 13216 24695
rect 13262 24692 13268 24704
rect 13320 24692 13326 24744
rect 13446 24732 13452 24744
rect 13407 24704 13452 24732
rect 13446 24692 13452 24704
rect 13504 24692 13510 24744
rect 14461 24735 14519 24741
rect 14461 24701 14473 24735
rect 14507 24732 14519 24735
rect 14921 24735 14979 24741
rect 14921 24732 14933 24735
rect 14507 24704 14933 24732
rect 14507 24701 14519 24704
rect 14461 24695 14519 24701
rect 14921 24701 14933 24704
rect 14967 24701 14979 24735
rect 16298 24732 16304 24744
rect 16259 24704 16304 24732
rect 14921 24695 14979 24701
rect 14476 24664 14504 24695
rect 16298 24692 16304 24704
rect 16356 24692 16362 24744
rect 16684 24741 16712 24772
rect 19797 24769 19809 24803
rect 19843 24800 19855 24803
rect 20165 24803 20223 24809
rect 20165 24800 20177 24803
rect 19843 24772 20177 24800
rect 19843 24769 19855 24772
rect 19797 24763 19855 24769
rect 20165 24769 20177 24772
rect 20211 24800 20223 24803
rect 20622 24800 20628 24812
rect 20211 24772 20628 24800
rect 20211 24769 20223 24772
rect 20165 24763 20223 24769
rect 20622 24760 20628 24772
rect 20680 24760 20686 24812
rect 21545 24803 21603 24809
rect 21545 24769 21557 24803
rect 21591 24800 21603 24803
rect 21910 24800 21916 24812
rect 21591 24772 21916 24800
rect 21591 24769 21603 24772
rect 21545 24763 21603 24769
rect 21910 24760 21916 24772
rect 21968 24800 21974 24812
rect 22189 24803 22247 24809
rect 22189 24800 22201 24803
rect 21968 24772 22201 24800
rect 21968 24760 21974 24772
rect 22189 24769 22201 24772
rect 22235 24769 22247 24803
rect 22189 24763 22247 24769
rect 24857 24803 24915 24809
rect 24857 24769 24869 24803
rect 24903 24800 24915 24803
rect 24903 24772 25360 24800
rect 24903 24769 24915 24772
rect 24857 24763 24915 24769
rect 16669 24735 16727 24741
rect 16669 24701 16681 24735
rect 16715 24701 16727 24735
rect 16669 24695 16727 24701
rect 16853 24735 16911 24741
rect 16853 24701 16865 24735
rect 16899 24732 16911 24735
rect 16942 24732 16948 24744
rect 16899 24704 16948 24732
rect 16899 24701 16911 24704
rect 16853 24695 16911 24701
rect 16942 24692 16948 24704
rect 17000 24692 17006 24744
rect 19886 24732 19892 24744
rect 19847 24704 19892 24732
rect 19886 24692 19892 24704
rect 19944 24692 19950 24744
rect 25332 24741 25360 24772
rect 25866 24760 25872 24812
rect 25924 24800 25930 24812
rect 27249 24803 27307 24809
rect 27249 24800 27261 24803
rect 25924 24772 27261 24800
rect 25924 24760 25930 24772
rect 27249 24769 27261 24772
rect 27295 24800 27307 24803
rect 28258 24800 28264 24812
rect 27295 24772 28264 24800
rect 27295 24769 27307 24772
rect 27249 24763 27307 24769
rect 28258 24760 28264 24772
rect 28316 24800 28322 24812
rect 29733 24803 29791 24809
rect 29733 24800 29745 24803
rect 28316 24772 29745 24800
rect 28316 24760 28322 24772
rect 29733 24769 29745 24772
rect 29779 24769 29791 24803
rect 29733 24763 29791 24769
rect 31205 24803 31263 24809
rect 31205 24769 31217 24803
rect 31251 24800 31263 24803
rect 31386 24800 31392 24812
rect 31251 24772 31392 24800
rect 31251 24769 31263 24772
rect 31205 24763 31263 24769
rect 31386 24760 31392 24772
rect 31444 24760 31450 24812
rect 24949 24735 25007 24741
rect 24949 24732 24961 24735
rect 24412 24704 24961 24732
rect 11848 24636 14504 24664
rect 11848 24624 11854 24636
rect 24412 24608 24440 24704
rect 24949 24701 24961 24704
rect 24995 24701 25007 24735
rect 24949 24695 25007 24701
rect 25317 24735 25375 24741
rect 25317 24701 25329 24735
rect 25363 24732 25375 24735
rect 25590 24732 25596 24744
rect 25363 24704 25596 24732
rect 25363 24701 25375 24704
rect 25317 24695 25375 24701
rect 25590 24692 25596 24704
rect 25648 24692 25654 24744
rect 25682 24692 25688 24744
rect 25740 24732 25746 24744
rect 26234 24732 26240 24744
rect 25740 24704 25785 24732
rect 26195 24704 26240 24732
rect 25740 24692 25746 24704
rect 26234 24692 26240 24704
rect 26292 24692 26298 24744
rect 27614 24732 27620 24744
rect 27575 24704 27620 24732
rect 27614 24692 27620 24704
rect 27672 24692 27678 24744
rect 27893 24735 27951 24741
rect 27893 24701 27905 24735
rect 27939 24701 27951 24735
rect 27893 24695 27951 24701
rect 29273 24735 29331 24741
rect 29273 24701 29285 24735
rect 29319 24732 29331 24735
rect 29362 24732 29368 24744
rect 29319 24704 29368 24732
rect 29319 24701 29331 24704
rect 29273 24695 29331 24701
rect 26145 24667 26203 24673
rect 26145 24633 26157 24667
rect 26191 24664 26203 24667
rect 26418 24664 26424 24676
rect 26191 24636 26424 24664
rect 26191 24633 26203 24636
rect 26145 24627 26203 24633
rect 26418 24624 26424 24636
rect 26476 24624 26482 24676
rect 27908 24664 27936 24695
rect 29362 24692 29368 24704
rect 29420 24692 29426 24744
rect 29454 24692 29460 24744
rect 29512 24732 29518 24744
rect 30101 24735 30159 24741
rect 30101 24732 30113 24735
rect 29512 24704 30113 24732
rect 29512 24692 29518 24704
rect 30101 24701 30113 24704
rect 30147 24701 30159 24735
rect 30101 24695 30159 24701
rect 30561 24735 30619 24741
rect 30561 24701 30573 24735
rect 30607 24732 30619 24735
rect 31478 24732 31484 24744
rect 30607 24704 31484 24732
rect 30607 24701 30619 24704
rect 30561 24695 30619 24701
rect 31478 24692 31484 24704
rect 31536 24692 31542 24744
rect 31588 24732 31616 24828
rect 32122 24760 32128 24812
rect 32180 24800 32186 24812
rect 35713 24803 35771 24809
rect 32180 24772 32628 24800
rect 32180 24760 32186 24772
rect 32600 24741 32628 24772
rect 35713 24769 35725 24803
rect 35759 24800 35771 24803
rect 36081 24803 36139 24809
rect 36081 24800 36093 24803
rect 35759 24772 36093 24800
rect 35759 24769 35771 24772
rect 35713 24763 35771 24769
rect 36081 24769 36093 24772
rect 36127 24800 36139 24803
rect 37182 24800 37188 24812
rect 36127 24772 37188 24800
rect 36127 24769 36139 24772
rect 36081 24763 36139 24769
rect 37182 24760 37188 24772
rect 37240 24760 37246 24812
rect 31665 24735 31723 24741
rect 31665 24732 31677 24735
rect 31588 24704 31677 24732
rect 31665 24701 31677 24704
rect 31711 24701 31723 24735
rect 31665 24695 31723 24701
rect 32585 24735 32643 24741
rect 32585 24701 32597 24735
rect 32631 24732 32643 24735
rect 32950 24732 32956 24744
rect 32631 24704 32956 24732
rect 32631 24701 32643 24704
rect 32585 24695 32643 24701
rect 32950 24692 32956 24704
rect 33008 24692 33014 24744
rect 35802 24732 35808 24744
rect 35763 24704 35808 24732
rect 35802 24692 35808 24704
rect 35860 24692 35866 24744
rect 28258 24664 28264 24676
rect 27540 24636 28264 24664
rect 5074 24596 5080 24608
rect 5035 24568 5080 24596
rect 5074 24556 5080 24568
rect 5132 24556 5138 24608
rect 6641 24599 6699 24605
rect 6641 24565 6653 24599
rect 6687 24596 6699 24599
rect 6914 24596 6920 24608
rect 6687 24568 6920 24596
rect 6687 24565 6699 24568
rect 6641 24559 6699 24565
rect 6914 24556 6920 24568
rect 6972 24596 6978 24608
rect 7009 24599 7067 24605
rect 7009 24596 7021 24599
rect 6972 24568 7021 24596
rect 6972 24556 6978 24568
rect 7009 24565 7021 24568
rect 7055 24565 7067 24599
rect 7834 24596 7840 24608
rect 7795 24568 7840 24596
rect 7009 24559 7067 24565
rect 7834 24556 7840 24568
rect 7892 24556 7898 24608
rect 11517 24599 11575 24605
rect 11517 24565 11529 24599
rect 11563 24596 11575 24599
rect 11606 24596 11612 24608
rect 11563 24568 11612 24596
rect 11563 24565 11575 24568
rect 11517 24559 11575 24565
rect 11606 24556 11612 24568
rect 11664 24556 11670 24608
rect 12250 24596 12256 24608
rect 12211 24568 12256 24596
rect 12250 24556 12256 24568
rect 12308 24556 12314 24608
rect 14645 24599 14703 24605
rect 14645 24565 14657 24599
rect 14691 24596 14703 24599
rect 15470 24596 15476 24608
rect 14691 24568 15476 24596
rect 14691 24565 14703 24568
rect 14645 24559 14703 24565
rect 15470 24556 15476 24568
rect 15528 24556 15534 24608
rect 15933 24599 15991 24605
rect 15933 24565 15945 24599
rect 15979 24596 15991 24599
rect 17034 24596 17040 24608
rect 15979 24568 17040 24596
rect 15979 24565 15991 24568
rect 15933 24559 15991 24565
rect 17034 24556 17040 24568
rect 17092 24556 17098 24608
rect 20254 24556 20260 24608
rect 20312 24596 20318 24608
rect 21726 24596 21732 24608
rect 20312 24568 21732 24596
rect 20312 24556 20318 24568
rect 21726 24556 21732 24568
rect 21784 24596 21790 24608
rect 21821 24599 21879 24605
rect 21821 24596 21833 24599
rect 21784 24568 21833 24596
rect 21784 24556 21790 24568
rect 21821 24565 21833 24568
rect 21867 24565 21879 24599
rect 24394 24596 24400 24608
rect 24355 24568 24400 24596
rect 21821 24559 21879 24565
rect 24394 24556 24400 24568
rect 24452 24556 24458 24608
rect 25958 24556 25964 24608
rect 26016 24596 26022 24608
rect 27540 24596 27568 24636
rect 28258 24624 28264 24636
rect 28316 24624 28322 24676
rect 28353 24667 28411 24673
rect 28353 24633 28365 24667
rect 28399 24664 28411 24667
rect 30006 24664 30012 24676
rect 28399 24636 30012 24664
rect 28399 24633 28411 24636
rect 28353 24627 28411 24633
rect 30006 24624 30012 24636
rect 30064 24624 30070 24676
rect 30653 24667 30711 24673
rect 30653 24633 30665 24667
rect 30699 24664 30711 24667
rect 31754 24664 31760 24676
rect 30699 24636 31760 24664
rect 30699 24633 30711 24636
rect 30653 24627 30711 24633
rect 31754 24624 31760 24636
rect 31812 24624 31818 24676
rect 26016 24568 27568 24596
rect 26016 24556 26022 24568
rect 27614 24556 27620 24608
rect 27672 24596 27678 24608
rect 28629 24599 28687 24605
rect 28629 24596 28641 24599
rect 27672 24568 28641 24596
rect 27672 24556 27678 24568
rect 28629 24565 28641 24568
rect 28675 24565 28687 24599
rect 28629 24559 28687 24565
rect 29457 24599 29515 24605
rect 29457 24565 29469 24599
rect 29503 24596 29515 24599
rect 29914 24596 29920 24608
rect 29503 24568 29920 24596
rect 29503 24565 29515 24568
rect 29457 24559 29515 24565
rect 29914 24556 29920 24568
rect 29972 24596 29978 24608
rect 30466 24596 30472 24608
rect 29972 24568 30472 24596
rect 29972 24556 29978 24568
rect 30466 24556 30472 24568
rect 30524 24556 30530 24608
rect 32214 24596 32220 24608
rect 32175 24568 32220 24596
rect 32214 24556 32220 24568
rect 32272 24556 32278 24608
rect 33502 24596 33508 24608
rect 33463 24568 33508 24596
rect 33502 24556 33508 24568
rect 33560 24556 33566 24608
rect 36078 24556 36084 24608
rect 36136 24596 36142 24608
rect 37185 24599 37243 24605
rect 37185 24596 37197 24599
rect 36136 24568 37197 24596
rect 36136 24556 36142 24568
rect 37185 24565 37197 24568
rect 37231 24565 37243 24599
rect 37185 24559 37243 24565
rect 1104 24506 38548 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 38548 24506
rect 1104 24432 38548 24454
rect 2961 24395 3019 24401
rect 2961 24361 2973 24395
rect 3007 24392 3019 24395
rect 3510 24392 3516 24404
rect 3007 24364 3516 24392
rect 3007 24361 3019 24364
rect 2961 24355 3019 24361
rect 3510 24352 3516 24364
rect 3568 24352 3574 24404
rect 7742 24392 7748 24404
rect 7703 24364 7748 24392
rect 7742 24352 7748 24364
rect 7800 24352 7806 24404
rect 16669 24395 16727 24401
rect 15120 24364 16620 24392
rect 4341 24327 4399 24333
rect 4341 24293 4353 24327
rect 4387 24324 4399 24327
rect 4890 24324 4896 24336
rect 4387 24296 4896 24324
rect 4387 24293 4399 24296
rect 4341 24287 4399 24293
rect 4890 24284 4896 24296
rect 4948 24284 4954 24336
rect 9677 24327 9735 24333
rect 9677 24293 9689 24327
rect 9723 24324 9735 24327
rect 11238 24324 11244 24336
rect 9723 24296 11244 24324
rect 9723 24293 9735 24296
rect 9677 24287 9735 24293
rect 11238 24284 11244 24296
rect 11296 24324 11302 24336
rect 11793 24327 11851 24333
rect 11793 24324 11805 24327
rect 11296 24296 11805 24324
rect 11296 24284 11302 24296
rect 11793 24293 11805 24296
rect 11839 24293 11851 24327
rect 11793 24287 11851 24293
rect 12894 24284 12900 24336
rect 12952 24324 12958 24336
rect 14645 24327 14703 24333
rect 14645 24324 14657 24327
rect 12952 24296 14657 24324
rect 12952 24284 12958 24296
rect 14645 24293 14657 24296
rect 14691 24293 14703 24327
rect 14645 24287 14703 24293
rect 1394 24256 1400 24268
rect 1355 24228 1400 24256
rect 1394 24216 1400 24228
rect 1452 24216 1458 24268
rect 4985 24259 5043 24265
rect 4985 24225 4997 24259
rect 5031 24256 5043 24259
rect 5258 24256 5264 24268
rect 5031 24228 5264 24256
rect 5031 24225 5043 24228
rect 4985 24219 5043 24225
rect 5258 24216 5264 24228
rect 5316 24216 5322 24268
rect 5353 24259 5411 24265
rect 5353 24225 5365 24259
rect 5399 24256 5411 24259
rect 5534 24256 5540 24268
rect 5399 24228 5540 24256
rect 5399 24225 5411 24228
rect 5353 24219 5411 24225
rect 5534 24216 5540 24228
rect 5592 24256 5598 24268
rect 6181 24259 6239 24265
rect 6181 24256 6193 24259
rect 5592 24228 6193 24256
rect 5592 24216 5598 24228
rect 6181 24225 6193 24228
rect 6227 24225 6239 24259
rect 6362 24256 6368 24268
rect 6323 24228 6368 24256
rect 6181 24219 6239 24225
rect 1578 24148 1584 24200
rect 1636 24188 1642 24200
rect 1673 24191 1731 24197
rect 1673 24188 1685 24191
rect 1636 24160 1685 24188
rect 1636 24148 1642 24160
rect 1673 24157 1685 24160
rect 1719 24157 1731 24191
rect 1673 24151 1731 24157
rect 4706 24148 4712 24200
rect 4764 24188 4770 24200
rect 4893 24191 4951 24197
rect 4893 24188 4905 24191
rect 4764 24160 4905 24188
rect 4764 24148 4770 24160
rect 4893 24157 4905 24160
rect 4939 24157 4951 24191
rect 4893 24151 4951 24157
rect 5166 24148 5172 24200
rect 5224 24188 5230 24200
rect 5445 24191 5503 24197
rect 5445 24188 5457 24191
rect 5224 24160 5457 24188
rect 5224 24148 5230 24160
rect 5445 24157 5457 24160
rect 5491 24157 5503 24191
rect 6196 24188 6224 24219
rect 6362 24216 6368 24228
rect 6420 24216 6426 24268
rect 7101 24259 7159 24265
rect 7101 24225 7113 24259
rect 7147 24256 7159 24259
rect 7282 24256 7288 24268
rect 7147 24228 7288 24256
rect 7147 24225 7159 24228
rect 7101 24219 7159 24225
rect 7282 24216 7288 24228
rect 7340 24216 7346 24268
rect 7377 24259 7435 24265
rect 7377 24225 7389 24259
rect 7423 24256 7435 24259
rect 7466 24256 7472 24268
rect 7423 24228 7472 24256
rect 7423 24225 7435 24228
rect 7377 24219 7435 24225
rect 7466 24216 7472 24228
rect 7524 24216 7530 24268
rect 7558 24216 7564 24268
rect 7616 24256 7622 24268
rect 8205 24259 8263 24265
rect 7616 24228 7661 24256
rect 7616 24216 7622 24228
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 8846 24256 8852 24268
rect 8251 24228 8852 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 8846 24216 8852 24228
rect 8904 24216 8910 24268
rect 10042 24256 10048 24268
rect 8956 24228 10048 24256
rect 8956 24197 8984 24228
rect 10042 24216 10048 24228
rect 10100 24216 10106 24268
rect 10226 24256 10232 24268
rect 10187 24228 10232 24256
rect 10226 24216 10232 24228
rect 10284 24216 10290 24268
rect 10321 24259 10379 24265
rect 10321 24225 10333 24259
rect 10367 24225 10379 24259
rect 10505 24259 10563 24265
rect 10505 24256 10517 24259
rect 10321 24219 10379 24225
rect 10428 24228 10517 24256
rect 8941 24191 8999 24197
rect 8941 24188 8953 24191
rect 6196 24160 8953 24188
rect 5445 24151 5503 24157
rect 8941 24157 8953 24160
rect 8987 24157 8999 24191
rect 8941 24151 8999 24157
rect 9858 24148 9864 24200
rect 9916 24188 9922 24200
rect 10336 24188 10364 24219
rect 9916 24160 10364 24188
rect 9916 24148 9922 24160
rect 3418 24080 3424 24132
rect 3476 24120 3482 24132
rect 5813 24123 5871 24129
rect 5813 24120 5825 24123
rect 3476 24092 5825 24120
rect 3476 24080 3482 24092
rect 5813 24089 5825 24092
rect 5859 24120 5871 24123
rect 7190 24120 7196 24132
rect 5859 24092 7196 24120
rect 5859 24089 5871 24092
rect 5813 24083 5871 24089
rect 6380 24064 6408 24092
rect 7190 24080 7196 24092
rect 7248 24120 7254 24132
rect 9309 24123 9367 24129
rect 9309 24120 9321 24123
rect 7248 24092 9321 24120
rect 7248 24080 7254 24092
rect 9309 24089 9321 24092
rect 9355 24089 9367 24123
rect 9309 24083 9367 24089
rect 9766 24080 9772 24132
rect 9824 24120 9830 24132
rect 10428 24120 10456 24228
rect 10505 24225 10517 24228
rect 10551 24225 10563 24259
rect 10505 24219 10563 24225
rect 12529 24259 12587 24265
rect 12529 24225 12541 24259
rect 12575 24256 12587 24259
rect 12912 24256 12940 24284
rect 13906 24256 13912 24268
rect 12575 24228 12940 24256
rect 13867 24228 13912 24256
rect 12575 24225 12587 24228
rect 12529 24219 12587 24225
rect 13906 24216 13912 24228
rect 13964 24216 13970 24268
rect 15120 24256 15148 24364
rect 15289 24327 15347 24333
rect 15289 24293 15301 24327
rect 15335 24324 15347 24327
rect 16206 24324 16212 24336
rect 15335 24296 16212 24324
rect 15335 24293 15347 24296
rect 15289 24287 15347 24293
rect 16206 24284 16212 24296
rect 16264 24284 16270 24336
rect 16592 24324 16620 24364
rect 16669 24361 16681 24395
rect 16715 24392 16727 24395
rect 16758 24392 16764 24404
rect 16715 24364 16764 24392
rect 16715 24361 16727 24364
rect 16669 24355 16727 24361
rect 16758 24352 16764 24364
rect 16816 24352 16822 24404
rect 17037 24395 17095 24401
rect 17037 24361 17049 24395
rect 17083 24392 17095 24395
rect 17494 24392 17500 24404
rect 17083 24364 17500 24392
rect 17083 24361 17095 24364
rect 17037 24355 17095 24361
rect 17494 24352 17500 24364
rect 17552 24352 17558 24404
rect 21177 24395 21235 24401
rect 21177 24361 21189 24395
rect 21223 24392 21235 24395
rect 21358 24392 21364 24404
rect 21223 24364 21364 24392
rect 21223 24361 21235 24364
rect 21177 24355 21235 24361
rect 21358 24352 21364 24364
rect 21416 24352 21422 24404
rect 24026 24392 24032 24404
rect 23987 24364 24032 24392
rect 24026 24352 24032 24364
rect 24084 24352 24090 24404
rect 25041 24395 25099 24401
rect 25041 24361 25053 24395
rect 25087 24392 25099 24395
rect 26234 24392 26240 24404
rect 25087 24364 26240 24392
rect 25087 24361 25099 24364
rect 25041 24355 25099 24361
rect 26234 24352 26240 24364
rect 26292 24352 26298 24404
rect 28258 24392 28264 24404
rect 28219 24364 28264 24392
rect 28258 24352 28264 24364
rect 28316 24392 28322 24404
rect 28316 24364 28764 24392
rect 28316 24352 28322 24364
rect 16942 24324 16948 24336
rect 16592 24296 16948 24324
rect 16942 24284 16948 24296
rect 17000 24324 17006 24336
rect 17313 24327 17371 24333
rect 17313 24324 17325 24327
rect 17000 24296 17325 24324
rect 17000 24284 17006 24296
rect 17313 24293 17325 24296
rect 17359 24324 17371 24327
rect 17402 24324 17408 24336
rect 17359 24296 17408 24324
rect 17359 24293 17371 24296
rect 17313 24287 17371 24293
rect 17402 24284 17408 24296
rect 17460 24284 17466 24336
rect 25958 24324 25964 24336
rect 25919 24296 25964 24324
rect 25958 24284 25964 24296
rect 26016 24284 26022 24336
rect 26878 24324 26884 24336
rect 26839 24296 26884 24324
rect 26878 24284 26884 24296
rect 26936 24284 26942 24336
rect 16114 24256 16120 24268
rect 14292 24228 15148 24256
rect 16075 24228 16120 24256
rect 10870 24188 10876 24200
rect 10831 24160 10876 24188
rect 10870 24148 10876 24160
rect 10928 24148 10934 24200
rect 11054 24188 11060 24200
rect 11015 24160 11060 24188
rect 11054 24148 11060 24160
rect 11112 24148 11118 24200
rect 12434 24148 12440 24200
rect 12492 24188 12498 24200
rect 12986 24188 12992 24200
rect 12492 24160 12537 24188
rect 12947 24160 12992 24188
rect 12492 24148 12498 24160
rect 12986 24148 12992 24160
rect 13044 24148 13050 24200
rect 13817 24191 13875 24197
rect 13817 24157 13829 24191
rect 13863 24188 13875 24191
rect 14090 24188 14096 24200
rect 13863 24160 14096 24188
rect 13863 24157 13875 24160
rect 13817 24151 13875 24157
rect 14090 24148 14096 24160
rect 14148 24188 14154 24200
rect 14292 24188 14320 24228
rect 16114 24216 16120 24228
rect 16172 24216 16178 24268
rect 17034 24216 17040 24268
rect 17092 24256 17098 24268
rect 17678 24256 17684 24268
rect 17092 24228 17684 24256
rect 17092 24216 17098 24228
rect 17678 24216 17684 24228
rect 17736 24256 17742 24268
rect 17865 24259 17923 24265
rect 17865 24256 17877 24259
rect 17736 24228 17877 24256
rect 17736 24216 17742 24228
rect 17865 24225 17877 24228
rect 17911 24225 17923 24259
rect 17865 24219 17923 24225
rect 22649 24259 22707 24265
rect 22649 24225 22661 24259
rect 22695 24256 22707 24259
rect 23198 24256 23204 24268
rect 22695 24228 23204 24256
rect 22695 24225 22707 24228
rect 22649 24219 22707 24225
rect 23198 24216 23204 24228
rect 23256 24216 23262 24268
rect 25409 24259 25467 24265
rect 25409 24225 25421 24259
rect 25455 24256 25467 24259
rect 25498 24256 25504 24268
rect 25455 24228 25504 24256
rect 25455 24225 25467 24228
rect 25409 24219 25467 24225
rect 25498 24216 25504 24228
rect 25556 24216 25562 24268
rect 27246 24256 27252 24268
rect 27207 24228 27252 24256
rect 27246 24216 27252 24228
rect 27304 24216 27310 24268
rect 28442 24256 28448 24268
rect 28403 24228 28448 24256
rect 28442 24216 28448 24228
rect 28500 24216 28506 24268
rect 28736 24265 28764 24364
rect 30926 24352 30932 24404
rect 30984 24392 30990 24404
rect 31205 24395 31263 24401
rect 31205 24392 31217 24395
rect 30984 24364 31217 24392
rect 30984 24352 30990 24364
rect 31205 24361 31217 24364
rect 31251 24361 31263 24395
rect 31205 24355 31263 24361
rect 31386 24352 31392 24404
rect 31444 24392 31450 24404
rect 31481 24395 31539 24401
rect 31481 24392 31493 24395
rect 31444 24364 31493 24392
rect 31444 24352 31450 24364
rect 31481 24361 31493 24364
rect 31527 24361 31539 24395
rect 32306 24392 32312 24404
rect 32267 24364 32312 24392
rect 31481 24355 31539 24361
rect 32306 24352 32312 24364
rect 32364 24352 32370 24404
rect 32582 24392 32588 24404
rect 32543 24364 32588 24392
rect 32582 24352 32588 24364
rect 32640 24352 32646 24404
rect 32950 24392 32956 24404
rect 32911 24364 32956 24392
rect 32950 24352 32956 24364
rect 33008 24352 33014 24404
rect 35802 24392 35808 24404
rect 35763 24364 35808 24392
rect 35802 24352 35808 24364
rect 35860 24352 35866 24404
rect 29178 24284 29184 24336
rect 29236 24324 29242 24336
rect 29638 24324 29644 24336
rect 29236 24296 29644 24324
rect 29236 24284 29242 24296
rect 29638 24284 29644 24296
rect 29696 24284 29702 24336
rect 28721 24259 28779 24265
rect 28721 24225 28733 24259
rect 28767 24225 28779 24259
rect 30006 24256 30012 24268
rect 29967 24228 30012 24256
rect 28721 24219 28779 24225
rect 30006 24216 30012 24228
rect 30064 24216 30070 24268
rect 31018 24256 31024 24268
rect 30931 24228 31024 24256
rect 31018 24216 31024 24228
rect 31076 24256 31082 24268
rect 31478 24256 31484 24268
rect 31076 24228 31484 24256
rect 31076 24216 31082 24228
rect 31478 24216 31484 24228
rect 31536 24216 31542 24268
rect 32125 24259 32183 24265
rect 32125 24225 32137 24259
rect 32171 24256 32183 24259
rect 32214 24256 32220 24268
rect 32171 24228 32220 24256
rect 32171 24225 32183 24228
rect 32125 24219 32183 24225
rect 32214 24216 32220 24228
rect 32272 24256 32278 24268
rect 32674 24256 32680 24268
rect 32272 24228 32680 24256
rect 32272 24216 32278 24228
rect 32674 24216 32680 24228
rect 32732 24216 32738 24268
rect 14148 24160 14320 24188
rect 14369 24191 14427 24197
rect 14148 24148 14154 24160
rect 14369 24157 14381 24191
rect 14415 24157 14427 24191
rect 14369 24151 14427 24157
rect 12342 24120 12348 24132
rect 9824 24092 10456 24120
rect 12303 24092 12348 24120
rect 9824 24080 9830 24092
rect 12342 24080 12348 24092
rect 12400 24080 12406 24132
rect 13538 24080 13544 24132
rect 13596 24080 13602 24132
rect 13722 24120 13728 24132
rect 13683 24092 13728 24120
rect 13722 24080 13728 24092
rect 13780 24080 13786 24132
rect 14384 24120 14412 24151
rect 15470 24148 15476 24200
rect 15528 24188 15534 24200
rect 15841 24191 15899 24197
rect 15841 24188 15853 24191
rect 15528 24160 15853 24188
rect 15528 24148 15534 24160
rect 15841 24157 15853 24160
rect 15887 24157 15899 24191
rect 15841 24151 15899 24157
rect 16301 24191 16359 24197
rect 16301 24157 16313 24191
rect 16347 24157 16359 24191
rect 16301 24151 16359 24157
rect 17589 24191 17647 24197
rect 17589 24157 17601 24191
rect 17635 24188 17647 24191
rect 17954 24188 17960 24200
rect 17635 24160 17960 24188
rect 17635 24157 17647 24160
rect 17589 24151 17647 24157
rect 15105 24123 15163 24129
rect 15105 24120 15117 24123
rect 14384 24092 15117 24120
rect 15105 24089 15117 24092
rect 15151 24120 15163 24123
rect 16316 24120 16344 24151
rect 17954 24148 17960 24160
rect 18012 24188 18018 24200
rect 18230 24188 18236 24200
rect 18012 24160 18236 24188
rect 18012 24148 18018 24160
rect 18230 24148 18236 24160
rect 18288 24148 18294 24200
rect 21082 24148 21088 24200
rect 21140 24188 21146 24200
rect 21453 24191 21511 24197
rect 21453 24188 21465 24191
rect 21140 24160 21465 24188
rect 21140 24148 21146 24160
rect 21453 24157 21465 24160
rect 21499 24157 21511 24191
rect 22922 24188 22928 24200
rect 22883 24160 22928 24188
rect 21453 24151 21511 24157
rect 22922 24148 22928 24160
rect 22980 24148 22986 24200
rect 27706 24148 27712 24200
rect 27764 24188 27770 24200
rect 28537 24191 28595 24197
rect 28537 24188 28549 24191
rect 27764 24160 28549 24188
rect 27764 24148 27770 24160
rect 28537 24157 28549 24160
rect 28583 24157 28595 24191
rect 29178 24188 29184 24200
rect 29139 24160 29184 24188
rect 28537 24151 28595 24157
rect 15151 24092 16344 24120
rect 20625 24123 20683 24129
rect 15151 24089 15163 24092
rect 15105 24083 15163 24089
rect 20625 24089 20637 24123
rect 20671 24120 20683 24123
rect 21542 24120 21548 24132
rect 20671 24092 21548 24120
rect 20671 24089 20683 24092
rect 20625 24083 20683 24089
rect 21542 24080 21548 24092
rect 21600 24080 21606 24132
rect 25593 24123 25651 24129
rect 25593 24089 25605 24123
rect 25639 24120 25651 24123
rect 26050 24120 26056 24132
rect 25639 24092 26056 24120
rect 25639 24089 25651 24092
rect 25593 24083 25651 24089
rect 26050 24080 26056 24092
rect 26108 24080 26114 24132
rect 3878 24052 3884 24064
rect 3839 24024 3884 24052
rect 3878 24012 3884 24024
rect 3936 24012 3942 24064
rect 6362 24012 6368 24064
rect 6420 24012 6426 24064
rect 8662 24052 8668 24064
rect 8623 24024 8668 24052
rect 8662 24012 8668 24024
rect 8720 24012 8726 24064
rect 11517 24055 11575 24061
rect 11517 24021 11529 24055
rect 11563 24052 11575 24055
rect 11606 24052 11612 24064
rect 11563 24024 11612 24052
rect 11563 24021 11575 24024
rect 11517 24015 11575 24021
rect 11606 24012 11612 24024
rect 11664 24052 11670 24064
rect 12158 24052 12164 24064
rect 11664 24024 12164 24052
rect 11664 24012 11670 24024
rect 12158 24012 12164 24024
rect 12216 24012 12222 24064
rect 12250 24012 12256 24064
rect 12308 24052 12314 24064
rect 13357 24055 13415 24061
rect 13357 24052 13369 24055
rect 12308 24024 13369 24052
rect 12308 24012 12314 24024
rect 13357 24021 13369 24024
rect 13403 24052 13415 24055
rect 13556 24052 13584 24080
rect 14366 24052 14372 24064
rect 13403 24024 14372 24052
rect 13403 24021 13415 24024
rect 13357 24015 13415 24021
rect 14366 24012 14372 24024
rect 14424 24012 14430 24064
rect 18690 24012 18696 24064
rect 18748 24052 18754 24064
rect 18969 24055 19027 24061
rect 18969 24052 18981 24055
rect 18748 24024 18981 24052
rect 18748 24012 18754 24024
rect 18969 24021 18981 24024
rect 19015 24021 19027 24055
rect 18969 24015 19027 24021
rect 19886 24012 19892 24064
rect 19944 24052 19950 24064
rect 19981 24055 20039 24061
rect 19981 24052 19993 24055
rect 19944 24024 19993 24052
rect 19944 24012 19950 24024
rect 19981 24021 19993 24024
rect 20027 24052 20039 24055
rect 20162 24052 20168 24064
rect 20027 24024 20168 24052
rect 20027 24021 20039 24024
rect 19981 24015 20039 24021
rect 20162 24012 20168 24024
rect 20220 24012 20226 24064
rect 27614 24012 27620 24064
rect 27672 24052 27678 24064
rect 27893 24055 27951 24061
rect 27893 24052 27905 24055
rect 27672 24024 27905 24052
rect 27672 24012 27678 24024
rect 27893 24021 27905 24024
rect 27939 24021 27951 24055
rect 28552 24052 28580 24151
rect 29178 24148 29184 24160
rect 29236 24148 29242 24200
rect 29270 24080 29276 24132
rect 29328 24120 29334 24132
rect 30193 24123 30251 24129
rect 30193 24120 30205 24123
rect 29328 24092 30205 24120
rect 29328 24080 29334 24092
rect 30193 24089 30205 24092
rect 30239 24120 30251 24123
rect 31570 24120 31576 24132
rect 30239 24092 31576 24120
rect 30239 24089 30251 24092
rect 30193 24083 30251 24089
rect 31570 24080 31576 24092
rect 31628 24080 31634 24132
rect 29362 24052 29368 24064
rect 28552 24024 29368 24052
rect 27893 24015 27951 24021
rect 29362 24012 29368 24024
rect 29420 24012 29426 24064
rect 29546 24052 29552 24064
rect 29507 24024 29552 24052
rect 29546 24012 29552 24024
rect 29604 24012 29610 24064
rect 30558 24012 30564 24064
rect 30616 24052 30622 24064
rect 30745 24055 30803 24061
rect 30745 24052 30757 24055
rect 30616 24024 30757 24052
rect 30616 24012 30622 24024
rect 30745 24021 30757 24024
rect 30791 24052 30803 24055
rect 30834 24052 30840 24064
rect 30791 24024 30840 24052
rect 30791 24021 30803 24024
rect 30745 24015 30803 24021
rect 30834 24012 30840 24024
rect 30892 24012 30898 24064
rect 1104 23962 38548 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 38548 23962
rect 1104 23888 38548 23910
rect 1578 23848 1584 23860
rect 1539 23820 1584 23848
rect 1578 23808 1584 23820
rect 1636 23808 1642 23860
rect 3786 23848 3792 23860
rect 3747 23820 3792 23848
rect 3786 23808 3792 23820
rect 3844 23808 3850 23860
rect 4706 23808 4712 23860
rect 4764 23848 4770 23860
rect 5169 23851 5227 23857
rect 5169 23848 5181 23851
rect 4764 23820 5181 23848
rect 4764 23808 4770 23820
rect 5169 23817 5181 23820
rect 5215 23817 5227 23851
rect 5169 23811 5227 23817
rect 5905 23851 5963 23857
rect 5905 23817 5917 23851
rect 5951 23817 5963 23851
rect 9766 23848 9772 23860
rect 9727 23820 9772 23848
rect 5905 23811 5963 23817
rect 1394 23740 1400 23792
rect 1452 23780 1458 23792
rect 1949 23783 2007 23789
rect 1949 23780 1961 23783
rect 1452 23752 1961 23780
rect 1452 23740 1458 23752
rect 1949 23749 1961 23752
rect 1995 23780 2007 23783
rect 2317 23783 2375 23789
rect 2317 23780 2329 23783
rect 1995 23752 2329 23780
rect 1995 23749 2007 23752
rect 1949 23743 2007 23749
rect 2317 23749 2329 23752
rect 2363 23749 2375 23783
rect 2317 23743 2375 23749
rect 4893 23783 4951 23789
rect 4893 23749 4905 23783
rect 4939 23780 4951 23783
rect 5534 23780 5540 23792
rect 4939 23752 5540 23780
rect 4939 23749 4951 23752
rect 4893 23743 4951 23749
rect 5534 23740 5540 23752
rect 5592 23780 5598 23792
rect 5920 23780 5948 23811
rect 9766 23808 9772 23820
rect 9824 23808 9830 23860
rect 10137 23851 10195 23857
rect 10137 23817 10149 23851
rect 10183 23848 10195 23851
rect 11054 23848 11060 23860
rect 10183 23820 11060 23848
rect 10183 23817 10195 23820
rect 10137 23811 10195 23817
rect 11054 23808 11060 23820
rect 11112 23808 11118 23860
rect 11422 23808 11428 23860
rect 11480 23848 11486 23860
rect 12161 23851 12219 23857
rect 12161 23848 12173 23851
rect 11480 23820 12173 23848
rect 11480 23808 11486 23820
rect 12161 23817 12173 23820
rect 12207 23848 12219 23851
rect 12434 23848 12440 23860
rect 12207 23820 12440 23848
rect 12207 23817 12219 23820
rect 12161 23811 12219 23817
rect 12434 23808 12440 23820
rect 12492 23808 12498 23860
rect 12710 23848 12716 23860
rect 12671 23820 12716 23848
rect 12710 23808 12716 23820
rect 12768 23848 12774 23860
rect 13998 23848 14004 23860
rect 12768 23820 14004 23848
rect 12768 23808 12774 23820
rect 13998 23808 14004 23820
rect 14056 23808 14062 23860
rect 15289 23851 15347 23857
rect 15289 23817 15301 23851
rect 15335 23848 15347 23851
rect 15930 23848 15936 23860
rect 15335 23820 15936 23848
rect 15335 23817 15347 23820
rect 15289 23811 15347 23817
rect 15930 23808 15936 23820
rect 15988 23808 15994 23860
rect 17402 23848 17408 23860
rect 17363 23820 17408 23848
rect 17402 23808 17408 23820
rect 17460 23808 17466 23860
rect 18874 23848 18880 23860
rect 18835 23820 18880 23848
rect 18874 23808 18880 23820
rect 18932 23808 18938 23860
rect 20254 23808 20260 23860
rect 20312 23848 20318 23860
rect 20349 23851 20407 23857
rect 20349 23848 20361 23851
rect 20312 23820 20361 23848
rect 20312 23808 20318 23820
rect 20349 23817 20361 23820
rect 20395 23817 20407 23851
rect 20349 23811 20407 23817
rect 23109 23851 23167 23857
rect 23109 23817 23121 23851
rect 23155 23848 23167 23851
rect 23198 23848 23204 23860
rect 23155 23820 23204 23848
rect 23155 23817 23167 23820
rect 23109 23811 23167 23817
rect 5592 23752 6868 23780
rect 5592 23740 5598 23752
rect 3418 23712 3424 23724
rect 3379 23684 3424 23712
rect 3418 23672 3424 23684
rect 3476 23672 3482 23724
rect 5902 23672 5908 23724
rect 5960 23712 5966 23724
rect 6840 23721 6868 23752
rect 13906 23740 13912 23792
rect 13964 23780 13970 23792
rect 14369 23783 14427 23789
rect 14369 23780 14381 23783
rect 13964 23752 14381 23780
rect 13964 23740 13970 23752
rect 14369 23749 14381 23752
rect 14415 23780 14427 23783
rect 15378 23780 15384 23792
rect 14415 23752 15384 23780
rect 14415 23749 14427 23752
rect 14369 23743 14427 23749
rect 15378 23740 15384 23752
rect 15436 23740 15442 23792
rect 6825 23715 6883 23721
rect 5960 23684 6684 23712
rect 5960 23672 5966 23684
rect 5721 23647 5779 23653
rect 5721 23613 5733 23647
rect 5767 23644 5779 23647
rect 6178 23644 6184 23656
rect 5767 23616 6184 23644
rect 5767 23613 5779 23616
rect 5721 23607 5779 23613
rect 6178 23604 6184 23616
rect 6236 23604 6242 23656
rect 6656 23653 6684 23684
rect 6825 23681 6837 23715
rect 6871 23681 6883 23715
rect 7558 23712 7564 23724
rect 7519 23684 7564 23712
rect 6825 23675 6883 23681
rect 7558 23672 7564 23684
rect 7616 23672 7622 23724
rect 10594 23672 10600 23724
rect 10652 23712 10658 23724
rect 11514 23712 11520 23724
rect 10652 23684 11100 23712
rect 11475 23684 11520 23712
rect 10652 23672 10658 23684
rect 6641 23647 6699 23653
rect 6641 23613 6653 23647
rect 6687 23644 6699 23647
rect 7101 23647 7159 23653
rect 7101 23644 7113 23647
rect 6687 23616 7113 23644
rect 6687 23613 6699 23616
rect 6641 23607 6699 23613
rect 7101 23613 7113 23616
rect 7147 23644 7159 23647
rect 7466 23644 7472 23656
rect 7147 23616 7472 23644
rect 7147 23613 7159 23616
rect 7101 23607 7159 23613
rect 7466 23604 7472 23616
rect 7524 23644 7530 23656
rect 8662 23644 8668 23656
rect 7524 23616 8668 23644
rect 7524 23604 7530 23616
rect 8662 23604 8668 23616
rect 8720 23644 8726 23656
rect 8849 23647 8907 23653
rect 8849 23644 8861 23647
rect 8720 23616 8861 23644
rect 8720 23604 8726 23616
rect 8849 23613 8861 23616
rect 8895 23613 8907 23647
rect 8849 23607 8907 23613
rect 9674 23604 9680 23656
rect 9732 23604 9738 23656
rect 10689 23647 10747 23653
rect 10689 23613 10701 23647
rect 10735 23644 10747 23647
rect 10778 23644 10784 23656
rect 10735 23616 10784 23644
rect 10735 23613 10747 23616
rect 10689 23607 10747 23613
rect 10778 23604 10784 23616
rect 10836 23604 10842 23656
rect 11072 23653 11100 23684
rect 11514 23672 11520 23684
rect 11572 23672 11578 23724
rect 14826 23712 14832 23724
rect 13924 23684 14832 23712
rect 11057 23647 11115 23653
rect 11057 23613 11069 23647
rect 11103 23644 11115 23647
rect 11330 23644 11336 23656
rect 11103 23616 11336 23644
rect 11103 23613 11115 23616
rect 11057 23607 11115 23613
rect 11330 23604 11336 23616
rect 11388 23604 11394 23656
rect 12342 23604 12348 23656
rect 12400 23644 12406 23656
rect 13541 23647 13599 23653
rect 13541 23644 13553 23647
rect 12400 23616 13553 23644
rect 12400 23604 12406 23616
rect 13541 23613 13553 23616
rect 13587 23613 13599 23647
rect 13541 23607 13599 23613
rect 13633 23647 13691 23653
rect 13633 23613 13645 23647
rect 13679 23613 13691 23647
rect 13633 23607 13691 23613
rect 3050 23576 3056 23588
rect 3011 23548 3056 23576
rect 3050 23536 3056 23548
rect 3108 23536 3114 23588
rect 4525 23579 4583 23585
rect 4525 23545 4537 23579
rect 4571 23576 4583 23579
rect 4798 23576 4804 23588
rect 4571 23548 4804 23576
rect 4571 23545 4583 23548
rect 4525 23539 4583 23545
rect 4798 23536 4804 23548
rect 4856 23536 4862 23588
rect 5629 23579 5687 23585
rect 5629 23545 5641 23579
rect 5675 23576 5687 23579
rect 7190 23576 7196 23588
rect 5675 23548 6500 23576
rect 7151 23548 7196 23576
rect 5675 23545 5687 23548
rect 5629 23539 5687 23545
rect 6472 23520 6500 23548
rect 7190 23536 7196 23548
rect 7248 23536 7254 23588
rect 8573 23579 8631 23585
rect 8573 23576 8585 23579
rect 8036 23548 8585 23576
rect 8036 23520 8064 23548
rect 8573 23545 8585 23548
rect 8619 23545 8631 23579
rect 8938 23576 8944 23588
rect 8899 23548 8944 23576
rect 8573 23539 8631 23545
rect 8938 23536 8944 23548
rect 8996 23536 9002 23588
rect 9309 23579 9367 23585
rect 9309 23545 9321 23579
rect 9355 23576 9367 23579
rect 9582 23576 9588 23588
rect 9355 23548 9588 23576
rect 9355 23545 9367 23548
rect 9309 23539 9367 23545
rect 9582 23536 9588 23548
rect 9640 23536 9646 23588
rect 9692 23576 9720 23604
rect 10965 23579 11023 23585
rect 10965 23576 10977 23579
rect 9692 23548 10977 23576
rect 10965 23545 10977 23548
rect 11011 23576 11023 23579
rect 11238 23576 11244 23588
rect 11011 23548 11244 23576
rect 11011 23545 11023 23548
rect 10965 23539 11023 23545
rect 11238 23536 11244 23548
rect 11296 23536 11302 23588
rect 12897 23579 12955 23585
rect 12897 23545 12909 23579
rect 12943 23576 12955 23579
rect 13354 23576 13360 23588
rect 12943 23548 13360 23576
rect 12943 23545 12955 23548
rect 12897 23539 12955 23545
rect 13354 23536 13360 23548
rect 13412 23536 13418 23588
rect 13648 23576 13676 23607
rect 13814 23604 13820 23656
rect 13872 23644 13878 23656
rect 13924 23653 13952 23684
rect 14826 23672 14832 23684
rect 14884 23672 14890 23724
rect 16574 23672 16580 23724
rect 16632 23712 16638 23724
rect 17129 23715 17187 23721
rect 17129 23712 17141 23715
rect 16632 23684 17141 23712
rect 16632 23672 16638 23684
rect 17129 23681 17141 23684
rect 17175 23712 17187 23715
rect 17773 23715 17831 23721
rect 17773 23712 17785 23715
rect 17175 23684 17785 23712
rect 17175 23681 17187 23684
rect 17129 23675 17187 23681
rect 17773 23681 17785 23684
rect 17819 23681 17831 23715
rect 17773 23675 17831 23681
rect 18509 23715 18567 23721
rect 18509 23681 18521 23715
rect 18555 23712 18567 23715
rect 20364 23712 20392 23811
rect 23198 23808 23204 23820
rect 23256 23808 23262 23860
rect 25866 23848 25872 23860
rect 25827 23820 25872 23848
rect 25866 23808 25872 23820
rect 25924 23808 25930 23860
rect 27157 23851 27215 23857
rect 27157 23848 27169 23851
rect 26804 23820 27169 23848
rect 24854 23780 24860 23792
rect 24815 23752 24860 23780
rect 24854 23740 24860 23752
rect 24912 23740 24918 23792
rect 25225 23783 25283 23789
rect 25225 23749 25237 23783
rect 25271 23780 25283 23783
rect 26804 23780 26832 23820
rect 27157 23817 27169 23820
rect 27203 23848 27215 23851
rect 27246 23848 27252 23860
rect 27203 23820 27252 23848
rect 27203 23817 27215 23820
rect 27157 23811 27215 23817
rect 27246 23808 27252 23820
rect 27304 23808 27310 23860
rect 28442 23808 28448 23860
rect 28500 23848 28506 23860
rect 28629 23851 28687 23857
rect 28629 23848 28641 23851
rect 28500 23820 28641 23848
rect 28500 23808 28506 23820
rect 28629 23817 28641 23820
rect 28675 23848 28687 23851
rect 29454 23848 29460 23860
rect 28675 23820 29460 23848
rect 28675 23817 28687 23820
rect 28629 23811 28687 23817
rect 29454 23808 29460 23820
rect 29512 23808 29518 23860
rect 30006 23808 30012 23860
rect 30064 23848 30070 23860
rect 30377 23851 30435 23857
rect 30377 23848 30389 23851
rect 30064 23820 30389 23848
rect 30064 23808 30070 23820
rect 30377 23817 30389 23820
rect 30423 23817 30435 23851
rect 30377 23811 30435 23817
rect 25271 23752 26832 23780
rect 25271 23749 25283 23752
rect 25225 23743 25283 23749
rect 26878 23740 26884 23792
rect 26936 23780 26942 23792
rect 27709 23783 27767 23789
rect 27709 23780 27721 23783
rect 26936 23752 27721 23780
rect 26936 23740 26942 23752
rect 27709 23749 27721 23752
rect 27755 23780 27767 23783
rect 27890 23780 27896 23792
rect 27755 23752 27896 23780
rect 27755 23749 27767 23752
rect 27709 23743 27767 23749
rect 27890 23740 27896 23752
rect 27948 23740 27954 23792
rect 21453 23715 21511 23721
rect 21453 23712 21465 23715
rect 18555 23684 18736 23712
rect 20364 23684 21465 23712
rect 18555 23681 18567 23684
rect 18509 23675 18567 23681
rect 18708 23656 18736 23684
rect 21453 23681 21465 23684
rect 21499 23712 21511 23715
rect 21726 23712 21732 23724
rect 21499 23684 21732 23712
rect 21499 23681 21511 23684
rect 21453 23675 21511 23681
rect 21726 23672 21732 23684
rect 21784 23672 21790 23724
rect 13909 23647 13967 23653
rect 13909 23644 13921 23647
rect 13872 23616 13921 23644
rect 13872 23604 13878 23616
rect 13909 23613 13921 23616
rect 13955 23613 13967 23647
rect 13909 23607 13967 23613
rect 13998 23604 14004 23656
rect 14056 23644 14062 23656
rect 14056 23616 14101 23644
rect 14056 23604 14062 23616
rect 14366 23604 14372 23656
rect 14424 23644 14430 23656
rect 15105 23647 15163 23653
rect 15105 23644 15117 23647
rect 14424 23616 15117 23644
rect 14424 23604 14430 23616
rect 15105 23613 15117 23616
rect 15151 23644 15163 23647
rect 15565 23647 15623 23653
rect 15565 23644 15577 23647
rect 15151 23616 15577 23644
rect 15151 23613 15163 23616
rect 15105 23607 15163 23613
rect 15565 23613 15577 23616
rect 15611 23613 15623 23647
rect 15565 23607 15623 23613
rect 16669 23647 16727 23653
rect 16669 23613 16681 23647
rect 16715 23644 16727 23647
rect 16758 23644 16764 23656
rect 16715 23616 16764 23644
rect 16715 23613 16727 23616
rect 16669 23607 16727 23613
rect 16758 23604 16764 23616
rect 16816 23604 16822 23656
rect 16945 23647 17003 23653
rect 16945 23613 16957 23647
rect 16991 23613 17003 23647
rect 18598 23644 18604 23656
rect 18559 23616 18604 23644
rect 16945 23607 17003 23613
rect 13722 23576 13728 23588
rect 13635 23548 13728 23576
rect 13722 23536 13728 23548
rect 13780 23576 13786 23588
rect 15013 23579 15071 23585
rect 15013 23576 15025 23579
rect 13780 23548 15025 23576
rect 13780 23536 13786 23548
rect 15013 23545 15025 23548
rect 15059 23576 15071 23579
rect 15470 23576 15476 23588
rect 15059 23548 15476 23576
rect 15059 23545 15071 23548
rect 15013 23539 15071 23545
rect 15470 23536 15476 23548
rect 15528 23536 15534 23588
rect 16114 23576 16120 23588
rect 16075 23548 16120 23576
rect 16114 23536 16120 23548
rect 16172 23536 16178 23588
rect 4157 23511 4215 23517
rect 4157 23477 4169 23511
rect 4203 23508 4215 23511
rect 5258 23508 5264 23520
rect 4203 23480 5264 23508
rect 4203 23477 4215 23480
rect 4157 23471 4215 23477
rect 5258 23468 5264 23480
rect 5316 23468 5322 23520
rect 6454 23468 6460 23520
rect 6512 23508 6518 23520
rect 7009 23511 7067 23517
rect 7009 23508 7021 23511
rect 6512 23480 7021 23508
rect 6512 23468 6518 23480
rect 7009 23477 7021 23480
rect 7055 23508 7067 23511
rect 7098 23508 7104 23520
rect 7055 23480 7104 23508
rect 7055 23477 7067 23480
rect 7009 23471 7067 23477
rect 7098 23468 7104 23480
rect 7156 23468 7162 23520
rect 8018 23508 8024 23520
rect 7979 23480 8024 23508
rect 8018 23468 8024 23480
rect 8076 23468 8082 23520
rect 8386 23508 8392 23520
rect 8347 23480 8392 23508
rect 8386 23468 8392 23480
rect 8444 23508 8450 23520
rect 8757 23511 8815 23517
rect 8757 23508 8769 23511
rect 8444 23480 8769 23508
rect 8444 23468 8450 23480
rect 8757 23477 8769 23480
rect 8803 23477 8815 23511
rect 8757 23471 8815 23477
rect 11054 23468 11060 23520
rect 11112 23508 11118 23520
rect 11793 23511 11851 23517
rect 11793 23508 11805 23511
rect 11112 23480 11805 23508
rect 11112 23468 11118 23480
rect 11793 23477 11805 23480
rect 11839 23477 11851 23511
rect 11793 23471 11851 23477
rect 15102 23468 15108 23520
rect 15160 23508 15166 23520
rect 16025 23511 16083 23517
rect 16025 23508 16037 23511
rect 15160 23480 16037 23508
rect 15160 23468 15166 23480
rect 16025 23477 16037 23480
rect 16071 23508 16083 23511
rect 16960 23508 16988 23607
rect 18598 23604 18604 23616
rect 18656 23604 18662 23656
rect 18690 23604 18696 23656
rect 18748 23644 18754 23656
rect 20993 23647 21051 23653
rect 20993 23644 21005 23647
rect 18748 23616 18793 23644
rect 19996 23616 21005 23644
rect 18748 23604 18754 23616
rect 18616 23576 18644 23604
rect 19429 23579 19487 23585
rect 19429 23576 19441 23579
rect 18616 23548 19441 23576
rect 19429 23545 19441 23548
rect 19475 23545 19487 23579
rect 19429 23539 19487 23545
rect 19886 23536 19892 23588
rect 19944 23576 19950 23588
rect 19996 23585 20024 23616
rect 20993 23613 21005 23616
rect 21039 23613 21051 23647
rect 20993 23607 21051 23613
rect 21082 23604 21088 23656
rect 21140 23644 21146 23656
rect 21177 23647 21235 23653
rect 21177 23644 21189 23647
rect 21140 23616 21189 23644
rect 21140 23604 21146 23616
rect 21177 23613 21189 23616
rect 21223 23613 21235 23647
rect 21542 23644 21548 23656
rect 21503 23616 21548 23644
rect 21177 23607 21235 23613
rect 21542 23604 21548 23616
rect 21600 23604 21606 23656
rect 24872 23644 24900 23740
rect 29086 23712 29092 23724
rect 27448 23684 27936 23712
rect 28999 23684 29092 23712
rect 25041 23647 25099 23653
rect 25041 23644 25053 23647
rect 24872 23616 25053 23644
rect 25041 23613 25053 23616
rect 25087 23613 25099 23647
rect 25041 23607 25099 23613
rect 25866 23604 25872 23656
rect 25924 23644 25930 23656
rect 27448 23653 27476 23684
rect 26145 23647 26203 23653
rect 26145 23644 26157 23647
rect 25924 23616 26157 23644
rect 25924 23604 25930 23616
rect 26145 23613 26157 23616
rect 26191 23644 26203 23647
rect 27433 23647 27491 23653
rect 27433 23644 27445 23647
rect 26191 23616 27445 23644
rect 26191 23613 26203 23616
rect 26145 23607 26203 23613
rect 27433 23613 27445 23616
rect 27479 23613 27491 23647
rect 27614 23644 27620 23656
rect 27575 23616 27620 23644
rect 27433 23607 27491 23613
rect 27614 23604 27620 23616
rect 27672 23604 27678 23656
rect 27908 23653 27936 23684
rect 29086 23672 29092 23684
rect 29144 23712 29150 23724
rect 30101 23715 30159 23721
rect 29144 23684 29684 23712
rect 29144 23672 29150 23684
rect 27893 23647 27951 23653
rect 27893 23613 27905 23647
rect 27939 23613 27951 23647
rect 29546 23644 29552 23656
rect 29459 23616 29552 23644
rect 27893 23607 27951 23613
rect 29546 23604 29552 23616
rect 29604 23604 29610 23656
rect 29656 23653 29684 23684
rect 30101 23681 30113 23715
rect 30147 23712 30159 23715
rect 30926 23712 30932 23724
rect 30147 23684 30932 23712
rect 30147 23681 30159 23684
rect 30101 23675 30159 23681
rect 30926 23672 30932 23684
rect 30984 23672 30990 23724
rect 31110 23712 31116 23724
rect 31071 23684 31116 23712
rect 31110 23672 31116 23684
rect 31168 23672 31174 23724
rect 35713 23715 35771 23721
rect 35713 23681 35725 23715
rect 35759 23712 35771 23715
rect 36078 23712 36084 23724
rect 35759 23684 36084 23712
rect 35759 23681 35771 23684
rect 35713 23675 35771 23681
rect 36078 23672 36084 23684
rect 36136 23672 36142 23724
rect 29641 23647 29699 23653
rect 29641 23613 29653 23647
rect 29687 23613 29699 23647
rect 29641 23607 29699 23613
rect 30837 23647 30895 23653
rect 30837 23613 30849 23647
rect 30883 23644 30895 23647
rect 31481 23647 31539 23653
rect 31481 23644 31493 23647
rect 30883 23616 31493 23644
rect 30883 23613 30895 23616
rect 30837 23607 30895 23613
rect 31481 23613 31493 23616
rect 31527 23644 31539 23647
rect 31570 23644 31576 23656
rect 31527 23616 31576 23644
rect 31527 23613 31539 23616
rect 31481 23607 31539 23613
rect 31570 23604 31576 23616
rect 31628 23604 31634 23656
rect 31754 23604 31760 23656
rect 31812 23644 31818 23656
rect 35802 23644 35808 23656
rect 31812 23616 31857 23644
rect 35763 23616 35808 23644
rect 31812 23604 31818 23616
rect 35802 23604 35808 23616
rect 35860 23604 35866 23656
rect 19981 23579 20039 23585
rect 19981 23576 19993 23579
rect 19944 23548 19993 23576
rect 19944 23536 19950 23548
rect 19981 23545 19993 23548
rect 20027 23545 20039 23579
rect 19981 23539 20039 23545
rect 22741 23579 22799 23585
rect 22741 23545 22753 23579
rect 22787 23576 22799 23579
rect 22922 23576 22928 23588
rect 22787 23548 22928 23576
rect 22787 23545 22799 23548
rect 22741 23539 22799 23545
rect 22922 23536 22928 23548
rect 22980 23576 22986 23588
rect 23382 23576 23388 23588
rect 22980 23548 23388 23576
rect 22980 23536 22986 23548
rect 23382 23536 23388 23548
rect 23440 23536 23446 23588
rect 26789 23579 26847 23585
rect 26789 23545 26801 23579
rect 26835 23576 26847 23579
rect 26878 23576 26884 23588
rect 26835 23548 26884 23576
rect 26835 23545 26847 23548
rect 26789 23539 26847 23545
rect 26878 23536 26884 23548
rect 26936 23536 26942 23588
rect 28353 23579 28411 23585
rect 28353 23545 28365 23579
rect 28399 23576 28411 23579
rect 28810 23576 28816 23588
rect 28399 23548 28816 23576
rect 28399 23545 28411 23548
rect 28353 23539 28411 23545
rect 28810 23536 28816 23548
rect 28868 23576 28874 23588
rect 29564 23576 29592 23604
rect 28868 23548 29592 23576
rect 32033 23579 32091 23585
rect 28868 23536 28874 23548
rect 32033 23545 32045 23579
rect 32079 23576 32091 23579
rect 32858 23576 32864 23588
rect 32079 23548 32864 23576
rect 32079 23545 32091 23548
rect 32033 23539 32091 23545
rect 32858 23536 32864 23548
rect 32916 23536 32922 23588
rect 16071 23480 16988 23508
rect 20809 23511 20867 23517
rect 16071 23477 16083 23480
rect 16025 23471 16083 23477
rect 20809 23477 20821 23511
rect 20855 23508 20867 23511
rect 25314 23508 25320 23520
rect 20855 23480 25320 23508
rect 20855 23477 20867 23480
rect 20809 23471 20867 23477
rect 25314 23468 25320 23480
rect 25372 23468 25378 23520
rect 25498 23508 25504 23520
rect 25459 23480 25504 23508
rect 25498 23468 25504 23480
rect 25556 23468 25562 23520
rect 32401 23511 32459 23517
rect 32401 23477 32413 23511
rect 32447 23508 32459 23511
rect 32674 23508 32680 23520
rect 32447 23480 32680 23508
rect 32447 23477 32459 23480
rect 32401 23471 32459 23477
rect 32674 23468 32680 23480
rect 32732 23468 32738 23520
rect 37366 23508 37372 23520
rect 37327 23480 37372 23508
rect 37366 23468 37372 23480
rect 37424 23468 37430 23520
rect 1104 23418 38548 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 38548 23418
rect 1104 23344 38548 23366
rect 3878 23304 3884 23316
rect 3839 23276 3884 23304
rect 3878 23264 3884 23276
rect 3936 23264 3942 23316
rect 6089 23307 6147 23313
rect 6089 23273 6101 23307
rect 6135 23304 6147 23307
rect 6454 23304 6460 23316
rect 6135 23276 6460 23304
rect 6135 23273 6147 23276
rect 6089 23267 6147 23273
rect 6454 23264 6460 23276
rect 6512 23264 6518 23316
rect 8294 23264 8300 23316
rect 8352 23304 8358 23316
rect 9033 23307 9091 23313
rect 9033 23304 9045 23307
rect 8352 23276 9045 23304
rect 8352 23264 8358 23276
rect 9033 23273 9045 23276
rect 9079 23273 9091 23307
rect 9858 23304 9864 23316
rect 9819 23276 9864 23304
rect 9033 23267 9091 23273
rect 9858 23264 9864 23276
rect 9916 23304 9922 23316
rect 10137 23307 10195 23313
rect 10137 23304 10149 23307
rect 9916 23276 10149 23304
rect 9916 23264 9922 23276
rect 10137 23273 10149 23276
rect 10183 23273 10195 23307
rect 10137 23267 10195 23273
rect 10226 23264 10232 23316
rect 10284 23304 10290 23316
rect 10505 23307 10563 23313
rect 10505 23304 10517 23307
rect 10284 23276 10517 23304
rect 10284 23264 10290 23276
rect 10505 23273 10517 23276
rect 10551 23273 10563 23307
rect 14642 23304 14648 23316
rect 14603 23276 14648 23304
rect 10505 23267 10563 23273
rect 14642 23264 14648 23276
rect 14700 23264 14706 23316
rect 15654 23304 15660 23316
rect 15615 23276 15660 23304
rect 15654 23264 15660 23276
rect 15712 23264 15718 23316
rect 16758 23264 16764 23316
rect 16816 23304 16822 23316
rect 16853 23307 16911 23313
rect 16853 23304 16865 23307
rect 16816 23276 16865 23304
rect 16816 23264 16822 23276
rect 16853 23273 16865 23276
rect 16899 23304 16911 23307
rect 17034 23304 17040 23316
rect 16899 23276 17040 23304
rect 16899 23273 16911 23276
rect 16853 23267 16911 23273
rect 17034 23264 17040 23276
rect 17092 23264 17098 23316
rect 17678 23304 17684 23316
rect 17639 23276 17684 23304
rect 17678 23264 17684 23276
rect 17736 23304 17742 23316
rect 21085 23307 21143 23313
rect 17736 23276 19104 23304
rect 17736 23264 17742 23276
rect 6178 23196 6184 23248
rect 6236 23236 6242 23248
rect 6273 23239 6331 23245
rect 6273 23236 6285 23239
rect 6236 23208 6285 23236
rect 6236 23196 6242 23208
rect 6273 23205 6285 23208
rect 6319 23205 6331 23239
rect 6638 23236 6644 23248
rect 6599 23208 6644 23236
rect 6273 23199 6331 23205
rect 6638 23196 6644 23208
rect 6696 23196 6702 23248
rect 7006 23236 7012 23248
rect 6967 23208 7012 23236
rect 7006 23196 7012 23208
rect 7064 23196 7070 23248
rect 7558 23196 7564 23248
rect 7616 23236 7622 23248
rect 8389 23239 8447 23245
rect 7616 23208 8340 23236
rect 7616 23196 7622 23208
rect 1394 23128 1400 23180
rect 1452 23168 1458 23180
rect 1489 23171 1547 23177
rect 1489 23168 1501 23171
rect 1452 23140 1501 23168
rect 1452 23128 1458 23140
rect 1489 23137 1501 23140
rect 1535 23137 1547 23171
rect 1489 23131 1547 23137
rect 4249 23171 4307 23177
rect 4249 23137 4261 23171
rect 4295 23168 4307 23171
rect 4614 23168 4620 23180
rect 4295 23140 4620 23168
rect 4295 23137 4307 23140
rect 4249 23131 4307 23137
rect 4614 23128 4620 23140
rect 4672 23168 4678 23180
rect 4801 23171 4859 23177
rect 4801 23168 4813 23171
rect 4672 23140 4813 23168
rect 4672 23128 4678 23140
rect 4801 23137 4813 23140
rect 4847 23137 4859 23171
rect 4801 23131 4859 23137
rect 4985 23171 5043 23177
rect 4985 23137 4997 23171
rect 5031 23168 5043 23171
rect 5442 23168 5448 23180
rect 5031 23140 5448 23168
rect 5031 23137 5043 23140
rect 4985 23131 5043 23137
rect 5442 23128 5448 23140
rect 5500 23168 5506 23180
rect 5626 23168 5632 23180
rect 5500 23140 5632 23168
rect 5500 23128 5506 23140
rect 5626 23128 5632 23140
rect 5684 23128 5690 23180
rect 6546 23168 6552 23180
rect 6507 23140 6552 23168
rect 6546 23128 6552 23140
rect 6604 23128 6610 23180
rect 8202 23168 8208 23180
rect 8163 23140 8208 23168
rect 8202 23128 8208 23140
rect 8260 23128 8266 23180
rect 8312 23177 8340 23208
rect 8389 23205 8401 23239
rect 8435 23236 8447 23239
rect 8662 23236 8668 23248
rect 8435 23208 8668 23236
rect 8435 23205 8447 23208
rect 8389 23199 8447 23205
rect 8662 23196 8668 23208
rect 8720 23196 8726 23248
rect 12069 23239 12127 23245
rect 12069 23205 12081 23239
rect 12115 23236 12127 23239
rect 12342 23236 12348 23248
rect 12115 23208 12348 23236
rect 12115 23205 12127 23208
rect 12069 23199 12127 23205
rect 12342 23196 12348 23208
rect 12400 23196 12406 23248
rect 12802 23196 12808 23248
rect 12860 23236 12866 23248
rect 12897 23239 12955 23245
rect 12897 23236 12909 23239
rect 12860 23208 12909 23236
rect 12860 23196 12866 23208
rect 12897 23205 12909 23208
rect 12943 23205 12955 23239
rect 12897 23199 12955 23205
rect 15930 23196 15936 23248
rect 15988 23236 15994 23248
rect 17954 23236 17960 23248
rect 15988 23208 16436 23236
rect 17915 23208 17960 23236
rect 15988 23196 15994 23208
rect 8297 23171 8355 23177
rect 8297 23137 8309 23171
rect 8343 23137 8355 23171
rect 8297 23131 8355 23137
rect 9677 23171 9735 23177
rect 9677 23137 9689 23171
rect 9723 23168 9735 23171
rect 9766 23168 9772 23180
rect 9723 23140 9772 23168
rect 9723 23137 9735 23140
rect 9677 23131 9735 23137
rect 9766 23128 9772 23140
rect 9824 23128 9830 23180
rect 11514 23168 11520 23180
rect 11475 23140 11520 23168
rect 11514 23128 11520 23140
rect 11572 23128 11578 23180
rect 11606 23128 11612 23180
rect 11664 23168 11670 23180
rect 13354 23168 13360 23180
rect 11664 23140 11709 23168
rect 13315 23140 13360 23168
rect 11664 23128 11670 23140
rect 13354 23128 13360 23140
rect 13412 23128 13418 23180
rect 13538 23168 13544 23180
rect 13499 23140 13544 23168
rect 13538 23128 13544 23140
rect 13596 23128 13602 23180
rect 13817 23171 13875 23177
rect 13817 23137 13829 23171
rect 13863 23168 13875 23171
rect 14366 23168 14372 23180
rect 13863 23140 14372 23168
rect 13863 23137 13875 23140
rect 13817 23131 13875 23137
rect 14366 23128 14372 23140
rect 14424 23128 14430 23180
rect 15105 23171 15163 23177
rect 15105 23137 15117 23171
rect 15151 23168 15163 23171
rect 16025 23171 16083 23177
rect 16025 23168 16037 23171
rect 15151 23140 16037 23168
rect 15151 23137 15163 23140
rect 15105 23131 15163 23137
rect 16025 23137 16037 23140
rect 16071 23168 16083 23171
rect 16114 23168 16120 23180
rect 16071 23140 16120 23168
rect 16071 23137 16083 23140
rect 16025 23131 16083 23137
rect 16114 23128 16120 23140
rect 16172 23128 16178 23180
rect 16408 23177 16436 23208
rect 17954 23196 17960 23208
rect 18012 23196 18018 23248
rect 19076 23236 19104 23276
rect 21085 23273 21097 23307
rect 21131 23304 21143 23307
rect 21358 23304 21364 23316
rect 21131 23276 21364 23304
rect 21131 23273 21143 23276
rect 21085 23267 21143 23273
rect 21358 23264 21364 23276
rect 21416 23264 21422 23316
rect 23474 23264 23480 23316
rect 23532 23304 23538 23316
rect 23845 23307 23903 23313
rect 23845 23304 23857 23307
rect 23532 23276 23857 23304
rect 23532 23264 23538 23276
rect 23845 23273 23857 23276
rect 23891 23273 23903 23307
rect 25590 23304 25596 23316
rect 25551 23276 25596 23304
rect 23845 23267 23903 23273
rect 25590 23264 25596 23276
rect 25648 23264 25654 23316
rect 26234 23304 26240 23316
rect 26195 23276 26240 23304
rect 26234 23264 26240 23276
rect 26292 23264 26298 23316
rect 27062 23264 27068 23316
rect 27120 23304 27126 23316
rect 27614 23304 27620 23316
rect 27120 23276 27620 23304
rect 27120 23264 27126 23276
rect 27614 23264 27620 23276
rect 27672 23264 27678 23316
rect 27890 23264 27896 23316
rect 27948 23304 27954 23316
rect 27985 23307 28043 23313
rect 27985 23304 27997 23307
rect 27948 23276 27997 23304
rect 27948 23264 27954 23276
rect 27985 23273 27997 23276
rect 28031 23273 28043 23307
rect 27985 23267 28043 23273
rect 19610 23236 19616 23248
rect 19076 23208 19616 23236
rect 16393 23171 16451 23177
rect 16393 23137 16405 23171
rect 16439 23137 16451 23171
rect 18874 23168 18880 23180
rect 18835 23140 18880 23168
rect 16393 23131 16451 23137
rect 18874 23128 18880 23140
rect 18932 23128 18938 23180
rect 19076 23177 19104 23208
rect 19610 23196 19616 23208
rect 19668 23196 19674 23248
rect 26252 23236 26280 23264
rect 26513 23239 26571 23245
rect 26513 23236 26525 23239
rect 26252 23208 26525 23236
rect 26513 23205 26525 23208
rect 26559 23205 26571 23239
rect 28000 23236 28028 23267
rect 28258 23264 28264 23316
rect 28316 23304 28322 23316
rect 28353 23307 28411 23313
rect 28353 23304 28365 23307
rect 28316 23276 28365 23304
rect 28316 23264 28322 23276
rect 28353 23273 28365 23276
rect 28399 23273 28411 23307
rect 28353 23267 28411 23273
rect 29362 23264 29368 23316
rect 29420 23304 29426 23316
rect 29825 23307 29883 23313
rect 29825 23304 29837 23307
rect 29420 23276 29837 23304
rect 29420 23264 29426 23276
rect 29825 23273 29837 23276
rect 29871 23273 29883 23307
rect 31018 23304 31024 23316
rect 30979 23276 31024 23304
rect 29825 23267 29883 23273
rect 31018 23264 31024 23276
rect 31076 23264 31082 23316
rect 31110 23264 31116 23316
rect 31168 23304 31174 23316
rect 31389 23307 31447 23313
rect 31389 23304 31401 23307
rect 31168 23276 31401 23304
rect 31168 23264 31174 23276
rect 31389 23273 31401 23276
rect 31435 23273 31447 23307
rect 31389 23267 31447 23273
rect 31754 23264 31760 23316
rect 31812 23304 31818 23316
rect 31941 23307 31999 23313
rect 31941 23304 31953 23307
rect 31812 23276 31953 23304
rect 31812 23264 31818 23276
rect 31941 23273 31953 23276
rect 31987 23273 31999 23307
rect 35802 23304 35808 23316
rect 35763 23276 35808 23304
rect 31941 23267 31999 23273
rect 35802 23264 35808 23276
rect 35860 23264 35866 23316
rect 28718 23236 28724 23248
rect 28000 23208 28724 23236
rect 26513 23199 26571 23205
rect 28718 23196 28724 23208
rect 28776 23236 28782 23248
rect 28776 23208 29592 23236
rect 28776 23196 28782 23208
rect 19061 23171 19119 23177
rect 19061 23137 19073 23171
rect 19107 23137 19119 23171
rect 19061 23131 19119 23137
rect 19245 23171 19303 23177
rect 19245 23137 19257 23171
rect 19291 23137 19303 23171
rect 19245 23131 19303 23137
rect 1670 23060 1676 23112
rect 1728 23100 1734 23112
rect 1765 23103 1823 23109
rect 1765 23100 1777 23103
rect 1728 23072 1777 23100
rect 1728 23060 1734 23072
rect 1765 23069 1777 23072
rect 1811 23100 1823 23103
rect 3510 23100 3516 23112
rect 1811 23072 3516 23100
rect 1811 23069 1823 23072
rect 1765 23063 1823 23069
rect 3510 23060 3516 23072
rect 3568 23060 3574 23112
rect 4157 23103 4215 23109
rect 4157 23069 4169 23103
rect 4203 23069 4215 23103
rect 4157 23063 4215 23069
rect 4172 23032 4200 23063
rect 7282 23060 7288 23112
rect 7340 23100 7346 23112
rect 7653 23103 7711 23109
rect 7653 23100 7665 23103
rect 7340 23072 7665 23100
rect 7340 23060 7346 23072
rect 7653 23069 7665 23072
rect 7699 23069 7711 23103
rect 8018 23100 8024 23112
rect 7979 23072 8024 23100
rect 7653 23063 7711 23069
rect 8018 23060 8024 23072
rect 8076 23060 8082 23112
rect 8757 23103 8815 23109
rect 8757 23069 8769 23103
rect 8803 23100 8815 23103
rect 10962 23100 10968 23112
rect 8803 23072 10968 23100
rect 8803 23069 8815 23072
rect 8757 23063 8815 23069
rect 10962 23060 10968 23072
rect 11020 23060 11026 23112
rect 14185 23103 14243 23109
rect 14185 23069 14197 23103
rect 14231 23069 14243 23103
rect 14185 23063 14243 23069
rect 5166 23032 5172 23044
rect 4172 23004 4936 23032
rect 5127 23004 5172 23032
rect 4908 22976 4936 23004
rect 5166 22992 5172 23004
rect 5224 22992 5230 23044
rect 10870 23032 10876 23044
rect 10831 23004 10876 23032
rect 10870 22992 10876 23004
rect 10928 22992 10934 23044
rect 14200 23032 14228 23063
rect 14274 23060 14280 23112
rect 14332 23100 14338 23112
rect 15838 23100 15844 23112
rect 14332 23072 14377 23100
rect 15799 23072 15844 23100
rect 14332 23060 14338 23072
rect 15838 23060 15844 23072
rect 15896 23060 15902 23112
rect 16298 23100 16304 23112
rect 16259 23072 16304 23100
rect 16298 23060 16304 23072
rect 16356 23060 16362 23112
rect 16758 23060 16764 23112
rect 16816 23100 16822 23112
rect 17221 23103 17279 23109
rect 17221 23100 17233 23103
rect 16816 23072 17233 23100
rect 16816 23060 16822 23072
rect 17221 23069 17233 23072
rect 17267 23069 17279 23103
rect 17221 23063 17279 23069
rect 18414 23060 18420 23112
rect 18472 23100 18478 23112
rect 19260 23100 19288 23131
rect 20070 23128 20076 23180
rect 20128 23168 20134 23180
rect 20714 23168 20720 23180
rect 20128 23140 20720 23168
rect 20128 23128 20134 23140
rect 20714 23128 20720 23140
rect 20772 23168 20778 23180
rect 20901 23171 20959 23177
rect 20901 23168 20913 23171
rect 20772 23140 20913 23168
rect 20772 23128 20778 23140
rect 20901 23137 20913 23140
rect 20947 23168 20959 23171
rect 21361 23171 21419 23177
rect 21361 23168 21373 23171
rect 20947 23140 21373 23168
rect 20947 23137 20959 23140
rect 20901 23131 20959 23137
rect 21361 23137 21373 23140
rect 21407 23137 21419 23171
rect 21361 23131 21419 23137
rect 22554 23128 22560 23180
rect 22612 23168 22618 23180
rect 22741 23171 22799 23177
rect 22741 23168 22753 23171
rect 22612 23140 22753 23168
rect 22612 23128 22618 23140
rect 22741 23137 22753 23140
rect 22787 23168 22799 23171
rect 25409 23171 25467 23177
rect 25409 23168 25421 23171
rect 22787 23140 25421 23168
rect 22787 23137 22799 23140
rect 22741 23131 22799 23137
rect 25409 23137 25421 23140
rect 25455 23168 25467 23171
rect 25958 23168 25964 23180
rect 25455 23140 25964 23168
rect 25455 23137 25467 23140
rect 25409 23131 25467 23137
rect 25958 23128 25964 23140
rect 26016 23128 26022 23180
rect 29089 23171 29147 23177
rect 29089 23137 29101 23171
rect 29135 23168 29147 23171
rect 29270 23168 29276 23180
rect 29135 23140 29276 23168
rect 29135 23137 29147 23140
rect 29089 23131 29147 23137
rect 29270 23128 29276 23140
rect 29328 23128 29334 23180
rect 29365 23171 29423 23177
rect 29365 23137 29377 23171
rect 29411 23168 29423 23171
rect 29454 23168 29460 23180
rect 29411 23140 29460 23168
rect 29411 23137 29423 23140
rect 29365 23131 29423 23137
rect 29454 23128 29460 23140
rect 29512 23128 29518 23180
rect 29564 23177 29592 23208
rect 29549 23171 29607 23177
rect 29549 23137 29561 23171
rect 29595 23137 29607 23171
rect 32309 23171 32367 23177
rect 32309 23168 32321 23171
rect 29549 23131 29607 23137
rect 31772 23140 32321 23168
rect 31772 23112 31800 23140
rect 32309 23137 32321 23140
rect 32355 23137 32367 23171
rect 32309 23131 32367 23137
rect 32950 23128 32956 23180
rect 33008 23168 33014 23180
rect 33045 23171 33103 23177
rect 33045 23168 33057 23171
rect 33008 23140 33057 23168
rect 33008 23128 33014 23140
rect 33045 23137 33057 23140
rect 33091 23137 33103 23171
rect 33045 23131 33103 23137
rect 18472 23072 19288 23100
rect 22465 23103 22523 23109
rect 18472 23060 18478 23072
rect 22465 23069 22477 23103
rect 22511 23100 22523 23103
rect 23198 23100 23204 23112
rect 22511 23072 23204 23100
rect 22511 23069 22523 23072
rect 22465 23063 22523 23069
rect 23198 23060 23204 23072
rect 23256 23060 23262 23112
rect 26878 23100 26884 23112
rect 26839 23072 26884 23100
rect 26878 23060 26884 23072
rect 26936 23060 26942 23112
rect 28534 23100 28540 23112
rect 28495 23072 28540 23100
rect 28534 23060 28540 23072
rect 28592 23060 28598 23112
rect 31754 23060 31760 23112
rect 31812 23060 31818 23112
rect 31941 23103 31999 23109
rect 31941 23069 31953 23103
rect 31987 23100 31999 23103
rect 32122 23100 32128 23112
rect 31987 23072 32128 23100
rect 31987 23069 31999 23072
rect 31941 23063 31999 23069
rect 32122 23060 32128 23072
rect 32180 23100 32186 23112
rect 32217 23103 32275 23109
rect 32217 23100 32229 23103
rect 32180 23072 32229 23100
rect 32180 23060 32186 23072
rect 32217 23069 32229 23072
rect 32263 23069 32275 23103
rect 32217 23063 32275 23069
rect 32490 23060 32496 23112
rect 32548 23100 32554 23112
rect 33137 23103 33195 23109
rect 33137 23100 33149 23103
rect 32548 23072 33149 23100
rect 32548 23060 32554 23072
rect 33137 23069 33149 23072
rect 33183 23069 33195 23103
rect 33137 23063 33195 23069
rect 18690 23032 18696 23044
rect 14200 23004 14320 23032
rect 18651 23004 18696 23032
rect 3053 22967 3111 22973
rect 3053 22933 3065 22967
rect 3099 22964 3111 22967
rect 3234 22964 3240 22976
rect 3099 22936 3240 22964
rect 3099 22933 3111 22936
rect 3053 22927 3111 22933
rect 3234 22924 3240 22936
rect 3292 22924 3298 22976
rect 3326 22924 3332 22976
rect 3384 22964 3390 22976
rect 3513 22967 3571 22973
rect 3513 22964 3525 22967
rect 3384 22936 3525 22964
rect 3384 22924 3390 22936
rect 3513 22933 3525 22936
rect 3559 22964 3571 22967
rect 3694 22964 3700 22976
rect 3559 22936 3700 22964
rect 3559 22933 3571 22936
rect 3513 22927 3571 22933
rect 3694 22924 3700 22936
rect 3752 22924 3758 22976
rect 4890 22924 4896 22976
rect 4948 22964 4954 22976
rect 5350 22964 5356 22976
rect 4948 22936 5356 22964
rect 4948 22924 4954 22936
rect 5350 22924 5356 22936
rect 5408 22964 5414 22976
rect 5721 22967 5779 22973
rect 5721 22964 5733 22967
rect 5408 22936 5733 22964
rect 5408 22924 5414 22936
rect 5721 22933 5733 22936
rect 5767 22933 5779 22967
rect 5721 22927 5779 22933
rect 7098 22924 7104 22976
rect 7156 22964 7162 22976
rect 7285 22967 7343 22973
rect 7285 22964 7297 22967
rect 7156 22936 7297 22964
rect 7156 22924 7162 22936
rect 7285 22933 7297 22936
rect 7331 22933 7343 22967
rect 9398 22964 9404 22976
rect 9359 22936 9404 22964
rect 7285 22927 7343 22933
rect 9398 22924 9404 22936
rect 9456 22924 9462 22976
rect 10778 22924 10784 22976
rect 10836 22964 10842 22976
rect 11333 22967 11391 22973
rect 11333 22964 11345 22967
rect 10836 22936 11345 22964
rect 10836 22924 10842 22936
rect 11333 22933 11345 22936
rect 11379 22964 11391 22967
rect 11422 22964 11428 22976
rect 11379 22936 11428 22964
rect 11379 22933 11391 22936
rect 11333 22927 11391 22933
rect 11422 22924 11428 22936
rect 11480 22924 11486 22976
rect 12434 22924 12440 22976
rect 12492 22964 12498 22976
rect 12802 22964 12808 22976
rect 12492 22936 12537 22964
rect 12763 22936 12808 22964
rect 12492 22924 12498 22936
rect 12802 22924 12808 22936
rect 12860 22924 12866 22976
rect 14292 22964 14320 23004
rect 18690 22992 18696 23004
rect 18748 22992 18754 23044
rect 26789 23035 26847 23041
rect 26789 23001 26801 23035
rect 26835 23032 26847 23035
rect 27246 23032 27252 23044
rect 26835 23004 27252 23032
rect 26835 23001 26847 23004
rect 26789 22995 26847 23001
rect 27246 22992 27252 23004
rect 27304 22992 27310 23044
rect 14550 22964 14556 22976
rect 14292 22936 14556 22964
rect 14550 22924 14556 22936
rect 14608 22964 14614 22976
rect 17402 22964 17408 22976
rect 14608 22936 17408 22964
rect 14608 22924 14614 22936
rect 17402 22924 17408 22936
rect 17460 22924 17466 22976
rect 18230 22924 18236 22976
rect 18288 22964 18294 22976
rect 20533 22967 20591 22973
rect 20533 22964 20545 22967
rect 18288 22936 20545 22964
rect 18288 22924 18294 22936
rect 20533 22933 20545 22936
rect 20579 22964 20591 22967
rect 20990 22964 20996 22976
rect 20579 22936 20996 22964
rect 20579 22933 20591 22936
rect 20533 22927 20591 22933
rect 20990 22924 20996 22936
rect 21048 22924 21054 22976
rect 25958 22964 25964 22976
rect 25919 22936 25964 22964
rect 25958 22924 25964 22936
rect 26016 22924 26022 22976
rect 26050 22924 26056 22976
rect 26108 22964 26114 22976
rect 26326 22964 26332 22976
rect 26108 22936 26332 22964
rect 26108 22924 26114 22936
rect 26326 22924 26332 22936
rect 26384 22964 26390 22976
rect 26651 22967 26709 22973
rect 26651 22964 26663 22967
rect 26384 22936 26663 22964
rect 26384 22924 26390 22936
rect 26651 22933 26663 22936
rect 26697 22933 26709 22967
rect 27154 22964 27160 22976
rect 27115 22936 27160 22964
rect 26651 22927 26709 22933
rect 27154 22924 27160 22936
rect 27212 22924 27218 22976
rect 30282 22964 30288 22976
rect 30243 22936 30288 22964
rect 30282 22924 30288 22936
rect 30340 22924 30346 22976
rect 1104 22874 38548 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 38548 22874
rect 1104 22800 38548 22822
rect 1670 22760 1676 22772
rect 1631 22732 1676 22760
rect 1670 22720 1676 22732
rect 1728 22720 1734 22772
rect 4157 22763 4215 22769
rect 4157 22729 4169 22763
rect 4203 22760 4215 22763
rect 4525 22763 4583 22769
rect 4525 22760 4537 22763
rect 4203 22732 4537 22760
rect 4203 22729 4215 22732
rect 4157 22723 4215 22729
rect 4525 22729 4537 22732
rect 4571 22760 4583 22763
rect 4614 22760 4620 22772
rect 4571 22732 4620 22760
rect 4571 22729 4583 22732
rect 4525 22723 4583 22729
rect 4614 22720 4620 22732
rect 4672 22720 4678 22772
rect 5169 22763 5227 22769
rect 5169 22729 5181 22763
rect 5215 22760 5227 22763
rect 5258 22760 5264 22772
rect 5215 22732 5264 22760
rect 5215 22729 5227 22732
rect 5169 22723 5227 22729
rect 5258 22720 5264 22732
rect 5316 22720 5322 22772
rect 10578 22763 10636 22769
rect 10578 22729 10590 22763
rect 10624 22760 10636 22763
rect 10962 22760 10968 22772
rect 10624 22732 10968 22760
rect 10624 22729 10636 22732
rect 10578 22723 10636 22729
rect 10962 22720 10968 22732
rect 11020 22720 11026 22772
rect 11057 22763 11115 22769
rect 11057 22729 11069 22763
rect 11103 22760 11115 22763
rect 11146 22760 11152 22772
rect 11103 22732 11152 22760
rect 11103 22729 11115 22732
rect 11057 22723 11115 22729
rect 11146 22720 11152 22732
rect 11204 22760 11210 22772
rect 11606 22760 11612 22772
rect 11204 22732 11612 22760
rect 11204 22720 11210 22732
rect 11606 22720 11612 22732
rect 11664 22720 11670 22772
rect 12250 22760 12256 22772
rect 12211 22732 12256 22760
rect 12250 22720 12256 22732
rect 12308 22720 12314 22772
rect 12526 22720 12532 22772
rect 12584 22760 12590 22772
rect 13538 22760 13544 22772
rect 12584 22732 13544 22760
rect 12584 22720 12590 22732
rect 13538 22720 13544 22732
rect 13596 22760 13602 22772
rect 13633 22763 13691 22769
rect 13633 22760 13645 22763
rect 13596 22732 13645 22760
rect 13596 22720 13602 22732
rect 13633 22729 13645 22732
rect 13679 22729 13691 22763
rect 13633 22723 13691 22729
rect 15194 22720 15200 22772
rect 15252 22760 15258 22772
rect 15933 22763 15991 22769
rect 15933 22760 15945 22763
rect 15252 22732 15945 22760
rect 15252 22720 15258 22732
rect 15933 22729 15945 22732
rect 15979 22760 15991 22763
rect 16942 22760 16948 22772
rect 15979 22732 16948 22760
rect 15979 22729 15991 22732
rect 15933 22723 15991 22729
rect 16942 22720 16948 22732
rect 17000 22720 17006 22772
rect 17402 22760 17408 22772
rect 17363 22732 17408 22760
rect 17402 22720 17408 22732
rect 17460 22720 17466 22772
rect 18230 22760 18236 22772
rect 18191 22732 18236 22760
rect 18230 22720 18236 22732
rect 18288 22720 18294 22772
rect 18598 22760 18604 22772
rect 18559 22732 18604 22760
rect 18598 22720 18604 22732
rect 18656 22720 18662 22772
rect 18874 22720 18880 22772
rect 18932 22760 18938 22772
rect 19245 22763 19303 22769
rect 19245 22760 19257 22763
rect 18932 22732 19257 22760
rect 18932 22720 18938 22732
rect 19245 22729 19257 22732
rect 19291 22729 19303 22763
rect 19610 22760 19616 22772
rect 19571 22732 19616 22760
rect 19245 22723 19303 22729
rect 19610 22720 19616 22732
rect 19668 22720 19674 22772
rect 19886 22720 19892 22772
rect 19944 22760 19950 22772
rect 19981 22763 20039 22769
rect 19981 22760 19993 22763
rect 19944 22732 19993 22760
rect 19944 22720 19950 22732
rect 19981 22729 19993 22732
rect 20027 22729 20039 22763
rect 21542 22760 21548 22772
rect 21503 22732 21548 22760
rect 19981 22723 20039 22729
rect 3142 22652 3148 22704
rect 3200 22692 3206 22704
rect 3200 22664 3372 22692
rect 3200 22652 3206 22664
rect 3344 22633 3372 22664
rect 6914 22652 6920 22704
rect 6972 22692 6978 22704
rect 8202 22692 8208 22704
rect 6972 22664 8208 22692
rect 6972 22652 6978 22664
rect 8202 22652 8208 22664
rect 8260 22692 8266 22704
rect 8297 22695 8355 22701
rect 8297 22692 8309 22695
rect 8260 22664 8309 22692
rect 8260 22652 8266 22664
rect 8297 22661 8309 22664
rect 8343 22692 8355 22695
rect 8665 22695 8723 22701
rect 8665 22692 8677 22695
rect 8343 22664 8677 22692
rect 8343 22661 8355 22664
rect 8297 22655 8355 22661
rect 8665 22661 8677 22664
rect 8711 22692 8723 22695
rect 9766 22692 9772 22704
rect 8711 22664 9772 22692
rect 8711 22661 8723 22664
rect 8665 22655 8723 22661
rect 2133 22627 2191 22633
rect 2133 22593 2145 22627
rect 2179 22624 2191 22627
rect 3329 22627 3387 22633
rect 2179 22596 3280 22624
rect 2179 22593 2191 22596
rect 2133 22587 2191 22593
rect 3252 22568 3280 22596
rect 3329 22593 3341 22627
rect 3375 22593 3387 22627
rect 3329 22587 3387 22593
rect 3510 22584 3516 22636
rect 3568 22624 3574 22636
rect 5166 22624 5172 22636
rect 3568 22596 5172 22624
rect 3568 22584 3574 22596
rect 2501 22559 2559 22565
rect 2501 22525 2513 22559
rect 2547 22556 2559 22559
rect 3050 22556 3056 22568
rect 2547 22528 3056 22556
rect 2547 22525 2559 22528
rect 2501 22519 2559 22525
rect 3050 22516 3056 22528
rect 3108 22516 3114 22568
rect 3234 22556 3240 22568
rect 3195 22528 3240 22556
rect 3234 22516 3240 22528
rect 3292 22516 3298 22568
rect 3620 22565 3648 22596
rect 5166 22584 5172 22596
rect 5224 22584 5230 22636
rect 7098 22584 7104 22636
rect 7156 22624 7162 22636
rect 7156 22596 7512 22624
rect 7156 22584 7162 22596
rect 3605 22559 3663 22565
rect 3605 22525 3617 22559
rect 3651 22525 3663 22559
rect 3786 22556 3792 22568
rect 3699 22528 3792 22556
rect 3605 22519 3663 22525
rect 3786 22516 3792 22528
rect 3844 22556 3850 22568
rect 4062 22556 4068 22568
rect 3844 22528 4068 22556
rect 3844 22516 3850 22528
rect 4062 22516 4068 22528
rect 4120 22516 4126 22568
rect 4890 22556 4896 22568
rect 4851 22528 4896 22556
rect 4890 22516 4896 22528
rect 4948 22516 4954 22568
rect 4985 22559 5043 22565
rect 4985 22525 4997 22559
rect 5031 22556 5043 22559
rect 5721 22559 5779 22565
rect 5721 22556 5733 22559
rect 5031 22528 5733 22556
rect 5031 22525 5043 22528
rect 4985 22519 5043 22525
rect 5721 22525 5733 22528
rect 5767 22556 5779 22559
rect 6638 22556 6644 22568
rect 5767 22528 6644 22556
rect 5767 22525 5779 22528
rect 5721 22519 5779 22525
rect 6638 22516 6644 22528
rect 6696 22516 6702 22568
rect 7484 22565 7512 22596
rect 8018 22584 8024 22636
rect 8076 22624 8082 22636
rect 8754 22624 8760 22636
rect 8076 22596 8760 22624
rect 8076 22584 8082 22596
rect 8754 22584 8760 22596
rect 8812 22624 8818 22636
rect 8849 22627 8907 22633
rect 8849 22624 8861 22627
rect 8812 22596 8861 22624
rect 8812 22584 8818 22596
rect 8849 22593 8861 22596
rect 8895 22593 8907 22627
rect 8849 22587 8907 22593
rect 7469 22559 7527 22565
rect 7469 22525 7481 22559
rect 7515 22525 7527 22559
rect 8956 22556 8984 22664
rect 9766 22652 9772 22664
rect 9824 22692 9830 22704
rect 9861 22695 9919 22701
rect 9861 22692 9873 22695
rect 9824 22664 9873 22692
rect 9824 22652 9830 22664
rect 9861 22661 9873 22664
rect 9907 22661 9919 22695
rect 10686 22692 10692 22704
rect 10647 22664 10692 22692
rect 9861 22655 9919 22661
rect 10686 22652 10692 22664
rect 10744 22652 10750 22704
rect 11422 22692 11428 22704
rect 11383 22664 11428 22692
rect 11422 22652 11428 22664
rect 11480 22652 11486 22704
rect 12618 22652 12624 22704
rect 12676 22692 12682 22704
rect 13081 22695 13139 22701
rect 13081 22692 13093 22695
rect 12676 22664 13093 22692
rect 12676 22652 12682 22664
rect 13081 22661 13093 22664
rect 13127 22692 13139 22695
rect 13311 22695 13369 22701
rect 13311 22692 13323 22695
rect 13127 22664 13323 22692
rect 13127 22661 13139 22664
rect 13081 22655 13139 22661
rect 13311 22661 13323 22664
rect 13357 22661 13369 22695
rect 17034 22692 17040 22704
rect 13311 22655 13369 22661
rect 16684 22664 17040 22692
rect 9674 22584 9680 22636
rect 9732 22624 9738 22636
rect 10781 22627 10839 22633
rect 10781 22624 10793 22627
rect 9732 22596 10793 22624
rect 9732 22584 9738 22596
rect 10781 22593 10793 22596
rect 10827 22624 10839 22627
rect 11054 22624 11060 22636
rect 10827 22596 11060 22624
rect 10827 22593 10839 22596
rect 10781 22587 10839 22593
rect 11054 22584 11060 22596
rect 11112 22584 11118 22636
rect 12713 22627 12771 22633
rect 12713 22593 12725 22627
rect 12759 22624 12771 22627
rect 13538 22624 13544 22636
rect 12759 22596 13544 22624
rect 12759 22593 12771 22596
rect 12713 22587 12771 22593
rect 13538 22584 13544 22596
rect 13596 22584 13602 22636
rect 14274 22624 14280 22636
rect 14187 22596 14280 22624
rect 14274 22584 14280 22596
rect 14332 22624 14338 22636
rect 14918 22624 14924 22636
rect 14332 22596 14924 22624
rect 14332 22584 14338 22596
rect 14918 22584 14924 22596
rect 14976 22584 14982 22636
rect 16684 22633 16712 22664
rect 17034 22652 17040 22664
rect 17092 22692 17098 22704
rect 17678 22692 17684 22704
rect 17092 22664 17684 22692
rect 17092 22652 17098 22664
rect 17678 22652 17684 22664
rect 17736 22652 17742 22704
rect 16669 22627 16727 22633
rect 16669 22593 16681 22627
rect 16715 22593 16727 22627
rect 16669 22587 16727 22593
rect 16758 22584 16764 22636
rect 16816 22624 16822 22636
rect 17129 22627 17187 22633
rect 17129 22624 17141 22627
rect 16816 22596 17141 22624
rect 16816 22584 16822 22596
rect 17129 22593 17141 22596
rect 17175 22593 17187 22627
rect 17129 22587 17187 22593
rect 18414 22584 18420 22636
rect 18472 22624 18478 22636
rect 18877 22627 18935 22633
rect 18877 22624 18889 22627
rect 18472 22596 18889 22624
rect 18472 22584 18478 22596
rect 18877 22593 18889 22596
rect 18923 22593 18935 22627
rect 18877 22587 18935 22593
rect 9033 22559 9091 22565
rect 9033 22556 9045 22559
rect 8956 22528 9045 22556
rect 7469 22519 7527 22525
rect 9033 22525 9045 22528
rect 9079 22525 9091 22559
rect 9033 22519 9091 22525
rect 12986 22516 12992 22568
rect 13044 22556 13050 22568
rect 13403 22559 13461 22565
rect 13403 22556 13415 22559
rect 13044 22528 13415 22556
rect 13044 22516 13050 22528
rect 13403 22525 13415 22528
rect 13449 22556 13461 22559
rect 13906 22556 13912 22568
rect 13449 22528 13912 22556
rect 13449 22525 13461 22528
rect 13403 22519 13461 22525
rect 13906 22516 13912 22528
rect 13964 22516 13970 22568
rect 13998 22516 14004 22568
rect 14056 22556 14062 22568
rect 14645 22559 14703 22565
rect 14645 22556 14657 22559
rect 14056 22528 14657 22556
rect 14056 22516 14062 22528
rect 14645 22525 14657 22528
rect 14691 22556 14703 22559
rect 14737 22559 14795 22565
rect 14737 22556 14749 22559
rect 14691 22528 14749 22556
rect 14691 22525 14703 22528
rect 14645 22519 14703 22525
rect 14737 22525 14749 22528
rect 14783 22525 14795 22559
rect 14737 22519 14795 22525
rect 14829 22559 14887 22565
rect 14829 22525 14841 22559
rect 14875 22556 14887 22559
rect 15102 22556 15108 22568
rect 14875 22528 15108 22556
rect 14875 22525 14887 22528
rect 14829 22519 14887 22525
rect 15102 22516 15108 22528
rect 15160 22556 15166 22568
rect 15565 22559 15623 22565
rect 15565 22556 15577 22559
rect 15160 22528 15577 22556
rect 15160 22516 15166 22528
rect 15565 22525 15577 22528
rect 15611 22525 15623 22559
rect 16942 22556 16948 22568
rect 16903 22528 16948 22556
rect 15565 22519 15623 22525
rect 16942 22516 16948 22528
rect 17000 22516 17006 22568
rect 18049 22559 18107 22565
rect 18049 22525 18061 22559
rect 18095 22556 18107 22559
rect 18598 22556 18604 22568
rect 18095 22528 18604 22556
rect 18095 22525 18107 22528
rect 18049 22519 18107 22525
rect 18598 22516 18604 22528
rect 18656 22516 18662 22568
rect 19996 22556 20024 22723
rect 21542 22720 21548 22732
rect 21600 22720 21606 22772
rect 22554 22760 22560 22772
rect 22515 22732 22560 22760
rect 22554 22720 22560 22732
rect 22612 22720 22618 22772
rect 22925 22763 22983 22769
rect 22925 22729 22937 22763
rect 22971 22760 22983 22763
rect 23198 22760 23204 22772
rect 22971 22732 23204 22760
rect 22971 22729 22983 22732
rect 22925 22723 22983 22729
rect 20162 22584 20168 22636
rect 20220 22633 20226 22636
rect 20220 22624 20230 22633
rect 22940 22624 22968 22723
rect 23198 22720 23204 22732
rect 23256 22720 23262 22772
rect 25869 22763 25927 22769
rect 25869 22729 25881 22763
rect 25915 22760 25927 22763
rect 26878 22760 26884 22772
rect 25915 22732 26884 22760
rect 25915 22729 25927 22732
rect 25869 22723 25927 22729
rect 26878 22720 26884 22732
rect 26936 22720 26942 22772
rect 26973 22763 27031 22769
rect 26973 22729 26985 22763
rect 27019 22760 27031 22763
rect 27246 22760 27252 22772
rect 27019 22732 27252 22760
rect 27019 22729 27031 22732
rect 26973 22723 27031 22729
rect 25590 22652 25596 22704
rect 25648 22692 25654 22704
rect 26145 22695 26203 22701
rect 26145 22692 26157 22695
rect 25648 22664 26157 22692
rect 25648 22652 25654 22664
rect 26145 22661 26157 22664
rect 26191 22661 26203 22695
rect 26145 22655 26203 22661
rect 25498 22624 25504 22636
rect 20220 22596 22968 22624
rect 25459 22596 25504 22624
rect 20220 22587 20230 22596
rect 20220 22584 20226 22587
rect 25498 22584 25504 22596
rect 25556 22584 25562 22636
rect 20441 22559 20499 22565
rect 20441 22556 20453 22559
rect 19996 22528 20453 22556
rect 20441 22525 20453 22528
rect 20487 22525 20499 22559
rect 20441 22519 20499 22525
rect 24673 22559 24731 22565
rect 24673 22525 24685 22559
rect 24719 22556 24731 22559
rect 25409 22559 25467 22565
rect 25409 22556 25421 22559
rect 24719 22528 25421 22556
rect 24719 22525 24731 22528
rect 24673 22519 24731 22525
rect 25409 22525 25421 22528
rect 25455 22556 25467 22559
rect 25958 22556 25964 22568
rect 25455 22528 25964 22556
rect 25455 22525 25467 22528
rect 25409 22519 25467 22525
rect 25958 22516 25964 22528
rect 26016 22516 26022 22568
rect 26160 22556 26188 22655
rect 26896 22624 26924 22720
rect 27172 22701 27200 22732
rect 27246 22720 27252 22732
rect 27304 22720 27310 22772
rect 28629 22763 28687 22769
rect 28629 22729 28641 22763
rect 28675 22760 28687 22763
rect 29270 22760 29276 22772
rect 28675 22732 29276 22760
rect 28675 22729 28687 22732
rect 28629 22723 28687 22729
rect 29270 22720 29276 22732
rect 29328 22720 29334 22772
rect 32122 22760 32128 22772
rect 32083 22732 32128 22760
rect 32122 22720 32128 22732
rect 32180 22720 32186 22772
rect 32490 22760 32496 22772
rect 32451 22732 32496 22760
rect 32490 22720 32496 22732
rect 32548 22720 32554 22772
rect 27157 22695 27215 22701
rect 27157 22661 27169 22695
rect 27203 22692 27215 22695
rect 27203 22664 27237 22692
rect 27203 22661 27215 22664
rect 27157 22655 27215 22661
rect 28718 22652 28724 22704
rect 28776 22692 28782 22704
rect 28905 22695 28963 22701
rect 28905 22692 28917 22695
rect 28776 22664 28917 22692
rect 28776 22652 28782 22664
rect 28905 22661 28917 22664
rect 28951 22661 28963 22695
rect 28905 22655 28963 22661
rect 29457 22695 29515 22701
rect 29457 22661 29469 22695
rect 29503 22692 29515 22695
rect 29546 22692 29552 22704
rect 29503 22664 29552 22692
rect 29503 22661 29515 22664
rect 29457 22655 29515 22661
rect 29546 22652 29552 22664
rect 29604 22652 29610 22704
rect 32950 22692 32956 22704
rect 32911 22664 32956 22692
rect 32950 22652 32956 22664
rect 33008 22652 33014 22704
rect 28077 22627 28135 22633
rect 28077 22624 28089 22627
rect 26896 22596 28089 22624
rect 27062 22556 27068 22568
rect 26160 22528 27068 22556
rect 27062 22516 27068 22528
rect 27120 22516 27126 22568
rect 27356 22565 27384 22596
rect 28077 22593 28089 22596
rect 28123 22593 28135 22627
rect 29564 22624 29592 22652
rect 30282 22624 30288 22636
rect 29564 22596 30288 22624
rect 28077 22587 28135 22593
rect 30282 22584 30288 22596
rect 30340 22624 30346 22636
rect 35713 22627 35771 22633
rect 30340 22596 30420 22624
rect 30340 22584 30346 22596
rect 27341 22559 27399 22565
rect 27341 22525 27353 22559
rect 27387 22525 27399 22559
rect 27341 22519 27399 22525
rect 27801 22559 27859 22565
rect 27801 22525 27813 22559
rect 27847 22556 27859 22559
rect 28442 22556 28448 22568
rect 27847 22528 28448 22556
rect 27847 22525 27859 22528
rect 27801 22519 27859 22525
rect 28442 22516 28448 22528
rect 28500 22556 28506 22568
rect 29086 22556 29092 22568
rect 28500 22528 29092 22556
rect 28500 22516 28506 22528
rect 29086 22516 29092 22528
rect 29144 22516 29150 22568
rect 29178 22516 29184 22568
rect 29236 22556 29242 22568
rect 30392 22565 30420 22596
rect 35713 22593 35725 22627
rect 35759 22624 35771 22627
rect 37274 22624 37280 22636
rect 35759 22596 36124 22624
rect 37235 22596 37280 22624
rect 35759 22593 35771 22596
rect 35713 22587 35771 22593
rect 36096 22568 36124 22596
rect 37274 22584 37280 22596
rect 37332 22584 37338 22636
rect 29273 22559 29331 22565
rect 29273 22556 29285 22559
rect 29236 22528 29285 22556
rect 29236 22516 29242 22528
rect 29273 22525 29285 22528
rect 29319 22556 29331 22559
rect 30101 22559 30159 22565
rect 30101 22556 30113 22559
rect 29319 22528 30113 22556
rect 29319 22525 29331 22528
rect 29273 22519 29331 22525
rect 30101 22525 30113 22528
rect 30147 22525 30159 22559
rect 30101 22519 30159 22525
rect 30377 22559 30435 22565
rect 30377 22525 30389 22559
rect 30423 22525 30435 22559
rect 35802 22556 35808 22568
rect 35763 22528 35808 22556
rect 30377 22519 30435 22525
rect 35802 22516 35808 22528
rect 35860 22516 35866 22568
rect 36078 22556 36084 22568
rect 36039 22528 36084 22556
rect 36078 22516 36084 22528
rect 36136 22516 36142 22568
rect 2590 22488 2596 22500
rect 2551 22460 2596 22488
rect 2590 22448 2596 22460
rect 2648 22448 2654 22500
rect 7282 22488 7288 22500
rect 7243 22460 7288 22488
rect 7282 22448 7288 22460
rect 7340 22448 7346 22500
rect 7653 22491 7711 22497
rect 7653 22488 7665 22491
rect 7484 22460 7665 22488
rect 6365 22423 6423 22429
rect 6365 22389 6377 22423
rect 6411 22420 6423 22423
rect 6546 22420 6552 22432
rect 6411 22392 6552 22420
rect 6411 22389 6423 22392
rect 6365 22383 6423 22389
rect 6546 22380 6552 22392
rect 6604 22380 6610 22432
rect 7193 22423 7251 22429
rect 7193 22389 7205 22423
rect 7239 22420 7251 22423
rect 7484 22420 7512 22460
rect 7653 22457 7665 22460
rect 7699 22488 7711 22491
rect 7834 22488 7840 22500
rect 7699 22460 7840 22488
rect 7699 22457 7711 22460
rect 7653 22451 7711 22457
rect 7834 22448 7840 22460
rect 7892 22448 7898 22500
rect 8021 22491 8079 22497
rect 8021 22457 8033 22491
rect 8067 22488 8079 22491
rect 8294 22488 8300 22500
rect 8067 22460 8300 22488
rect 8067 22457 8079 22460
rect 8021 22451 8079 22457
rect 8294 22448 8300 22460
rect 8352 22448 8358 22500
rect 9214 22488 9220 22500
rect 9175 22460 9220 22488
rect 9214 22448 9220 22460
rect 9272 22448 9278 22500
rect 9582 22488 9588 22500
rect 9543 22460 9588 22488
rect 9582 22448 9588 22460
rect 9640 22448 9646 22500
rect 10413 22491 10471 22497
rect 10413 22457 10425 22491
rect 10459 22488 10471 22491
rect 10778 22488 10784 22500
rect 10459 22460 10784 22488
rect 10459 22457 10471 22460
rect 10413 22451 10471 22457
rect 10778 22448 10784 22460
rect 10836 22448 10842 22500
rect 11514 22448 11520 22500
rect 11572 22488 11578 22500
rect 11885 22491 11943 22497
rect 11885 22488 11897 22491
rect 11572 22460 11897 22488
rect 11572 22448 11578 22460
rect 11885 22457 11897 22460
rect 11931 22488 11943 22491
rect 12342 22488 12348 22500
rect 11931 22460 12348 22488
rect 11931 22457 11943 22460
rect 11885 22451 11943 22457
rect 12342 22448 12348 22460
rect 12400 22448 12406 22500
rect 12802 22448 12808 22500
rect 12860 22488 12866 22500
rect 13173 22491 13231 22497
rect 13173 22488 13185 22491
rect 12860 22460 13185 22488
rect 12860 22448 12866 22460
rect 13173 22457 13185 22460
rect 13219 22488 13231 22491
rect 15289 22491 15347 22497
rect 15289 22488 15301 22491
rect 13219 22460 15301 22488
rect 13219 22457 13231 22460
rect 13173 22451 13231 22457
rect 15289 22457 15301 22460
rect 15335 22457 15347 22491
rect 15289 22451 15347 22457
rect 16117 22491 16175 22497
rect 16117 22457 16129 22491
rect 16163 22488 16175 22491
rect 16206 22488 16212 22500
rect 16163 22460 16212 22488
rect 16163 22457 16175 22460
rect 16117 22451 16175 22457
rect 16206 22448 16212 22460
rect 16264 22448 16270 22500
rect 16298 22448 16304 22500
rect 16356 22488 16362 22500
rect 17773 22491 17831 22497
rect 17773 22488 17785 22491
rect 16356 22460 17785 22488
rect 16356 22448 16362 22460
rect 17773 22457 17785 22460
rect 17819 22457 17831 22491
rect 17773 22451 17831 22457
rect 26605 22491 26663 22497
rect 26605 22457 26617 22491
rect 26651 22488 26663 22491
rect 27246 22488 27252 22500
rect 26651 22460 27252 22488
rect 26651 22457 26663 22460
rect 26605 22451 26663 22457
rect 27246 22448 27252 22460
rect 27304 22448 27310 22500
rect 29454 22448 29460 22500
rect 29512 22488 29518 22500
rect 29733 22491 29791 22497
rect 29733 22488 29745 22491
rect 29512 22460 29745 22488
rect 29512 22448 29518 22460
rect 29733 22457 29745 22460
rect 29779 22457 29791 22491
rect 29733 22451 29791 22457
rect 30834 22448 30840 22500
rect 30892 22488 30898 22500
rect 31021 22491 31079 22497
rect 31021 22488 31033 22491
rect 30892 22460 31033 22488
rect 30892 22448 30898 22460
rect 31021 22457 31033 22460
rect 31067 22488 31079 22491
rect 31570 22488 31576 22500
rect 31067 22460 31576 22488
rect 31067 22457 31079 22460
rect 31021 22451 31079 22457
rect 31570 22448 31576 22460
rect 31628 22448 31634 22500
rect 7239 22392 7512 22420
rect 7239 22389 7251 22392
rect 7193 22383 7251 22389
rect 7558 22380 7564 22432
rect 7616 22420 7622 22432
rect 9125 22423 9183 22429
rect 9125 22420 9137 22423
rect 7616 22392 9137 22420
rect 7616 22380 7622 22392
rect 9125 22389 9137 22392
rect 9171 22420 9183 22423
rect 9398 22420 9404 22432
rect 9171 22392 9404 22420
rect 9171 22389 9183 22392
rect 9125 22383 9183 22389
rect 9398 22380 9404 22392
rect 9456 22420 9462 22432
rect 10229 22423 10287 22429
rect 10229 22420 10241 22423
rect 9456 22392 10241 22420
rect 9456 22380 9462 22392
rect 10229 22389 10241 22392
rect 10275 22420 10287 22423
rect 10502 22420 10508 22432
rect 10275 22392 10508 22420
rect 10275 22389 10287 22392
rect 10229 22383 10287 22389
rect 10502 22380 10508 22392
rect 10560 22380 10566 22432
rect 1104 22330 38548 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 38548 22330
rect 1104 22256 38548 22278
rect 3053 22219 3111 22225
rect 3053 22185 3065 22219
rect 3099 22216 3111 22219
rect 3510 22216 3516 22228
rect 3099 22188 3516 22216
rect 3099 22185 3111 22188
rect 3053 22179 3111 22185
rect 3510 22176 3516 22188
rect 3568 22176 3574 22228
rect 3881 22219 3939 22225
rect 3881 22185 3893 22219
rect 3927 22216 3939 22219
rect 3970 22216 3976 22228
rect 3927 22188 3976 22216
rect 3927 22185 3939 22188
rect 3881 22179 3939 22185
rect 3786 22148 3792 22160
rect 2792 22120 3792 22148
rect 2685 22083 2743 22089
rect 2685 22049 2697 22083
rect 2731 22080 2743 22083
rect 2792 22080 2820 22120
rect 3786 22108 3792 22120
rect 3844 22108 3850 22160
rect 2731 22052 2820 22080
rect 2731 22049 2743 22052
rect 2685 22043 2743 22049
rect 2866 22040 2872 22092
rect 2924 22080 2930 22092
rect 3896 22080 3924 22179
rect 3970 22176 3976 22188
rect 4028 22176 4034 22228
rect 5353 22219 5411 22225
rect 5353 22185 5365 22219
rect 5399 22216 5411 22219
rect 5721 22219 5779 22225
rect 5721 22216 5733 22219
rect 5399 22188 5733 22216
rect 5399 22185 5411 22188
rect 5353 22179 5411 22185
rect 5721 22185 5733 22188
rect 5767 22216 5779 22219
rect 5902 22216 5908 22228
rect 5767 22188 5908 22216
rect 5767 22185 5779 22188
rect 5721 22179 5779 22185
rect 5902 22176 5908 22188
rect 5960 22176 5966 22228
rect 6178 22176 6184 22228
rect 6236 22216 6242 22228
rect 6457 22219 6515 22225
rect 6457 22216 6469 22219
rect 6236 22188 6469 22216
rect 6236 22176 6242 22188
rect 6457 22185 6469 22188
rect 6503 22185 6515 22219
rect 6457 22179 6515 22185
rect 4614 22108 4620 22160
rect 4672 22148 4678 22160
rect 5813 22151 5871 22157
rect 5813 22148 5825 22151
rect 4672 22120 5825 22148
rect 4672 22108 4678 22120
rect 5813 22117 5825 22120
rect 5859 22148 5871 22151
rect 6086 22148 6092 22160
rect 5859 22120 6092 22148
rect 5859 22117 5871 22120
rect 5813 22111 5871 22117
rect 6086 22108 6092 22120
rect 6144 22108 6150 22160
rect 6472 22148 6500 22179
rect 7282 22176 7288 22228
rect 7340 22216 7346 22228
rect 8754 22216 8760 22228
rect 7340 22188 8156 22216
rect 8715 22188 8760 22216
rect 7340 22176 7346 22188
rect 8018 22148 8024 22160
rect 6472 22120 8024 22148
rect 8018 22108 8024 22120
rect 8076 22108 8082 22160
rect 8128 22148 8156 22188
rect 8754 22176 8760 22188
rect 8812 22216 8818 22228
rect 9033 22219 9091 22225
rect 9033 22216 9045 22219
rect 8812 22188 9045 22216
rect 8812 22176 8818 22188
rect 9033 22185 9045 22188
rect 9079 22185 9091 22219
rect 9398 22216 9404 22228
rect 9359 22188 9404 22216
rect 9033 22179 9091 22185
rect 9398 22176 9404 22188
rect 9456 22216 9462 22228
rect 9953 22219 10011 22225
rect 9953 22216 9965 22219
rect 9456 22188 9965 22216
rect 9456 22176 9462 22188
rect 9953 22185 9965 22188
rect 9999 22185 10011 22219
rect 9953 22179 10011 22185
rect 13354 22176 13360 22228
rect 13412 22216 13418 22228
rect 15838 22216 15844 22228
rect 13412 22188 13768 22216
rect 15799 22188 15844 22216
rect 13412 22176 13418 22188
rect 10042 22148 10048 22160
rect 8128 22120 8340 22148
rect 10003 22120 10048 22148
rect 2924 22052 3924 22080
rect 4433 22083 4491 22089
rect 2924 22040 2930 22052
rect 4433 22049 4445 22083
rect 4479 22080 4491 22083
rect 4706 22080 4712 22092
rect 4479 22052 4712 22080
rect 4479 22049 4491 22052
rect 4433 22043 4491 22049
rect 4706 22040 4712 22052
rect 4764 22040 4770 22092
rect 4985 22083 5043 22089
rect 4985 22049 4997 22083
rect 5031 22080 5043 22083
rect 5077 22083 5135 22089
rect 5077 22080 5089 22083
rect 5031 22052 5089 22080
rect 5031 22049 5043 22052
rect 4985 22043 5043 22049
rect 5077 22049 5089 22052
rect 5123 22080 5135 22083
rect 5258 22080 5264 22092
rect 5123 22052 5264 22080
rect 5123 22049 5135 22052
rect 5077 22043 5135 22049
rect 5258 22040 5264 22052
rect 5316 22040 5322 22092
rect 5445 22083 5503 22089
rect 5445 22049 5457 22083
rect 5491 22080 5503 22083
rect 5534 22080 5540 22092
rect 5491 22052 5540 22080
rect 5491 22049 5503 22052
rect 5445 22043 5503 22049
rect 1673 22015 1731 22021
rect 1673 21981 1685 22015
rect 1719 22012 1731 22015
rect 1854 22012 1860 22024
rect 1719 21984 1860 22012
rect 1719 21981 1731 21984
rect 1673 21975 1731 21981
rect 1854 21972 1860 21984
rect 1912 22012 1918 22024
rect 2884 22012 2912 22040
rect 1912 21984 2912 22012
rect 4341 22015 4399 22021
rect 1912 21972 1918 21984
rect 4341 21981 4353 22015
rect 4387 22012 4399 22015
rect 5169 22015 5227 22021
rect 5169 22012 5181 22015
rect 4387 21984 5181 22012
rect 4387 21981 4399 21984
rect 4341 21975 4399 21981
rect 5169 21981 5181 21984
rect 5215 21981 5227 22015
rect 5169 21975 5227 21981
rect 4617 21947 4675 21953
rect 4617 21913 4629 21947
rect 4663 21944 4675 21947
rect 5460 21944 5488 22043
rect 5534 22040 5540 22052
rect 5592 22040 5598 22092
rect 5629 22083 5687 22089
rect 5629 22049 5641 22083
rect 5675 22080 5687 22083
rect 6454 22080 6460 22092
rect 5675 22052 6460 22080
rect 5675 22049 5687 22052
rect 5629 22043 5687 22049
rect 6454 22040 6460 22052
rect 6512 22080 6518 22092
rect 6822 22080 6828 22092
rect 6512 22052 6828 22080
rect 6512 22040 6518 22052
rect 6822 22040 6828 22052
rect 6880 22040 6886 22092
rect 7006 22080 7012 22092
rect 6967 22052 7012 22080
rect 7006 22040 7012 22052
rect 7064 22040 7070 22092
rect 7156 22083 7214 22089
rect 7156 22049 7168 22083
rect 7202 22080 7214 22083
rect 8202 22080 8208 22092
rect 7202 22052 8208 22080
rect 7202 22049 7214 22052
rect 7156 22043 7214 22049
rect 8202 22040 8208 22052
rect 8260 22040 8266 22092
rect 8312 22080 8340 22120
rect 10042 22108 10048 22120
rect 10100 22108 10106 22160
rect 10502 22108 10508 22160
rect 10560 22148 10566 22160
rect 10689 22151 10747 22157
rect 10689 22148 10701 22151
rect 10560 22120 10701 22148
rect 10560 22108 10566 22120
rect 10689 22117 10701 22120
rect 10735 22117 10747 22151
rect 12526 22148 12532 22160
rect 12487 22120 12532 22148
rect 10689 22111 10747 22117
rect 12526 22108 12532 22120
rect 12584 22108 12590 22160
rect 8573 22083 8631 22089
rect 8573 22080 8585 22083
rect 8312 22052 8585 22080
rect 8404 22024 8432 22052
rect 8573 22049 8585 22052
rect 8619 22049 8631 22083
rect 8573 22043 8631 22049
rect 9214 22040 9220 22092
rect 9272 22080 9278 22092
rect 9861 22083 9919 22089
rect 9861 22080 9873 22083
rect 9272 22052 9873 22080
rect 9272 22040 9278 22052
rect 9861 22049 9873 22052
rect 9907 22049 9919 22083
rect 11054 22080 11060 22092
rect 11015 22052 11060 22080
rect 9861 22043 9919 22049
rect 11054 22040 11060 22052
rect 11112 22040 11118 22092
rect 11241 22083 11299 22089
rect 11241 22049 11253 22083
rect 11287 22080 11299 22083
rect 11330 22080 11336 22092
rect 11287 22052 11336 22080
rect 11287 22049 11299 22052
rect 11241 22043 11299 22049
rect 11330 22040 11336 22052
rect 11388 22040 11394 22092
rect 11425 22083 11483 22089
rect 11425 22049 11437 22083
rect 11471 22080 11483 22083
rect 11882 22080 11888 22092
rect 11471 22052 11888 22080
rect 11471 22049 11483 22052
rect 11425 22043 11483 22049
rect 11882 22040 11888 22052
rect 11940 22080 11946 22092
rect 12250 22080 12256 22092
rect 11940 22052 12256 22080
rect 11940 22040 11946 22052
rect 12250 22040 12256 22052
rect 12308 22040 12314 22092
rect 12621 22083 12679 22089
rect 12621 22049 12633 22083
rect 12667 22080 12679 22083
rect 12710 22080 12716 22092
rect 12667 22052 12716 22080
rect 12667 22049 12679 22052
rect 12621 22043 12679 22049
rect 12710 22040 12716 22052
rect 12768 22040 12774 22092
rect 12802 22040 12808 22092
rect 12860 22080 12866 22092
rect 12860 22052 12905 22080
rect 12860 22040 12866 22052
rect 6181 22015 6239 22021
rect 6181 21981 6193 22015
rect 6227 22012 6239 22015
rect 6270 22012 6276 22024
rect 6227 21984 6276 22012
rect 6227 21981 6239 21984
rect 6181 21975 6239 21981
rect 6270 21972 6276 21984
rect 6328 21972 6334 22024
rect 7374 22012 7380 22024
rect 7335 21984 7380 22012
rect 7374 21972 7380 21984
rect 7432 21972 7438 22024
rect 7650 22012 7656 22024
rect 7611 21984 7656 22012
rect 7650 21972 7656 21984
rect 7708 21972 7714 22024
rect 8386 21972 8392 22024
rect 8444 21972 8450 22024
rect 9674 22012 9680 22024
rect 9635 21984 9680 22012
rect 9674 21972 9680 21984
rect 9732 21972 9738 22024
rect 10413 22015 10471 22021
rect 10413 21981 10425 22015
rect 10459 22012 10471 22015
rect 10686 22012 10692 22024
rect 10459 21984 10692 22012
rect 10459 21981 10471 21984
rect 10413 21975 10471 21981
rect 10686 21972 10692 21984
rect 10744 22012 10750 22024
rect 12069 22015 12127 22021
rect 12069 22012 12081 22015
rect 10744 21984 12081 22012
rect 10744 21972 10750 21984
rect 12069 21981 12081 21984
rect 12115 21981 12127 22015
rect 13740 22012 13768 22188
rect 15838 22176 15844 22188
rect 15896 22176 15902 22228
rect 16022 22176 16028 22228
rect 16080 22216 16086 22228
rect 16209 22219 16267 22225
rect 16209 22216 16221 22219
rect 16080 22188 16221 22216
rect 16080 22176 16086 22188
rect 16209 22185 16221 22188
rect 16255 22185 16267 22219
rect 16209 22179 16267 22185
rect 19426 22176 19432 22228
rect 19484 22216 19490 22228
rect 19521 22219 19579 22225
rect 19521 22216 19533 22219
rect 19484 22188 19533 22216
rect 19484 22176 19490 22188
rect 19521 22185 19533 22188
rect 19567 22216 19579 22219
rect 20162 22216 20168 22228
rect 19567 22188 20168 22216
rect 19567 22185 19579 22188
rect 19521 22179 19579 22185
rect 20162 22176 20168 22188
rect 20220 22176 20226 22228
rect 26326 22216 26332 22228
rect 26287 22188 26332 22216
rect 26326 22176 26332 22188
rect 26384 22176 26390 22228
rect 29454 22176 29460 22228
rect 29512 22216 29518 22228
rect 29822 22216 29828 22228
rect 29512 22188 29828 22216
rect 29512 22176 29518 22188
rect 29822 22176 29828 22188
rect 29880 22176 29886 22228
rect 35802 22216 35808 22228
rect 35763 22188 35808 22216
rect 35802 22176 35808 22188
rect 35860 22176 35866 22228
rect 15565 22151 15623 22157
rect 15565 22117 15577 22151
rect 15611 22148 15623 22151
rect 15930 22148 15936 22160
rect 15611 22120 15936 22148
rect 15611 22117 15623 22120
rect 15565 22111 15623 22117
rect 15930 22108 15936 22120
rect 15988 22148 15994 22160
rect 15988 22120 16896 22148
rect 15988 22108 15994 22120
rect 13906 22080 13912 22092
rect 13867 22052 13912 22080
rect 13906 22040 13912 22052
rect 13964 22040 13970 22092
rect 14642 22080 14648 22092
rect 14603 22052 14648 22080
rect 14642 22040 14648 22052
rect 14700 22040 14706 22092
rect 16761 22083 16819 22089
rect 16761 22080 16773 22083
rect 16408 22052 16773 22080
rect 14277 22015 14335 22021
rect 14277 22012 14289 22015
rect 13740 21984 14289 22012
rect 12069 21975 12127 21981
rect 14277 21981 14289 21984
rect 14323 21981 14335 22015
rect 14277 21975 14335 21981
rect 16022 21972 16028 22024
rect 16080 22012 16086 22024
rect 16206 22012 16212 22024
rect 16080 21984 16212 22012
rect 16080 21972 16086 21984
rect 16206 21972 16212 21984
rect 16264 22012 16270 22024
rect 16408 22012 16436 22052
rect 16761 22049 16773 22052
rect 16807 22049 16819 22083
rect 16868 22080 16896 22120
rect 17129 22083 17187 22089
rect 17129 22080 17141 22083
rect 16868 22052 17141 22080
rect 16761 22043 16819 22049
rect 17129 22049 17141 22052
rect 17175 22080 17187 22083
rect 17402 22080 17408 22092
rect 17175 22052 17408 22080
rect 17175 22049 17187 22052
rect 17129 22043 17187 22049
rect 17402 22040 17408 22052
rect 17460 22040 17466 22092
rect 18598 22040 18604 22092
rect 18656 22080 18662 22092
rect 18969 22083 19027 22089
rect 18969 22080 18981 22083
rect 18656 22052 18981 22080
rect 18656 22040 18662 22052
rect 18969 22049 18981 22052
rect 19015 22049 19027 22083
rect 21266 22080 21272 22092
rect 21227 22052 21272 22080
rect 18969 22043 19027 22049
rect 21266 22040 21272 22052
rect 21324 22040 21330 22092
rect 22085 22083 22143 22089
rect 22085 22049 22097 22083
rect 22131 22080 22143 22083
rect 22278 22080 22284 22092
rect 22131 22052 22284 22080
rect 22131 22049 22143 22052
rect 22085 22043 22143 22049
rect 22278 22040 22284 22052
rect 22336 22040 22342 22092
rect 23661 22083 23719 22089
rect 23661 22049 23673 22083
rect 23707 22049 23719 22083
rect 23661 22043 23719 22049
rect 24029 22083 24087 22089
rect 24029 22049 24041 22083
rect 24075 22080 24087 22083
rect 24486 22080 24492 22092
rect 24075 22052 24492 22080
rect 24075 22049 24087 22052
rect 24029 22043 24087 22049
rect 16574 22012 16580 22024
rect 16264 21984 16436 22012
rect 16535 21984 16580 22012
rect 16264 21972 16270 21984
rect 16574 21972 16580 21984
rect 16632 21972 16638 22024
rect 17037 22015 17095 22021
rect 17037 21981 17049 22015
rect 17083 21981 17095 22015
rect 17037 21975 17095 21981
rect 4663 21916 5488 21944
rect 4663 21913 4675 21916
rect 4617 21907 4675 21913
rect 8662 21904 8668 21956
rect 8720 21944 8726 21956
rect 16298 21944 16304 21956
rect 8720 21916 16304 21944
rect 8720 21904 8726 21916
rect 16298 21904 16304 21916
rect 16356 21944 16362 21956
rect 17052 21944 17080 21975
rect 17218 21972 17224 22024
rect 17276 22012 17282 22024
rect 18141 22015 18199 22021
rect 18141 22012 18153 22015
rect 17276 21984 18153 22012
rect 17276 21972 17282 21984
rect 18141 21981 18153 21984
rect 18187 21981 18199 22015
rect 18141 21975 18199 21981
rect 18693 22015 18751 22021
rect 18693 21981 18705 22015
rect 18739 21981 18751 22015
rect 18693 21975 18751 21981
rect 17589 21947 17647 21953
rect 17589 21944 17601 21947
rect 16356 21916 17601 21944
rect 16356 21904 16362 21916
rect 17589 21913 17601 21916
rect 17635 21913 17647 21947
rect 17589 21907 17647 21913
rect 17678 21904 17684 21956
rect 17736 21944 17742 21956
rect 18708 21944 18736 21975
rect 18782 21972 18788 22024
rect 18840 22012 18846 22024
rect 19153 22015 19211 22021
rect 19153 22012 19165 22015
rect 18840 21984 19165 22012
rect 18840 21972 18846 21984
rect 19153 21981 19165 21984
rect 19199 21981 19211 22015
rect 21358 22012 21364 22024
rect 21319 21984 21364 22012
rect 19153 21975 19211 21981
rect 21358 21972 21364 21984
rect 21416 21972 21422 22024
rect 22189 22015 22247 22021
rect 22189 21981 22201 22015
rect 22235 22012 22247 22015
rect 22370 22012 22376 22024
rect 22235 21984 22376 22012
rect 22235 21981 22247 21984
rect 22189 21975 22247 21981
rect 22370 21972 22376 21984
rect 22428 21972 22434 22024
rect 23290 22012 23296 22024
rect 23251 21984 23296 22012
rect 23290 21972 23296 21984
rect 23348 21972 23354 22024
rect 23676 22012 23704 22043
rect 24486 22040 24492 22052
rect 24544 22040 24550 22092
rect 27338 22080 27344 22092
rect 27299 22052 27344 22080
rect 27338 22040 27344 22052
rect 27396 22040 27402 22092
rect 28810 22080 28816 22092
rect 28771 22052 28816 22080
rect 28810 22040 28816 22052
rect 28868 22040 28874 22092
rect 30466 22080 30472 22092
rect 30427 22052 30472 22080
rect 30466 22040 30472 22052
rect 30524 22040 30530 22092
rect 31021 22083 31079 22089
rect 31021 22049 31033 22083
rect 31067 22080 31079 22083
rect 31294 22080 31300 22092
rect 31067 22052 31300 22080
rect 31067 22049 31079 22052
rect 31021 22043 31079 22049
rect 31294 22040 31300 22052
rect 31352 22040 31358 22092
rect 32677 22083 32735 22089
rect 32677 22049 32689 22083
rect 32723 22080 32735 22083
rect 33042 22080 33048 22092
rect 32723 22052 33048 22080
rect 32723 22049 32735 22052
rect 32677 22043 32735 22049
rect 33042 22040 33048 22052
rect 33100 22080 33106 22092
rect 35250 22080 35256 22092
rect 33100 22052 35256 22080
rect 33100 22040 33106 22052
rect 35250 22040 35256 22052
rect 35308 22080 35314 22092
rect 35820 22080 35848 22176
rect 35308 22052 35848 22080
rect 35308 22040 35314 22052
rect 26513 22015 26571 22021
rect 26513 22012 26525 22015
rect 23676 21984 24072 22012
rect 24044 21956 24072 21984
rect 25884 21984 26525 22012
rect 17736 21916 18736 21944
rect 17736 21904 17742 21916
rect 23658 21904 23664 21956
rect 23716 21944 23722 21956
rect 23937 21947 23995 21953
rect 23937 21944 23949 21947
rect 23716 21916 23949 21944
rect 23716 21904 23722 21916
rect 23937 21913 23949 21916
rect 23983 21913 23995 21947
rect 23937 21907 23995 21913
rect 24026 21904 24032 21956
rect 24084 21904 24090 21956
rect 25884 21888 25912 21984
rect 26513 21981 26525 21984
rect 26559 21981 26571 22015
rect 26513 21975 26571 21981
rect 27065 22015 27123 22021
rect 27065 21981 27077 22015
rect 27111 21981 27123 22015
rect 27065 21975 27123 21981
rect 27080 21944 27108 21975
rect 27154 21972 27160 22024
rect 27212 22012 27218 22024
rect 27525 22015 27583 22021
rect 27525 22012 27537 22015
rect 27212 21984 27537 22012
rect 27212 21972 27218 21984
rect 27525 21981 27537 21984
rect 27571 21981 27583 22015
rect 30282 22012 30288 22024
rect 30243 21984 30288 22012
rect 27525 21975 27583 21981
rect 30282 21972 30288 21984
rect 30340 21972 30346 22024
rect 30650 21972 30656 22024
rect 30708 22012 30714 22024
rect 30929 22015 30987 22021
rect 30929 22012 30941 22015
rect 30708 21984 30941 22012
rect 30708 21972 30714 21984
rect 30929 21981 30941 21984
rect 30975 21981 30987 22015
rect 32950 22012 32956 22024
rect 32911 21984 32956 22012
rect 30929 21975 30987 21981
rect 32950 21972 32956 21984
rect 33008 21972 33014 22024
rect 27614 21944 27620 21956
rect 27080 21916 27620 21944
rect 27614 21904 27620 21916
rect 27672 21904 27678 21956
rect 2038 21876 2044 21888
rect 1999 21848 2044 21876
rect 2038 21836 2044 21848
rect 2096 21836 2102 21888
rect 3510 21876 3516 21888
rect 3471 21848 3516 21876
rect 3510 21836 3516 21848
rect 3568 21836 3574 21888
rect 5074 21876 5080 21888
rect 5035 21848 5080 21876
rect 5074 21836 5080 21848
rect 5132 21836 5138 21888
rect 5169 21879 5227 21885
rect 5169 21845 5181 21879
rect 5215 21876 5227 21879
rect 5442 21876 5448 21888
rect 5215 21848 5448 21876
rect 5215 21845 5227 21848
rect 5169 21839 5227 21845
rect 5442 21836 5448 21848
rect 5500 21876 5506 21888
rect 5626 21876 5632 21888
rect 5500 21848 5632 21876
rect 5500 21836 5506 21848
rect 5626 21836 5632 21848
rect 5684 21836 5690 21888
rect 6917 21879 6975 21885
rect 6917 21845 6929 21879
rect 6963 21876 6975 21879
rect 7190 21876 7196 21888
rect 6963 21848 7196 21876
rect 6963 21845 6975 21848
rect 6917 21839 6975 21845
rect 7190 21836 7196 21848
rect 7248 21836 7254 21888
rect 7285 21879 7343 21885
rect 7285 21845 7297 21879
rect 7331 21876 7343 21879
rect 7558 21876 7564 21888
rect 7331 21848 7564 21876
rect 7331 21845 7343 21848
rect 7285 21839 7343 21845
rect 7558 21836 7564 21848
rect 7616 21836 7622 21888
rect 8481 21879 8539 21885
rect 8481 21845 8493 21879
rect 8527 21876 8539 21879
rect 8570 21876 8576 21888
rect 8527 21848 8576 21876
rect 8527 21845 8539 21848
rect 8481 21839 8539 21845
rect 8570 21836 8576 21848
rect 8628 21836 8634 21888
rect 9122 21836 9128 21888
rect 9180 21876 9186 21888
rect 9582 21876 9588 21888
rect 9180 21848 9588 21876
rect 9180 21836 9186 21848
rect 9582 21836 9588 21848
rect 9640 21836 9646 21888
rect 11238 21836 11244 21888
rect 11296 21876 11302 21888
rect 11517 21879 11575 21885
rect 11517 21876 11529 21879
rect 11296 21848 11529 21876
rect 11296 21836 11302 21848
rect 11517 21845 11529 21848
rect 11563 21845 11575 21879
rect 11517 21839 11575 21845
rect 12434 21836 12440 21888
rect 12492 21876 12498 21888
rect 12897 21879 12955 21885
rect 12897 21876 12909 21879
rect 12492 21848 12909 21876
rect 12492 21836 12498 21848
rect 12897 21845 12909 21848
rect 12943 21845 12955 21879
rect 12897 21839 12955 21845
rect 13262 21836 13268 21888
rect 13320 21876 13326 21888
rect 13541 21879 13599 21885
rect 13541 21876 13553 21879
rect 13320 21848 13553 21876
rect 13320 21836 13326 21848
rect 13541 21845 13553 21848
rect 13587 21845 13599 21879
rect 15010 21876 15016 21888
rect 14971 21848 15016 21876
rect 13541 21839 13599 21845
rect 15010 21836 15016 21848
rect 15068 21836 15074 21888
rect 17954 21876 17960 21888
rect 17915 21848 17960 21876
rect 17954 21836 17960 21848
rect 18012 21836 18018 21888
rect 25685 21879 25743 21885
rect 25685 21845 25697 21879
rect 25731 21876 25743 21879
rect 25866 21876 25872 21888
rect 25731 21848 25872 21876
rect 25731 21845 25743 21848
rect 25685 21839 25743 21845
rect 25866 21836 25872 21848
rect 25924 21836 25930 21888
rect 28626 21876 28632 21888
rect 28587 21848 28632 21876
rect 28626 21836 28632 21848
rect 28684 21836 28690 21888
rect 31573 21879 31631 21885
rect 31573 21845 31585 21879
rect 31619 21876 31631 21879
rect 31662 21876 31668 21888
rect 31619 21848 31668 21876
rect 31619 21845 31631 21848
rect 31573 21839 31631 21845
rect 31662 21836 31668 21848
rect 31720 21836 31726 21888
rect 34054 21876 34060 21888
rect 34015 21848 34060 21876
rect 34054 21836 34060 21848
rect 34112 21836 34118 21888
rect 1104 21786 38548 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 38548 21786
rect 1104 21712 38548 21734
rect 3878 21632 3884 21684
rect 3936 21672 3942 21684
rect 4065 21675 4123 21681
rect 4065 21672 4077 21675
rect 3936 21644 4077 21672
rect 3936 21632 3942 21644
rect 4065 21641 4077 21644
rect 4111 21641 4123 21675
rect 5534 21672 5540 21684
rect 5495 21644 5540 21672
rect 4065 21635 4123 21641
rect 1857 21607 1915 21613
rect 1857 21573 1869 21607
rect 1903 21604 1915 21607
rect 1903 21576 3096 21604
rect 1903 21573 1915 21576
rect 1857 21567 1915 21573
rect 1946 21536 1952 21548
rect 1907 21508 1952 21536
rect 1946 21496 1952 21508
rect 2004 21496 2010 21548
rect 2685 21539 2743 21545
rect 2685 21505 2697 21539
rect 2731 21536 2743 21539
rect 2866 21536 2872 21548
rect 2731 21508 2872 21536
rect 2731 21505 2743 21508
rect 2685 21499 2743 21505
rect 2866 21496 2872 21508
rect 2924 21496 2930 21548
rect 2038 21428 2044 21480
rect 2096 21468 2102 21480
rect 3068 21477 3096 21576
rect 2593 21471 2651 21477
rect 2593 21468 2605 21471
rect 2096 21440 2605 21468
rect 2096 21428 2102 21440
rect 2593 21437 2605 21440
rect 2639 21437 2651 21471
rect 2593 21431 2651 21437
rect 2961 21471 3019 21477
rect 2961 21437 2973 21471
rect 3007 21437 3019 21471
rect 2961 21431 3019 21437
rect 3053 21471 3111 21477
rect 3053 21437 3065 21471
rect 3099 21468 3111 21471
rect 3234 21468 3240 21480
rect 3099 21440 3240 21468
rect 3099 21437 3111 21440
rect 3053 21431 3111 21437
rect 2608 21332 2636 21431
rect 2976 21400 3004 21431
rect 3234 21428 3240 21440
rect 3292 21428 3298 21480
rect 4080 21468 4108 21635
rect 5534 21632 5540 21644
rect 5592 21632 5598 21684
rect 5905 21675 5963 21681
rect 5905 21641 5917 21675
rect 5951 21672 5963 21675
rect 6454 21672 6460 21684
rect 5951 21644 6460 21672
rect 5951 21641 5963 21644
rect 5905 21635 5963 21641
rect 5169 21607 5227 21613
rect 5169 21573 5181 21607
rect 5215 21604 5227 21607
rect 5920 21604 5948 21635
rect 6454 21632 6460 21644
rect 6512 21632 6518 21684
rect 9214 21632 9220 21684
rect 9272 21672 9278 21684
rect 9401 21675 9459 21681
rect 9401 21672 9413 21675
rect 9272 21644 9413 21672
rect 9272 21632 9278 21644
rect 9401 21641 9413 21644
rect 9447 21641 9459 21675
rect 9401 21635 9459 21641
rect 9750 21675 9808 21681
rect 9750 21641 9762 21675
rect 9796 21672 9808 21675
rect 9950 21672 9956 21684
rect 9796 21644 9956 21672
rect 9796 21641 9808 21644
rect 9750 21635 9808 21641
rect 9950 21632 9956 21644
rect 10008 21632 10014 21684
rect 10229 21675 10287 21681
rect 10229 21641 10241 21675
rect 10275 21672 10287 21675
rect 10594 21672 10600 21684
rect 10275 21644 10600 21672
rect 10275 21641 10287 21644
rect 10229 21635 10287 21641
rect 10594 21632 10600 21644
rect 10652 21632 10658 21684
rect 11146 21632 11152 21684
rect 11204 21672 11210 21684
rect 11977 21675 12035 21681
rect 11977 21672 11989 21675
rect 11204 21644 11989 21672
rect 11204 21632 11210 21644
rect 11977 21641 11989 21644
rect 12023 21641 12035 21675
rect 13998 21672 14004 21684
rect 11977 21635 12035 21641
rect 12452 21644 14004 21672
rect 5215 21576 5948 21604
rect 5215 21573 5227 21576
rect 5169 21567 5227 21573
rect 8570 21564 8576 21616
rect 8628 21564 8634 21616
rect 9125 21607 9183 21613
rect 9125 21573 9137 21607
rect 9171 21604 9183 21607
rect 9582 21604 9588 21616
rect 9171 21576 9588 21604
rect 9171 21573 9183 21576
rect 9125 21567 9183 21573
rect 4706 21496 4712 21548
rect 4764 21536 4770 21548
rect 4801 21539 4859 21545
rect 4801 21536 4813 21539
rect 4764 21508 4813 21536
rect 4764 21496 4770 21508
rect 4801 21505 4813 21508
rect 4847 21536 4859 21539
rect 6641 21539 6699 21545
rect 6641 21536 6653 21539
rect 4847 21508 6653 21536
rect 4847 21505 4859 21508
rect 4801 21499 4859 21505
rect 6641 21505 6653 21508
rect 6687 21536 6699 21539
rect 6825 21539 6883 21545
rect 6825 21536 6837 21539
rect 6687 21508 6837 21536
rect 6687 21505 6699 21508
rect 6641 21499 6699 21505
rect 6825 21505 6837 21508
rect 6871 21536 6883 21539
rect 7098 21536 7104 21548
rect 6871 21508 7104 21536
rect 6871 21505 6883 21508
rect 6825 21499 6883 21505
rect 7098 21496 7104 21508
rect 7156 21496 7162 21548
rect 7190 21496 7196 21548
rect 7248 21496 7254 21548
rect 7742 21536 7748 21548
rect 7300 21508 7748 21536
rect 4249 21471 4307 21477
rect 4249 21468 4261 21471
rect 4080 21440 4261 21468
rect 4249 21437 4261 21440
rect 4295 21437 4307 21471
rect 4249 21431 4307 21437
rect 5721 21471 5779 21477
rect 5721 21437 5733 21471
rect 5767 21468 5779 21471
rect 6181 21471 6239 21477
rect 6181 21468 6193 21471
rect 5767 21440 6193 21468
rect 5767 21437 5779 21440
rect 5721 21431 5779 21437
rect 6181 21437 6193 21440
rect 6227 21468 6239 21471
rect 6914 21468 6920 21480
rect 6227 21440 6920 21468
rect 6227 21437 6239 21440
rect 6181 21431 6239 21437
rect 6914 21428 6920 21440
rect 6972 21468 6978 21480
rect 7009 21471 7067 21477
rect 7009 21468 7021 21471
rect 6972 21440 7021 21468
rect 6972 21428 6978 21440
rect 7009 21437 7021 21440
rect 7055 21437 7067 21471
rect 7208 21468 7236 21496
rect 7009 21431 7067 21437
rect 7116 21440 7236 21468
rect 3142 21400 3148 21412
rect 2976 21372 3148 21400
rect 3142 21360 3148 21372
rect 3200 21400 3206 21412
rect 7116 21409 7144 21440
rect 3421 21403 3479 21409
rect 3421 21400 3433 21403
rect 3200 21372 3433 21400
rect 3200 21360 3206 21372
rect 3421 21369 3433 21372
rect 3467 21369 3479 21403
rect 3421 21363 3479 21369
rect 7101 21403 7159 21409
rect 7101 21369 7113 21403
rect 7147 21369 7159 21403
rect 7101 21363 7159 21369
rect 7193 21403 7251 21409
rect 7193 21369 7205 21403
rect 7239 21400 7251 21403
rect 7300 21400 7328 21508
rect 7742 21496 7748 21508
rect 7800 21536 7806 21548
rect 8588 21536 8616 21564
rect 7800 21508 8616 21536
rect 7800 21496 7806 21508
rect 7374 21428 7380 21480
rect 7432 21468 7438 21480
rect 8573 21471 8631 21477
rect 7432 21440 7972 21468
rect 7432 21428 7438 21440
rect 7558 21400 7564 21412
rect 7239 21372 7328 21400
rect 7519 21372 7564 21400
rect 7239 21369 7251 21372
rect 7193 21363 7251 21369
rect 7558 21360 7564 21372
rect 7616 21360 7622 21412
rect 7944 21409 7972 21440
rect 8573 21437 8585 21471
rect 8619 21468 8631 21471
rect 9140 21468 9168 21567
rect 9582 21564 9588 21576
rect 9640 21564 9646 21616
rect 9861 21607 9919 21613
rect 9861 21573 9873 21607
rect 9907 21604 9919 21607
rect 10502 21604 10508 21616
rect 9907 21576 10508 21604
rect 9907 21573 9919 21576
rect 9861 21567 9919 21573
rect 10502 21564 10508 21576
rect 10560 21564 10566 21616
rect 11057 21607 11115 21613
rect 11057 21573 11069 21607
rect 11103 21604 11115 21607
rect 11790 21604 11796 21616
rect 11103 21576 11796 21604
rect 11103 21573 11115 21576
rect 11057 21567 11115 21573
rect 9950 21536 9956 21548
rect 9911 21508 9956 21536
rect 9950 21496 9956 21508
rect 10008 21496 10014 21548
rect 10042 21496 10048 21548
rect 10100 21536 10106 21548
rect 11072 21536 11100 21567
rect 11790 21564 11796 21576
rect 11848 21604 11854 21616
rect 12452 21604 12480 21644
rect 13998 21632 14004 21644
rect 14056 21632 14062 21684
rect 15930 21632 15936 21684
rect 15988 21672 15994 21684
rect 16209 21675 16267 21681
rect 16209 21672 16221 21675
rect 15988 21644 16221 21672
rect 15988 21632 15994 21644
rect 16209 21641 16221 21644
rect 16255 21641 16267 21675
rect 16209 21635 16267 21641
rect 17678 21632 17684 21684
rect 17736 21672 17742 21684
rect 17773 21675 17831 21681
rect 17773 21672 17785 21675
rect 17736 21644 17785 21672
rect 17736 21632 17742 21644
rect 17773 21641 17785 21644
rect 17819 21641 17831 21675
rect 20165 21675 20223 21681
rect 20165 21672 20177 21675
rect 17773 21635 17831 21641
rect 19720 21644 20177 21672
rect 11848 21576 12480 21604
rect 11848 21564 11854 21576
rect 12710 21564 12716 21616
rect 12768 21604 12774 21616
rect 13357 21607 13415 21613
rect 13357 21604 13369 21607
rect 12768 21576 13369 21604
rect 12768 21564 12774 21576
rect 13357 21573 13369 21576
rect 13403 21573 13415 21607
rect 13357 21567 13415 21573
rect 10100 21508 11100 21536
rect 10100 21496 10106 21508
rect 12986 21496 12992 21548
rect 13044 21536 13050 21548
rect 13446 21536 13452 21548
rect 13044 21508 13452 21536
rect 13044 21496 13050 21508
rect 13446 21496 13452 21508
rect 13504 21496 13510 21548
rect 14093 21539 14151 21545
rect 14093 21505 14105 21539
rect 14139 21536 14151 21539
rect 15010 21536 15016 21548
rect 14139 21508 15016 21536
rect 14139 21505 14151 21508
rect 14093 21499 14151 21505
rect 15010 21496 15016 21508
rect 15068 21536 15074 21548
rect 15933 21539 15991 21545
rect 15933 21536 15945 21539
rect 15068 21508 15945 21536
rect 15068 21496 15074 21508
rect 15933 21505 15945 21508
rect 15979 21505 15991 21539
rect 15933 21499 15991 21505
rect 18693 21539 18751 21545
rect 18693 21505 18705 21539
rect 18739 21536 18751 21539
rect 18739 21508 19104 21536
rect 18739 21505 18751 21508
rect 18693 21499 18751 21505
rect 19076 21480 19104 21508
rect 8619 21440 9168 21468
rect 9585 21471 9643 21477
rect 8619 21437 8631 21440
rect 8573 21431 8631 21437
rect 9585 21437 9597 21471
rect 9631 21468 9643 21471
rect 9631 21440 9720 21468
rect 9631 21437 9643 21440
rect 9585 21431 9643 21437
rect 7929 21403 7987 21409
rect 7929 21369 7941 21403
rect 7975 21400 7987 21403
rect 9692 21400 9720 21440
rect 9766 21428 9772 21480
rect 9824 21468 9830 21480
rect 10597 21471 10655 21477
rect 10597 21468 10609 21471
rect 9824 21440 10609 21468
rect 9824 21428 9830 21440
rect 10597 21437 10609 21440
rect 10643 21437 10655 21471
rect 10597 21431 10655 21437
rect 11149 21471 11207 21477
rect 11149 21437 11161 21471
rect 11195 21468 11207 21471
rect 11238 21468 11244 21480
rect 11195 21440 11244 21468
rect 11195 21437 11207 21440
rect 11149 21431 11207 21437
rect 11238 21428 11244 21440
rect 11296 21428 11302 21480
rect 12529 21471 12587 21477
rect 12529 21437 12541 21471
rect 12575 21468 12587 21471
rect 12575 21440 13124 21468
rect 12575 21437 12587 21440
rect 12529 21431 12587 21437
rect 10042 21400 10048 21412
rect 7975 21372 8800 21400
rect 9692 21372 10048 21400
rect 7975 21369 7987 21372
rect 7929 21363 7987 21369
rect 3050 21332 3056 21344
rect 2608 21304 3056 21332
rect 3050 21292 3056 21304
rect 3108 21332 3114 21344
rect 4433 21335 4491 21341
rect 4433 21332 4445 21335
rect 3108 21304 4445 21332
rect 3108 21292 3114 21304
rect 4433 21301 4445 21304
rect 4479 21301 4491 21335
rect 4433 21295 4491 21301
rect 6638 21292 6644 21344
rect 6696 21332 6702 21344
rect 8018 21332 8024 21344
rect 6696 21304 8024 21332
rect 6696 21292 6702 21304
rect 8018 21292 8024 21304
rect 8076 21292 8082 21344
rect 8386 21332 8392 21344
rect 8347 21304 8392 21332
rect 8386 21292 8392 21304
rect 8444 21292 8450 21344
rect 8772 21341 8800 21372
rect 10042 21360 10048 21372
rect 10100 21360 10106 21412
rect 8757 21335 8815 21341
rect 8757 21301 8769 21335
rect 8803 21332 8815 21335
rect 8846 21332 8852 21344
rect 8803 21304 8852 21332
rect 8803 21301 8815 21304
rect 8757 21295 8815 21301
rect 8846 21292 8852 21304
rect 8904 21292 8910 21344
rect 11330 21332 11336 21344
rect 11291 21304 11336 21332
rect 11330 21292 11336 21304
rect 11388 21292 11394 21344
rect 11422 21292 11428 21344
rect 11480 21332 11486 21344
rect 11609 21335 11667 21341
rect 11609 21332 11621 21335
rect 11480 21304 11621 21332
rect 11480 21292 11486 21304
rect 11609 21301 11621 21304
rect 11655 21332 11667 21335
rect 12710 21332 12716 21344
rect 11655 21304 12716 21332
rect 11655 21301 11667 21304
rect 11609 21295 11667 21301
rect 12710 21292 12716 21304
rect 12768 21292 12774 21344
rect 13096 21341 13124 21440
rect 13262 21428 13268 21480
rect 13320 21468 13326 21480
rect 13541 21471 13599 21477
rect 13541 21468 13553 21471
rect 13320 21440 13553 21468
rect 13320 21428 13326 21440
rect 13541 21437 13553 21440
rect 13587 21437 13599 21471
rect 13541 21431 13599 21437
rect 13633 21471 13691 21477
rect 13633 21437 13645 21471
rect 13679 21437 13691 21471
rect 13633 21431 13691 21437
rect 13648 21400 13676 21431
rect 13906 21428 13912 21480
rect 13964 21468 13970 21480
rect 14829 21471 14887 21477
rect 14829 21468 14841 21471
rect 13964 21440 14841 21468
rect 13964 21428 13970 21440
rect 14829 21437 14841 21440
rect 14875 21468 14887 21471
rect 15470 21468 15476 21480
rect 14875 21440 15476 21468
rect 14875 21437 14887 21440
rect 14829 21431 14887 21437
rect 15470 21428 15476 21440
rect 15528 21428 15534 21480
rect 15654 21428 15660 21480
rect 15712 21468 15718 21480
rect 15749 21471 15807 21477
rect 15749 21468 15761 21471
rect 15712 21440 15761 21468
rect 15712 21428 15718 21440
rect 15749 21437 15761 21440
rect 15795 21468 15807 21471
rect 16577 21471 16635 21477
rect 16577 21468 16589 21471
rect 15795 21440 16589 21468
rect 15795 21437 15807 21440
rect 15749 21431 15807 21437
rect 16577 21437 16589 21440
rect 16623 21437 16635 21471
rect 16577 21431 16635 21437
rect 18785 21471 18843 21477
rect 18785 21437 18797 21471
rect 18831 21437 18843 21471
rect 19058 21468 19064 21480
rect 19019 21440 19064 21468
rect 18785 21431 18843 21437
rect 14921 21403 14979 21409
rect 13648 21372 14136 21400
rect 14108 21344 14136 21372
rect 14921 21369 14933 21403
rect 14967 21400 14979 21403
rect 15838 21400 15844 21412
rect 14967 21372 15844 21400
rect 14967 21369 14979 21372
rect 14921 21363 14979 21369
rect 15838 21360 15844 21372
rect 15896 21360 15902 21412
rect 13081 21335 13139 21341
rect 13081 21301 13093 21335
rect 13127 21332 13139 21335
rect 13446 21332 13452 21344
rect 13127 21304 13452 21332
rect 13127 21301 13139 21304
rect 13081 21295 13139 21301
rect 13446 21292 13452 21304
rect 13504 21292 13510 21344
rect 14090 21292 14096 21344
rect 14148 21332 14154 21344
rect 14369 21335 14427 21341
rect 14369 21332 14381 21335
rect 14148 21304 14381 21332
rect 14148 21292 14154 21304
rect 14369 21301 14381 21304
rect 14415 21332 14427 21335
rect 15102 21332 15108 21344
rect 14415 21304 15108 21332
rect 14415 21301 14427 21304
rect 14369 21295 14427 21301
rect 15102 21292 15108 21304
rect 15160 21292 15166 21344
rect 15930 21292 15936 21344
rect 15988 21332 15994 21344
rect 16574 21332 16580 21344
rect 15988 21304 16580 21332
rect 15988 21292 15994 21304
rect 16574 21292 16580 21304
rect 16632 21332 16638 21344
rect 16945 21335 17003 21341
rect 16945 21332 16957 21335
rect 16632 21304 16957 21332
rect 16632 21292 16638 21304
rect 16945 21301 16957 21304
rect 16991 21301 17003 21335
rect 17310 21332 17316 21344
rect 17271 21304 17316 21332
rect 16945 21295 17003 21301
rect 17310 21292 17316 21304
rect 17368 21292 17374 21344
rect 18138 21292 18144 21344
rect 18196 21332 18202 21344
rect 18233 21335 18291 21341
rect 18233 21332 18245 21335
rect 18196 21304 18245 21332
rect 18196 21292 18202 21304
rect 18233 21301 18245 21304
rect 18279 21332 18291 21335
rect 18598 21332 18604 21344
rect 18279 21304 18604 21332
rect 18279 21301 18291 21304
rect 18233 21295 18291 21301
rect 18598 21292 18604 21304
rect 18656 21292 18662 21344
rect 18800 21332 18828 21431
rect 19058 21428 19064 21440
rect 19116 21428 19122 21480
rect 19334 21428 19340 21480
rect 19392 21468 19398 21480
rect 19720 21468 19748 21644
rect 20165 21641 20177 21644
rect 20211 21672 20223 21675
rect 20254 21672 20260 21684
rect 20211 21644 20260 21672
rect 20211 21641 20223 21644
rect 20165 21635 20223 21641
rect 20254 21632 20260 21644
rect 20312 21632 20318 21684
rect 21177 21675 21235 21681
rect 21177 21641 21189 21675
rect 21223 21672 21235 21675
rect 21266 21672 21272 21684
rect 21223 21644 21272 21672
rect 21223 21641 21235 21644
rect 21177 21635 21235 21641
rect 21266 21632 21272 21644
rect 21324 21632 21330 21684
rect 26050 21632 26056 21684
rect 26108 21672 26114 21684
rect 27065 21675 27123 21681
rect 27065 21672 27077 21675
rect 26108 21644 27077 21672
rect 26108 21632 26114 21644
rect 27065 21641 27077 21644
rect 27111 21672 27123 21675
rect 27338 21672 27344 21684
rect 27111 21644 27344 21672
rect 27111 21641 27123 21644
rect 27065 21635 27123 21641
rect 27338 21632 27344 21644
rect 27396 21632 27402 21684
rect 28537 21675 28595 21681
rect 28537 21641 28549 21675
rect 28583 21672 28595 21675
rect 28810 21672 28816 21684
rect 28583 21644 28816 21672
rect 28583 21641 28595 21644
rect 28537 21635 28595 21641
rect 28810 21632 28816 21644
rect 28868 21632 28874 21684
rect 32769 21675 32827 21681
rect 32769 21641 32781 21675
rect 32815 21672 32827 21675
rect 32950 21672 32956 21684
rect 32815 21644 32956 21672
rect 32815 21641 32827 21644
rect 32769 21635 32827 21641
rect 32950 21632 32956 21644
rect 33008 21632 33014 21684
rect 33042 21632 33048 21684
rect 33100 21672 33106 21684
rect 35250 21672 35256 21684
rect 33100 21644 33145 21672
rect 35211 21644 35256 21672
rect 33100 21632 33106 21644
rect 35250 21632 35256 21644
rect 35308 21632 35314 21684
rect 35342 21632 35348 21684
rect 35400 21672 35406 21684
rect 37185 21675 37243 21681
rect 37185 21672 37197 21675
rect 35400 21644 37197 21672
rect 35400 21632 35406 21644
rect 37185 21641 37197 21644
rect 37231 21641 37243 21675
rect 37185 21635 37243 21641
rect 20809 21607 20867 21613
rect 20809 21573 20821 21607
rect 20855 21604 20867 21607
rect 22370 21604 22376 21616
rect 20855 21576 22376 21604
rect 20855 21573 20867 21576
rect 20809 21567 20867 21573
rect 22370 21564 22376 21576
rect 22428 21564 22434 21616
rect 23566 21564 23572 21616
rect 23624 21604 23630 21616
rect 24489 21607 24547 21613
rect 24489 21604 24501 21607
rect 23624 21576 24501 21604
rect 23624 21564 23630 21576
rect 24489 21573 24501 21576
rect 24535 21573 24547 21607
rect 26510 21604 26516 21616
rect 26471 21576 26516 21604
rect 24489 21567 24547 21573
rect 26510 21564 26516 21576
rect 26568 21564 26574 21616
rect 28169 21607 28227 21613
rect 28169 21573 28181 21607
rect 28215 21604 28227 21607
rect 29178 21604 29184 21616
rect 28215 21576 29184 21604
rect 28215 21573 28227 21576
rect 28169 21567 28227 21573
rect 29178 21564 29184 21576
rect 29236 21604 29242 21616
rect 29454 21604 29460 21616
rect 29236 21576 29460 21604
rect 29236 21564 29242 21576
rect 29454 21564 29460 21576
rect 29512 21564 29518 21616
rect 29638 21564 29644 21616
rect 29696 21604 29702 21616
rect 29914 21604 29920 21616
rect 29696 21576 29920 21604
rect 29696 21564 29702 21576
rect 29914 21564 29920 21576
rect 29972 21564 29978 21616
rect 30193 21607 30251 21613
rect 30193 21573 30205 21607
rect 30239 21604 30251 21607
rect 30282 21604 30288 21616
rect 30239 21576 30288 21604
rect 30239 21573 30251 21576
rect 30193 21567 30251 21573
rect 30282 21564 30288 21576
rect 30340 21604 30346 21616
rect 30469 21607 30527 21613
rect 30469 21604 30481 21607
rect 30340 21576 30481 21604
rect 30340 21564 30346 21576
rect 30469 21573 30481 21576
rect 30515 21604 30527 21607
rect 30515 21576 31248 21604
rect 30515 21573 30527 21576
rect 30469 21567 30527 21573
rect 23477 21539 23535 21545
rect 23477 21505 23489 21539
rect 23523 21536 23535 21539
rect 23842 21536 23848 21548
rect 23523 21508 23848 21536
rect 23523 21505 23535 21508
rect 23477 21499 23535 21505
rect 23842 21496 23848 21508
rect 23900 21496 23906 21548
rect 25866 21496 25872 21548
rect 25924 21536 25930 21548
rect 28258 21536 28264 21548
rect 25924 21508 26464 21536
rect 25924 21496 25930 21508
rect 21634 21468 21640 21480
rect 19392 21440 19748 21468
rect 21595 21440 21640 21468
rect 19392 21428 19398 21440
rect 21634 21428 21640 21440
rect 21692 21428 21698 21480
rect 24026 21468 24032 21480
rect 23987 21440 24032 21468
rect 24026 21428 24032 21440
rect 24084 21428 24090 21480
rect 24486 21468 24492 21480
rect 24447 21440 24492 21468
rect 24486 21428 24492 21440
rect 24544 21428 24550 21480
rect 25498 21468 25504 21480
rect 25459 21440 25504 21468
rect 25498 21428 25504 21440
rect 25556 21468 25562 21480
rect 25593 21471 25651 21477
rect 25593 21468 25605 21471
rect 25556 21440 25605 21468
rect 25556 21428 25562 21440
rect 25593 21437 25605 21440
rect 25639 21437 25651 21471
rect 25958 21468 25964 21480
rect 25919 21440 25964 21468
rect 25593 21431 25651 21437
rect 25958 21428 25964 21440
rect 26016 21428 26022 21480
rect 26436 21477 26464 21508
rect 28000 21508 28264 21536
rect 28000 21477 28028 21508
rect 28258 21496 28264 21508
rect 28316 21536 28322 21548
rect 28626 21536 28632 21548
rect 28316 21508 28632 21536
rect 28316 21496 28322 21508
rect 28626 21496 28632 21508
rect 28684 21536 28690 21548
rect 28813 21539 28871 21545
rect 28813 21536 28825 21539
rect 28684 21508 28825 21536
rect 28684 21496 28690 21508
rect 28813 21505 28825 21508
rect 28859 21505 28871 21539
rect 28813 21499 28871 21505
rect 26421 21471 26479 21477
rect 26421 21437 26433 21471
rect 26467 21437 26479 21471
rect 26421 21431 26479 21437
rect 27985 21471 28043 21477
rect 27985 21437 27997 21471
rect 28031 21437 28043 21471
rect 27985 21431 28043 21437
rect 29273 21471 29331 21477
rect 29273 21437 29285 21471
rect 29319 21468 29331 21471
rect 29546 21468 29552 21480
rect 29319 21440 29552 21468
rect 29319 21437 29331 21440
rect 29273 21431 29331 21437
rect 29546 21428 29552 21440
rect 29604 21468 29610 21480
rect 29604 21440 29868 21468
rect 29604 21428 29610 21440
rect 21266 21400 21272 21412
rect 21227 21372 21272 21400
rect 21266 21360 21272 21372
rect 21324 21360 21330 21412
rect 29840 21344 29868 21440
rect 29914 21428 29920 21480
rect 29972 21468 29978 21480
rect 30285 21471 30343 21477
rect 30285 21468 30297 21471
rect 29972 21440 30297 21468
rect 29972 21428 29978 21440
rect 30285 21437 30297 21440
rect 30331 21468 30343 21471
rect 30374 21468 30380 21480
rect 30331 21440 30380 21468
rect 30331 21437 30343 21440
rect 30285 21431 30343 21437
rect 30374 21428 30380 21440
rect 30432 21468 30438 21480
rect 31220 21477 31248 21576
rect 31294 21496 31300 21548
rect 31352 21536 31358 21548
rect 32401 21539 32459 21545
rect 31352 21508 32168 21536
rect 31352 21496 31358 21508
rect 30745 21471 30803 21477
rect 30745 21468 30757 21471
rect 30432 21440 30757 21468
rect 30432 21428 30438 21440
rect 30745 21437 30757 21440
rect 30791 21437 30803 21471
rect 30745 21431 30803 21437
rect 31205 21471 31263 21477
rect 31205 21437 31217 21471
rect 31251 21468 31263 21471
rect 31386 21468 31392 21480
rect 31251 21440 31392 21468
rect 31251 21437 31263 21440
rect 31205 21431 31263 21437
rect 31386 21428 31392 21440
rect 31444 21428 31450 21480
rect 31662 21468 31668 21480
rect 31623 21440 31668 21468
rect 31662 21428 31668 21440
rect 31720 21428 31726 21480
rect 32140 21477 32168 21508
rect 32401 21505 32413 21539
rect 32447 21536 32459 21539
rect 32766 21536 32772 21548
rect 32447 21508 32772 21536
rect 32447 21505 32459 21508
rect 32401 21499 32459 21505
rect 32766 21496 32772 21508
rect 32824 21496 32830 21548
rect 36081 21539 36139 21545
rect 36081 21536 36093 21539
rect 35728 21508 36093 21536
rect 35728 21480 35756 21508
rect 36081 21505 36093 21508
rect 36127 21505 36139 21539
rect 36081 21499 36139 21505
rect 32125 21471 32183 21477
rect 32125 21437 32137 21471
rect 32171 21437 32183 21471
rect 35710 21468 35716 21480
rect 35671 21440 35716 21468
rect 32125 21431 32183 21437
rect 35710 21428 35716 21440
rect 35768 21428 35774 21480
rect 35802 21428 35808 21480
rect 35860 21468 35866 21480
rect 35860 21440 35905 21468
rect 35860 21428 35866 21440
rect 19150 21332 19156 21344
rect 18800 21304 19156 21332
rect 19150 21292 19156 21304
rect 19208 21332 19214 21344
rect 19426 21332 19432 21344
rect 19208 21304 19432 21332
rect 19208 21292 19214 21304
rect 19426 21292 19432 21304
rect 19484 21292 19490 21344
rect 22370 21332 22376 21344
rect 22331 21304 22376 21332
rect 22370 21292 22376 21304
rect 22428 21292 22434 21344
rect 22646 21332 22652 21344
rect 22607 21304 22652 21332
rect 22646 21292 22652 21304
rect 22704 21292 22710 21344
rect 23109 21335 23167 21341
rect 23109 21301 23121 21335
rect 23155 21332 23167 21335
rect 23290 21332 23296 21344
rect 23155 21304 23296 21332
rect 23155 21301 23167 21304
rect 23109 21295 23167 21301
rect 23290 21292 23296 21304
rect 23348 21292 23354 21344
rect 27154 21292 27160 21344
rect 27212 21332 27218 21344
rect 27341 21335 27399 21341
rect 27341 21332 27353 21335
rect 27212 21304 27353 21332
rect 27212 21292 27218 21304
rect 27341 21301 27353 21304
rect 27387 21301 27399 21335
rect 27341 21295 27399 21301
rect 27614 21292 27620 21344
rect 27672 21332 27678 21344
rect 27709 21335 27767 21341
rect 27709 21332 27721 21335
rect 27672 21304 27721 21332
rect 27672 21292 27678 21304
rect 27709 21301 27721 21304
rect 27755 21301 27767 21335
rect 27709 21295 27767 21301
rect 29457 21335 29515 21341
rect 29457 21301 29469 21335
rect 29503 21332 29515 21335
rect 29546 21332 29552 21344
rect 29503 21304 29552 21332
rect 29503 21301 29515 21304
rect 29457 21295 29515 21301
rect 29546 21292 29552 21304
rect 29604 21292 29610 21344
rect 29822 21332 29828 21344
rect 29783 21304 29828 21332
rect 29822 21292 29828 21304
rect 29880 21292 29886 21344
rect 1104 21242 38548 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 38548 21242
rect 1104 21168 38548 21190
rect 3878 21128 3884 21140
rect 3839 21100 3884 21128
rect 3878 21088 3884 21100
rect 3936 21088 3942 21140
rect 4062 21088 4068 21140
rect 4120 21128 4126 21140
rect 4341 21131 4399 21137
rect 4341 21128 4353 21131
rect 4120 21100 4353 21128
rect 4120 21088 4126 21100
rect 4341 21097 4353 21100
rect 4387 21128 4399 21131
rect 4522 21128 4528 21140
rect 4387 21100 4528 21128
rect 4387 21097 4399 21100
rect 4341 21091 4399 21097
rect 4522 21088 4528 21100
rect 4580 21088 4586 21140
rect 5994 21128 6000 21140
rect 5955 21100 6000 21128
rect 5994 21088 6000 21100
rect 6052 21088 6058 21140
rect 6914 21128 6920 21140
rect 6875 21100 6920 21128
rect 6914 21088 6920 21100
rect 6972 21128 6978 21140
rect 7285 21131 7343 21137
rect 7285 21128 7297 21131
rect 6972 21100 7297 21128
rect 6972 21088 6978 21100
rect 7285 21097 7297 21100
rect 7331 21097 7343 21131
rect 7285 21091 7343 21097
rect 7558 21088 7564 21140
rect 7616 21128 7622 21140
rect 9125 21131 9183 21137
rect 9125 21128 9137 21131
rect 7616 21100 9137 21128
rect 7616 21088 7622 21100
rect 9125 21097 9137 21100
rect 9171 21097 9183 21131
rect 9125 21091 9183 21097
rect 9398 21088 9404 21140
rect 9456 21128 9462 21140
rect 9953 21131 10011 21137
rect 9953 21128 9965 21131
rect 9456 21100 9965 21128
rect 9456 21088 9462 21100
rect 9953 21097 9965 21100
rect 9999 21128 10011 21131
rect 10689 21131 10747 21137
rect 10689 21128 10701 21131
rect 9999 21100 10701 21128
rect 9999 21097 10011 21100
rect 9953 21091 10011 21097
rect 10689 21097 10701 21100
rect 10735 21097 10747 21131
rect 12618 21128 12624 21140
rect 12579 21100 12624 21128
rect 10689 21091 10747 21097
rect 12618 21088 12624 21100
rect 12676 21088 12682 21140
rect 14826 21088 14832 21140
rect 14884 21128 14890 21140
rect 15102 21128 15108 21140
rect 14884 21100 15108 21128
rect 14884 21088 14890 21100
rect 15102 21088 15108 21100
rect 15160 21088 15166 21140
rect 15378 21088 15384 21140
rect 15436 21128 15442 21140
rect 15473 21131 15531 21137
rect 15473 21128 15485 21131
rect 15436 21100 15485 21128
rect 15436 21088 15442 21100
rect 15473 21097 15485 21100
rect 15519 21097 15531 21131
rect 15473 21091 15531 21097
rect 16022 21088 16028 21140
rect 16080 21128 16086 21140
rect 16117 21131 16175 21137
rect 16117 21128 16129 21131
rect 16080 21100 16129 21128
rect 16080 21088 16086 21100
rect 16117 21097 16129 21100
rect 16163 21097 16175 21131
rect 16117 21091 16175 21097
rect 16758 21088 16764 21140
rect 16816 21128 16822 21140
rect 16853 21131 16911 21137
rect 16853 21128 16865 21131
rect 16816 21100 16865 21128
rect 16816 21088 16822 21100
rect 16853 21097 16865 21100
rect 16899 21097 16911 21131
rect 16853 21091 16911 21097
rect 22370 21088 22376 21140
rect 22428 21128 22434 21140
rect 24029 21131 24087 21137
rect 24029 21128 24041 21131
rect 22428 21100 24041 21128
rect 22428 21088 22434 21100
rect 24029 21097 24041 21100
rect 24075 21128 24087 21131
rect 24486 21128 24492 21140
rect 24075 21100 24492 21128
rect 24075 21097 24087 21100
rect 24029 21091 24087 21097
rect 3142 21060 3148 21072
rect 3103 21032 3148 21060
rect 3142 21020 3148 21032
rect 3200 21020 3206 21072
rect 6270 21060 6276 21072
rect 5552 21032 6276 21060
rect 1765 20995 1823 21001
rect 1765 20961 1777 20995
rect 1811 20992 1823 20995
rect 1854 20992 1860 21004
rect 1811 20964 1860 20992
rect 1811 20961 1823 20964
rect 1765 20955 1823 20961
rect 1854 20952 1860 20964
rect 1912 20952 1918 21004
rect 4801 20995 4859 21001
rect 4801 20961 4813 20995
rect 4847 20961 4859 20995
rect 4801 20955 4859 20961
rect 1489 20927 1547 20933
rect 1489 20893 1501 20927
rect 1535 20924 1547 20927
rect 1946 20924 1952 20936
rect 1535 20896 1952 20924
rect 1535 20893 1547 20896
rect 1489 20887 1547 20893
rect 1946 20884 1952 20896
rect 2004 20884 2010 20936
rect 4816 20924 4844 20955
rect 4890 20952 4896 21004
rect 4948 20992 4954 21004
rect 5552 21001 5580 21032
rect 6270 21020 6276 21032
rect 6328 21020 6334 21072
rect 7469 21063 7527 21069
rect 7469 21029 7481 21063
rect 7515 21060 7527 21063
rect 8202 21060 8208 21072
rect 7515 21032 8208 21060
rect 7515 21029 7527 21032
rect 7469 21023 7527 21029
rect 8202 21020 8208 21032
rect 8260 21020 8266 21072
rect 9214 21020 9220 21072
rect 9272 21060 9278 21072
rect 9858 21060 9864 21072
rect 9272 21032 9864 21060
rect 9272 21020 9278 21032
rect 9858 21020 9864 21032
rect 9916 21020 9922 21072
rect 10045 21063 10103 21069
rect 10045 21029 10057 21063
rect 10091 21060 10103 21063
rect 10318 21060 10324 21072
rect 10091 21032 10324 21060
rect 10091 21029 10103 21032
rect 10045 21023 10103 21029
rect 10318 21020 10324 21032
rect 10376 21020 10382 21072
rect 10413 21063 10471 21069
rect 10413 21029 10425 21063
rect 10459 21060 10471 21063
rect 10502 21060 10508 21072
rect 10459 21032 10508 21060
rect 10459 21029 10471 21032
rect 10413 21023 10471 21029
rect 10502 21020 10508 21032
rect 10560 21020 10566 21072
rect 14642 21060 14648 21072
rect 14603 21032 14648 21060
rect 14642 21020 14648 21032
rect 14700 21020 14706 21072
rect 24228 21069 24256 21100
rect 24486 21088 24492 21100
rect 24544 21088 24550 21140
rect 25685 21131 25743 21137
rect 25685 21097 25697 21131
rect 25731 21128 25743 21131
rect 25958 21128 25964 21140
rect 25731 21100 25964 21128
rect 25731 21097 25743 21100
rect 25685 21091 25743 21097
rect 25958 21088 25964 21100
rect 26016 21128 26022 21140
rect 26694 21128 26700 21140
rect 26016 21100 26700 21128
rect 26016 21088 26022 21100
rect 26694 21088 26700 21100
rect 26752 21088 26758 21140
rect 30193 21131 30251 21137
rect 30193 21097 30205 21131
rect 30239 21128 30251 21131
rect 30466 21128 30472 21140
rect 30239 21100 30472 21128
rect 30239 21097 30251 21100
rect 30193 21091 30251 21097
rect 30466 21088 30472 21100
rect 30524 21088 30530 21140
rect 35250 21128 35256 21140
rect 34900 21100 35256 21128
rect 24213 21063 24271 21069
rect 24213 21029 24225 21063
rect 24259 21029 24271 21063
rect 24213 21023 24271 21029
rect 27617 21063 27675 21069
rect 27617 21029 27629 21063
rect 27663 21060 27675 21063
rect 28810 21060 28816 21072
rect 27663 21032 28816 21060
rect 27663 21029 27675 21032
rect 27617 21023 27675 21029
rect 28810 21020 28816 21032
rect 28868 21020 28874 21072
rect 33318 21060 33324 21072
rect 33279 21032 33324 21060
rect 33318 21020 33324 21032
rect 33376 21020 33382 21072
rect 5537 20995 5595 21001
rect 5537 20992 5549 20995
rect 4948 20964 5549 20992
rect 4948 20952 4954 20964
rect 5537 20961 5549 20964
rect 5583 20961 5595 20995
rect 5537 20955 5595 20961
rect 5626 20952 5632 21004
rect 5684 20992 5690 21004
rect 6178 20992 6184 21004
rect 5684 20964 5729 20992
rect 6139 20964 6184 20992
rect 5684 20952 5690 20964
rect 6178 20952 6184 20964
rect 6236 20952 6242 21004
rect 7377 20995 7435 21001
rect 7377 20961 7389 20995
rect 7423 20992 7435 20995
rect 7650 20992 7656 21004
rect 7423 20964 7656 20992
rect 7423 20961 7435 20964
rect 7377 20955 7435 20961
rect 7650 20952 7656 20964
rect 7708 20952 7714 21004
rect 11054 20952 11060 21004
rect 11112 20992 11118 21004
rect 11241 20995 11299 21001
rect 11241 20992 11253 20995
rect 11112 20964 11253 20992
rect 11112 20952 11118 20964
rect 11241 20961 11253 20964
rect 11287 20961 11299 20995
rect 11422 20992 11428 21004
rect 11383 20964 11428 20992
rect 11241 20955 11299 20961
rect 11422 20952 11428 20964
rect 11480 20952 11486 21004
rect 13906 20992 13912 21004
rect 13867 20964 13912 20992
rect 13906 20952 13912 20964
rect 13964 20952 13970 21004
rect 14182 20992 14188 21004
rect 14143 20964 14188 20992
rect 14182 20952 14188 20964
rect 14240 20952 14246 21004
rect 15289 20995 15347 21001
rect 15289 20961 15301 20995
rect 15335 20992 15347 20995
rect 15378 20992 15384 21004
rect 15335 20964 15384 20992
rect 15335 20961 15347 20964
rect 15289 20955 15347 20961
rect 15378 20952 15384 20964
rect 15436 20952 15442 21004
rect 17218 20992 17224 21004
rect 17179 20964 17224 20992
rect 17218 20952 17224 20964
rect 17276 20952 17282 21004
rect 17586 20992 17592 21004
rect 17547 20964 17592 20992
rect 17586 20952 17592 20964
rect 17644 20952 17650 21004
rect 17773 20995 17831 21001
rect 17773 20961 17785 20995
rect 17819 20992 17831 20995
rect 18322 20992 18328 21004
rect 17819 20964 18328 20992
rect 17819 20961 17831 20964
rect 17773 20955 17831 20961
rect 18322 20952 18328 20964
rect 18380 20952 18386 21004
rect 18598 20992 18604 21004
rect 18559 20964 18604 20992
rect 18598 20952 18604 20964
rect 18656 20952 18662 21004
rect 20441 20995 20499 21001
rect 20441 20961 20453 20995
rect 20487 20992 20499 20995
rect 20622 20992 20628 21004
rect 20487 20964 20628 20992
rect 20487 20961 20499 20964
rect 20441 20955 20499 20961
rect 20622 20952 20628 20964
rect 20680 20952 20686 21004
rect 22646 20992 22652 21004
rect 22607 20964 22652 20992
rect 22646 20952 22652 20964
rect 22704 20952 22710 21004
rect 23014 20952 23020 21004
rect 23072 20992 23078 21004
rect 23109 20995 23167 21001
rect 23109 20992 23121 20995
rect 23072 20964 23121 20992
rect 23072 20952 23078 20964
rect 23109 20961 23121 20964
rect 23155 20961 23167 20995
rect 23109 20955 23167 20961
rect 24670 20952 24676 21004
rect 24728 20992 24734 21004
rect 25041 20995 25099 21001
rect 25041 20992 25053 20995
rect 24728 20964 25053 20992
rect 24728 20952 24734 20964
rect 25041 20961 25053 20964
rect 25087 20961 25099 20995
rect 25041 20955 25099 20961
rect 26418 20952 26424 21004
rect 26476 20992 26482 21004
rect 26513 20995 26571 21001
rect 26513 20992 26525 20995
rect 26476 20964 26525 20992
rect 26476 20952 26482 20964
rect 26513 20961 26525 20964
rect 26559 20961 26571 20995
rect 28442 20992 28448 21004
rect 28403 20964 28448 20992
rect 26513 20955 26571 20961
rect 28442 20952 28448 20964
rect 28500 20952 28506 21004
rect 28534 20952 28540 21004
rect 28592 20992 28598 21004
rect 28905 20995 28963 21001
rect 28905 20992 28917 20995
rect 28592 20964 28917 20992
rect 28592 20952 28598 20964
rect 28905 20961 28917 20964
rect 28951 20992 28963 20995
rect 29086 20992 29092 21004
rect 28951 20964 29092 20992
rect 28951 20961 28963 20964
rect 28905 20955 28963 20961
rect 29086 20952 29092 20964
rect 29144 20992 29150 21004
rect 29457 20995 29515 21001
rect 29457 20992 29469 20995
rect 29144 20964 29469 20992
rect 29144 20952 29150 20964
rect 29457 20961 29469 20964
rect 29503 20961 29515 20995
rect 29457 20955 29515 20961
rect 29822 20952 29828 21004
rect 29880 20992 29886 21004
rect 30285 20995 30343 21001
rect 30285 20992 30297 20995
rect 29880 20964 30297 20992
rect 29880 20952 29886 20964
rect 30285 20961 30297 20964
rect 30331 20992 30343 20995
rect 30650 20992 30656 21004
rect 30331 20964 30656 20992
rect 30331 20961 30343 20964
rect 30285 20955 30343 20961
rect 30650 20952 30656 20964
rect 30708 20952 30714 21004
rect 32490 20952 32496 21004
rect 32548 20992 32554 21004
rect 32585 20995 32643 21001
rect 32585 20992 32597 20995
rect 32548 20964 32597 20992
rect 32548 20952 32554 20964
rect 32585 20961 32597 20964
rect 32631 20961 32643 20995
rect 33042 20992 33048 21004
rect 33003 20964 33048 20992
rect 32585 20955 32643 20961
rect 33042 20952 33048 20964
rect 33100 20952 33106 21004
rect 34900 21001 34928 21100
rect 35250 21088 35256 21100
rect 35308 21088 35314 21140
rect 36262 21128 36268 21140
rect 36223 21100 36268 21128
rect 36262 21088 36268 21100
rect 36320 21088 36326 21140
rect 34885 20995 34943 21001
rect 34885 20961 34897 20995
rect 34931 20961 34943 20995
rect 34885 20955 34943 20961
rect 5258 20924 5264 20936
rect 4816 20896 5264 20924
rect 5258 20884 5264 20896
rect 5316 20884 5322 20936
rect 7098 20924 7104 20936
rect 7059 20896 7104 20924
rect 7098 20884 7104 20896
rect 7156 20884 7162 20936
rect 7837 20927 7895 20933
rect 7837 20893 7849 20927
rect 7883 20893 7895 20927
rect 7837 20887 7895 20893
rect 4709 20859 4767 20865
rect 4709 20825 4721 20859
rect 4755 20856 4767 20859
rect 7006 20856 7012 20868
rect 4755 20828 7012 20856
rect 4755 20825 4767 20828
rect 4709 20819 4767 20825
rect 7006 20816 7012 20828
rect 7064 20856 7070 20868
rect 7852 20856 7880 20887
rect 9122 20884 9128 20936
rect 9180 20924 9186 20936
rect 9398 20924 9404 20936
rect 9180 20896 9404 20924
rect 9180 20884 9186 20896
rect 9398 20884 9404 20896
rect 9456 20924 9462 20936
rect 9677 20927 9735 20933
rect 9677 20924 9689 20927
rect 9456 20896 9689 20924
rect 9456 20884 9462 20896
rect 9677 20893 9689 20896
rect 9723 20893 9735 20927
rect 9677 20887 9735 20893
rect 10502 20884 10508 20936
rect 10560 20924 10566 20936
rect 12253 20927 12311 20933
rect 12253 20924 12265 20927
rect 10560 20896 12265 20924
rect 10560 20884 10566 20896
rect 12253 20893 12265 20896
rect 12299 20893 12311 20927
rect 13354 20924 13360 20936
rect 13315 20896 13360 20924
rect 12253 20887 12311 20893
rect 13354 20884 13360 20896
rect 13412 20884 13418 20936
rect 14369 20927 14427 20933
rect 14369 20893 14381 20927
rect 14415 20924 14427 20927
rect 14734 20924 14740 20936
rect 14415 20896 14740 20924
rect 14415 20893 14427 20896
rect 14369 20887 14427 20893
rect 7064 20828 7880 20856
rect 7064 20816 7070 20828
rect 13814 20816 13820 20868
rect 13872 20856 13878 20868
rect 14384 20856 14412 20887
rect 14734 20884 14740 20896
rect 14792 20884 14798 20936
rect 16942 20884 16948 20936
rect 17000 20924 17006 20936
rect 17037 20927 17095 20933
rect 17037 20924 17049 20927
rect 17000 20896 17049 20924
rect 17000 20884 17006 20896
rect 17037 20893 17049 20896
rect 17083 20893 17095 20927
rect 21634 20924 21640 20936
rect 21595 20896 21640 20924
rect 17037 20887 17095 20893
rect 21634 20884 21640 20896
rect 21692 20884 21698 20936
rect 22370 20924 22376 20936
rect 22331 20896 22376 20924
rect 22370 20884 22376 20896
rect 22428 20884 22434 20936
rect 22664 20924 22692 20952
rect 23661 20927 23719 20933
rect 23661 20924 23673 20927
rect 22664 20896 23673 20924
rect 23661 20893 23673 20896
rect 23707 20924 23719 20927
rect 24026 20924 24032 20936
rect 23707 20896 24032 20924
rect 23707 20893 23719 20896
rect 23661 20887 23719 20893
rect 24026 20884 24032 20896
rect 24084 20884 24090 20936
rect 24762 20924 24768 20936
rect 24723 20896 24768 20924
rect 24762 20884 24768 20896
rect 24820 20884 24826 20936
rect 25222 20924 25228 20936
rect 25183 20896 25228 20924
rect 25222 20884 25228 20896
rect 25280 20884 25286 20936
rect 28169 20927 28227 20933
rect 28169 20924 28181 20927
rect 27908 20896 28181 20924
rect 13872 20828 14412 20856
rect 13872 20816 13878 20828
rect 20254 20816 20260 20868
rect 20312 20856 20318 20868
rect 20625 20859 20683 20865
rect 20625 20856 20637 20859
rect 20312 20828 20637 20856
rect 20312 20816 20318 20828
rect 20625 20825 20637 20828
rect 20671 20825 20683 20859
rect 23106 20856 23112 20868
rect 23067 20828 23112 20856
rect 20625 20819 20683 20825
rect 23106 20816 23112 20828
rect 23164 20816 23170 20868
rect 27157 20859 27215 20865
rect 27157 20825 27169 20859
rect 27203 20856 27215 20859
rect 27614 20856 27620 20868
rect 27203 20828 27620 20856
rect 27203 20825 27215 20828
rect 27157 20819 27215 20825
rect 27614 20816 27620 20828
rect 27672 20816 27678 20868
rect 5442 20748 5448 20800
rect 5500 20788 5506 20800
rect 5810 20788 5816 20800
rect 5500 20760 5816 20788
rect 5500 20748 5506 20760
rect 5810 20748 5816 20760
rect 5868 20748 5874 20800
rect 7282 20748 7288 20800
rect 7340 20788 7346 20800
rect 8113 20791 8171 20797
rect 8113 20788 8125 20791
rect 7340 20760 8125 20788
rect 7340 20748 7346 20760
rect 8113 20757 8125 20760
rect 8159 20788 8171 20791
rect 8386 20788 8392 20800
rect 8159 20760 8392 20788
rect 8159 20757 8171 20760
rect 8113 20751 8171 20757
rect 8386 20748 8392 20760
rect 8444 20748 8450 20800
rect 8849 20791 8907 20797
rect 8849 20757 8861 20791
rect 8895 20788 8907 20791
rect 9122 20788 9128 20800
rect 8895 20760 9128 20788
rect 8895 20757 8907 20760
rect 8849 20751 8907 20757
rect 9122 20748 9128 20760
rect 9180 20748 9186 20800
rect 10318 20748 10324 20800
rect 10376 20788 10382 20800
rect 11057 20791 11115 20797
rect 11057 20788 11069 20791
rect 10376 20760 11069 20788
rect 10376 20748 10382 20760
rect 11057 20757 11069 20760
rect 11103 20757 11115 20791
rect 11057 20751 11115 20757
rect 12158 20748 12164 20800
rect 12216 20788 12222 20800
rect 13265 20791 13323 20797
rect 13265 20788 13277 20791
rect 12216 20760 13277 20788
rect 12216 20748 12222 20760
rect 13265 20757 13277 20760
rect 13311 20788 13323 20791
rect 13354 20788 13360 20800
rect 13311 20760 13360 20788
rect 13311 20757 13323 20760
rect 13265 20751 13323 20757
rect 13354 20748 13360 20760
rect 13412 20748 13418 20800
rect 13538 20748 13544 20800
rect 13596 20788 13602 20800
rect 15013 20791 15071 20797
rect 15013 20788 15025 20791
rect 13596 20760 15025 20788
rect 13596 20748 13602 20760
rect 15013 20757 15025 20760
rect 15059 20757 15071 20791
rect 15838 20788 15844 20800
rect 15799 20760 15844 20788
rect 15013 20751 15071 20757
rect 15838 20748 15844 20760
rect 15896 20748 15902 20800
rect 18233 20791 18291 20797
rect 18233 20757 18245 20791
rect 18279 20788 18291 20791
rect 18782 20788 18788 20800
rect 18279 20760 18788 20788
rect 18279 20757 18291 20760
rect 18233 20751 18291 20757
rect 18782 20748 18788 20760
rect 18840 20788 18846 20800
rect 19058 20788 19064 20800
rect 18840 20760 19064 20788
rect 18840 20748 18846 20760
rect 19058 20748 19064 20760
rect 19116 20748 19122 20800
rect 20070 20788 20076 20800
rect 20031 20760 20076 20788
rect 20070 20748 20076 20760
rect 20128 20788 20134 20800
rect 20438 20788 20444 20800
rect 20128 20760 20444 20788
rect 20128 20748 20134 20760
rect 20438 20748 20444 20760
rect 20496 20748 20502 20800
rect 21269 20791 21327 20797
rect 21269 20757 21281 20791
rect 21315 20788 21327 20791
rect 22278 20788 22284 20800
rect 21315 20760 22284 20788
rect 21315 20757 21327 20760
rect 21269 20751 21327 20757
rect 22278 20748 22284 20760
rect 22336 20748 22342 20800
rect 25682 20748 25688 20800
rect 25740 20788 25746 20800
rect 25961 20791 26019 20797
rect 25961 20788 25973 20791
rect 25740 20760 25973 20788
rect 25740 20748 25746 20760
rect 25961 20757 25973 20760
rect 26007 20757 26019 20791
rect 25961 20751 26019 20757
rect 27798 20748 27804 20800
rect 27856 20788 27862 20800
rect 27908 20797 27936 20896
rect 28169 20893 28181 20896
rect 28215 20893 28227 20927
rect 32306 20924 32312 20936
rect 32267 20896 32312 20924
rect 28169 20887 28227 20893
rect 32306 20884 32312 20896
rect 32364 20884 32370 20936
rect 35161 20927 35219 20933
rect 35161 20893 35173 20927
rect 35207 20924 35219 20927
rect 35250 20924 35256 20936
rect 35207 20896 35256 20924
rect 35207 20893 35219 20896
rect 35161 20887 35219 20893
rect 35250 20884 35256 20896
rect 35308 20884 35314 20936
rect 28718 20816 28724 20868
rect 28776 20856 28782 20868
rect 28997 20859 29055 20865
rect 28997 20856 29009 20859
rect 28776 20828 29009 20856
rect 28776 20816 28782 20828
rect 28997 20825 29009 20828
rect 29043 20825 29055 20859
rect 28997 20819 29055 20825
rect 27893 20791 27951 20797
rect 27893 20788 27905 20791
rect 27856 20760 27905 20788
rect 27856 20748 27862 20760
rect 27893 20757 27905 20760
rect 27939 20757 27951 20791
rect 30466 20788 30472 20800
rect 30427 20760 30472 20788
rect 27893 20751 27951 20757
rect 30466 20748 30472 20760
rect 30524 20748 30530 20800
rect 30837 20791 30895 20797
rect 30837 20757 30849 20791
rect 30883 20788 30895 20791
rect 31294 20788 31300 20800
rect 30883 20760 31300 20788
rect 30883 20757 30895 20760
rect 30837 20751 30895 20757
rect 31294 20748 31300 20760
rect 31352 20748 31358 20800
rect 31757 20791 31815 20797
rect 31757 20757 31769 20791
rect 31803 20788 31815 20791
rect 32122 20788 32128 20800
rect 31803 20760 32128 20788
rect 31803 20757 31815 20760
rect 31757 20751 31815 20757
rect 32122 20748 32128 20760
rect 32180 20748 32186 20800
rect 1104 20698 38548 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 38548 20698
rect 1104 20624 38548 20646
rect 3510 20584 3516 20596
rect 3160 20556 3516 20584
rect 3160 20460 3188 20556
rect 3510 20544 3516 20556
rect 3568 20544 3574 20596
rect 4614 20584 4620 20596
rect 4575 20556 4620 20584
rect 4614 20544 4620 20556
rect 4672 20544 4678 20596
rect 5258 20584 5264 20596
rect 5219 20556 5264 20584
rect 5258 20544 5264 20556
rect 5316 20544 5322 20596
rect 5997 20587 6055 20593
rect 5997 20553 6009 20587
rect 6043 20584 6055 20587
rect 6086 20584 6092 20596
rect 6043 20556 6092 20584
rect 6043 20553 6055 20556
rect 5997 20547 6055 20553
rect 4341 20519 4399 20525
rect 4341 20485 4353 20519
rect 4387 20516 4399 20519
rect 4890 20516 4896 20528
rect 4387 20488 4896 20516
rect 4387 20485 4399 20488
rect 4341 20479 4399 20485
rect 4890 20476 4896 20488
rect 4948 20476 4954 20528
rect 2406 20448 2412 20460
rect 2367 20420 2412 20448
rect 2406 20408 2412 20420
rect 2464 20408 2470 20460
rect 3142 20448 3148 20460
rect 3055 20420 3148 20448
rect 3142 20408 3148 20420
rect 3200 20408 3206 20460
rect 3234 20408 3240 20460
rect 3292 20448 3298 20460
rect 3329 20451 3387 20457
rect 3329 20448 3341 20451
rect 3292 20420 3341 20448
rect 3292 20408 3298 20420
rect 3329 20417 3341 20420
rect 3375 20417 3387 20451
rect 3329 20411 3387 20417
rect 3510 20408 3516 20460
rect 3568 20448 3574 20460
rect 5813 20451 5871 20457
rect 5813 20448 5825 20451
rect 3568 20420 5825 20448
rect 3568 20408 3574 20420
rect 5813 20417 5825 20420
rect 5859 20417 5871 20451
rect 5813 20411 5871 20417
rect 3050 20380 3056 20392
rect 3011 20352 3056 20380
rect 3050 20340 3056 20352
rect 3108 20340 3114 20392
rect 3421 20383 3479 20389
rect 3421 20349 3433 20383
rect 3467 20349 3479 20383
rect 3421 20343 3479 20349
rect 4433 20383 4491 20389
rect 4433 20349 4445 20383
rect 4479 20380 4491 20383
rect 4479 20352 4844 20380
rect 4479 20349 4491 20352
rect 4433 20343 4491 20349
rect 1949 20315 2007 20321
rect 1949 20281 1961 20315
rect 1995 20312 2007 20315
rect 3436 20312 3464 20343
rect 3694 20312 3700 20324
rect 1995 20284 3700 20312
rect 1995 20281 2007 20284
rect 1949 20275 2007 20281
rect 3694 20272 3700 20284
rect 3752 20272 3758 20324
rect 4816 20256 4844 20352
rect 4890 20340 4896 20392
rect 4948 20380 4954 20392
rect 5445 20383 5503 20389
rect 5445 20380 5457 20383
rect 4948 20352 5457 20380
rect 4948 20340 4954 20352
rect 5445 20349 5457 20352
rect 5491 20380 5503 20383
rect 6012 20380 6040 20547
rect 6086 20544 6092 20556
rect 6144 20544 6150 20596
rect 6641 20587 6699 20593
rect 6641 20553 6653 20587
rect 6687 20584 6699 20587
rect 6914 20584 6920 20596
rect 6687 20556 6920 20584
rect 6687 20553 6699 20556
rect 6641 20547 6699 20553
rect 6914 20544 6920 20556
rect 6972 20544 6978 20596
rect 7098 20584 7104 20596
rect 7011 20556 7104 20584
rect 7098 20544 7104 20556
rect 7156 20584 7162 20596
rect 9398 20584 9404 20596
rect 7156 20556 9404 20584
rect 7156 20544 7162 20556
rect 9398 20544 9404 20556
rect 9456 20544 9462 20596
rect 9858 20584 9864 20596
rect 9819 20556 9864 20584
rect 9858 20544 9864 20556
rect 9916 20544 9922 20596
rect 10486 20587 10544 20593
rect 10486 20553 10498 20587
rect 10532 20584 10544 20587
rect 12434 20584 12440 20596
rect 10532 20556 12440 20584
rect 10532 20553 10544 20556
rect 10486 20547 10544 20553
rect 12434 20544 12440 20556
rect 12492 20584 12498 20596
rect 12621 20587 12679 20593
rect 12621 20584 12633 20587
rect 12492 20556 12633 20584
rect 12492 20544 12498 20556
rect 12621 20553 12633 20556
rect 12667 20553 12679 20587
rect 12621 20547 12679 20553
rect 12710 20544 12716 20596
rect 12768 20584 12774 20596
rect 13081 20587 13139 20593
rect 13081 20584 13093 20587
rect 12768 20556 13093 20584
rect 12768 20544 12774 20556
rect 13081 20553 13093 20556
rect 13127 20584 13139 20587
rect 13814 20584 13820 20596
rect 13127 20556 13820 20584
rect 13127 20553 13139 20556
rect 13081 20547 13139 20553
rect 13814 20544 13820 20556
rect 13872 20544 13878 20596
rect 16942 20544 16948 20596
rect 17000 20584 17006 20596
rect 17037 20587 17095 20593
rect 17037 20584 17049 20587
rect 17000 20556 17049 20584
rect 17000 20544 17006 20556
rect 17037 20553 17049 20556
rect 17083 20553 17095 20587
rect 17037 20547 17095 20553
rect 17218 20544 17224 20596
rect 17276 20584 17282 20596
rect 17405 20587 17463 20593
rect 17405 20584 17417 20587
rect 17276 20556 17417 20584
rect 17276 20544 17282 20556
rect 17405 20553 17417 20556
rect 17451 20553 17463 20587
rect 18966 20584 18972 20596
rect 18927 20556 18972 20584
rect 17405 20547 17463 20553
rect 18966 20544 18972 20556
rect 19024 20544 19030 20596
rect 22370 20584 22376 20596
rect 22283 20556 22376 20584
rect 22370 20544 22376 20556
rect 22428 20584 22434 20596
rect 22738 20584 22744 20596
rect 22428 20556 22744 20584
rect 22428 20544 22434 20556
rect 22738 20544 22744 20556
rect 22796 20584 22802 20596
rect 24670 20584 24676 20596
rect 22796 20556 24676 20584
rect 22796 20544 22802 20556
rect 24670 20544 24676 20556
rect 24728 20544 24734 20596
rect 26418 20544 26424 20596
rect 26476 20584 26482 20596
rect 26513 20587 26571 20593
rect 26513 20584 26525 20587
rect 26476 20556 26525 20584
rect 26476 20544 26482 20556
rect 26513 20553 26525 20556
rect 26559 20553 26571 20587
rect 28442 20584 28448 20596
rect 28403 20556 28448 20584
rect 26513 20547 26571 20553
rect 28442 20544 28448 20556
rect 28500 20584 28506 20596
rect 28997 20587 29055 20593
rect 28997 20584 29009 20587
rect 28500 20556 29009 20584
rect 28500 20544 28506 20556
rect 28997 20553 29009 20556
rect 29043 20553 29055 20587
rect 30650 20584 30656 20596
rect 30611 20556 30656 20584
rect 28997 20547 29055 20553
rect 8662 20516 8668 20528
rect 8623 20488 8668 20516
rect 8662 20476 8668 20488
rect 8720 20516 8726 20528
rect 8720 20488 8800 20516
rect 8720 20476 8726 20488
rect 7926 20448 7932 20460
rect 7887 20420 7932 20448
rect 7926 20408 7932 20420
rect 7984 20408 7990 20460
rect 8772 20457 8800 20488
rect 9582 20476 9588 20528
rect 9640 20516 9646 20528
rect 10594 20516 10600 20528
rect 9640 20488 10600 20516
rect 9640 20476 9646 20488
rect 10594 20476 10600 20488
rect 10652 20476 10658 20528
rect 10778 20516 10784 20528
rect 10739 20488 10784 20516
rect 10778 20476 10784 20488
rect 10836 20476 10842 20528
rect 11422 20516 11428 20528
rect 11383 20488 11428 20516
rect 11422 20476 11428 20488
rect 11480 20476 11486 20528
rect 11793 20519 11851 20525
rect 11793 20485 11805 20519
rect 11839 20516 11851 20519
rect 11882 20516 11888 20528
rect 11839 20488 11888 20516
rect 11839 20485 11851 20488
rect 11793 20479 11851 20485
rect 11882 20476 11888 20488
rect 11940 20476 11946 20528
rect 13449 20519 13507 20525
rect 13449 20485 13461 20519
rect 13495 20516 13507 20519
rect 14182 20516 14188 20528
rect 13495 20488 14188 20516
rect 13495 20485 13507 20488
rect 13449 20479 13507 20485
rect 14182 20476 14188 20488
rect 14240 20516 14246 20528
rect 14461 20519 14519 20525
rect 14461 20516 14473 20519
rect 14240 20488 14473 20516
rect 14240 20476 14246 20488
rect 14461 20485 14473 20488
rect 14507 20485 14519 20519
rect 15654 20516 15660 20528
rect 15615 20488 15660 20516
rect 14461 20479 14519 20485
rect 15654 20476 15660 20488
rect 15712 20476 15718 20528
rect 16761 20519 16819 20525
rect 16761 20485 16773 20519
rect 16807 20516 16819 20519
rect 17586 20516 17592 20528
rect 16807 20488 17592 20516
rect 16807 20485 16819 20488
rect 16761 20479 16819 20485
rect 17586 20476 17592 20488
rect 17644 20476 17650 20528
rect 8757 20451 8815 20457
rect 8757 20417 8769 20451
rect 8803 20417 8815 20451
rect 8757 20411 8815 20417
rect 9674 20408 9680 20460
rect 9732 20448 9738 20460
rect 10137 20451 10195 20457
rect 10137 20448 10149 20451
rect 9732 20420 10149 20448
rect 9732 20408 9738 20420
rect 10137 20417 10149 20420
rect 10183 20448 10195 20451
rect 10689 20451 10747 20457
rect 10689 20448 10701 20451
rect 10183 20420 10701 20448
rect 10183 20417 10195 20420
rect 10137 20411 10195 20417
rect 10689 20417 10701 20420
rect 10735 20448 10747 20451
rect 11054 20448 11060 20460
rect 10735 20420 11060 20448
rect 10735 20417 10747 20420
rect 10689 20411 10747 20417
rect 11054 20408 11060 20420
rect 11112 20408 11118 20460
rect 17218 20448 17224 20460
rect 16040 20420 17224 20448
rect 16040 20392 16068 20420
rect 17218 20408 17224 20420
rect 17276 20448 17282 20460
rect 17773 20451 17831 20457
rect 17773 20448 17785 20451
rect 17276 20420 17785 20448
rect 17276 20408 17282 20420
rect 17773 20417 17785 20420
rect 17819 20417 17831 20451
rect 18984 20448 19012 20544
rect 25958 20516 25964 20528
rect 25919 20488 25964 20516
rect 25958 20476 25964 20488
rect 26016 20476 26022 20528
rect 19429 20451 19487 20457
rect 19429 20448 19441 20451
rect 18984 20420 19441 20448
rect 17773 20411 17831 20417
rect 19429 20417 19441 20420
rect 19475 20417 19487 20451
rect 19429 20411 19487 20417
rect 25590 20408 25596 20460
rect 25648 20448 25654 20460
rect 26973 20451 27031 20457
rect 26973 20448 26985 20451
rect 25648 20420 26985 20448
rect 25648 20408 25654 20420
rect 26973 20417 26985 20420
rect 27019 20448 27031 20451
rect 29012 20448 29040 20547
rect 30650 20544 30656 20556
rect 30708 20544 30714 20596
rect 35342 20544 35348 20596
rect 35400 20584 35406 20596
rect 35437 20587 35495 20593
rect 35437 20584 35449 20587
rect 35400 20556 35449 20584
rect 35400 20544 35406 20556
rect 35437 20553 35449 20556
rect 35483 20553 35495 20587
rect 35437 20547 35495 20553
rect 29822 20476 29828 20528
rect 29880 20516 29886 20528
rect 30101 20519 30159 20525
rect 30101 20516 30113 20519
rect 29880 20488 30113 20516
rect 29880 20476 29886 20488
rect 30101 20485 30113 20488
rect 30147 20485 30159 20519
rect 30101 20479 30159 20485
rect 31846 20476 31852 20528
rect 31904 20516 31910 20528
rect 32033 20519 32091 20525
rect 32033 20516 32045 20519
rect 31904 20488 32045 20516
rect 31904 20476 31910 20488
rect 32033 20485 32045 20488
rect 32079 20485 32091 20519
rect 32033 20479 32091 20485
rect 32490 20448 32496 20460
rect 27019 20420 27936 20448
rect 29012 20420 29684 20448
rect 27019 20417 27031 20420
rect 26973 20411 27031 20417
rect 27908 20392 27936 20420
rect 5491 20352 6040 20380
rect 5491 20349 5503 20352
rect 5445 20343 5503 20349
rect 6914 20340 6920 20392
rect 6972 20380 6978 20392
rect 7377 20383 7435 20389
rect 7377 20380 7389 20383
rect 6972 20352 7389 20380
rect 6972 20340 6978 20352
rect 7377 20349 7389 20352
rect 7423 20349 7435 20383
rect 7377 20343 7435 20349
rect 7466 20340 7472 20392
rect 7524 20380 7530 20392
rect 8941 20383 8999 20389
rect 7524 20352 7569 20380
rect 7524 20340 7530 20352
rect 8941 20349 8953 20383
rect 8987 20380 8999 20383
rect 9030 20380 9036 20392
rect 8987 20352 9036 20380
rect 8987 20349 8999 20352
rect 8941 20343 8999 20349
rect 9030 20340 9036 20352
rect 9088 20340 9094 20392
rect 9493 20383 9551 20389
rect 9493 20349 9505 20383
rect 9539 20380 9551 20383
rect 10321 20383 10379 20389
rect 10321 20380 10333 20383
rect 9539 20352 10333 20380
rect 9539 20349 9551 20352
rect 9493 20343 9551 20349
rect 10321 20349 10333 20352
rect 10367 20380 10379 20383
rect 10502 20380 10508 20392
rect 10367 20352 10508 20380
rect 10367 20349 10379 20352
rect 10321 20343 10379 20349
rect 10502 20340 10508 20352
rect 10560 20340 10566 20392
rect 13078 20340 13084 20392
rect 13136 20380 13142 20392
rect 13633 20383 13691 20389
rect 13633 20380 13645 20383
rect 13136 20352 13645 20380
rect 13136 20340 13142 20352
rect 13633 20349 13645 20352
rect 13679 20349 13691 20383
rect 13633 20343 13691 20349
rect 13817 20383 13875 20389
rect 13817 20349 13829 20383
rect 13863 20380 13875 20383
rect 13906 20380 13912 20392
rect 13863 20352 13912 20380
rect 13863 20349 13875 20352
rect 13817 20343 13875 20349
rect 13906 20340 13912 20352
rect 13964 20340 13970 20392
rect 14001 20383 14059 20389
rect 14001 20349 14013 20383
rect 14047 20349 14059 20383
rect 15838 20380 15844 20392
rect 15799 20352 15844 20380
rect 14001 20343 14059 20349
rect 7098 20312 7104 20324
rect 5644 20284 7104 20312
rect 2317 20247 2375 20253
rect 2317 20213 2329 20247
rect 2363 20244 2375 20247
rect 3234 20244 3240 20256
rect 2363 20216 3240 20244
rect 2363 20213 2375 20216
rect 2317 20207 2375 20213
rect 3234 20204 3240 20216
rect 3292 20204 3298 20256
rect 3970 20244 3976 20256
rect 3931 20216 3976 20244
rect 3970 20204 3976 20216
rect 4028 20204 4034 20256
rect 4798 20204 4804 20256
rect 4856 20244 4862 20256
rect 5644 20253 5672 20284
rect 7098 20272 7104 20284
rect 7156 20272 7162 20324
rect 7193 20315 7251 20321
rect 7193 20281 7205 20315
rect 7239 20312 7251 20315
rect 7282 20312 7288 20324
rect 7239 20284 7288 20312
rect 7239 20281 7251 20284
rect 7193 20275 7251 20281
rect 7282 20272 7288 20284
rect 7340 20272 7346 20324
rect 7553 20315 7611 20321
rect 7553 20312 7565 20315
rect 7392 20284 7565 20312
rect 7392 20256 7420 20284
rect 7553 20281 7565 20284
rect 7599 20281 7611 20315
rect 7553 20275 7611 20281
rect 7834 20272 7840 20324
rect 7892 20312 7898 20324
rect 9122 20312 9128 20324
rect 7892 20284 8340 20312
rect 9083 20284 9128 20312
rect 7892 20272 7898 20284
rect 4893 20247 4951 20253
rect 4893 20244 4905 20247
rect 4856 20216 4905 20244
rect 4856 20204 4862 20216
rect 4893 20213 4905 20216
rect 4939 20213 4951 20247
rect 4893 20207 4951 20213
rect 5629 20247 5687 20253
rect 5629 20213 5641 20247
rect 5675 20213 5687 20247
rect 5629 20207 5687 20213
rect 5813 20247 5871 20253
rect 5813 20213 5825 20247
rect 5859 20244 5871 20247
rect 7374 20244 7380 20256
rect 5859 20216 7380 20244
rect 5859 20213 5871 20216
rect 5813 20207 5871 20213
rect 7374 20204 7380 20216
rect 7432 20204 7438 20256
rect 7650 20204 7656 20256
rect 7708 20244 7714 20256
rect 8205 20247 8263 20253
rect 8205 20244 8217 20247
rect 7708 20216 8217 20244
rect 7708 20204 7714 20216
rect 8205 20213 8217 20216
rect 8251 20213 8263 20247
rect 8312 20244 8340 20284
rect 9122 20272 9128 20284
rect 9180 20272 9186 20324
rect 10594 20272 10600 20324
rect 10652 20312 10658 20324
rect 12069 20315 12127 20321
rect 12069 20312 12081 20315
rect 10652 20284 12081 20312
rect 10652 20272 10658 20284
rect 12069 20281 12081 20284
rect 12115 20281 12127 20315
rect 12069 20275 12127 20281
rect 13354 20272 13360 20324
rect 13412 20312 13418 20324
rect 14016 20312 14044 20343
rect 15838 20340 15844 20352
rect 15896 20340 15902 20392
rect 16022 20380 16028 20392
rect 15983 20352 16028 20380
rect 16022 20340 16028 20352
rect 16080 20340 16086 20392
rect 16209 20383 16267 20389
rect 16209 20349 16221 20383
rect 16255 20380 16267 20383
rect 17126 20380 17132 20392
rect 16255 20352 17132 20380
rect 16255 20349 16267 20352
rect 16209 20343 16267 20349
rect 14921 20315 14979 20321
rect 14921 20312 14933 20315
rect 13412 20284 14933 20312
rect 13412 20272 13418 20284
rect 14921 20281 14933 20284
rect 14967 20312 14979 20315
rect 16224 20312 16252 20343
rect 17126 20340 17132 20352
rect 17184 20340 17190 20392
rect 19150 20380 19156 20392
rect 19111 20352 19156 20380
rect 19150 20340 19156 20352
rect 19208 20340 19214 20392
rect 25041 20383 25099 20389
rect 25041 20349 25053 20383
rect 25087 20380 25099 20383
rect 25133 20383 25191 20389
rect 25133 20380 25145 20383
rect 25087 20352 25145 20380
rect 25087 20349 25099 20352
rect 25041 20343 25099 20349
rect 25133 20349 25145 20352
rect 25179 20349 25191 20383
rect 25682 20380 25688 20392
rect 25643 20352 25688 20380
rect 25133 20343 25191 20349
rect 20806 20312 20812 20324
rect 14967 20284 16252 20312
rect 20767 20284 20812 20312
rect 14967 20281 14979 20284
rect 14921 20275 14979 20281
rect 20806 20272 20812 20284
rect 20864 20272 20870 20324
rect 22554 20272 22560 20324
rect 22612 20312 22618 20324
rect 23014 20312 23020 20324
rect 22612 20284 23020 20312
rect 22612 20272 22618 20284
rect 23014 20272 23020 20284
rect 23072 20272 23078 20324
rect 23937 20315 23995 20321
rect 23937 20281 23949 20315
rect 23983 20312 23995 20315
rect 24762 20312 24768 20324
rect 23983 20284 24768 20312
rect 23983 20281 23995 20284
rect 23937 20275 23995 20281
rect 24762 20272 24768 20284
rect 24820 20272 24826 20324
rect 25148 20312 25176 20343
rect 25682 20340 25688 20352
rect 25740 20340 25746 20392
rect 25958 20380 25964 20392
rect 25919 20352 25964 20380
rect 25958 20340 25964 20352
rect 26016 20340 26022 20392
rect 27614 20380 27620 20392
rect 27575 20352 27620 20380
rect 27614 20340 27620 20352
rect 27672 20340 27678 20392
rect 27890 20380 27896 20392
rect 27851 20352 27896 20380
rect 27890 20340 27896 20352
rect 27948 20340 27954 20392
rect 28074 20380 28080 20392
rect 27987 20352 28080 20380
rect 28074 20340 28080 20352
rect 28132 20340 28138 20392
rect 29362 20380 29368 20392
rect 29323 20352 29368 20380
rect 29362 20340 29368 20352
rect 29420 20340 29426 20392
rect 29656 20389 29684 20420
rect 31588 20420 32496 20448
rect 29641 20383 29699 20389
rect 29641 20349 29653 20383
rect 29687 20349 29699 20383
rect 29641 20343 29699 20349
rect 30101 20383 30159 20389
rect 30101 20349 30113 20383
rect 30147 20349 30159 20383
rect 30101 20343 30159 20349
rect 31205 20383 31263 20389
rect 31205 20349 31217 20383
rect 31251 20349 31263 20383
rect 31205 20343 31263 20349
rect 26142 20312 26148 20324
rect 25148 20284 26148 20312
rect 26142 20272 26148 20284
rect 26200 20272 26206 20324
rect 26326 20272 26332 20324
rect 26384 20312 26390 20324
rect 27065 20315 27123 20321
rect 27065 20312 27077 20315
rect 26384 20284 27077 20312
rect 26384 20272 26390 20284
rect 27065 20281 27077 20284
rect 27111 20281 27123 20315
rect 27065 20275 27123 20281
rect 27154 20272 27160 20324
rect 27212 20312 27218 20324
rect 28092 20312 28120 20340
rect 27212 20284 28120 20312
rect 27212 20272 27218 20284
rect 29086 20272 29092 20324
rect 29144 20312 29150 20324
rect 30116 20312 30144 20343
rect 29144 20284 30144 20312
rect 29144 20272 29150 20284
rect 9033 20247 9091 20253
rect 9033 20244 9045 20247
rect 8312 20216 9045 20244
rect 8205 20207 8263 20213
rect 9033 20213 9045 20216
rect 9079 20244 9091 20247
rect 9306 20244 9312 20256
rect 9079 20216 9312 20244
rect 9079 20213 9091 20216
rect 9033 20207 9091 20213
rect 9306 20204 9312 20216
rect 9364 20204 9370 20256
rect 10962 20204 10968 20256
rect 11020 20244 11026 20256
rect 11146 20244 11152 20256
rect 11020 20216 11152 20244
rect 11020 20204 11026 20216
rect 11146 20204 11152 20216
rect 11204 20244 11210 20256
rect 11882 20244 11888 20256
rect 11204 20216 11888 20244
rect 11204 20204 11210 20216
rect 11882 20204 11888 20216
rect 11940 20204 11946 20256
rect 15289 20247 15347 20253
rect 15289 20213 15301 20247
rect 15335 20244 15347 20247
rect 15378 20244 15384 20256
rect 15335 20216 15384 20244
rect 15335 20213 15347 20216
rect 15289 20207 15347 20213
rect 15378 20204 15384 20216
rect 15436 20204 15442 20256
rect 18322 20244 18328 20256
rect 18283 20216 18328 20244
rect 18322 20204 18328 20216
rect 18380 20204 18386 20256
rect 18598 20244 18604 20256
rect 18559 20216 18604 20244
rect 18598 20204 18604 20216
rect 18656 20204 18662 20256
rect 20714 20204 20720 20256
rect 20772 20244 20778 20256
rect 21085 20247 21143 20253
rect 21085 20244 21097 20247
rect 20772 20216 21097 20244
rect 20772 20204 20778 20216
rect 21085 20213 21097 20216
rect 21131 20213 21143 20247
rect 21085 20207 21143 20213
rect 22094 20204 22100 20256
rect 22152 20244 22158 20256
rect 22646 20244 22652 20256
rect 22152 20216 22652 20244
rect 22152 20204 22158 20216
rect 22646 20204 22652 20216
rect 22704 20204 22710 20256
rect 24305 20247 24363 20253
rect 24305 20213 24317 20247
rect 24351 20244 24363 20247
rect 24486 20244 24492 20256
rect 24351 20216 24492 20244
rect 24351 20213 24363 20216
rect 24305 20207 24363 20213
rect 24486 20204 24492 20216
rect 24544 20204 24550 20256
rect 31110 20244 31116 20256
rect 31071 20216 31116 20244
rect 31110 20204 31116 20216
rect 31168 20244 31174 20256
rect 31220 20244 31248 20343
rect 31478 20340 31484 20392
rect 31536 20380 31542 20392
rect 31588 20389 31616 20420
rect 32490 20408 32496 20420
rect 32548 20408 32554 20460
rect 31573 20383 31631 20389
rect 31573 20380 31585 20383
rect 31536 20352 31585 20380
rect 31536 20340 31542 20352
rect 31573 20349 31585 20352
rect 31619 20349 31631 20383
rect 32122 20380 32128 20392
rect 32083 20352 32128 20380
rect 31573 20343 31631 20349
rect 32122 20340 32128 20352
rect 32180 20340 32186 20392
rect 32490 20272 32496 20324
rect 32548 20312 32554 20324
rect 32953 20315 33011 20321
rect 32953 20312 32965 20315
rect 32548 20284 32965 20312
rect 32548 20272 32554 20284
rect 32953 20281 32965 20284
rect 32999 20281 33011 20315
rect 32953 20275 33011 20281
rect 31168 20216 31248 20244
rect 31168 20204 31174 20216
rect 32306 20204 32312 20256
rect 32364 20244 32370 20256
rect 32585 20247 32643 20253
rect 32585 20244 32597 20247
rect 32364 20216 32597 20244
rect 32364 20204 32370 20216
rect 32585 20213 32597 20216
rect 32631 20213 32643 20247
rect 35158 20244 35164 20256
rect 35119 20216 35164 20244
rect 32585 20207 32643 20213
rect 35158 20204 35164 20216
rect 35216 20204 35222 20256
rect 1104 20154 38548 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 38548 20154
rect 1104 20080 38548 20102
rect 1946 20040 1952 20052
rect 1907 20012 1952 20040
rect 1946 20000 1952 20012
rect 2004 20000 2010 20052
rect 2501 20043 2559 20049
rect 2501 20009 2513 20043
rect 2547 20040 2559 20043
rect 2682 20040 2688 20052
rect 2547 20012 2688 20040
rect 2547 20009 2559 20012
rect 2501 20003 2559 20009
rect 2682 20000 2688 20012
rect 2740 20040 2746 20052
rect 3050 20040 3056 20052
rect 2740 20012 3056 20040
rect 2740 20000 2746 20012
rect 3050 20000 3056 20012
rect 3108 20000 3114 20052
rect 3510 20040 3516 20052
rect 3471 20012 3516 20040
rect 3510 20000 3516 20012
rect 3568 20000 3574 20052
rect 4614 20040 4620 20052
rect 4575 20012 4620 20040
rect 4614 20000 4620 20012
rect 4672 20000 4678 20052
rect 4893 20043 4951 20049
rect 4893 20009 4905 20043
rect 4939 20040 4951 20043
rect 5166 20040 5172 20052
rect 4939 20012 5172 20040
rect 4939 20009 4951 20012
rect 4893 20003 4951 20009
rect 5166 20000 5172 20012
rect 5224 20000 5230 20052
rect 6178 20040 6184 20052
rect 6139 20012 6184 20040
rect 6178 20000 6184 20012
rect 6236 20000 6242 20052
rect 6914 20000 6920 20052
rect 6972 20040 6978 20052
rect 7101 20043 7159 20049
rect 7101 20040 7113 20043
rect 6972 20012 7113 20040
rect 6972 20000 6978 20012
rect 7101 20009 7113 20012
rect 7147 20040 7159 20043
rect 7469 20043 7527 20049
rect 7469 20040 7481 20043
rect 7147 20012 7481 20040
rect 7147 20009 7159 20012
rect 7101 20003 7159 20009
rect 7469 20009 7481 20012
rect 7515 20040 7527 20043
rect 7834 20040 7840 20052
rect 7515 20012 7840 20040
rect 7515 20009 7527 20012
rect 7469 20003 7527 20009
rect 7834 20000 7840 20012
rect 7892 20000 7898 20052
rect 8294 20040 8300 20052
rect 8255 20012 8300 20040
rect 8294 20000 8300 20012
rect 8352 20000 8358 20052
rect 9398 20040 9404 20052
rect 9359 20012 9404 20040
rect 9398 20000 9404 20012
rect 9456 20000 9462 20052
rect 10042 20000 10048 20052
rect 10100 20040 10106 20052
rect 10597 20043 10655 20049
rect 10597 20040 10609 20043
rect 10100 20012 10609 20040
rect 10100 20000 10106 20012
rect 10597 20009 10609 20012
rect 10643 20040 10655 20043
rect 13538 20040 13544 20052
rect 10643 20012 13544 20040
rect 10643 20009 10655 20012
rect 10597 20003 10655 20009
rect 13538 20000 13544 20012
rect 13596 20000 13602 20052
rect 13633 20043 13691 20049
rect 13633 20009 13645 20043
rect 13679 20040 13691 20043
rect 13814 20040 13820 20052
rect 13679 20012 13820 20040
rect 13679 20009 13691 20012
rect 13633 20003 13691 20009
rect 13814 20000 13820 20012
rect 13872 20000 13878 20052
rect 19150 20040 19156 20052
rect 19111 20012 19156 20040
rect 19150 20000 19156 20012
rect 19208 20000 19214 20052
rect 24394 20000 24400 20052
rect 24452 20040 24458 20052
rect 24670 20040 24676 20052
rect 24452 20012 24676 20040
rect 24452 20000 24458 20012
rect 24670 20000 24676 20012
rect 24728 20000 24734 20052
rect 25225 20043 25283 20049
rect 25225 20009 25237 20043
rect 25271 20040 25283 20043
rect 25958 20040 25964 20052
rect 25271 20012 25964 20040
rect 25271 20009 25283 20012
rect 25225 20003 25283 20009
rect 25958 20000 25964 20012
rect 26016 20000 26022 20052
rect 26326 20040 26332 20052
rect 26287 20012 26332 20040
rect 26326 20000 26332 20012
rect 26384 20000 26390 20052
rect 27614 20040 27620 20052
rect 27575 20012 27620 20040
rect 27614 20000 27620 20012
rect 27672 20000 27678 20052
rect 28997 20043 29055 20049
rect 28997 20009 29009 20043
rect 29043 20040 29055 20043
rect 29086 20040 29092 20052
rect 29043 20012 29092 20040
rect 29043 20009 29055 20012
rect 28997 20003 29055 20009
rect 29086 20000 29092 20012
rect 29144 20000 29150 20052
rect 31478 20040 31484 20052
rect 31439 20012 31484 20040
rect 31478 20000 31484 20012
rect 31536 20000 31542 20052
rect 1673 19975 1731 19981
rect 1673 19941 1685 19975
rect 1719 19972 1731 19975
rect 1854 19972 1860 19984
rect 1719 19944 1860 19972
rect 1719 19941 1731 19944
rect 1673 19935 1731 19941
rect 1854 19932 1860 19944
rect 1912 19932 1918 19984
rect 2869 19975 2927 19981
rect 2869 19941 2881 19975
rect 2915 19972 2927 19975
rect 3142 19972 3148 19984
rect 2915 19944 3148 19972
rect 2915 19941 2927 19944
rect 2869 19935 2927 19941
rect 3142 19932 3148 19944
rect 3200 19932 3206 19984
rect 5258 19972 5264 19984
rect 5219 19944 5264 19972
rect 5258 19932 5264 19944
rect 5316 19932 5322 19984
rect 5902 19932 5908 19984
rect 5960 19972 5966 19984
rect 6825 19975 6883 19981
rect 6825 19972 6837 19975
rect 5960 19944 6837 19972
rect 5960 19932 5966 19944
rect 6825 19941 6837 19944
rect 6871 19972 6883 19975
rect 7374 19972 7380 19984
rect 6871 19944 7380 19972
rect 6871 19941 6883 19944
rect 6825 19935 6883 19941
rect 7374 19932 7380 19944
rect 7432 19932 7438 19984
rect 7653 19975 7711 19981
rect 7653 19941 7665 19975
rect 7699 19972 7711 19975
rect 7926 19972 7932 19984
rect 7699 19944 7932 19972
rect 7699 19941 7711 19944
rect 7653 19935 7711 19941
rect 7926 19932 7932 19944
rect 7984 19932 7990 19984
rect 11606 19972 11612 19984
rect 11567 19944 11612 19972
rect 11606 19932 11612 19944
rect 11664 19932 11670 19984
rect 15838 19972 15844 19984
rect 15799 19944 15844 19972
rect 15838 19932 15844 19944
rect 15896 19932 15902 19984
rect 25682 19932 25688 19984
rect 25740 19972 25746 19984
rect 25869 19975 25927 19981
rect 25869 19972 25881 19975
rect 25740 19944 25881 19972
rect 25740 19932 25746 19944
rect 25869 19941 25881 19944
rect 25915 19941 25927 19975
rect 25869 19935 25927 19941
rect 27816 19944 30144 19972
rect 4709 19907 4767 19913
rect 4709 19873 4721 19907
rect 4755 19904 4767 19907
rect 4755 19876 5304 19904
rect 4755 19873 4767 19876
rect 4709 19867 4767 19873
rect 5276 19712 5304 19876
rect 5534 19864 5540 19916
rect 5592 19904 5598 19916
rect 5721 19907 5779 19913
rect 5721 19904 5733 19907
rect 5592 19876 5733 19904
rect 5592 19864 5598 19876
rect 5721 19873 5733 19876
rect 5767 19873 5779 19907
rect 5721 19867 5779 19873
rect 5997 19907 6055 19913
rect 5997 19873 6009 19907
rect 6043 19904 6055 19907
rect 6178 19904 6184 19916
rect 6043 19876 6184 19904
rect 6043 19873 6055 19876
rect 5997 19867 6055 19873
rect 6178 19864 6184 19876
rect 6236 19904 6242 19916
rect 7558 19904 7564 19916
rect 6236 19876 7420 19904
rect 7519 19876 7564 19904
rect 6236 19864 6242 19876
rect 7282 19836 7288 19848
rect 7243 19808 7288 19836
rect 7282 19796 7288 19808
rect 7340 19796 7346 19848
rect 7392 19836 7420 19876
rect 7558 19864 7564 19876
rect 7616 19864 7622 19916
rect 9953 19907 10011 19913
rect 9953 19873 9965 19907
rect 9999 19904 10011 19907
rect 10778 19904 10784 19916
rect 9999 19876 10784 19904
rect 9999 19873 10011 19876
rect 9953 19867 10011 19873
rect 10778 19864 10784 19876
rect 10836 19864 10842 19916
rect 12342 19864 12348 19916
rect 12400 19904 12406 19916
rect 12437 19907 12495 19913
rect 12437 19904 12449 19907
rect 12400 19876 12449 19904
rect 12400 19864 12406 19876
rect 12437 19873 12449 19876
rect 12483 19904 12495 19907
rect 12710 19904 12716 19916
rect 12483 19876 12716 19904
rect 12483 19873 12495 19876
rect 12437 19867 12495 19873
rect 12710 19864 12716 19876
rect 12768 19864 12774 19916
rect 13906 19904 13912 19916
rect 13867 19876 13912 19904
rect 13906 19864 13912 19876
rect 13964 19864 13970 19916
rect 15378 19904 15384 19916
rect 15339 19876 15384 19904
rect 15378 19864 15384 19876
rect 15436 19864 15442 19916
rect 16942 19904 16948 19916
rect 16903 19876 16948 19904
rect 16942 19864 16948 19876
rect 17000 19864 17006 19916
rect 17037 19907 17095 19913
rect 17037 19873 17049 19907
rect 17083 19904 17095 19907
rect 17126 19904 17132 19916
rect 17083 19876 17132 19904
rect 17083 19873 17095 19876
rect 17037 19867 17095 19873
rect 17126 19864 17132 19876
rect 17184 19864 17190 19916
rect 17402 19904 17408 19916
rect 17363 19876 17408 19904
rect 17402 19864 17408 19876
rect 17460 19864 17466 19916
rect 17497 19907 17555 19913
rect 17497 19873 17509 19907
rect 17543 19904 17555 19907
rect 17586 19904 17592 19916
rect 17543 19876 17592 19904
rect 17543 19873 17555 19876
rect 17497 19867 17555 19873
rect 17586 19864 17592 19876
rect 17644 19864 17650 19916
rect 22094 19864 22100 19916
rect 22152 19904 22158 19916
rect 22373 19907 22431 19913
rect 22152 19876 22197 19904
rect 22152 19864 22158 19876
rect 22373 19873 22385 19907
rect 22419 19904 22431 19907
rect 22554 19904 22560 19916
rect 22419 19876 22560 19904
rect 22419 19873 22431 19876
rect 22373 19867 22431 19873
rect 22554 19864 22560 19876
rect 22612 19864 22618 19916
rect 24026 19904 24032 19916
rect 23987 19876 24032 19904
rect 24026 19864 24032 19876
rect 24084 19864 24090 19916
rect 24394 19904 24400 19916
rect 24355 19876 24400 19904
rect 24394 19864 24400 19876
rect 24452 19864 24458 19916
rect 25222 19864 25228 19916
rect 25280 19904 25286 19916
rect 25409 19907 25467 19913
rect 25409 19904 25421 19907
rect 25280 19876 25421 19904
rect 25280 19864 25286 19876
rect 25409 19873 25421 19876
rect 25455 19873 25467 19907
rect 25409 19867 25467 19873
rect 27430 19864 27436 19916
rect 27488 19904 27494 19916
rect 27816 19913 27844 19944
rect 30116 19916 30144 19944
rect 32490 19932 32496 19984
rect 32548 19972 32554 19984
rect 34241 19975 34299 19981
rect 32548 19944 33548 19972
rect 32548 19932 32554 19944
rect 27801 19907 27859 19913
rect 27801 19904 27813 19907
rect 27488 19876 27813 19904
rect 27488 19864 27494 19876
rect 27801 19873 27813 19876
rect 27847 19873 27859 19907
rect 27801 19867 27859 19873
rect 28353 19907 28411 19913
rect 28353 19873 28365 19907
rect 28399 19873 28411 19907
rect 28353 19867 28411 19873
rect 28537 19907 28595 19913
rect 28537 19873 28549 19907
rect 28583 19904 28595 19907
rect 28810 19904 28816 19916
rect 28583 19876 28816 19904
rect 28583 19873 28595 19876
rect 28537 19867 28595 19873
rect 8021 19839 8079 19845
rect 8021 19836 8033 19839
rect 7392 19808 8033 19836
rect 8021 19805 8033 19808
rect 8067 19805 8079 19839
rect 8021 19799 8079 19805
rect 10134 19796 10140 19848
rect 10192 19836 10198 19848
rect 10321 19839 10379 19845
rect 10192 19808 10272 19836
rect 10192 19796 10198 19808
rect 5813 19771 5871 19777
rect 5813 19737 5825 19771
rect 5859 19768 5871 19771
rect 6454 19768 6460 19780
rect 5859 19740 6460 19768
rect 5859 19737 5871 19740
rect 5813 19731 5871 19737
rect 6454 19728 6460 19740
rect 6512 19728 6518 19780
rect 10244 19777 10272 19808
rect 10321 19805 10333 19839
rect 10367 19836 10379 19839
rect 10502 19836 10508 19848
rect 10367 19808 10508 19836
rect 10367 19805 10379 19808
rect 10321 19799 10379 19805
rect 10502 19796 10508 19808
rect 10560 19836 10566 19848
rect 11333 19839 11391 19845
rect 11333 19836 11345 19839
rect 10560 19808 11345 19836
rect 10560 19796 10566 19808
rect 11333 19805 11345 19808
rect 11379 19805 11391 19839
rect 12158 19836 12164 19848
rect 12119 19808 12164 19836
rect 11333 19799 11391 19805
rect 12158 19796 12164 19808
rect 12216 19796 12222 19848
rect 12526 19796 12532 19848
rect 12584 19836 12590 19848
rect 12621 19839 12679 19845
rect 12621 19836 12633 19839
rect 12584 19808 12633 19836
rect 12584 19796 12590 19808
rect 12621 19805 12633 19808
rect 12667 19805 12679 19839
rect 12621 19799 12679 19805
rect 13817 19839 13875 19845
rect 13817 19805 13829 19839
rect 13863 19836 13875 19839
rect 14550 19836 14556 19848
rect 13863 19808 14556 19836
rect 13863 19805 13875 19808
rect 13817 19799 13875 19805
rect 14550 19796 14556 19808
rect 14608 19796 14614 19848
rect 15286 19836 15292 19848
rect 15247 19808 15292 19836
rect 15286 19796 15292 19808
rect 15344 19836 15350 19848
rect 21726 19836 21732 19848
rect 15344 19808 16528 19836
rect 21687 19808 21732 19836
rect 15344 19796 15350 19808
rect 10229 19771 10287 19777
rect 10229 19737 10241 19771
rect 10275 19737 10287 19771
rect 10229 19731 10287 19737
rect 12802 19728 12808 19780
rect 12860 19768 12866 19780
rect 15105 19771 15163 19777
rect 15105 19768 15117 19771
rect 12860 19740 15117 19768
rect 12860 19728 12866 19740
rect 15105 19737 15117 19740
rect 15151 19768 15163 19771
rect 15654 19768 15660 19780
rect 15151 19740 15660 19768
rect 15151 19737 15163 19740
rect 15105 19731 15163 19737
rect 15654 19728 15660 19740
rect 15712 19728 15718 19780
rect 3878 19700 3884 19712
rect 3839 19672 3884 19700
rect 3878 19660 3884 19672
rect 3936 19660 3942 19712
rect 5258 19660 5264 19712
rect 5316 19700 5322 19712
rect 5629 19703 5687 19709
rect 5629 19700 5641 19703
rect 5316 19672 5641 19700
rect 5316 19660 5322 19672
rect 5629 19669 5641 19672
rect 5675 19700 5687 19703
rect 7190 19700 7196 19712
rect 5675 19672 7196 19700
rect 5675 19669 5687 19672
rect 5629 19663 5687 19669
rect 7190 19660 7196 19672
rect 7248 19660 7254 19712
rect 8849 19703 8907 19709
rect 8849 19669 8861 19703
rect 8895 19700 8907 19703
rect 9030 19700 9036 19712
rect 8895 19672 9036 19700
rect 8895 19669 8907 19672
rect 8849 19663 8907 19669
rect 9030 19660 9036 19672
rect 9088 19660 9094 19712
rect 9858 19660 9864 19712
rect 9916 19700 9922 19712
rect 10091 19703 10149 19709
rect 10091 19700 10103 19703
rect 9916 19672 10103 19700
rect 9916 19660 9922 19672
rect 10091 19669 10103 19672
rect 10137 19669 10149 19703
rect 11054 19700 11060 19712
rect 11015 19672 11060 19700
rect 10091 19663 10149 19669
rect 11054 19660 11060 19672
rect 11112 19660 11118 19712
rect 13078 19660 13084 19712
rect 13136 19700 13142 19712
rect 13173 19703 13231 19709
rect 13173 19700 13185 19703
rect 13136 19672 13185 19700
rect 13136 19660 13142 19672
rect 13173 19669 13185 19672
rect 13219 19669 13231 19703
rect 13173 19663 13231 19669
rect 13630 19660 13636 19712
rect 13688 19700 13694 19712
rect 14093 19703 14151 19709
rect 14093 19700 14105 19703
rect 13688 19672 14105 19700
rect 13688 19660 13694 19672
rect 14093 19669 14105 19672
rect 14139 19669 14151 19703
rect 14642 19700 14648 19712
rect 14603 19672 14648 19700
rect 14093 19663 14151 19669
rect 14642 19660 14648 19672
rect 14700 19660 14706 19712
rect 15470 19660 15476 19712
rect 15528 19700 15534 19712
rect 16206 19700 16212 19712
rect 15528 19672 16212 19700
rect 15528 19660 15534 19672
rect 16206 19660 16212 19672
rect 16264 19660 16270 19712
rect 16500 19700 16528 19808
rect 21726 19796 21732 19808
rect 21784 19796 21790 19848
rect 23661 19839 23719 19845
rect 23661 19805 23673 19839
rect 23707 19836 23719 19839
rect 23934 19836 23940 19848
rect 23707 19808 23940 19836
rect 23707 19805 23719 19808
rect 23661 19799 23719 19805
rect 23934 19796 23940 19808
rect 23992 19796 23998 19848
rect 28368 19836 28396 19867
rect 28810 19864 28816 19876
rect 28868 19864 28874 19916
rect 29733 19907 29791 19913
rect 29733 19873 29745 19907
rect 29779 19904 29791 19907
rect 30006 19904 30012 19916
rect 29779 19876 30012 19904
rect 29779 19873 29791 19876
rect 29733 19867 29791 19873
rect 30006 19864 30012 19876
rect 30064 19864 30070 19916
rect 30098 19864 30104 19916
rect 30156 19904 30162 19916
rect 30285 19907 30343 19913
rect 30156 19876 30201 19904
rect 30156 19864 30162 19876
rect 30285 19873 30297 19907
rect 30331 19873 30343 19907
rect 33134 19904 33140 19916
rect 33095 19876 33140 19904
rect 30285 19867 30343 19873
rect 28718 19836 28724 19848
rect 28368 19808 28724 19836
rect 28718 19796 28724 19808
rect 28776 19796 28782 19848
rect 30190 19796 30196 19848
rect 30248 19836 30254 19848
rect 30300 19836 30328 19867
rect 33134 19864 33140 19876
rect 33192 19864 33198 19916
rect 33520 19913 33548 19944
rect 34241 19941 34253 19975
rect 34287 19972 34299 19975
rect 34422 19972 34428 19984
rect 34287 19944 34428 19972
rect 34287 19941 34299 19944
rect 34241 19935 34299 19941
rect 34422 19932 34428 19944
rect 34480 19932 34486 19984
rect 33505 19907 33563 19913
rect 33505 19873 33517 19907
rect 33551 19873 33563 19907
rect 33962 19904 33968 19916
rect 33923 19876 33968 19904
rect 33505 19867 33563 19873
rect 33962 19864 33968 19876
rect 34020 19864 34026 19916
rect 35894 19904 35900 19916
rect 35855 19876 35900 19904
rect 35894 19864 35900 19876
rect 35952 19864 35958 19916
rect 30248 19808 30328 19836
rect 30248 19796 30254 19808
rect 32122 19796 32128 19848
rect 32180 19836 32186 19848
rect 32401 19839 32459 19845
rect 32401 19836 32413 19839
rect 32180 19808 32413 19836
rect 32180 19796 32186 19808
rect 32401 19805 32413 19808
rect 32447 19836 32459 19839
rect 33042 19836 33048 19848
rect 32447 19808 33048 19836
rect 32447 19805 32459 19808
rect 32401 19799 32459 19805
rect 33042 19796 33048 19808
rect 33100 19836 33106 19848
rect 35069 19839 35127 19845
rect 35069 19836 35081 19839
rect 33100 19808 35081 19836
rect 33100 19796 33106 19808
rect 35069 19805 35081 19808
rect 35115 19805 35127 19839
rect 35618 19836 35624 19848
rect 35579 19808 35624 19836
rect 35069 19799 35127 19805
rect 35618 19796 35624 19808
rect 35676 19796 35682 19848
rect 36078 19836 36084 19848
rect 36039 19808 36084 19836
rect 36078 19796 36084 19808
rect 36136 19796 36142 19848
rect 16577 19771 16635 19777
rect 16577 19737 16589 19771
rect 16623 19768 16635 19771
rect 17310 19768 17316 19780
rect 16623 19740 17316 19768
rect 16623 19737 16635 19740
rect 16577 19731 16635 19737
rect 17310 19728 17316 19740
rect 17368 19768 17374 19780
rect 17865 19771 17923 19777
rect 17865 19768 17877 19771
rect 17368 19740 17877 19768
rect 17368 19728 17374 19740
rect 17865 19737 17877 19740
rect 17911 19737 17923 19771
rect 17865 19731 17923 19737
rect 22002 19728 22008 19780
rect 22060 19768 22066 19780
rect 22373 19771 22431 19777
rect 22373 19768 22385 19771
rect 22060 19740 22385 19768
rect 22060 19728 22066 19740
rect 22373 19737 22385 19740
rect 22419 19737 22431 19771
rect 24302 19768 24308 19780
rect 24263 19740 24308 19768
rect 22373 19731 22431 19737
rect 24302 19728 24308 19740
rect 24360 19728 24366 19780
rect 25593 19771 25651 19777
rect 25593 19737 25605 19771
rect 25639 19768 25651 19771
rect 26050 19768 26056 19780
rect 25639 19740 26056 19768
rect 25639 19737 25651 19740
rect 25593 19731 25651 19737
rect 26050 19728 26056 19740
rect 26108 19728 26114 19780
rect 30282 19768 30288 19780
rect 30243 19740 30288 19768
rect 30282 19728 30288 19740
rect 30340 19728 30346 19780
rect 17402 19700 17408 19712
rect 16500 19672 17408 19700
rect 17402 19660 17408 19672
rect 17460 19660 17466 19712
rect 18414 19700 18420 19712
rect 18375 19672 18420 19700
rect 18414 19660 18420 19672
rect 18472 19660 18478 19712
rect 19797 19703 19855 19709
rect 19797 19669 19809 19703
rect 19843 19700 19855 19703
rect 19886 19700 19892 19712
rect 19843 19672 19892 19700
rect 19843 19669 19855 19672
rect 19797 19663 19855 19669
rect 19886 19660 19892 19672
rect 19944 19660 19950 19712
rect 26786 19700 26792 19712
rect 26747 19672 26792 19700
rect 26786 19660 26792 19672
rect 26844 19660 26850 19712
rect 27062 19700 27068 19712
rect 27023 19672 27068 19700
rect 27062 19660 27068 19672
rect 27120 19660 27126 19712
rect 29362 19700 29368 19712
rect 29323 19672 29368 19700
rect 29362 19660 29368 19672
rect 29420 19660 29426 19712
rect 31113 19703 31171 19709
rect 31113 19669 31125 19703
rect 31159 19700 31171 19703
rect 31478 19700 31484 19712
rect 31159 19672 31484 19700
rect 31159 19669 31171 19672
rect 31113 19663 31171 19669
rect 31478 19660 31484 19672
rect 31536 19660 31542 19712
rect 33042 19700 33048 19712
rect 33003 19672 33048 19700
rect 33042 19660 33048 19672
rect 33100 19660 33106 19712
rect 1104 19610 38548 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 38548 19610
rect 1104 19536 38548 19558
rect 1857 19499 1915 19505
rect 1857 19465 1869 19499
rect 1903 19496 1915 19499
rect 1946 19496 1952 19508
rect 1903 19468 1952 19496
rect 1903 19465 1915 19468
rect 1857 19459 1915 19465
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 3694 19496 3700 19508
rect 3655 19468 3700 19496
rect 3694 19456 3700 19468
rect 3752 19456 3758 19508
rect 7834 19496 7840 19508
rect 7795 19468 7840 19496
rect 7834 19456 7840 19468
rect 7892 19456 7898 19508
rect 8662 19456 8668 19508
rect 8720 19496 8726 19508
rect 8941 19499 8999 19505
rect 8941 19496 8953 19499
rect 8720 19468 8953 19496
rect 8720 19456 8726 19468
rect 8941 19465 8953 19468
rect 8987 19465 8999 19499
rect 10134 19496 10140 19508
rect 10095 19468 10140 19496
rect 8941 19459 8999 19465
rect 1964 19360 1992 19456
rect 2317 19363 2375 19369
rect 2317 19360 2329 19363
rect 1964 19332 2329 19360
rect 2317 19329 2329 19332
rect 2363 19329 2375 19363
rect 3418 19360 3424 19372
rect 2317 19323 2375 19329
rect 2792 19332 3424 19360
rect 2593 19295 2651 19301
rect 2593 19292 2605 19295
rect 2424 19264 2605 19292
rect 2225 19227 2283 19233
rect 2225 19193 2237 19227
rect 2271 19224 2283 19227
rect 2424 19224 2452 19264
rect 2593 19261 2605 19264
rect 2639 19292 2651 19295
rect 2792 19292 2820 19332
rect 3418 19320 3424 19332
rect 3476 19320 3482 19372
rect 4709 19363 4767 19369
rect 4709 19329 4721 19363
rect 4755 19360 4767 19363
rect 5258 19360 5264 19372
rect 4755 19332 5264 19360
rect 4755 19329 4767 19332
rect 4709 19323 4767 19329
rect 5258 19320 5264 19332
rect 5316 19320 5322 19372
rect 5534 19320 5540 19372
rect 5592 19360 5598 19372
rect 5905 19363 5963 19369
rect 5905 19360 5917 19363
rect 5592 19332 5917 19360
rect 5592 19320 5598 19332
rect 5905 19329 5917 19332
rect 5951 19329 5963 19363
rect 5905 19323 5963 19329
rect 6454 19320 6460 19372
rect 6512 19360 6518 19372
rect 7561 19363 7619 19369
rect 7561 19360 7573 19363
rect 6512 19332 7573 19360
rect 6512 19320 6518 19332
rect 7561 19329 7573 19332
rect 7607 19329 7619 19363
rect 8956 19360 8984 19459
rect 10134 19456 10140 19468
rect 10192 19456 10198 19508
rect 12710 19456 12716 19508
rect 12768 19496 12774 19508
rect 13078 19496 13084 19508
rect 12768 19468 13084 19496
rect 12768 19456 12774 19468
rect 13078 19456 13084 19468
rect 13136 19456 13142 19508
rect 16206 19456 16212 19508
rect 16264 19496 16270 19508
rect 17497 19499 17555 19505
rect 16264 19468 16712 19496
rect 16264 19456 16270 19468
rect 11422 19388 11428 19440
rect 11480 19428 11486 19440
rect 12066 19428 12072 19440
rect 11480 19400 12072 19428
rect 11480 19388 11486 19400
rect 12066 19388 12072 19400
rect 12124 19388 12130 19440
rect 16022 19388 16028 19440
rect 16080 19428 16086 19440
rect 16298 19428 16304 19440
rect 16080 19400 16304 19428
rect 16080 19388 16086 19400
rect 16298 19388 16304 19400
rect 16356 19388 16362 19440
rect 9125 19363 9183 19369
rect 9125 19360 9137 19363
rect 7561 19323 7619 19329
rect 7668 19332 8248 19360
rect 8956 19332 9137 19360
rect 2639 19264 2820 19292
rect 4341 19295 4399 19301
rect 2639 19261 2651 19264
rect 2593 19255 2651 19261
rect 4341 19261 4353 19295
rect 4387 19292 4399 19295
rect 5074 19292 5080 19304
rect 4387 19264 5080 19292
rect 4387 19261 4399 19264
rect 4341 19255 4399 19261
rect 5074 19252 5080 19264
rect 5132 19292 5138 19304
rect 6273 19295 6331 19301
rect 5132 19264 5580 19292
rect 5132 19252 5138 19264
rect 2271 19196 2452 19224
rect 2271 19193 2283 19196
rect 2225 19187 2283 19193
rect 4890 19184 4896 19236
rect 4948 19224 4954 19236
rect 5166 19224 5172 19236
rect 4948 19196 5172 19224
rect 4948 19184 4954 19196
rect 5166 19184 5172 19196
rect 5224 19184 5230 19236
rect 5258 19184 5264 19236
rect 5316 19224 5322 19236
rect 5552 19233 5580 19264
rect 6273 19261 6285 19295
rect 6319 19292 6331 19295
rect 6825 19295 6883 19301
rect 6825 19292 6837 19295
rect 6319 19264 6837 19292
rect 6319 19261 6331 19264
rect 6273 19255 6331 19261
rect 6825 19261 6837 19264
rect 6871 19292 6883 19295
rect 7282 19292 7288 19304
rect 6871 19264 7288 19292
rect 6871 19261 6883 19264
rect 6825 19255 6883 19261
rect 7282 19252 7288 19264
rect 7340 19292 7346 19304
rect 7668 19292 7696 19332
rect 7340 19264 7696 19292
rect 8220 19292 8248 19332
rect 9125 19329 9137 19332
rect 9171 19329 9183 19363
rect 9125 19323 9183 19329
rect 11517 19363 11575 19369
rect 11517 19329 11529 19363
rect 11563 19360 11575 19363
rect 12434 19360 12440 19372
rect 11563 19332 12440 19360
rect 11563 19329 11575 19332
rect 11517 19323 11575 19329
rect 12434 19320 12440 19332
rect 12492 19320 12498 19372
rect 15930 19320 15936 19372
rect 15988 19360 15994 19372
rect 16117 19363 16175 19369
rect 16117 19360 16129 19363
rect 15988 19332 16129 19360
rect 15988 19320 15994 19332
rect 16117 19329 16129 19332
rect 16163 19329 16175 19363
rect 16117 19323 16175 19329
rect 8220 19264 8340 19292
rect 7340 19252 7346 19264
rect 8312 19236 8340 19264
rect 9030 19252 9036 19304
rect 9088 19292 9094 19304
rect 9309 19295 9367 19301
rect 9309 19292 9321 19295
rect 9088 19264 9321 19292
rect 9088 19252 9094 19264
rect 9309 19261 9321 19264
rect 9355 19261 9367 19295
rect 9309 19255 9367 19261
rect 10781 19295 10839 19301
rect 10781 19261 10793 19295
rect 10827 19292 10839 19295
rect 11330 19292 11336 19304
rect 10827 19264 11336 19292
rect 10827 19261 10839 19264
rect 10781 19255 10839 19261
rect 11330 19252 11336 19264
rect 11388 19252 11394 19304
rect 12253 19295 12311 19301
rect 12253 19261 12265 19295
rect 12299 19292 12311 19295
rect 12342 19292 12348 19304
rect 12299 19264 12348 19292
rect 12299 19261 12311 19264
rect 12253 19255 12311 19261
rect 12342 19252 12348 19264
rect 12400 19252 12406 19304
rect 12618 19252 12624 19304
rect 12676 19292 12682 19304
rect 12802 19292 12808 19304
rect 12676 19264 12808 19292
rect 12676 19252 12682 19264
rect 12802 19252 12808 19264
rect 12860 19252 12866 19304
rect 12894 19252 12900 19304
rect 12952 19292 12958 19304
rect 14182 19292 14188 19304
rect 12952 19264 12997 19292
rect 14143 19264 14188 19292
rect 12952 19252 12958 19264
rect 14182 19252 14188 19264
rect 14240 19252 14246 19304
rect 14277 19295 14335 19301
rect 14277 19261 14289 19295
rect 14323 19261 14335 19295
rect 14734 19292 14740 19304
rect 14695 19264 14740 19292
rect 14277 19255 14335 19261
rect 5445 19227 5503 19233
rect 5445 19224 5457 19227
rect 5316 19196 5457 19224
rect 5316 19184 5322 19196
rect 5445 19193 5457 19196
rect 5491 19193 5503 19227
rect 5445 19187 5503 19193
rect 5537 19227 5595 19233
rect 5537 19193 5549 19227
rect 5583 19193 5595 19227
rect 7190 19224 7196 19236
rect 7151 19196 7196 19224
rect 5537 19187 5595 19193
rect 7190 19184 7196 19196
rect 7248 19184 7254 19236
rect 8294 19224 8300 19236
rect 8255 19196 8300 19224
rect 8294 19184 8300 19196
rect 8352 19184 8358 19236
rect 9214 19184 9220 19236
rect 9272 19224 9278 19236
rect 9493 19227 9551 19233
rect 9493 19224 9505 19227
rect 9272 19196 9505 19224
rect 9272 19184 9278 19196
rect 9493 19193 9505 19196
rect 9539 19193 9551 19227
rect 9858 19224 9864 19236
rect 9819 19196 9864 19224
rect 9493 19187 9551 19193
rect 9858 19184 9864 19196
rect 9916 19184 9922 19236
rect 11149 19227 11207 19233
rect 11149 19193 11161 19227
rect 11195 19224 11207 19227
rect 11606 19224 11612 19236
rect 11195 19196 11612 19224
rect 11195 19193 11207 19196
rect 11149 19187 11207 19193
rect 11606 19184 11612 19196
rect 11664 19184 11670 19236
rect 11885 19227 11943 19233
rect 11885 19193 11897 19227
rect 11931 19224 11943 19227
rect 12526 19224 12532 19236
rect 11931 19196 12532 19224
rect 11931 19193 11943 19196
rect 11885 19187 11943 19193
rect 12526 19184 12532 19196
rect 12584 19184 12590 19236
rect 12713 19227 12771 19233
rect 12713 19193 12725 19227
rect 12759 19224 12771 19227
rect 12912 19224 12940 19252
rect 12759 19196 12940 19224
rect 12759 19193 12771 19196
rect 12713 19187 12771 19193
rect 4798 19116 4804 19168
rect 4856 19156 4862 19168
rect 5077 19159 5135 19165
rect 5077 19156 5089 19159
rect 4856 19128 5089 19156
rect 4856 19116 4862 19128
rect 5077 19125 5089 19128
rect 5123 19156 5135 19159
rect 5353 19159 5411 19165
rect 5353 19156 5365 19159
rect 5123 19128 5365 19156
rect 5123 19125 5135 19128
rect 5077 19119 5135 19125
rect 5353 19125 5365 19128
rect 5399 19125 5411 19159
rect 5353 19119 5411 19125
rect 6641 19159 6699 19165
rect 6641 19125 6653 19159
rect 6687 19156 6699 19159
rect 7006 19156 7012 19168
rect 6687 19128 7012 19156
rect 6687 19125 6699 19128
rect 6641 19119 6699 19125
rect 7006 19116 7012 19128
rect 7064 19116 7070 19168
rect 7098 19116 7104 19168
rect 7156 19156 7162 19168
rect 8573 19159 8631 19165
rect 8573 19156 8585 19159
rect 7156 19128 8585 19156
rect 7156 19116 7162 19128
rect 8573 19125 8585 19128
rect 8619 19125 8631 19159
rect 9398 19156 9404 19168
rect 9359 19128 9404 19156
rect 8573 19119 8631 19125
rect 9398 19116 9404 19128
rect 9456 19116 9462 19168
rect 10686 19156 10692 19168
rect 10647 19128 10692 19156
rect 10686 19116 10692 19128
rect 10744 19156 10750 19168
rect 10965 19159 11023 19165
rect 10965 19156 10977 19159
rect 10744 19128 10977 19156
rect 10744 19116 10750 19128
rect 10965 19125 10977 19128
rect 11011 19125 11023 19159
rect 10965 19119 11023 19125
rect 11054 19116 11060 19168
rect 11112 19156 11118 19168
rect 11112 19128 11157 19156
rect 11112 19116 11118 19128
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 12728 19156 12756 19187
rect 14090 19184 14096 19236
rect 14148 19224 14154 19236
rect 14292 19224 14320 19255
rect 14734 19252 14740 19264
rect 14792 19252 14798 19304
rect 16684 19301 16712 19468
rect 17497 19465 17509 19499
rect 17543 19496 17555 19499
rect 17586 19496 17592 19508
rect 17543 19468 17592 19496
rect 17543 19465 17555 19468
rect 17497 19459 17555 19465
rect 17586 19456 17592 19468
rect 17644 19456 17650 19508
rect 21726 19496 21732 19508
rect 21687 19468 21732 19496
rect 21726 19456 21732 19468
rect 21784 19456 21790 19508
rect 23290 19456 23296 19508
rect 23348 19496 23354 19508
rect 23934 19496 23940 19508
rect 23348 19468 23940 19496
rect 23348 19456 23354 19468
rect 23934 19456 23940 19468
rect 23992 19456 23998 19508
rect 16942 19388 16948 19440
rect 17000 19428 17006 19440
rect 23477 19431 23535 19437
rect 17000 19400 17356 19428
rect 17000 19388 17006 19400
rect 17328 19369 17356 19400
rect 23477 19397 23489 19431
rect 23523 19428 23535 19431
rect 24026 19428 24032 19440
rect 23523 19400 24032 19428
rect 23523 19397 23535 19400
rect 23477 19391 23535 19397
rect 24026 19388 24032 19400
rect 24084 19428 24090 19440
rect 24489 19431 24547 19437
rect 24489 19428 24501 19431
rect 24084 19400 24501 19428
rect 24084 19388 24090 19400
rect 24489 19397 24501 19400
rect 24535 19428 24547 19431
rect 25682 19428 25688 19440
rect 24535 19400 25688 19428
rect 24535 19397 24547 19400
rect 24489 19391 24547 19397
rect 25682 19388 25688 19400
rect 25740 19388 25746 19440
rect 25774 19388 25780 19440
rect 25832 19428 25838 19440
rect 26145 19431 26203 19437
rect 26145 19428 26157 19431
rect 25832 19400 26157 19428
rect 25832 19388 25838 19400
rect 26145 19397 26157 19400
rect 26191 19397 26203 19431
rect 26145 19391 26203 19397
rect 31478 19388 31484 19440
rect 31536 19428 31542 19440
rect 33962 19428 33968 19440
rect 31536 19400 31800 19428
rect 31536 19388 31542 19400
rect 17313 19363 17371 19369
rect 17313 19329 17325 19363
rect 17359 19360 17371 19363
rect 17773 19363 17831 19369
rect 17773 19360 17785 19363
rect 17359 19332 17785 19360
rect 17359 19329 17371 19332
rect 17313 19323 17371 19329
rect 17773 19329 17785 19332
rect 17819 19329 17831 19363
rect 17773 19323 17831 19329
rect 19705 19363 19763 19369
rect 19705 19329 19717 19363
rect 19751 19360 19763 19363
rect 19886 19360 19892 19372
rect 19751 19332 19892 19360
rect 19751 19329 19763 19332
rect 19705 19323 19763 19329
rect 19886 19320 19892 19332
rect 19944 19320 19950 19372
rect 26326 19360 26332 19372
rect 26160 19332 26332 19360
rect 16669 19295 16727 19301
rect 16669 19261 16681 19295
rect 16715 19261 16727 19295
rect 16942 19292 16948 19304
rect 16903 19264 16948 19292
rect 16669 19255 16727 19261
rect 16942 19252 16948 19264
rect 17000 19252 17006 19304
rect 17129 19295 17187 19301
rect 17129 19261 17141 19295
rect 17175 19292 17187 19295
rect 17221 19295 17279 19301
rect 17221 19292 17233 19295
rect 17175 19264 17233 19292
rect 17175 19261 17187 19264
rect 17129 19255 17187 19261
rect 17221 19261 17233 19264
rect 17267 19261 17279 19295
rect 17221 19255 17279 19261
rect 17402 19252 17408 19304
rect 17460 19252 17466 19304
rect 19978 19292 19984 19304
rect 19812 19264 19984 19292
rect 15013 19227 15071 19233
rect 15013 19224 15025 19227
rect 14148 19196 15025 19224
rect 14148 19184 14154 19196
rect 15013 19193 15025 19196
rect 15059 19193 15071 19227
rect 17310 19224 17316 19236
rect 17271 19196 17316 19224
rect 15013 19187 15071 19193
rect 17310 19184 17316 19196
rect 17368 19184 17374 19236
rect 17420 19224 17448 19252
rect 18782 19224 18788 19236
rect 17420 19196 18788 19224
rect 18782 19184 18788 19196
rect 18840 19184 18846 19236
rect 19613 19227 19671 19233
rect 19613 19193 19625 19227
rect 19659 19224 19671 19227
rect 19812 19224 19840 19264
rect 19978 19252 19984 19264
rect 20036 19252 20042 19304
rect 24302 19292 24308 19304
rect 24263 19264 24308 19292
rect 24302 19252 24308 19264
rect 24360 19252 24366 19304
rect 25133 19295 25191 19301
rect 25133 19261 25145 19295
rect 25179 19292 25191 19295
rect 25314 19292 25320 19304
rect 25179 19264 25320 19292
rect 25179 19261 25191 19264
rect 25133 19255 25191 19261
rect 25314 19252 25320 19264
rect 25372 19252 25378 19304
rect 25682 19292 25688 19304
rect 25643 19264 25688 19292
rect 25682 19252 25688 19264
rect 25740 19252 25746 19304
rect 26050 19252 26056 19304
rect 26108 19292 26114 19304
rect 26160 19301 26188 19332
rect 26326 19320 26332 19332
rect 26384 19320 26390 19372
rect 26786 19360 26792 19372
rect 26699 19332 26792 19360
rect 26786 19320 26792 19332
rect 26844 19360 26850 19372
rect 28718 19360 28724 19372
rect 26844 19332 28724 19360
rect 26844 19320 26850 19332
rect 26145 19295 26203 19301
rect 26145 19292 26157 19295
rect 26108 19264 26157 19292
rect 26108 19252 26114 19264
rect 26145 19261 26157 19264
rect 26191 19261 26203 19295
rect 26145 19255 26203 19261
rect 27157 19295 27215 19301
rect 27157 19261 27169 19295
rect 27203 19292 27215 19295
rect 27430 19292 27436 19304
rect 27203 19264 27436 19292
rect 27203 19261 27215 19264
rect 27157 19255 27215 19261
rect 27430 19252 27436 19264
rect 27488 19252 27494 19304
rect 28092 19301 28120 19332
rect 28718 19320 28724 19332
rect 28776 19320 28782 19372
rect 30006 19320 30012 19372
rect 30064 19360 30070 19372
rect 30285 19363 30343 19369
rect 30285 19360 30297 19363
rect 30064 19332 30297 19360
rect 30064 19320 30070 19332
rect 30285 19329 30297 19332
rect 30331 19329 30343 19363
rect 30285 19323 30343 19329
rect 27525 19295 27583 19301
rect 27525 19261 27537 19295
rect 27571 19261 27583 19295
rect 27525 19255 27583 19261
rect 28077 19295 28135 19301
rect 28077 19261 28089 19295
rect 28123 19261 28135 19295
rect 28077 19255 28135 19261
rect 21358 19224 21364 19236
rect 19659 19196 19840 19224
rect 21319 19196 21364 19224
rect 19659 19193 19671 19196
rect 19613 19187 19671 19193
rect 21358 19184 21364 19196
rect 21416 19184 21422 19236
rect 24857 19227 24915 19233
rect 24857 19193 24869 19227
rect 24903 19224 24915 19227
rect 25222 19224 25228 19236
rect 24903 19196 25228 19224
rect 24903 19193 24915 19196
rect 24857 19187 24915 19193
rect 25222 19184 25228 19196
rect 25280 19184 25286 19236
rect 27540 19224 27568 19255
rect 28166 19252 28172 19304
rect 28224 19292 28230 19304
rect 28261 19295 28319 19301
rect 28261 19292 28273 19295
rect 28224 19264 28273 19292
rect 28224 19252 28230 19264
rect 28261 19261 28273 19264
rect 28307 19261 28319 19295
rect 29270 19292 29276 19304
rect 29231 19264 29276 19292
rect 28261 19255 28319 19261
rect 29270 19252 29276 19264
rect 29328 19252 29334 19304
rect 29549 19295 29607 19301
rect 29549 19292 29561 19295
rect 29380 19264 29561 19292
rect 29089 19227 29147 19233
rect 27540 19196 28120 19224
rect 28092 19168 28120 19196
rect 29089 19193 29101 19227
rect 29135 19224 29147 19227
rect 29178 19224 29184 19236
rect 29135 19196 29184 19224
rect 29135 19193 29147 19196
rect 29089 19187 29147 19193
rect 29178 19184 29184 19196
rect 29236 19224 29242 19236
rect 29380 19224 29408 19264
rect 29549 19261 29561 19264
rect 29595 19261 29607 19295
rect 31021 19295 31079 19301
rect 31021 19292 31033 19295
rect 29549 19255 29607 19261
rect 30944 19264 31033 19292
rect 29236 19196 29408 19224
rect 29469 19227 29527 19233
rect 29236 19184 29242 19196
rect 29469 19193 29481 19227
rect 29515 19224 29527 19227
rect 30009 19227 30067 19233
rect 29515 19196 29592 19224
rect 29515 19193 29527 19196
rect 29469 19187 29527 19193
rect 13814 19156 13820 19168
rect 12492 19128 12756 19156
rect 13775 19128 13820 19156
rect 12492 19116 12498 19128
rect 13814 19116 13820 19128
rect 13872 19116 13878 19168
rect 15470 19156 15476 19168
rect 15431 19128 15476 19156
rect 15470 19116 15476 19128
rect 15528 19116 15534 19168
rect 16025 19159 16083 19165
rect 16025 19125 16037 19159
rect 16071 19156 16083 19159
rect 17126 19156 17132 19168
rect 16071 19128 17132 19156
rect 16071 19125 16083 19128
rect 16025 19119 16083 19125
rect 17126 19116 17132 19128
rect 17184 19156 17190 19168
rect 17221 19159 17279 19165
rect 17221 19156 17233 19159
rect 17184 19128 17233 19156
rect 17184 19116 17190 19128
rect 17221 19125 17233 19128
rect 17267 19125 17279 19159
rect 17221 19119 17279 19125
rect 17402 19116 17408 19168
rect 17460 19156 17466 19168
rect 17589 19159 17647 19165
rect 17589 19156 17601 19159
rect 17460 19128 17601 19156
rect 17460 19116 17466 19128
rect 17589 19125 17601 19128
rect 17635 19125 17647 19159
rect 17589 19119 17647 19125
rect 18138 19116 18144 19168
rect 18196 19156 18202 19168
rect 18233 19159 18291 19165
rect 18233 19156 18245 19159
rect 18196 19128 18245 19156
rect 18196 19116 18202 19128
rect 18233 19125 18245 19128
rect 18279 19125 18291 19159
rect 18233 19119 18291 19125
rect 18322 19116 18328 19168
rect 18380 19156 18386 19168
rect 18601 19159 18659 19165
rect 18601 19156 18613 19159
rect 18380 19128 18613 19156
rect 18380 19116 18386 19128
rect 18601 19125 18613 19128
rect 18647 19125 18659 19159
rect 18601 19119 18659 19125
rect 22094 19116 22100 19168
rect 22152 19156 22158 19168
rect 22465 19159 22523 19165
rect 22152 19128 22197 19156
rect 22152 19116 22158 19128
rect 22465 19125 22477 19159
rect 22511 19156 22523 19159
rect 22554 19156 22560 19168
rect 22511 19128 22560 19156
rect 22511 19125 22523 19128
rect 22465 19119 22523 19125
rect 22554 19116 22560 19128
rect 22612 19116 22618 19168
rect 23106 19156 23112 19168
rect 23067 19128 23112 19156
rect 23106 19116 23112 19128
rect 23164 19116 23170 19168
rect 25958 19116 25964 19168
rect 26016 19156 26022 19168
rect 27341 19159 27399 19165
rect 27341 19156 27353 19159
rect 26016 19128 27353 19156
rect 26016 19116 26022 19128
rect 27341 19125 27353 19128
rect 27387 19125 27399 19159
rect 27341 19119 27399 19125
rect 28074 19116 28080 19168
rect 28132 19116 28138 19168
rect 28626 19156 28632 19168
rect 28587 19128 28632 19156
rect 28626 19116 28632 19128
rect 28684 19156 28690 19168
rect 29270 19156 29276 19168
rect 28684 19128 29276 19156
rect 28684 19116 28690 19128
rect 29270 19116 29276 19128
rect 29328 19116 29334 19168
rect 29564 19156 29592 19196
rect 30009 19193 30021 19227
rect 30055 19224 30067 19227
rect 30098 19224 30104 19236
rect 30055 19196 30104 19224
rect 30055 19193 30067 19196
rect 30009 19187 30067 19193
rect 30098 19184 30104 19196
rect 30156 19184 30162 19236
rect 30944 19168 30972 19264
rect 31021 19261 31033 19264
rect 31067 19261 31079 19295
rect 31021 19255 31079 19261
rect 31573 19295 31631 19301
rect 31573 19261 31585 19295
rect 31619 19261 31631 19295
rect 31772 19292 31800 19400
rect 32968 19400 33968 19428
rect 32968 19372 32996 19400
rect 33962 19388 33968 19400
rect 34020 19388 34026 19440
rect 32030 19360 32036 19372
rect 31991 19332 32036 19360
rect 32030 19320 32036 19332
rect 32088 19320 32094 19372
rect 32950 19360 32956 19372
rect 32863 19332 32956 19360
rect 32950 19320 32956 19332
rect 33008 19320 33014 19372
rect 33134 19360 33140 19372
rect 33060 19332 33140 19360
rect 31849 19295 31907 19301
rect 31849 19292 31861 19295
rect 31772 19264 31861 19292
rect 31573 19255 31631 19261
rect 31849 19261 31861 19264
rect 31895 19261 31907 19295
rect 31849 19255 31907 19261
rect 31588 19224 31616 19255
rect 31662 19224 31668 19236
rect 31588 19196 31668 19224
rect 31662 19184 31668 19196
rect 31720 19184 31726 19236
rect 30282 19156 30288 19168
rect 29564 19128 30288 19156
rect 30282 19116 30288 19128
rect 30340 19116 30346 19168
rect 30926 19156 30932 19168
rect 30887 19128 30932 19156
rect 30926 19116 30932 19128
rect 30984 19116 30990 19168
rect 32490 19156 32496 19168
rect 32451 19128 32496 19156
rect 32490 19116 32496 19128
rect 32548 19116 32554 19168
rect 32582 19116 32588 19168
rect 32640 19156 32646 19168
rect 32769 19159 32827 19165
rect 32769 19156 32781 19159
rect 32640 19128 32781 19156
rect 32640 19116 32646 19128
rect 32769 19125 32781 19128
rect 32815 19156 32827 19159
rect 33060 19156 33088 19332
rect 33134 19320 33140 19332
rect 33192 19320 33198 19372
rect 36078 19360 36084 19372
rect 35912 19332 36084 19360
rect 33502 19292 33508 19304
rect 33463 19264 33508 19292
rect 33502 19252 33508 19264
rect 33560 19252 33566 19304
rect 33778 19292 33784 19304
rect 33739 19264 33784 19292
rect 33778 19252 33784 19264
rect 33836 19252 33842 19304
rect 33870 19252 33876 19304
rect 33928 19292 33934 19304
rect 33965 19295 34023 19301
rect 33965 19292 33977 19295
rect 33928 19264 33977 19292
rect 33928 19252 33934 19264
rect 33965 19261 33977 19264
rect 34011 19292 34023 19295
rect 34241 19295 34299 19301
rect 34241 19292 34253 19295
rect 34011 19264 34253 19292
rect 34011 19261 34023 19264
rect 33965 19255 34023 19261
rect 34241 19261 34253 19264
rect 34287 19292 34299 19295
rect 35437 19295 35495 19301
rect 35437 19292 35449 19295
rect 34287 19264 35449 19292
rect 34287 19261 34299 19264
rect 34241 19255 34299 19261
rect 35437 19261 35449 19264
rect 35483 19292 35495 19295
rect 35912 19292 35940 19332
rect 36078 19320 36084 19332
rect 36136 19320 36142 19372
rect 35483 19264 35940 19292
rect 35483 19261 35495 19264
rect 35437 19255 35495 19261
rect 33520 19224 33548 19252
rect 34609 19227 34667 19233
rect 34609 19224 34621 19227
rect 33520 19196 34621 19224
rect 34609 19193 34621 19196
rect 34655 19224 34667 19227
rect 35618 19224 35624 19236
rect 34655 19196 35624 19224
rect 34655 19193 34667 19196
rect 34609 19187 34667 19193
rect 35618 19184 35624 19196
rect 35676 19224 35682 19236
rect 35805 19227 35863 19233
rect 35805 19224 35817 19227
rect 35676 19196 35817 19224
rect 35676 19184 35682 19196
rect 35805 19193 35817 19196
rect 35851 19193 35863 19227
rect 35805 19187 35863 19193
rect 32815 19128 33088 19156
rect 32815 19125 32827 19128
rect 32769 19119 32827 19125
rect 33134 19116 33140 19168
rect 33192 19156 33198 19168
rect 33778 19156 33784 19168
rect 33192 19128 33784 19156
rect 33192 19116 33198 19128
rect 33778 19116 33784 19128
rect 33836 19156 33842 19168
rect 34422 19156 34428 19168
rect 33836 19128 34428 19156
rect 33836 19116 33842 19128
rect 34422 19116 34428 19128
rect 34480 19116 34486 19168
rect 35066 19156 35072 19168
rect 35027 19128 35072 19156
rect 35066 19116 35072 19128
rect 35124 19156 35130 19168
rect 35894 19156 35900 19168
rect 35124 19128 35900 19156
rect 35124 19116 35130 19128
rect 35894 19116 35900 19128
rect 35952 19116 35958 19168
rect 1104 19066 38548 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 38548 19066
rect 1104 18992 38548 19014
rect 3510 18952 3516 18964
rect 3471 18924 3516 18952
rect 3510 18912 3516 18924
rect 3568 18912 3574 18964
rect 4893 18955 4951 18961
rect 4893 18921 4905 18955
rect 4939 18952 4951 18955
rect 5442 18952 5448 18964
rect 4939 18924 5448 18952
rect 4939 18921 4951 18924
rect 4893 18915 4951 18921
rect 5442 18912 5448 18924
rect 5500 18912 5506 18964
rect 6178 18952 6184 18964
rect 6139 18924 6184 18952
rect 6178 18912 6184 18924
rect 6236 18912 6242 18964
rect 6454 18952 6460 18964
rect 6415 18924 6460 18952
rect 6454 18912 6460 18924
rect 6512 18912 6518 18964
rect 6825 18955 6883 18961
rect 6825 18921 6837 18955
rect 6871 18952 6883 18955
rect 6914 18952 6920 18964
rect 6871 18924 6920 18952
rect 6871 18921 6883 18924
rect 6825 18915 6883 18921
rect 6914 18912 6920 18924
rect 6972 18912 6978 18964
rect 8754 18952 8760 18964
rect 8715 18924 8760 18952
rect 8754 18912 8760 18924
rect 8812 18912 8818 18964
rect 11054 18952 11060 18964
rect 10336 18924 11060 18952
rect 5166 18884 5172 18896
rect 5127 18856 5172 18884
rect 5166 18844 5172 18856
rect 5224 18844 5230 18896
rect 7466 18844 7472 18896
rect 7524 18884 7530 18896
rect 7837 18887 7895 18893
rect 7837 18884 7849 18887
rect 7524 18856 7849 18884
rect 7524 18844 7530 18856
rect 7837 18853 7849 18856
rect 7883 18853 7895 18887
rect 7837 18847 7895 18853
rect 10042 18844 10048 18896
rect 10100 18884 10106 18896
rect 10336 18893 10364 18924
rect 11054 18912 11060 18924
rect 11112 18912 11118 18964
rect 11698 18952 11704 18964
rect 11611 18924 11704 18952
rect 11698 18912 11704 18924
rect 11756 18952 11762 18964
rect 12158 18952 12164 18964
rect 11756 18924 12164 18952
rect 11756 18912 11762 18924
rect 12158 18912 12164 18924
rect 12216 18912 12222 18964
rect 13449 18955 13507 18961
rect 13449 18921 13461 18955
rect 13495 18952 13507 18955
rect 13630 18952 13636 18964
rect 13495 18924 13636 18952
rect 13495 18921 13507 18924
rect 13449 18915 13507 18921
rect 13630 18912 13636 18924
rect 13688 18912 13694 18964
rect 14642 18952 14648 18964
rect 14603 18924 14648 18952
rect 14642 18912 14648 18924
rect 14700 18912 14706 18964
rect 16022 18912 16028 18964
rect 16080 18912 16086 18964
rect 16206 18952 16212 18964
rect 16167 18924 16212 18952
rect 16206 18912 16212 18924
rect 16264 18912 16270 18964
rect 17221 18955 17279 18961
rect 17221 18921 17233 18955
rect 17267 18952 17279 18955
rect 17586 18952 17592 18964
rect 17267 18924 17592 18952
rect 17267 18921 17279 18924
rect 17221 18915 17279 18921
rect 17586 18912 17592 18924
rect 17644 18912 17650 18964
rect 17678 18912 17684 18964
rect 17736 18952 17742 18964
rect 18509 18955 18567 18961
rect 18509 18952 18521 18955
rect 17736 18924 18521 18952
rect 17736 18912 17742 18924
rect 18509 18921 18521 18924
rect 18555 18921 18567 18955
rect 18509 18915 18567 18921
rect 18598 18912 18604 18964
rect 18656 18952 18662 18964
rect 18877 18955 18935 18961
rect 18877 18952 18889 18955
rect 18656 18924 18889 18952
rect 18656 18912 18662 18924
rect 18877 18921 18889 18924
rect 18923 18921 18935 18955
rect 18877 18915 18935 18921
rect 21358 18912 21364 18964
rect 21416 18952 21422 18964
rect 22557 18955 22615 18961
rect 22557 18952 22569 18955
rect 21416 18924 22569 18952
rect 21416 18912 21422 18924
rect 22557 18921 22569 18924
rect 22603 18952 22615 18955
rect 23474 18952 23480 18964
rect 22603 18924 23480 18952
rect 22603 18921 22615 18924
rect 22557 18915 22615 18921
rect 23474 18912 23480 18924
rect 23532 18912 23538 18964
rect 24302 18912 24308 18964
rect 24360 18952 24366 18964
rect 24489 18955 24547 18961
rect 24489 18952 24501 18955
rect 24360 18924 24501 18952
rect 24360 18912 24366 18924
rect 24489 18921 24501 18924
rect 24535 18921 24547 18955
rect 24489 18915 24547 18921
rect 25041 18955 25099 18961
rect 25041 18921 25053 18955
rect 25087 18952 25099 18955
rect 26050 18952 26056 18964
rect 25087 18924 26056 18952
rect 25087 18921 25099 18924
rect 25041 18915 25099 18921
rect 26050 18912 26056 18924
rect 26108 18912 26114 18964
rect 26234 18912 26240 18964
rect 26292 18952 26298 18964
rect 26970 18952 26976 18964
rect 26292 18924 26976 18952
rect 26292 18912 26298 18924
rect 26970 18912 26976 18924
rect 27028 18912 27034 18964
rect 27706 18912 27712 18964
rect 27764 18952 27770 18964
rect 28261 18955 28319 18961
rect 28261 18952 28273 18955
rect 27764 18924 28273 18952
rect 27764 18912 27770 18924
rect 28261 18921 28273 18924
rect 28307 18921 28319 18955
rect 28261 18915 28319 18921
rect 30009 18955 30067 18961
rect 30009 18921 30021 18955
rect 30055 18952 30067 18955
rect 30098 18952 30104 18964
rect 30055 18924 30104 18952
rect 30055 18921 30067 18924
rect 30009 18915 30067 18921
rect 30098 18912 30104 18924
rect 30156 18912 30162 18964
rect 30190 18912 30196 18964
rect 30248 18952 30254 18964
rect 30285 18955 30343 18961
rect 30285 18952 30297 18955
rect 30248 18924 30297 18952
rect 30248 18912 30254 18924
rect 30285 18921 30297 18924
rect 30331 18921 30343 18955
rect 30285 18915 30343 18921
rect 31202 18912 31208 18964
rect 31260 18952 31266 18964
rect 31389 18955 31447 18961
rect 31389 18952 31401 18955
rect 31260 18924 31401 18952
rect 31260 18912 31266 18924
rect 31389 18921 31401 18924
rect 31435 18921 31447 18955
rect 31389 18915 31447 18921
rect 32861 18955 32919 18961
rect 32861 18921 32873 18955
rect 32907 18952 32919 18955
rect 32950 18952 32956 18964
rect 32907 18924 32956 18952
rect 32907 18921 32919 18924
rect 32861 18915 32919 18921
rect 32950 18912 32956 18924
rect 33008 18912 33014 18964
rect 10321 18887 10379 18893
rect 10321 18884 10333 18887
rect 10100 18856 10333 18884
rect 10100 18844 10106 18856
rect 10321 18853 10333 18856
rect 10367 18853 10379 18887
rect 10321 18847 10379 18853
rect 10413 18887 10471 18893
rect 10413 18853 10425 18887
rect 10459 18884 10471 18887
rect 10594 18884 10600 18896
rect 10459 18856 10600 18884
rect 10459 18853 10471 18856
rect 10413 18847 10471 18853
rect 10594 18844 10600 18856
rect 10652 18844 10658 18896
rect 10778 18884 10784 18896
rect 10739 18856 10784 18884
rect 10778 18844 10784 18856
rect 10836 18844 10842 18896
rect 15838 18844 15844 18896
rect 15896 18884 15902 18896
rect 15933 18887 15991 18893
rect 15933 18884 15945 18887
rect 15896 18856 15945 18884
rect 15896 18844 15902 18856
rect 15933 18853 15945 18856
rect 15979 18853 15991 18887
rect 16040 18884 16068 18912
rect 23017 18887 23075 18893
rect 16040 18856 17356 18884
rect 15933 18847 15991 18853
rect 1670 18816 1676 18828
rect 1631 18788 1676 18816
rect 1670 18776 1676 18788
rect 1728 18776 1734 18828
rect 1946 18776 1952 18828
rect 2004 18776 2010 18828
rect 5626 18816 5632 18828
rect 5587 18788 5632 18816
rect 5626 18776 5632 18788
rect 5684 18776 5690 18828
rect 6641 18819 6699 18825
rect 6641 18785 6653 18819
rect 6687 18816 6699 18819
rect 7006 18816 7012 18828
rect 6687 18788 7012 18816
rect 6687 18785 6699 18788
rect 6641 18779 6699 18785
rect 7006 18776 7012 18788
rect 7064 18776 7070 18828
rect 7374 18776 7380 18828
rect 7432 18816 7438 18828
rect 7653 18819 7711 18825
rect 7653 18816 7665 18819
rect 7432 18788 7665 18816
rect 7432 18776 7438 18788
rect 7653 18785 7665 18788
rect 7699 18785 7711 18819
rect 7926 18816 7932 18828
rect 7887 18788 7932 18816
rect 7653 18779 7711 18785
rect 7926 18776 7932 18788
rect 7984 18776 7990 18828
rect 10229 18819 10287 18825
rect 10229 18785 10241 18819
rect 10275 18816 10287 18819
rect 10686 18816 10692 18828
rect 10275 18788 10692 18816
rect 10275 18785 10287 18788
rect 10229 18779 10287 18785
rect 10686 18776 10692 18788
rect 10744 18776 10750 18828
rect 12253 18819 12311 18825
rect 12253 18785 12265 18819
rect 12299 18785 12311 18819
rect 12253 18779 12311 18785
rect 1397 18751 1455 18757
rect 1397 18717 1409 18751
rect 1443 18748 1455 18751
rect 1964 18748 1992 18776
rect 1443 18720 1992 18748
rect 1443 18717 1455 18720
rect 1397 18711 1455 18717
rect 8662 18708 8668 18760
rect 8720 18748 8726 18760
rect 9214 18748 9220 18760
rect 8720 18720 9220 18748
rect 8720 18708 8726 18720
rect 9214 18708 9220 18720
rect 9272 18708 9278 18760
rect 9490 18708 9496 18760
rect 9548 18748 9554 18760
rect 10045 18751 10103 18757
rect 10045 18748 10057 18751
rect 9548 18720 10057 18748
rect 9548 18708 9554 18720
rect 10045 18717 10057 18720
rect 10091 18748 10103 18751
rect 12268 18748 12296 18779
rect 12434 18776 12440 18828
rect 12492 18816 12498 18828
rect 12492 18788 12537 18816
rect 12492 18776 12498 18788
rect 12710 18776 12716 18828
rect 12768 18816 12774 18828
rect 12805 18819 12863 18825
rect 12805 18816 12817 18819
rect 12768 18788 12817 18816
rect 12768 18776 12774 18788
rect 12805 18785 12817 18788
rect 12851 18785 12863 18819
rect 12805 18779 12863 18785
rect 14185 18819 14243 18825
rect 14185 18785 14197 18819
rect 14231 18816 14243 18819
rect 14274 18816 14280 18828
rect 14231 18788 14280 18816
rect 14231 18785 14243 18788
rect 14185 18779 14243 18785
rect 14274 18776 14280 18788
rect 14332 18776 14338 18828
rect 16022 18776 16028 18828
rect 16080 18816 16086 18828
rect 17328 18825 17356 18856
rect 23017 18853 23029 18887
rect 23063 18884 23075 18887
rect 23106 18884 23112 18896
rect 23063 18856 23112 18884
rect 23063 18853 23075 18856
rect 23017 18847 23075 18853
rect 23106 18844 23112 18856
rect 23164 18884 23170 18896
rect 23164 18856 24072 18884
rect 23164 18844 23170 18856
rect 16117 18819 16175 18825
rect 16117 18816 16129 18819
rect 16080 18788 16129 18816
rect 16080 18776 16086 18788
rect 16117 18785 16129 18788
rect 16163 18785 16175 18819
rect 16117 18779 16175 18785
rect 17313 18819 17371 18825
rect 17313 18785 17325 18819
rect 17359 18785 17371 18819
rect 17313 18779 17371 18785
rect 17405 18819 17463 18825
rect 17405 18785 17417 18819
rect 17451 18816 17463 18819
rect 17954 18816 17960 18828
rect 17451 18788 17960 18816
rect 17451 18785 17463 18788
rect 17405 18779 17463 18785
rect 12526 18748 12532 18760
rect 10091 18720 11192 18748
rect 12268 18720 12532 18748
rect 10091 18717 10103 18720
rect 10045 18711 10103 18717
rect 4430 18680 4436 18692
rect 4391 18652 4436 18680
rect 4430 18640 4436 18652
rect 4488 18640 4494 18692
rect 5442 18640 5448 18692
rect 5500 18680 5506 18692
rect 5813 18683 5871 18689
rect 5813 18680 5825 18683
rect 5500 18652 5825 18680
rect 5500 18640 5506 18652
rect 5813 18649 5825 18652
rect 5859 18680 5871 18683
rect 6546 18680 6552 18692
rect 5859 18652 6552 18680
rect 5859 18649 5871 18652
rect 5813 18643 5871 18649
rect 6546 18640 6552 18652
rect 6604 18680 6610 18692
rect 7190 18680 7196 18692
rect 6604 18652 7196 18680
rect 6604 18640 6610 18652
rect 7190 18640 7196 18652
rect 7248 18640 7254 18692
rect 8938 18640 8944 18692
rect 8996 18680 9002 18692
rect 9398 18680 9404 18692
rect 8996 18652 9404 18680
rect 8996 18640 9002 18652
rect 9398 18640 9404 18652
rect 9456 18680 9462 18692
rect 9861 18683 9919 18689
rect 9861 18680 9873 18683
rect 9456 18652 9873 18680
rect 9456 18640 9462 18652
rect 9861 18649 9873 18652
rect 9907 18649 9919 18683
rect 9861 18643 9919 18649
rect 9950 18640 9956 18692
rect 10008 18680 10014 18692
rect 10594 18680 10600 18692
rect 10008 18652 10600 18680
rect 10008 18640 10014 18652
rect 10594 18640 10600 18652
rect 10652 18680 10658 18692
rect 10962 18680 10968 18692
rect 10652 18652 10968 18680
rect 10652 18640 10658 18652
rect 10962 18640 10968 18652
rect 11020 18640 11026 18692
rect 2590 18572 2596 18624
rect 2648 18612 2654 18624
rect 2777 18615 2835 18621
rect 2777 18612 2789 18615
rect 2648 18584 2789 18612
rect 2648 18572 2654 18584
rect 2777 18581 2789 18584
rect 2823 18581 2835 18615
rect 2777 18575 2835 18581
rect 3142 18572 3148 18624
rect 3200 18612 3206 18624
rect 3789 18615 3847 18621
rect 3789 18612 3801 18615
rect 3200 18584 3801 18612
rect 3200 18572 3206 18584
rect 3789 18581 3801 18584
rect 3835 18581 3847 18615
rect 3789 18575 3847 18581
rect 6454 18572 6460 18624
rect 6512 18612 6518 18624
rect 7285 18615 7343 18621
rect 7285 18612 7297 18615
rect 6512 18584 7297 18612
rect 6512 18572 6518 18584
rect 7285 18581 7297 18584
rect 7331 18612 7343 18615
rect 7558 18612 7564 18624
rect 7331 18584 7564 18612
rect 7331 18581 7343 18584
rect 7285 18575 7343 18581
rect 7558 18572 7564 18584
rect 7616 18572 7622 18624
rect 8110 18612 8116 18624
rect 8071 18584 8116 18612
rect 8110 18572 8116 18584
rect 8168 18572 8174 18624
rect 9030 18572 9036 18624
rect 9088 18612 9094 18624
rect 11164 18621 11192 18720
rect 12526 18708 12532 18720
rect 12584 18708 12590 18760
rect 17328 18748 17356 18779
rect 17954 18776 17960 18788
rect 18012 18816 18018 18828
rect 18693 18819 18751 18825
rect 18693 18816 18705 18819
rect 18012 18788 18705 18816
rect 18012 18776 18018 18788
rect 18693 18785 18705 18788
rect 18739 18785 18751 18819
rect 18693 18779 18751 18785
rect 23661 18819 23719 18825
rect 23661 18785 23673 18819
rect 23707 18816 23719 18819
rect 23934 18816 23940 18828
rect 23707 18788 23940 18816
rect 23707 18785 23719 18788
rect 23661 18779 23719 18785
rect 23934 18776 23940 18788
rect 23992 18776 23998 18828
rect 24044 18825 24072 18856
rect 25682 18844 25688 18896
rect 25740 18884 25746 18896
rect 25961 18887 26019 18893
rect 25961 18884 25973 18887
rect 25740 18856 25973 18884
rect 25740 18844 25746 18856
rect 25961 18853 25973 18856
rect 26007 18853 26019 18887
rect 25961 18847 26019 18853
rect 27430 18844 27436 18896
rect 27488 18884 27494 18896
rect 27798 18884 27804 18896
rect 27488 18856 27804 18884
rect 27488 18844 27494 18856
rect 27798 18844 27804 18856
rect 27856 18884 27862 18896
rect 29365 18887 29423 18893
rect 29365 18884 29377 18887
rect 27856 18856 29377 18884
rect 27856 18844 27862 18856
rect 29365 18853 29377 18856
rect 29411 18853 29423 18887
rect 29365 18847 29423 18853
rect 24029 18819 24087 18825
rect 24029 18785 24041 18819
rect 24075 18816 24087 18819
rect 24394 18816 24400 18828
rect 24075 18788 24400 18816
rect 24075 18785 24087 18788
rect 24029 18779 24087 18785
rect 24394 18776 24400 18788
rect 24452 18776 24458 18828
rect 25133 18819 25191 18825
rect 25133 18785 25145 18819
rect 25179 18816 25191 18819
rect 26789 18819 26847 18825
rect 25179 18788 25728 18816
rect 25179 18785 25191 18788
rect 25133 18779 25191 18785
rect 18414 18748 18420 18760
rect 17328 18720 18420 18748
rect 18414 18708 18420 18720
rect 18472 18708 18478 18760
rect 23198 18708 23204 18760
rect 23256 18748 23262 18760
rect 23293 18751 23351 18757
rect 23293 18748 23305 18751
rect 23256 18720 23305 18748
rect 23256 18708 23262 18720
rect 23293 18717 23305 18720
rect 23339 18748 23351 18751
rect 24302 18748 24308 18760
rect 23339 18720 24308 18748
rect 23339 18717 23351 18720
rect 23293 18711 23351 18717
rect 24302 18708 24308 18720
rect 24360 18708 24366 18760
rect 12802 18680 12808 18692
rect 12763 18652 12808 18680
rect 12802 18640 12808 18652
rect 12860 18640 12866 18692
rect 13998 18640 14004 18692
rect 14056 18680 14062 18692
rect 15013 18683 15071 18689
rect 15013 18680 15025 18683
rect 14056 18652 15025 18680
rect 14056 18640 14062 18652
rect 15013 18649 15025 18652
rect 15059 18649 15071 18683
rect 15013 18643 15071 18649
rect 16853 18683 16911 18689
rect 16853 18649 16865 18683
rect 16899 18680 16911 18683
rect 17494 18680 17500 18692
rect 16899 18652 17500 18680
rect 16899 18649 16911 18652
rect 16853 18643 16911 18649
rect 17494 18640 17500 18652
rect 17552 18640 17558 18692
rect 23934 18680 23940 18692
rect 23895 18652 23940 18680
rect 23934 18640 23940 18652
rect 23992 18640 23998 18692
rect 25317 18683 25375 18689
rect 25317 18649 25329 18683
rect 25363 18680 25375 18683
rect 25590 18680 25596 18692
rect 25363 18652 25596 18680
rect 25363 18649 25375 18652
rect 25317 18643 25375 18649
rect 25590 18640 25596 18652
rect 25648 18640 25654 18692
rect 25700 18689 25728 18788
rect 26789 18785 26801 18819
rect 26835 18816 26847 18819
rect 26970 18816 26976 18828
rect 26835 18788 26976 18816
rect 26835 18785 26847 18788
rect 26789 18779 26847 18785
rect 26970 18776 26976 18788
rect 27028 18776 27034 18828
rect 28166 18816 28172 18828
rect 28127 18788 28172 18816
rect 28166 18776 28172 18788
rect 28224 18776 28230 18828
rect 28718 18776 28724 18828
rect 28776 18816 28782 18828
rect 28997 18819 29055 18825
rect 28997 18816 29009 18819
rect 28776 18788 29009 18816
rect 28776 18776 28782 18788
rect 28997 18785 29009 18788
rect 29043 18816 29055 18819
rect 30208 18816 30236 18912
rect 34054 18884 34060 18896
rect 34015 18856 34060 18884
rect 34054 18844 34060 18856
rect 34112 18844 34118 18896
rect 33502 18816 33508 18828
rect 29043 18788 30236 18816
rect 33463 18788 33508 18816
rect 29043 18785 29055 18788
rect 28997 18779 29055 18785
rect 33502 18776 33508 18788
rect 33560 18776 33566 18828
rect 33778 18816 33784 18828
rect 33739 18788 33784 18816
rect 33778 18776 33784 18788
rect 33836 18776 33842 18828
rect 29086 18748 29092 18760
rect 29047 18720 29092 18748
rect 29086 18708 29092 18720
rect 29144 18708 29150 18760
rect 33042 18748 33048 18760
rect 33003 18720 33048 18748
rect 33042 18708 33048 18720
rect 33100 18708 33106 18760
rect 25685 18683 25743 18689
rect 25685 18649 25697 18683
rect 25731 18680 25743 18683
rect 26142 18680 26148 18692
rect 25731 18652 26148 18680
rect 25731 18649 25743 18652
rect 25685 18643 25743 18649
rect 26142 18640 26148 18652
rect 26200 18640 26206 18692
rect 9125 18615 9183 18621
rect 9125 18612 9137 18615
rect 9088 18584 9137 18612
rect 9088 18572 9094 18584
rect 9125 18581 9137 18584
rect 9171 18581 9183 18615
rect 9125 18575 9183 18581
rect 11149 18615 11207 18621
rect 11149 18581 11161 18615
rect 11195 18612 11207 18615
rect 11330 18612 11336 18624
rect 11195 18584 11336 18612
rect 11195 18581 11207 18584
rect 11149 18575 11207 18581
rect 11330 18572 11336 18584
rect 11388 18572 11394 18624
rect 13538 18572 13544 18624
rect 13596 18612 13602 18624
rect 13725 18615 13783 18621
rect 13725 18612 13737 18615
rect 13596 18584 13737 18612
rect 13596 18572 13602 18584
rect 13725 18581 13737 18584
rect 13771 18581 13783 18615
rect 13725 18575 13783 18581
rect 13906 18572 13912 18624
rect 13964 18612 13970 18624
rect 14369 18615 14427 18621
rect 14369 18612 14381 18615
rect 13964 18584 14381 18612
rect 13964 18572 13970 18584
rect 14369 18581 14381 18584
rect 14415 18581 14427 18615
rect 14369 18575 14427 18581
rect 14550 18572 14556 18624
rect 14608 18612 14614 18624
rect 15378 18612 15384 18624
rect 14608 18584 15384 18612
rect 14608 18572 14614 18584
rect 15378 18572 15384 18584
rect 15436 18612 15442 18624
rect 15565 18615 15623 18621
rect 15565 18612 15577 18615
rect 15436 18584 15577 18612
rect 15436 18572 15442 18584
rect 15565 18581 15577 18584
rect 15611 18612 15623 18615
rect 16942 18612 16948 18624
rect 15611 18584 16948 18612
rect 15611 18581 15623 18584
rect 15565 18575 15623 18581
rect 16942 18572 16948 18584
rect 17000 18572 17006 18624
rect 17126 18572 17132 18624
rect 17184 18612 17190 18624
rect 17586 18612 17592 18624
rect 17184 18584 17592 18612
rect 17184 18572 17190 18584
rect 17586 18572 17592 18584
rect 17644 18572 17650 18624
rect 18233 18615 18291 18621
rect 18233 18581 18245 18615
rect 18279 18612 18291 18615
rect 18782 18612 18788 18624
rect 18279 18584 18788 18612
rect 18279 18581 18291 18584
rect 18233 18575 18291 18581
rect 18782 18572 18788 18584
rect 18840 18572 18846 18624
rect 19702 18612 19708 18624
rect 19663 18584 19708 18612
rect 19702 18572 19708 18584
rect 19760 18572 19766 18624
rect 27433 18615 27491 18621
rect 27433 18581 27445 18615
rect 27479 18612 27491 18615
rect 27614 18612 27620 18624
rect 27479 18584 27620 18612
rect 27479 18581 27491 18584
rect 27433 18575 27491 18581
rect 27614 18572 27620 18584
rect 27672 18572 27678 18624
rect 29365 18615 29423 18621
rect 29365 18581 29377 18615
rect 29411 18612 29423 18615
rect 29641 18615 29699 18621
rect 29641 18612 29653 18615
rect 29411 18584 29653 18612
rect 29411 18581 29423 18584
rect 29365 18575 29423 18581
rect 29641 18581 29653 18584
rect 29687 18612 29699 18615
rect 30282 18612 30288 18624
rect 29687 18584 30288 18612
rect 29687 18581 29699 18584
rect 29641 18575 29699 18581
rect 30282 18572 30288 18584
rect 30340 18572 30346 18624
rect 30650 18612 30656 18624
rect 30611 18584 30656 18612
rect 30650 18572 30656 18584
rect 30708 18572 30714 18624
rect 30926 18572 30932 18624
rect 30984 18612 30990 18624
rect 31021 18615 31079 18621
rect 31021 18612 31033 18615
rect 30984 18584 31033 18612
rect 30984 18572 30990 18584
rect 31021 18581 31033 18584
rect 31067 18612 31079 18615
rect 31662 18612 31668 18624
rect 31067 18584 31668 18612
rect 31067 18581 31079 18584
rect 31021 18575 31079 18581
rect 31662 18572 31668 18584
rect 31720 18612 31726 18624
rect 32582 18612 32588 18624
rect 31720 18584 32588 18612
rect 31720 18572 31726 18584
rect 32582 18572 32588 18584
rect 32640 18572 32646 18624
rect 1104 18522 38548 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 38548 18522
rect 1104 18448 38548 18470
rect 1670 18408 1676 18420
rect 1631 18380 1676 18408
rect 1670 18368 1676 18380
rect 1728 18368 1734 18420
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 4157 18411 4215 18417
rect 4157 18377 4169 18411
rect 4203 18408 4215 18411
rect 4614 18408 4620 18420
rect 4203 18380 4620 18408
rect 4203 18377 4215 18380
rect 4157 18371 4215 18377
rect 4614 18368 4620 18380
rect 4672 18368 4678 18420
rect 4890 18408 4896 18420
rect 4851 18380 4896 18408
rect 4890 18368 4896 18380
rect 4948 18368 4954 18420
rect 5258 18408 5264 18420
rect 5219 18380 5264 18408
rect 5258 18368 5264 18380
rect 5316 18368 5322 18420
rect 5626 18408 5632 18420
rect 5587 18380 5632 18408
rect 5626 18368 5632 18380
rect 5684 18368 5690 18420
rect 5902 18408 5908 18420
rect 5863 18380 5908 18408
rect 5902 18368 5908 18380
rect 5960 18368 5966 18420
rect 8570 18368 8576 18420
rect 8628 18408 8634 18420
rect 8665 18411 8723 18417
rect 8665 18408 8677 18411
rect 8628 18380 8677 18408
rect 8628 18368 8634 18380
rect 8665 18377 8677 18380
rect 8711 18408 8723 18411
rect 10686 18408 10692 18420
rect 8711 18380 8892 18408
rect 10647 18380 10692 18408
rect 8711 18377 8723 18380
rect 8665 18371 8723 18377
rect 5644 18340 5672 18368
rect 6914 18340 6920 18352
rect 5644 18312 6920 18340
rect 6914 18300 6920 18312
rect 6972 18300 6978 18352
rect 7006 18232 7012 18284
rect 7064 18272 7070 18284
rect 8864 18281 8892 18380
rect 10686 18368 10692 18380
rect 10744 18368 10750 18420
rect 13814 18368 13820 18420
rect 13872 18408 13878 18420
rect 15657 18411 15715 18417
rect 13872 18380 15608 18408
rect 13872 18368 13878 18380
rect 12526 18340 12532 18352
rect 12360 18312 12532 18340
rect 7101 18275 7159 18281
rect 7101 18272 7113 18275
rect 7064 18244 7113 18272
rect 7064 18232 7070 18244
rect 7101 18241 7113 18244
rect 7147 18272 7159 18275
rect 8481 18275 8539 18281
rect 8481 18272 8493 18275
rect 7147 18244 8493 18272
rect 7147 18241 7159 18244
rect 7101 18235 7159 18241
rect 8481 18241 8493 18244
rect 8527 18241 8539 18275
rect 8481 18235 8539 18241
rect 8849 18275 8907 18281
rect 8849 18241 8861 18275
rect 8895 18241 8907 18275
rect 9582 18272 9588 18284
rect 9543 18244 9588 18272
rect 8849 18235 8907 18241
rect 9582 18232 9588 18244
rect 9640 18232 9646 18284
rect 11330 18272 11336 18284
rect 11291 18244 11336 18272
rect 11330 18232 11336 18244
rect 11388 18232 11394 18284
rect 12069 18275 12127 18281
rect 12069 18241 12081 18275
rect 12115 18272 12127 18275
rect 12360 18272 12388 18312
rect 12526 18300 12532 18312
rect 12584 18340 12590 18352
rect 13173 18343 13231 18349
rect 13173 18340 13185 18343
rect 12584 18312 13185 18340
rect 12584 18300 12590 18312
rect 13173 18309 13185 18312
rect 13219 18340 13231 18343
rect 13219 18312 13308 18340
rect 13219 18309 13231 18312
rect 13173 18303 13231 18309
rect 12115 18244 12388 18272
rect 13280 18272 13308 18312
rect 13630 18300 13636 18352
rect 13688 18340 13694 18352
rect 15580 18340 15608 18380
rect 15657 18377 15669 18411
rect 15703 18408 15715 18411
rect 15838 18408 15844 18420
rect 15703 18380 15844 18408
rect 15703 18377 15715 18380
rect 15657 18371 15715 18377
rect 15838 18368 15844 18380
rect 15896 18368 15902 18420
rect 17310 18368 17316 18420
rect 17368 18408 17374 18420
rect 18322 18408 18328 18420
rect 17368 18380 18328 18408
rect 17368 18368 17374 18380
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 23198 18408 23204 18420
rect 23159 18380 23204 18408
rect 23198 18368 23204 18380
rect 23256 18368 23262 18420
rect 23937 18411 23995 18417
rect 23937 18377 23949 18411
rect 23983 18408 23995 18411
rect 24026 18408 24032 18420
rect 23983 18380 24032 18408
rect 23983 18377 23995 18380
rect 23937 18371 23995 18377
rect 24026 18368 24032 18380
rect 24084 18368 24090 18420
rect 24302 18408 24308 18420
rect 24263 18380 24308 18408
rect 24302 18368 24308 18380
rect 24360 18368 24366 18420
rect 28718 18408 28724 18420
rect 28679 18380 28724 18408
rect 28718 18368 28724 18380
rect 28776 18368 28782 18420
rect 29825 18411 29883 18417
rect 29825 18377 29837 18411
rect 29871 18408 29883 18411
rect 29914 18408 29920 18420
rect 29871 18380 29920 18408
rect 29871 18377 29883 18380
rect 29825 18371 29883 18377
rect 29914 18368 29920 18380
rect 29972 18408 29978 18420
rect 30466 18408 30472 18420
rect 29972 18380 30472 18408
rect 29972 18368 29978 18380
rect 30466 18368 30472 18380
rect 30524 18368 30530 18420
rect 33042 18368 33048 18420
rect 33100 18368 33106 18420
rect 16393 18343 16451 18349
rect 16393 18340 16405 18343
rect 13688 18312 14136 18340
rect 15580 18312 16405 18340
rect 13688 18300 13694 18312
rect 13280 18244 13952 18272
rect 12115 18241 12127 18244
rect 12069 18235 12127 18241
rect 13924 18216 13952 18244
rect 5721 18207 5779 18213
rect 5721 18173 5733 18207
rect 5767 18204 5779 18207
rect 6641 18207 6699 18213
rect 5767 18176 6040 18204
rect 5767 18173 5779 18176
rect 5721 18167 5779 18173
rect 6012 18080 6040 18176
rect 6641 18173 6653 18207
rect 6687 18204 6699 18207
rect 7190 18204 7196 18216
rect 6687 18176 7196 18204
rect 6687 18173 6699 18176
rect 6641 18167 6699 18173
rect 7190 18164 7196 18176
rect 7248 18164 7254 18216
rect 7377 18207 7435 18213
rect 7377 18173 7389 18207
rect 7423 18204 7435 18207
rect 8754 18204 8760 18216
rect 7423 18176 8760 18204
rect 7423 18173 7435 18176
rect 7377 18167 7435 18173
rect 8754 18164 8760 18176
rect 8812 18164 8818 18216
rect 8938 18164 8944 18216
rect 8996 18204 9002 18216
rect 9125 18207 9183 18213
rect 9125 18204 9137 18207
rect 8996 18176 9137 18204
rect 8996 18164 9002 18176
rect 9125 18173 9137 18176
rect 9171 18173 9183 18207
rect 9125 18167 9183 18173
rect 9766 18164 9772 18216
rect 9824 18204 9830 18216
rect 10413 18207 10471 18213
rect 10413 18204 10425 18207
rect 9824 18176 10425 18204
rect 9824 18164 9830 18176
rect 10413 18173 10425 18176
rect 10459 18173 10471 18207
rect 10413 18167 10471 18173
rect 10502 18164 10508 18216
rect 10560 18204 10566 18216
rect 11609 18207 11667 18213
rect 11609 18204 11621 18207
rect 10560 18176 11621 18204
rect 10560 18164 10566 18176
rect 11609 18173 11621 18176
rect 11655 18204 11667 18207
rect 11974 18204 11980 18216
rect 11655 18176 11980 18204
rect 11655 18173 11667 18176
rect 11609 18167 11667 18173
rect 11974 18164 11980 18176
rect 12032 18164 12038 18216
rect 13538 18204 13544 18216
rect 13499 18176 13544 18204
rect 13538 18164 13544 18176
rect 13596 18164 13602 18216
rect 13906 18204 13912 18216
rect 13867 18176 13912 18204
rect 13906 18164 13912 18176
rect 13964 18164 13970 18216
rect 14108 18213 14136 18312
rect 16393 18309 16405 18312
rect 16439 18340 16451 18343
rect 17954 18340 17960 18352
rect 16439 18312 17960 18340
rect 16439 18309 16451 18312
rect 16393 18303 16451 18309
rect 17954 18300 17960 18312
rect 18012 18340 18018 18352
rect 19061 18343 19119 18349
rect 19061 18340 19073 18343
rect 18012 18312 19073 18340
rect 18012 18300 18018 18312
rect 19061 18309 19073 18312
rect 19107 18309 19119 18343
rect 19061 18303 19119 18309
rect 22281 18343 22339 18349
rect 22281 18309 22293 18343
rect 22327 18340 22339 18343
rect 24210 18340 24216 18352
rect 22327 18312 24216 18340
rect 22327 18309 22339 18312
rect 22281 18303 22339 18309
rect 16577 18275 16635 18281
rect 16577 18241 16589 18275
rect 16623 18272 16635 18275
rect 17678 18272 17684 18284
rect 16623 18244 17684 18272
rect 16623 18241 16635 18244
rect 16577 18235 16635 18241
rect 17678 18232 17684 18244
rect 17736 18232 17742 18284
rect 19702 18272 19708 18284
rect 19615 18244 19708 18272
rect 19702 18232 19708 18244
rect 19760 18272 19766 18284
rect 20438 18272 20444 18284
rect 19760 18244 20444 18272
rect 19760 18232 19766 18244
rect 20438 18232 20444 18244
rect 20496 18232 20502 18284
rect 21818 18232 21824 18284
rect 21876 18272 21882 18284
rect 22388 18272 22416 18312
rect 24210 18300 24216 18312
rect 24268 18300 24274 18352
rect 31938 18300 31944 18352
rect 31996 18340 32002 18352
rect 32033 18343 32091 18349
rect 32033 18340 32045 18343
rect 31996 18312 32045 18340
rect 31996 18300 32002 18312
rect 32033 18309 32045 18312
rect 32079 18309 32091 18343
rect 32033 18303 32091 18309
rect 32677 18343 32735 18349
rect 32677 18309 32689 18343
rect 32723 18340 32735 18343
rect 32950 18340 32956 18352
rect 32723 18312 32956 18340
rect 32723 18309 32735 18312
rect 32677 18303 32735 18309
rect 32950 18300 32956 18312
rect 33008 18300 33014 18352
rect 21876 18244 22416 18272
rect 21876 18232 21882 18244
rect 14093 18207 14151 18213
rect 14093 18173 14105 18207
rect 14139 18173 14151 18207
rect 14734 18204 14740 18216
rect 14695 18176 14740 18204
rect 14093 18167 14151 18173
rect 14734 18164 14740 18176
rect 14792 18164 14798 18216
rect 14829 18207 14887 18213
rect 14829 18173 14841 18207
rect 14875 18173 14887 18207
rect 14829 18167 14887 18173
rect 16669 18207 16727 18213
rect 16669 18173 16681 18207
rect 16715 18204 16727 18207
rect 16942 18204 16948 18216
rect 16715 18176 16948 18204
rect 16715 18173 16727 18176
rect 16669 18167 16727 18173
rect 7561 18139 7619 18145
rect 7561 18105 7573 18139
rect 7607 18105 7619 18139
rect 7926 18136 7932 18148
rect 7887 18108 7932 18136
rect 7561 18099 7619 18105
rect 4522 18068 4528 18080
rect 4483 18040 4528 18068
rect 4522 18028 4528 18040
rect 4580 18028 4586 18080
rect 5994 18028 6000 18080
rect 6052 18068 6058 18080
rect 6181 18071 6239 18077
rect 6181 18068 6193 18071
rect 6052 18040 6193 18068
rect 6052 18028 6058 18040
rect 6181 18037 6193 18040
rect 6227 18068 6239 18071
rect 6454 18068 6460 18080
rect 6227 18040 6460 18068
rect 6227 18037 6239 18040
rect 6181 18031 6239 18037
rect 6454 18028 6460 18040
rect 6512 18028 6518 18080
rect 6914 18028 6920 18080
rect 6972 18068 6978 18080
rect 7469 18071 7527 18077
rect 7469 18068 7481 18071
rect 6972 18040 7481 18068
rect 6972 18028 6978 18040
rect 7469 18037 7481 18040
rect 7515 18037 7527 18071
rect 7576 18068 7604 18099
rect 7926 18096 7932 18108
rect 7984 18096 7990 18148
rect 8389 18139 8447 18145
rect 8389 18105 8401 18139
rect 8435 18136 8447 18139
rect 8481 18139 8539 18145
rect 8481 18136 8493 18139
rect 8435 18108 8493 18136
rect 8435 18105 8447 18108
rect 8389 18099 8447 18105
rect 8481 18105 8493 18108
rect 8527 18136 8539 18139
rect 9214 18136 9220 18148
rect 8527 18108 8800 18136
rect 9175 18108 9220 18136
rect 8527 18105 8539 18108
rect 8481 18099 8539 18105
rect 8202 18068 8208 18080
rect 7576 18040 8208 18068
rect 7469 18031 7527 18037
rect 8202 18028 8208 18040
rect 8260 18068 8266 18080
rect 8662 18068 8668 18080
rect 8260 18040 8668 18068
rect 8260 18028 8266 18040
rect 8662 18028 8668 18040
rect 8720 18028 8726 18080
rect 8772 18068 8800 18108
rect 9214 18096 9220 18108
rect 9272 18096 9278 18148
rect 10137 18139 10195 18145
rect 10137 18105 10149 18139
rect 10183 18136 10195 18139
rect 10778 18136 10784 18148
rect 10183 18108 10784 18136
rect 10183 18105 10195 18108
rect 10137 18099 10195 18105
rect 10778 18096 10784 18108
rect 10836 18096 10842 18148
rect 13262 18136 13268 18148
rect 13223 18108 13268 18136
rect 13262 18096 13268 18108
rect 13320 18096 13326 18148
rect 14182 18096 14188 18148
rect 14240 18136 14246 18148
rect 14844 18136 14872 18167
rect 16942 18164 16948 18176
rect 17000 18204 17006 18216
rect 17000 18176 17264 18204
rect 17000 18164 17006 18176
rect 17129 18139 17187 18145
rect 17129 18136 17141 18139
rect 14240 18108 14872 18136
rect 16040 18108 17141 18136
rect 14240 18096 14246 18108
rect 9030 18068 9036 18080
rect 8772 18040 9036 18068
rect 9030 18028 9036 18040
rect 9088 18068 9094 18080
rect 9582 18068 9588 18080
rect 9088 18040 9588 18068
rect 9088 18028 9094 18040
rect 9582 18028 9588 18040
rect 9640 18028 9646 18080
rect 10226 18028 10232 18080
rect 10284 18068 10290 18080
rect 10594 18068 10600 18080
rect 10284 18040 10600 18068
rect 10284 18028 10290 18040
rect 10594 18028 10600 18040
rect 10652 18028 10658 18080
rect 12805 18071 12863 18077
rect 12805 18037 12817 18071
rect 12851 18068 12863 18071
rect 14200 18068 14228 18096
rect 16040 18080 16068 18108
rect 17129 18105 17141 18108
rect 17175 18105 17187 18139
rect 17236 18136 17264 18176
rect 17402 18164 17408 18216
rect 17460 18204 17466 18216
rect 17589 18207 17647 18213
rect 17589 18204 17601 18207
rect 17460 18176 17601 18204
rect 17460 18164 17466 18176
rect 17589 18173 17601 18176
rect 17635 18204 17647 18207
rect 17773 18207 17831 18213
rect 17773 18204 17785 18207
rect 17635 18176 17785 18204
rect 17635 18173 17647 18176
rect 17589 18167 17647 18173
rect 17773 18173 17785 18176
rect 17819 18173 17831 18207
rect 17773 18167 17831 18173
rect 18141 18207 18199 18213
rect 18141 18173 18153 18207
rect 18187 18173 18199 18207
rect 19981 18207 20039 18213
rect 19981 18204 19993 18207
rect 18141 18167 18199 18173
rect 19536 18176 19993 18204
rect 17497 18139 17555 18145
rect 17497 18136 17509 18139
rect 17236 18108 17509 18136
rect 17129 18099 17187 18105
rect 17497 18105 17509 18108
rect 17543 18136 17555 18139
rect 18049 18139 18107 18145
rect 18049 18136 18061 18139
rect 17543 18108 18061 18136
rect 17543 18105 17555 18108
rect 17497 18099 17555 18105
rect 18049 18105 18061 18108
rect 18095 18105 18107 18139
rect 18049 18099 18107 18105
rect 16022 18068 16028 18080
rect 12851 18040 14228 18068
rect 15983 18040 16028 18068
rect 12851 18037 12863 18040
rect 12805 18031 12863 18037
rect 16022 18028 16028 18040
rect 16080 18028 16086 18080
rect 17589 18071 17647 18077
rect 17589 18037 17601 18071
rect 17635 18068 17647 18071
rect 17770 18068 17776 18080
rect 17635 18040 17776 18068
rect 17635 18037 17647 18040
rect 17589 18031 17647 18037
rect 17770 18028 17776 18040
rect 17828 18068 17834 18080
rect 18156 18068 18184 18167
rect 19242 18068 19248 18080
rect 17828 18040 19248 18068
rect 17828 18028 17834 18040
rect 19242 18028 19248 18040
rect 19300 18028 19306 18080
rect 19426 18028 19432 18080
rect 19484 18068 19490 18080
rect 19536 18077 19564 18176
rect 19981 18173 19993 18176
rect 20027 18204 20039 18207
rect 20622 18204 20628 18216
rect 20027 18176 20628 18204
rect 20027 18173 20039 18176
rect 19981 18167 20039 18173
rect 20622 18164 20628 18176
rect 20680 18164 20686 18216
rect 22388 18213 22416 18244
rect 25774 18232 25780 18284
rect 25832 18272 25838 18284
rect 25961 18275 26019 18281
rect 25961 18272 25973 18275
rect 25832 18244 25973 18272
rect 25832 18232 25838 18244
rect 25961 18241 25973 18244
rect 26007 18241 26019 18275
rect 28074 18272 28080 18284
rect 28035 18244 28080 18272
rect 25961 18235 26019 18241
rect 28074 18232 28080 18244
rect 28132 18232 28138 18284
rect 28166 18232 28172 18284
rect 28224 18272 28230 18284
rect 30101 18275 30159 18281
rect 30101 18272 30113 18275
rect 28224 18244 30113 18272
rect 28224 18232 28230 18244
rect 30101 18241 30113 18244
rect 30147 18241 30159 18275
rect 30101 18235 30159 18241
rect 30834 18232 30840 18284
rect 30892 18272 30898 18284
rect 31113 18275 31171 18281
rect 31113 18272 31125 18275
rect 30892 18244 31125 18272
rect 30892 18232 30898 18244
rect 31113 18241 31125 18244
rect 31159 18272 31171 18275
rect 31389 18275 31447 18281
rect 31389 18272 31401 18275
rect 31159 18244 31401 18272
rect 31159 18241 31171 18244
rect 31113 18235 31171 18241
rect 31389 18241 31401 18244
rect 31435 18272 31447 18275
rect 33060 18272 33088 18368
rect 33502 18300 33508 18352
rect 33560 18340 33566 18352
rect 33689 18343 33747 18349
rect 33689 18340 33701 18343
rect 33560 18312 33701 18340
rect 33560 18300 33566 18312
rect 33689 18309 33701 18312
rect 33735 18309 33747 18343
rect 33689 18303 33747 18309
rect 31435 18244 33088 18272
rect 31435 18241 31447 18244
rect 31389 18235 31447 18241
rect 22373 18207 22431 18213
rect 22373 18173 22385 18207
rect 22419 18173 22431 18207
rect 22373 18167 22431 18173
rect 24121 18207 24179 18213
rect 24121 18173 24133 18207
rect 24167 18204 24179 18207
rect 25041 18207 25099 18213
rect 24167 18176 24716 18204
rect 24167 18173 24179 18176
rect 24121 18167 24179 18173
rect 21361 18139 21419 18145
rect 21361 18105 21373 18139
rect 21407 18136 21419 18139
rect 21910 18136 21916 18148
rect 21407 18108 21916 18136
rect 21407 18105 21419 18108
rect 21361 18099 21419 18105
rect 21910 18096 21916 18108
rect 21968 18096 21974 18148
rect 19521 18071 19579 18077
rect 19521 18068 19533 18071
rect 19484 18040 19533 18068
rect 19484 18028 19490 18040
rect 19521 18037 19533 18040
rect 19567 18037 19579 18071
rect 19521 18031 19579 18037
rect 22002 18028 22008 18080
rect 22060 18068 22066 18080
rect 22094 18068 22100 18080
rect 22060 18040 22100 18068
rect 22060 18028 22066 18040
rect 22094 18028 22100 18040
rect 22152 18068 22158 18080
rect 22557 18071 22615 18077
rect 22557 18068 22569 18071
rect 22152 18040 22569 18068
rect 22152 18028 22158 18040
rect 22557 18037 22569 18040
rect 22603 18037 22615 18071
rect 22557 18031 22615 18037
rect 23658 18028 23664 18080
rect 23716 18068 23722 18080
rect 24486 18068 24492 18080
rect 23716 18040 24492 18068
rect 23716 18028 23722 18040
rect 24486 18028 24492 18040
rect 24544 18028 24550 18080
rect 24688 18077 24716 18176
rect 25041 18173 25053 18207
rect 25087 18204 25099 18207
rect 25130 18204 25136 18216
rect 25087 18176 25136 18204
rect 25087 18173 25099 18176
rect 25041 18167 25099 18173
rect 25130 18164 25136 18176
rect 25188 18164 25194 18216
rect 25682 18204 25688 18216
rect 25643 18176 25688 18204
rect 25682 18164 25688 18176
rect 25740 18164 25746 18216
rect 26050 18204 26056 18216
rect 26011 18176 26056 18204
rect 26050 18164 26056 18176
rect 26108 18164 26114 18216
rect 27341 18207 27399 18213
rect 27341 18173 27353 18207
rect 27387 18204 27399 18207
rect 27614 18204 27620 18216
rect 27387 18176 27620 18204
rect 27387 18173 27399 18176
rect 27341 18167 27399 18173
rect 27614 18164 27620 18176
rect 27672 18204 27678 18216
rect 28353 18207 28411 18213
rect 28353 18204 28365 18207
rect 27672 18176 28365 18204
rect 27672 18164 27678 18176
rect 28353 18173 28365 18176
rect 28399 18204 28411 18207
rect 28626 18204 28632 18216
rect 28399 18176 28632 18204
rect 28399 18173 28411 18176
rect 28353 18167 28411 18173
rect 28626 18164 28632 18176
rect 28684 18164 28690 18216
rect 29273 18207 29331 18213
rect 29273 18173 29285 18207
rect 29319 18204 29331 18207
rect 29914 18204 29920 18216
rect 29319 18176 29920 18204
rect 29319 18173 29331 18176
rect 29273 18167 29331 18173
rect 29914 18164 29920 18176
rect 29972 18164 29978 18216
rect 31202 18164 31208 18216
rect 31260 18204 31266 18216
rect 31573 18207 31631 18213
rect 31573 18204 31585 18207
rect 31260 18176 31585 18204
rect 31260 18164 31266 18176
rect 31573 18173 31585 18176
rect 31619 18204 31631 18207
rect 31754 18204 31760 18216
rect 31619 18176 31760 18204
rect 31619 18173 31631 18176
rect 31573 18167 31631 18173
rect 31754 18164 31760 18176
rect 31812 18164 31818 18216
rect 32033 18207 32091 18213
rect 32033 18173 32045 18207
rect 32079 18173 32091 18207
rect 32033 18167 32091 18173
rect 27249 18139 27307 18145
rect 27249 18105 27261 18139
rect 27295 18136 27307 18139
rect 27709 18139 27767 18145
rect 27709 18136 27721 18139
rect 27295 18108 27721 18136
rect 27295 18105 27307 18108
rect 27249 18099 27307 18105
rect 27709 18105 27721 18108
rect 27755 18136 27767 18139
rect 27798 18136 27804 18148
rect 27755 18108 27804 18136
rect 27755 18105 27767 18108
rect 27709 18099 27767 18105
rect 27798 18096 27804 18108
rect 27856 18096 27862 18148
rect 30745 18139 30803 18145
rect 30745 18105 30757 18139
rect 30791 18136 30803 18139
rect 32048 18136 32076 18167
rect 33060 18148 33088 18244
rect 32214 18136 32220 18148
rect 30791 18108 32220 18136
rect 30791 18105 30803 18108
rect 30745 18099 30803 18105
rect 32214 18096 32220 18108
rect 32272 18096 32278 18148
rect 33042 18136 33048 18148
rect 33003 18108 33048 18136
rect 33042 18096 33048 18108
rect 33100 18096 33106 18148
rect 24673 18071 24731 18077
rect 24673 18037 24685 18071
rect 24719 18068 24731 18071
rect 24762 18068 24768 18080
rect 24719 18040 24768 18068
rect 24719 18037 24731 18040
rect 24673 18031 24731 18037
rect 24762 18028 24768 18040
rect 24820 18028 24826 18080
rect 26881 18071 26939 18077
rect 26881 18037 26893 18071
rect 26927 18068 26939 18071
rect 26970 18068 26976 18080
rect 26927 18040 26976 18068
rect 26927 18037 26939 18040
rect 26881 18031 26939 18037
rect 26970 18028 26976 18040
rect 27028 18028 27034 18080
rect 27430 18028 27436 18080
rect 27488 18068 27494 18080
rect 27525 18071 27583 18077
rect 27525 18068 27537 18071
rect 27488 18040 27537 18068
rect 27488 18028 27494 18040
rect 27525 18037 27537 18040
rect 27571 18037 27583 18071
rect 27525 18031 27583 18037
rect 27617 18071 27675 18077
rect 27617 18037 27629 18071
rect 27663 18068 27675 18071
rect 27890 18068 27896 18080
rect 27663 18040 27896 18068
rect 27663 18037 27675 18040
rect 27617 18031 27675 18037
rect 27890 18028 27896 18040
rect 27948 18028 27954 18080
rect 29457 18071 29515 18077
rect 29457 18037 29469 18071
rect 29503 18068 29515 18071
rect 29638 18068 29644 18080
rect 29503 18040 29644 18068
rect 29503 18037 29515 18040
rect 29457 18031 29515 18037
rect 29638 18028 29644 18040
rect 29696 18028 29702 18080
rect 31478 18028 31484 18080
rect 31536 18068 31542 18080
rect 32766 18068 32772 18080
rect 31536 18040 32772 18068
rect 31536 18028 31542 18040
rect 32766 18028 32772 18040
rect 32824 18068 32830 18080
rect 33321 18071 33379 18077
rect 33321 18068 33333 18071
rect 32824 18040 33333 18068
rect 32824 18028 32830 18040
rect 33321 18037 33333 18040
rect 33367 18068 33379 18071
rect 33778 18068 33784 18080
rect 33367 18040 33784 18068
rect 33367 18037 33379 18040
rect 33321 18031 33379 18037
rect 33778 18028 33784 18040
rect 33836 18028 33842 18080
rect 1104 17978 38548 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 38548 17978
rect 1104 17904 38548 17926
rect 1854 17864 1860 17876
rect 1815 17836 1860 17864
rect 1854 17824 1860 17836
rect 1912 17824 1918 17876
rect 3326 17864 3332 17876
rect 2424 17836 3332 17864
rect 1946 17796 1952 17808
rect 1907 17768 1952 17796
rect 1946 17756 1952 17768
rect 2004 17756 2010 17808
rect 2424 17740 2452 17836
rect 3326 17824 3332 17836
rect 3384 17824 3390 17876
rect 4614 17864 4620 17876
rect 4575 17836 4620 17864
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 5166 17864 5172 17876
rect 5127 17836 5172 17864
rect 5166 17824 5172 17836
rect 5224 17824 5230 17876
rect 7006 17824 7012 17876
rect 7064 17864 7070 17876
rect 7193 17867 7251 17873
rect 7193 17864 7205 17867
rect 7064 17836 7205 17864
rect 7064 17824 7070 17836
rect 7193 17833 7205 17836
rect 7239 17833 7251 17867
rect 7193 17827 7251 17833
rect 4985 17799 5043 17805
rect 4985 17765 4997 17799
rect 5031 17796 5043 17799
rect 7208 17796 7236 17827
rect 7374 17824 7380 17876
rect 7432 17864 7438 17876
rect 7653 17867 7711 17873
rect 7653 17864 7665 17867
rect 7432 17836 7665 17864
rect 7432 17824 7438 17836
rect 7653 17833 7665 17836
rect 7699 17833 7711 17867
rect 7653 17827 7711 17833
rect 8478 17824 8484 17876
rect 8536 17864 8542 17876
rect 8665 17867 8723 17873
rect 8665 17864 8677 17867
rect 8536 17836 8677 17864
rect 8536 17824 8542 17836
rect 8665 17833 8677 17836
rect 8711 17833 8723 17867
rect 11514 17864 11520 17876
rect 11475 17836 11520 17864
rect 8665 17827 8723 17833
rect 11514 17824 11520 17836
rect 11572 17824 11578 17876
rect 11698 17824 11704 17876
rect 11756 17864 11762 17876
rect 12345 17867 12403 17873
rect 11756 17836 12112 17864
rect 11756 17824 11762 17836
rect 9122 17796 9128 17808
rect 5031 17768 5948 17796
rect 7208 17768 9128 17796
rect 5031 17765 5043 17768
rect 4985 17759 5043 17765
rect 5920 17740 5948 17768
rect 9122 17756 9128 17768
rect 9180 17796 9186 17808
rect 9398 17796 9404 17808
rect 9180 17768 9404 17796
rect 9180 17756 9186 17768
rect 9398 17756 9404 17768
rect 9456 17796 9462 17808
rect 10042 17796 10048 17808
rect 9456 17768 10048 17796
rect 9456 17756 9462 17768
rect 2406 17728 2412 17740
rect 2319 17700 2412 17728
rect 2406 17688 2412 17700
rect 2464 17688 2470 17740
rect 2498 17688 2504 17740
rect 2556 17728 2562 17740
rect 2593 17731 2651 17737
rect 2593 17728 2605 17731
rect 2556 17700 2605 17728
rect 2556 17688 2562 17700
rect 2593 17697 2605 17700
rect 2639 17728 2651 17731
rect 2682 17728 2688 17740
rect 2639 17700 2688 17728
rect 2639 17697 2651 17700
rect 2593 17691 2651 17697
rect 2682 17688 2688 17700
rect 2740 17688 2746 17740
rect 2961 17731 3019 17737
rect 2961 17697 2973 17731
rect 3007 17728 3019 17731
rect 3510 17728 3516 17740
rect 3007 17700 3516 17728
rect 3007 17697 3019 17700
rect 2961 17691 3019 17697
rect 3510 17688 3516 17700
rect 3568 17688 3574 17740
rect 5353 17731 5411 17737
rect 5353 17697 5365 17731
rect 5399 17697 5411 17731
rect 5534 17728 5540 17740
rect 5495 17700 5540 17728
rect 5353 17691 5411 17697
rect 2869 17663 2927 17669
rect 2869 17629 2881 17663
rect 2915 17660 2927 17663
rect 3234 17660 3240 17672
rect 2915 17632 3240 17660
rect 2915 17629 2927 17632
rect 2869 17623 2927 17629
rect 3234 17620 3240 17632
rect 3292 17620 3298 17672
rect 5368 17660 5396 17691
rect 5534 17688 5540 17700
rect 5592 17688 5598 17740
rect 5902 17728 5908 17740
rect 5863 17700 5908 17728
rect 5902 17688 5908 17700
rect 5960 17688 5966 17740
rect 6638 17688 6644 17740
rect 6696 17728 6702 17740
rect 7009 17731 7067 17737
rect 7009 17728 7021 17731
rect 6696 17700 7021 17728
rect 6696 17688 6702 17700
rect 7009 17697 7021 17700
rect 7055 17697 7067 17731
rect 8018 17728 8024 17740
rect 7979 17700 8024 17728
rect 7009 17691 7067 17697
rect 8018 17688 8024 17700
rect 8076 17728 8082 17740
rect 8202 17728 8208 17740
rect 8076 17700 8208 17728
rect 8076 17688 8082 17700
rect 8202 17688 8208 17700
rect 8260 17688 8266 17740
rect 9493 17731 9551 17737
rect 9493 17697 9505 17731
rect 9539 17728 9551 17731
rect 9674 17728 9680 17740
rect 9539 17700 9680 17728
rect 9539 17697 9551 17700
rect 9493 17691 9551 17697
rect 9674 17688 9680 17700
rect 9732 17688 9738 17740
rect 9968 17737 9996 17768
rect 10042 17756 10048 17768
rect 10100 17796 10106 17808
rect 10689 17799 10747 17805
rect 10689 17796 10701 17799
rect 10100 17768 10701 17796
rect 10100 17756 10106 17768
rect 10689 17765 10701 17768
rect 10735 17765 10747 17799
rect 11606 17796 11612 17808
rect 11567 17768 11612 17796
rect 10689 17759 10747 17765
rect 11606 17756 11612 17768
rect 11664 17756 11670 17808
rect 11974 17796 11980 17808
rect 11935 17768 11980 17796
rect 11974 17756 11980 17768
rect 12032 17756 12038 17808
rect 12084 17796 12112 17836
rect 12345 17833 12357 17867
rect 12391 17864 12403 17867
rect 12434 17864 12440 17876
rect 12391 17836 12440 17864
rect 12391 17833 12403 17836
rect 12345 17827 12403 17833
rect 12434 17824 12440 17836
rect 12492 17824 12498 17876
rect 12710 17864 12716 17876
rect 12671 17836 12716 17864
rect 12710 17824 12716 17836
rect 12768 17824 12774 17876
rect 15378 17864 15384 17876
rect 12820 17836 15384 17864
rect 12526 17796 12532 17808
rect 12084 17768 12532 17796
rect 12526 17756 12532 17768
rect 12584 17796 12590 17808
rect 12820 17796 12848 17836
rect 15378 17824 15384 17836
rect 15436 17864 15442 17876
rect 15473 17867 15531 17873
rect 15473 17864 15485 17867
rect 15436 17836 15485 17864
rect 15436 17824 15442 17836
rect 15473 17833 15485 17836
rect 15519 17833 15531 17867
rect 15473 17827 15531 17833
rect 17402 17824 17408 17876
rect 17460 17864 17466 17876
rect 17770 17864 17776 17876
rect 17460 17836 17776 17864
rect 17460 17824 17466 17836
rect 17770 17824 17776 17836
rect 17828 17824 17834 17876
rect 17954 17824 17960 17876
rect 18012 17864 18018 17876
rect 18049 17867 18107 17873
rect 18049 17864 18061 17867
rect 18012 17836 18061 17864
rect 18012 17824 18018 17836
rect 18049 17833 18061 17836
rect 18095 17833 18107 17867
rect 18414 17864 18420 17876
rect 18375 17836 18420 17864
rect 18049 17827 18107 17833
rect 18414 17824 18420 17836
rect 18472 17824 18478 17876
rect 20254 17824 20260 17876
rect 20312 17864 20318 17876
rect 20625 17867 20683 17873
rect 20625 17864 20637 17867
rect 20312 17836 20637 17864
rect 20312 17824 20318 17836
rect 20625 17833 20637 17836
rect 20671 17864 20683 17867
rect 20898 17864 20904 17876
rect 20671 17836 20904 17864
rect 20671 17833 20683 17836
rect 20625 17827 20683 17833
rect 20898 17824 20904 17836
rect 20956 17824 20962 17876
rect 21545 17867 21603 17873
rect 21545 17833 21557 17867
rect 21591 17864 21603 17867
rect 22002 17864 22008 17876
rect 21591 17836 22008 17864
rect 21591 17833 21603 17836
rect 21545 17827 21603 17833
rect 22002 17824 22008 17836
rect 22060 17824 22066 17876
rect 23937 17867 23995 17873
rect 23937 17833 23949 17867
rect 23983 17864 23995 17867
rect 25406 17864 25412 17876
rect 23983 17836 25412 17864
rect 23983 17833 23995 17836
rect 23937 17827 23995 17833
rect 25406 17824 25412 17836
rect 25464 17824 25470 17876
rect 26697 17867 26755 17873
rect 26697 17833 26709 17867
rect 26743 17864 26755 17867
rect 26743 17836 27476 17864
rect 26743 17833 26755 17836
rect 26697 17827 26755 17833
rect 12584 17768 12848 17796
rect 12584 17756 12590 17768
rect 13538 17756 13544 17808
rect 13596 17796 13602 17808
rect 13633 17799 13691 17805
rect 13633 17796 13645 17799
rect 13596 17768 13645 17796
rect 13596 17756 13602 17768
rect 13633 17765 13645 17768
rect 13679 17765 13691 17799
rect 17586 17796 17592 17808
rect 13633 17759 13691 17765
rect 16132 17768 17592 17796
rect 9953 17731 10011 17737
rect 9953 17697 9965 17731
rect 9999 17697 10011 17731
rect 9953 17691 10011 17697
rect 11146 17688 11152 17740
rect 11204 17728 11210 17740
rect 11241 17731 11299 17737
rect 11241 17728 11253 17731
rect 11204 17700 11253 17728
rect 11204 17688 11210 17700
rect 11241 17697 11253 17700
rect 11287 17697 11299 17731
rect 11241 17691 11299 17697
rect 11330 17688 11336 17740
rect 11388 17728 11394 17740
rect 11425 17731 11483 17737
rect 11425 17728 11437 17731
rect 11388 17700 11437 17728
rect 11388 17688 11394 17700
rect 11425 17697 11437 17700
rect 11471 17697 11483 17731
rect 11425 17691 11483 17697
rect 13173 17731 13231 17737
rect 13173 17697 13185 17731
rect 13219 17728 13231 17731
rect 13354 17728 13360 17740
rect 13219 17700 13360 17728
rect 13219 17697 13231 17700
rect 13173 17691 13231 17697
rect 13354 17688 13360 17700
rect 13412 17688 13418 17740
rect 16132 17737 16160 17768
rect 17586 17756 17592 17768
rect 17644 17756 17650 17808
rect 22554 17796 22560 17808
rect 22515 17768 22560 17796
rect 22554 17756 22560 17768
rect 22612 17756 22618 17808
rect 24394 17796 24400 17808
rect 24355 17768 24400 17796
rect 24394 17756 24400 17768
rect 24452 17756 24458 17808
rect 16117 17731 16175 17737
rect 16117 17697 16129 17731
rect 16163 17697 16175 17731
rect 16117 17691 16175 17697
rect 16485 17731 16543 17737
rect 16485 17697 16497 17731
rect 16531 17728 16543 17731
rect 16574 17728 16580 17740
rect 16531 17700 16580 17728
rect 16531 17697 16543 17700
rect 16485 17691 16543 17697
rect 16574 17688 16580 17700
rect 16632 17688 16638 17740
rect 16669 17731 16727 17737
rect 16669 17697 16681 17731
rect 16715 17697 16727 17731
rect 16669 17691 16727 17697
rect 17313 17731 17371 17737
rect 17313 17697 17325 17731
rect 17359 17728 17371 17731
rect 17770 17728 17776 17740
rect 17359 17700 17632 17728
rect 17731 17700 17776 17728
rect 17359 17697 17371 17700
rect 17313 17691 17371 17697
rect 5442 17660 5448 17672
rect 5368 17632 5448 17660
rect 5442 17620 5448 17632
rect 5500 17620 5506 17672
rect 5552 17660 5580 17688
rect 6457 17663 6515 17669
rect 6457 17660 6469 17663
rect 5552 17632 6469 17660
rect 6457 17629 6469 17632
rect 6503 17660 6515 17663
rect 6914 17660 6920 17672
rect 6503 17632 6920 17660
rect 6503 17629 6515 17632
rect 6457 17623 6515 17629
rect 6914 17620 6920 17632
rect 6972 17620 6978 17672
rect 8386 17660 8392 17672
rect 8347 17632 8392 17660
rect 8386 17620 8392 17632
rect 8444 17620 8450 17672
rect 10413 17663 10471 17669
rect 10413 17629 10425 17663
rect 10459 17660 10471 17663
rect 11054 17660 11060 17672
rect 10459 17632 11060 17660
rect 10459 17629 10471 17632
rect 10413 17623 10471 17629
rect 11054 17620 11060 17632
rect 11112 17620 11118 17672
rect 13078 17660 13084 17672
rect 12991 17632 13084 17660
rect 13078 17620 13084 17632
rect 13136 17660 13142 17672
rect 14645 17663 14703 17669
rect 14645 17660 14657 17663
rect 13136 17632 14657 17660
rect 13136 17620 13142 17632
rect 14645 17629 14657 17632
rect 14691 17660 14703 17663
rect 14734 17660 14740 17672
rect 14691 17632 14740 17660
rect 14691 17629 14703 17632
rect 14645 17623 14703 17629
rect 14734 17620 14740 17632
rect 14792 17620 14798 17672
rect 15838 17660 15844 17672
rect 15799 17632 15844 17660
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 16022 17620 16028 17672
rect 16080 17660 16086 17672
rect 16684 17660 16712 17691
rect 16080 17632 16712 17660
rect 16080 17620 16086 17632
rect 8294 17592 8300 17604
rect 8255 17564 8300 17592
rect 8294 17552 8300 17564
rect 8352 17552 8358 17604
rect 8570 17552 8576 17604
rect 8628 17592 8634 17604
rect 8628 17564 9260 17592
rect 8628 17552 8634 17564
rect 3878 17524 3884 17536
rect 3839 17496 3884 17524
rect 3878 17484 3884 17496
rect 3936 17484 3942 17536
rect 6917 17527 6975 17533
rect 6917 17493 6929 17527
rect 6963 17524 6975 17527
rect 7466 17524 7472 17536
rect 6963 17496 7472 17524
rect 6963 17493 6975 17496
rect 6917 17487 6975 17493
rect 7466 17484 7472 17496
rect 7524 17484 7530 17536
rect 8110 17484 8116 17536
rect 8168 17533 8174 17536
rect 8168 17527 8217 17533
rect 8168 17493 8171 17527
rect 8205 17493 8217 17527
rect 8168 17487 8217 17493
rect 8168 17484 8174 17487
rect 8938 17484 8944 17536
rect 8996 17524 9002 17536
rect 9033 17527 9091 17533
rect 9033 17524 9045 17527
rect 8996 17496 9045 17524
rect 8996 17484 9002 17496
rect 9033 17493 9045 17496
rect 9079 17493 9091 17527
rect 9232 17524 9260 17564
rect 9306 17552 9312 17604
rect 9364 17592 9370 17604
rect 9766 17592 9772 17604
rect 9364 17564 9772 17592
rect 9364 17552 9370 17564
rect 9766 17552 9772 17564
rect 9824 17592 9830 17604
rect 11149 17595 11207 17601
rect 11149 17592 11161 17595
rect 9824 17564 11161 17592
rect 9824 17552 9830 17564
rect 11149 17561 11161 17564
rect 11195 17561 11207 17595
rect 17604 17592 17632 17700
rect 17770 17688 17776 17700
rect 17828 17688 17834 17740
rect 19429 17731 19487 17737
rect 19429 17697 19441 17731
rect 19475 17728 19487 17731
rect 22097 17731 22155 17737
rect 19475 17700 19932 17728
rect 19475 17697 19487 17700
rect 19429 17691 19487 17697
rect 18690 17620 18696 17672
rect 18748 17660 18754 17672
rect 18785 17663 18843 17669
rect 18785 17660 18797 17663
rect 18748 17632 18797 17660
rect 18748 17620 18754 17632
rect 18785 17629 18797 17632
rect 18831 17629 18843 17663
rect 18785 17623 18843 17629
rect 17604 17564 18828 17592
rect 11149 17555 11207 17561
rect 18800 17536 18828 17564
rect 9582 17524 9588 17536
rect 9232 17496 9588 17524
rect 9033 17487 9091 17493
rect 9582 17484 9588 17496
rect 9640 17484 9646 17536
rect 14274 17524 14280 17536
rect 14235 17496 14280 17524
rect 14274 17484 14280 17496
rect 14332 17484 14338 17536
rect 14826 17484 14832 17536
rect 14884 17524 14890 17536
rect 15010 17524 15016 17536
rect 14884 17496 15016 17524
rect 14884 17484 14890 17496
rect 15010 17484 15016 17496
rect 15068 17484 15074 17536
rect 18782 17484 18788 17536
rect 18840 17484 18846 17536
rect 19904 17533 19932 17700
rect 22097 17697 22109 17731
rect 22143 17728 22155 17731
rect 23106 17728 23112 17740
rect 22143 17700 23112 17728
rect 22143 17697 22155 17700
rect 22097 17691 22155 17697
rect 23106 17688 23112 17700
rect 23164 17688 23170 17740
rect 23198 17688 23204 17740
rect 23256 17728 23262 17740
rect 23385 17731 23443 17737
rect 23385 17728 23397 17731
rect 23256 17700 23397 17728
rect 23256 17688 23262 17700
rect 23385 17697 23397 17700
rect 23431 17697 23443 17731
rect 23385 17691 23443 17697
rect 23569 17731 23627 17737
rect 23569 17697 23581 17731
rect 23615 17728 23627 17731
rect 23658 17728 23664 17740
rect 23615 17700 23664 17728
rect 23615 17697 23627 17700
rect 23569 17691 23627 17697
rect 22922 17620 22928 17672
rect 22980 17660 22986 17672
rect 23584 17660 23612 17691
rect 23658 17688 23664 17700
rect 23716 17728 23722 17740
rect 23934 17728 23940 17740
rect 23716 17700 23940 17728
rect 23716 17688 23722 17700
rect 23934 17688 23940 17700
rect 23992 17688 23998 17740
rect 25225 17731 25283 17737
rect 25225 17728 25237 17731
rect 24228 17700 25237 17728
rect 22980 17632 23612 17660
rect 22980 17620 22986 17632
rect 24228 17604 24256 17700
rect 25225 17697 25237 17700
rect 25271 17697 25283 17731
rect 25958 17728 25964 17740
rect 25225 17691 25283 17697
rect 25332 17700 25964 17728
rect 24949 17663 25007 17669
rect 24949 17629 24961 17663
rect 24995 17660 25007 17663
rect 25332 17660 25360 17700
rect 25958 17688 25964 17700
rect 26016 17688 26022 17740
rect 26510 17728 26516 17740
rect 26471 17700 26516 17728
rect 26510 17688 26516 17700
rect 26568 17688 26574 17740
rect 24995 17632 25360 17660
rect 24995 17629 25007 17632
rect 24949 17623 25007 17629
rect 22465 17595 22523 17601
rect 22465 17561 22477 17595
rect 22511 17592 22523 17595
rect 24210 17592 24216 17604
rect 22511 17564 24072 17592
rect 24171 17564 24216 17592
rect 22511 17561 22523 17564
rect 22465 17555 22523 17561
rect 19889 17527 19947 17533
rect 19889 17493 19901 17527
rect 19935 17524 19947 17527
rect 19978 17524 19984 17536
rect 19935 17496 19984 17524
rect 19935 17493 19947 17496
rect 19889 17487 19947 17493
rect 19978 17484 19984 17496
rect 20036 17524 20042 17536
rect 20165 17527 20223 17533
rect 20165 17524 20177 17527
rect 20036 17496 20177 17524
rect 20036 17484 20042 17496
rect 20165 17493 20177 17496
rect 20211 17493 20223 17527
rect 24044 17524 24072 17564
rect 24210 17552 24216 17564
rect 24268 17552 24274 17604
rect 24964 17524 24992 17623
rect 25406 17620 25412 17672
rect 25464 17660 25470 17672
rect 27448 17669 27476 17836
rect 29178 17824 29184 17876
rect 29236 17864 29242 17876
rect 29730 17864 29736 17876
rect 29236 17836 29736 17864
rect 29236 17824 29242 17836
rect 29730 17824 29736 17836
rect 29788 17824 29794 17876
rect 30834 17864 30840 17876
rect 30795 17836 30840 17864
rect 30834 17824 30840 17836
rect 30892 17824 30898 17876
rect 29362 17796 29368 17808
rect 28184 17768 29368 17796
rect 27614 17688 27620 17740
rect 27672 17728 27678 17740
rect 27985 17731 28043 17737
rect 27985 17728 27997 17731
rect 27672 17700 27997 17728
rect 27672 17688 27678 17700
rect 27985 17697 27997 17700
rect 28031 17697 28043 17731
rect 27985 17691 28043 17697
rect 28074 17688 28080 17740
rect 28132 17728 28138 17740
rect 28184 17737 28212 17768
rect 29362 17756 29368 17768
rect 29420 17756 29426 17808
rect 30374 17796 30380 17808
rect 30335 17768 30380 17796
rect 30374 17756 30380 17768
rect 30432 17756 30438 17808
rect 28169 17731 28227 17737
rect 28169 17728 28181 17731
rect 28132 17700 28181 17728
rect 28132 17688 28138 17700
rect 28169 17697 28181 17700
rect 28215 17697 28227 17731
rect 28169 17691 28227 17697
rect 28258 17688 28264 17740
rect 28316 17728 28322 17740
rect 29546 17728 29552 17740
rect 28316 17700 28361 17728
rect 29507 17700 29552 17728
rect 28316 17688 28322 17700
rect 29546 17688 29552 17700
rect 29604 17688 29610 17740
rect 30466 17688 30472 17740
rect 30524 17728 30530 17740
rect 30653 17731 30711 17737
rect 30653 17728 30665 17731
rect 30524 17700 30665 17728
rect 30524 17688 30530 17700
rect 30653 17697 30665 17700
rect 30699 17697 30711 17731
rect 30653 17691 30711 17697
rect 32401 17731 32459 17737
rect 32401 17697 32413 17731
rect 32447 17728 32459 17731
rect 32490 17728 32496 17740
rect 32447 17700 32496 17728
rect 32447 17697 32459 17700
rect 32401 17691 32459 17697
rect 32490 17688 32496 17700
rect 32548 17728 32554 17740
rect 32861 17731 32919 17737
rect 32861 17728 32873 17731
rect 32548 17700 32873 17728
rect 32548 17688 32554 17700
rect 32861 17697 32873 17700
rect 32907 17697 32919 17731
rect 32861 17691 32919 17697
rect 33134 17688 33140 17740
rect 33192 17728 33198 17740
rect 33321 17731 33379 17737
rect 33321 17728 33333 17731
rect 33192 17700 33333 17728
rect 33192 17688 33198 17700
rect 33321 17697 33333 17700
rect 33367 17697 33379 17731
rect 34514 17728 34520 17740
rect 34475 17700 34520 17728
rect 33321 17691 33379 17697
rect 34514 17688 34520 17700
rect 34572 17688 34578 17740
rect 34790 17728 34796 17740
rect 34751 17700 34796 17728
rect 34790 17688 34796 17700
rect 34848 17688 34854 17740
rect 35250 17728 35256 17740
rect 35211 17700 35256 17728
rect 35250 17688 35256 17700
rect 35308 17688 35314 17740
rect 35526 17728 35532 17740
rect 35487 17700 35532 17728
rect 35526 17688 35532 17700
rect 35584 17688 35590 17740
rect 27433 17663 27491 17669
rect 25464 17632 25509 17660
rect 25464 17620 25470 17632
rect 27433 17629 27445 17663
rect 27479 17660 27491 17663
rect 27890 17660 27896 17672
rect 27479 17632 27896 17660
rect 27479 17629 27491 17632
rect 27433 17623 27491 17629
rect 27890 17620 27896 17632
rect 27948 17620 27954 17672
rect 29730 17620 29736 17672
rect 29788 17660 29794 17672
rect 30009 17663 30067 17669
rect 30009 17660 30021 17663
rect 29788 17632 30021 17660
rect 29788 17620 29794 17632
rect 30009 17629 30021 17632
rect 30055 17629 30067 17663
rect 30009 17623 30067 17629
rect 32582 17620 32588 17672
rect 32640 17660 32646 17672
rect 32677 17663 32735 17669
rect 32677 17660 32689 17663
rect 32640 17632 32689 17660
rect 32640 17620 32646 17632
rect 32677 17629 32689 17632
rect 32723 17660 32735 17663
rect 33502 17660 33508 17672
rect 32723 17632 33508 17660
rect 32723 17629 32735 17632
rect 32677 17623 32735 17629
rect 33502 17620 33508 17632
rect 33560 17620 33566 17672
rect 33597 17663 33655 17669
rect 33597 17629 33609 17663
rect 33643 17660 33655 17663
rect 33962 17660 33968 17672
rect 33643 17632 33968 17660
rect 33643 17629 33655 17632
rect 33597 17623 33655 17629
rect 33962 17620 33968 17632
rect 34020 17620 34026 17672
rect 26329 17595 26387 17601
rect 26329 17561 26341 17595
rect 26375 17592 26387 17595
rect 28166 17592 28172 17604
rect 26375 17564 28172 17592
rect 26375 17561 26387 17564
rect 26329 17555 26387 17561
rect 28166 17552 28172 17564
rect 28224 17592 28230 17604
rect 28224 17564 28488 17592
rect 28224 17552 28230 17564
rect 25958 17524 25964 17536
rect 24044 17496 24992 17524
rect 25919 17496 25964 17524
rect 20165 17487 20223 17493
rect 25958 17484 25964 17496
rect 26016 17484 26022 17536
rect 27062 17524 27068 17536
rect 27023 17496 27068 17524
rect 27062 17484 27068 17496
rect 27120 17484 27126 17536
rect 27706 17524 27712 17536
rect 27667 17496 27712 17524
rect 27706 17484 27712 17496
rect 27764 17484 27770 17536
rect 28460 17533 28488 17564
rect 28445 17527 28503 17533
rect 28445 17493 28457 17527
rect 28491 17493 28503 17527
rect 29362 17524 29368 17536
rect 29323 17496 29368 17524
rect 28445 17487 28503 17493
rect 29362 17484 29368 17496
rect 29420 17484 29426 17536
rect 29733 17527 29791 17533
rect 29733 17493 29745 17527
rect 29779 17524 29791 17527
rect 29914 17524 29920 17536
rect 29779 17496 29920 17524
rect 29779 17493 29791 17496
rect 29733 17487 29791 17493
rect 29914 17484 29920 17496
rect 29972 17484 29978 17536
rect 31202 17524 31208 17536
rect 31163 17496 31208 17524
rect 31202 17484 31208 17496
rect 31260 17484 31266 17536
rect 31573 17527 31631 17533
rect 31573 17493 31585 17527
rect 31619 17524 31631 17527
rect 31662 17524 31668 17536
rect 31619 17496 31668 17524
rect 31619 17493 31631 17496
rect 31573 17487 31631 17493
rect 31662 17484 31668 17496
rect 31720 17484 31726 17536
rect 1104 17434 38548 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 38548 17434
rect 1104 17360 38548 17382
rect 2041 17323 2099 17329
rect 2041 17289 2053 17323
rect 2087 17320 2099 17323
rect 3234 17320 3240 17332
rect 2087 17292 3240 17320
rect 2087 17289 2099 17292
rect 2041 17283 2099 17289
rect 3234 17280 3240 17292
rect 3292 17280 3298 17332
rect 3510 17320 3516 17332
rect 3471 17292 3516 17320
rect 3510 17280 3516 17292
rect 3568 17280 3574 17332
rect 4433 17323 4491 17329
rect 4433 17289 4445 17323
rect 4479 17320 4491 17323
rect 5534 17320 5540 17332
rect 4479 17292 5540 17320
rect 4479 17289 4491 17292
rect 4433 17283 4491 17289
rect 5534 17280 5540 17292
rect 5592 17280 5598 17332
rect 5629 17323 5687 17329
rect 5629 17289 5641 17323
rect 5675 17320 5687 17323
rect 5718 17320 5724 17332
rect 5675 17292 5724 17320
rect 5675 17289 5687 17292
rect 5629 17283 5687 17289
rect 5718 17280 5724 17292
rect 5776 17280 5782 17332
rect 8113 17323 8171 17329
rect 8113 17289 8125 17323
rect 8159 17320 8171 17323
rect 8386 17320 8392 17332
rect 8159 17292 8392 17320
rect 8159 17289 8171 17292
rect 8113 17283 8171 17289
rect 8386 17280 8392 17292
rect 8444 17280 8450 17332
rect 8662 17280 8668 17332
rect 8720 17320 8726 17332
rect 8757 17323 8815 17329
rect 8757 17320 8769 17323
rect 8720 17292 8769 17320
rect 8720 17280 8726 17292
rect 8757 17289 8769 17292
rect 8803 17289 8815 17323
rect 8757 17283 8815 17289
rect 9125 17323 9183 17329
rect 9125 17289 9137 17323
rect 9171 17320 9183 17323
rect 9490 17320 9496 17332
rect 9171 17292 9496 17320
rect 9171 17289 9183 17292
rect 9125 17283 9183 17289
rect 5169 17255 5227 17261
rect 5169 17221 5181 17255
rect 5215 17252 5227 17255
rect 5442 17252 5448 17264
rect 5215 17224 5448 17252
rect 5215 17221 5227 17224
rect 5169 17215 5227 17221
rect 5442 17212 5448 17224
rect 5500 17212 5506 17264
rect 5994 17212 6000 17264
rect 6052 17252 6058 17264
rect 6730 17252 6736 17264
rect 6052 17224 6736 17252
rect 6052 17212 6058 17224
rect 6730 17212 6736 17224
rect 6788 17212 6794 17264
rect 2406 17184 2412 17196
rect 2367 17156 2412 17184
rect 2406 17144 2412 17156
rect 2464 17144 2470 17196
rect 5353 17187 5411 17193
rect 5353 17153 5365 17187
rect 5399 17184 5411 17187
rect 6270 17184 6276 17196
rect 5399 17156 6276 17184
rect 5399 17153 5411 17156
rect 5353 17147 5411 17153
rect 6270 17144 6276 17156
rect 6328 17144 6334 17196
rect 7009 17187 7067 17193
rect 7009 17153 7021 17187
rect 7055 17184 7067 17187
rect 7098 17184 7104 17196
rect 7055 17156 7104 17184
rect 7055 17153 7067 17156
rect 7009 17147 7067 17153
rect 7098 17144 7104 17156
rect 7156 17144 7162 17196
rect 9140 17184 9168 17283
rect 9490 17280 9496 17292
rect 9548 17280 9554 17332
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 12713 17323 12771 17329
rect 12713 17320 12725 17323
rect 12492 17292 12725 17320
rect 12492 17280 12498 17292
rect 12713 17289 12725 17292
rect 12759 17289 12771 17323
rect 14182 17320 14188 17332
rect 14143 17292 14188 17320
rect 12713 17283 12771 17289
rect 14182 17280 14188 17292
rect 14240 17280 14246 17332
rect 14274 17280 14280 17332
rect 14332 17320 14338 17332
rect 15289 17323 15347 17329
rect 15289 17320 15301 17323
rect 14332 17292 15301 17320
rect 14332 17280 14338 17292
rect 15289 17289 15301 17292
rect 15335 17289 15347 17323
rect 15289 17283 15347 17289
rect 16574 17280 16580 17332
rect 16632 17320 16638 17332
rect 16669 17323 16727 17329
rect 16669 17320 16681 17323
rect 16632 17292 16681 17320
rect 16632 17280 16638 17292
rect 16669 17289 16681 17292
rect 16715 17289 16727 17323
rect 17586 17320 17592 17332
rect 17547 17292 17592 17320
rect 16669 17283 16727 17289
rect 17586 17280 17592 17292
rect 17644 17280 17650 17332
rect 17770 17280 17776 17332
rect 17828 17320 17834 17332
rect 18233 17323 18291 17329
rect 18233 17320 18245 17323
rect 17828 17292 18245 17320
rect 17828 17280 17834 17292
rect 18233 17289 18245 17292
rect 18279 17289 18291 17323
rect 18233 17283 18291 17289
rect 18782 17280 18788 17332
rect 18840 17320 18846 17332
rect 18877 17323 18935 17329
rect 18877 17320 18889 17323
rect 18840 17292 18889 17320
rect 18840 17280 18846 17292
rect 18877 17289 18889 17292
rect 18923 17289 18935 17323
rect 18877 17283 18935 17289
rect 19334 17280 19340 17332
rect 19392 17320 19398 17332
rect 20257 17323 20315 17329
rect 20257 17320 20269 17323
rect 19392 17292 20269 17320
rect 19392 17280 19398 17292
rect 20257 17289 20269 17292
rect 20303 17289 20315 17323
rect 22922 17320 22928 17332
rect 22883 17292 22928 17320
rect 20257 17283 20315 17289
rect 22922 17280 22928 17292
rect 22980 17280 22986 17332
rect 25866 17280 25872 17332
rect 25924 17320 25930 17332
rect 26145 17323 26203 17329
rect 26145 17320 26157 17323
rect 25924 17292 26157 17320
rect 25924 17280 25930 17292
rect 26145 17289 26157 17292
rect 26191 17289 26203 17323
rect 26145 17283 26203 17289
rect 26513 17323 26571 17329
rect 26513 17289 26525 17323
rect 26559 17320 26571 17323
rect 27430 17320 27436 17332
rect 26559 17292 27436 17320
rect 26559 17289 26571 17292
rect 26513 17283 26571 17289
rect 27430 17280 27436 17292
rect 27488 17280 27494 17332
rect 28258 17280 28264 17332
rect 28316 17320 28322 17332
rect 28629 17323 28687 17329
rect 28629 17320 28641 17323
rect 28316 17292 28641 17320
rect 28316 17280 28322 17292
rect 28629 17289 28641 17292
rect 28675 17289 28687 17323
rect 28629 17283 28687 17289
rect 29546 17280 29552 17332
rect 29604 17320 29610 17332
rect 30285 17323 30343 17329
rect 30285 17320 30297 17323
rect 29604 17292 30297 17320
rect 29604 17280 29610 17292
rect 30285 17289 30297 17292
rect 30331 17289 30343 17323
rect 30285 17283 30343 17289
rect 30466 17280 30472 17332
rect 30524 17320 30530 17332
rect 30653 17323 30711 17329
rect 30653 17320 30665 17323
rect 30524 17292 30665 17320
rect 30524 17280 30530 17292
rect 30653 17289 30665 17292
rect 30699 17289 30711 17323
rect 32582 17320 32588 17332
rect 32543 17292 32588 17320
rect 30653 17283 30711 17289
rect 32582 17280 32588 17292
rect 32640 17280 32646 17332
rect 34330 17280 34336 17332
rect 34388 17320 34394 17332
rect 34514 17320 34520 17332
rect 34388 17292 34520 17320
rect 34388 17280 34394 17292
rect 34514 17280 34520 17292
rect 34572 17320 34578 17332
rect 35069 17323 35127 17329
rect 35069 17320 35081 17323
rect 34572 17292 35081 17320
rect 34572 17280 34578 17292
rect 35069 17289 35081 17292
rect 35115 17289 35127 17323
rect 35069 17283 35127 17289
rect 11698 17212 11704 17264
rect 11756 17252 11762 17264
rect 12250 17252 12256 17264
rect 11756 17224 12256 17252
rect 11756 17212 11762 17224
rect 12250 17212 12256 17224
rect 12308 17252 12314 17264
rect 14734 17252 14740 17264
rect 12308 17224 14740 17252
rect 12308 17212 12314 17224
rect 14734 17212 14740 17224
rect 14792 17212 14798 17264
rect 16301 17255 16359 17261
rect 16301 17221 16313 17255
rect 16347 17252 16359 17255
rect 17788 17252 17816 17280
rect 16347 17224 17816 17252
rect 16347 17221 16359 17224
rect 16301 17215 16359 17221
rect 8588 17156 9168 17184
rect 1854 17076 1860 17128
rect 1912 17116 1918 17128
rect 2133 17119 2191 17125
rect 2133 17116 2145 17119
rect 1912 17088 2145 17116
rect 1912 17076 1918 17088
rect 2133 17085 2145 17088
rect 2179 17085 2191 17119
rect 2498 17116 2504 17128
rect 2133 17079 2191 17085
rect 2240 17088 2504 17116
rect 1673 17051 1731 17057
rect 1673 17017 1685 17051
rect 1719 17048 1731 17051
rect 2240 17048 2268 17088
rect 2498 17076 2504 17088
rect 2556 17076 2562 17128
rect 5442 17076 5448 17128
rect 5500 17116 5506 17128
rect 7193 17119 7251 17125
rect 5500 17088 5545 17116
rect 5500 17076 5506 17088
rect 7193 17085 7205 17119
rect 7239 17116 7251 17119
rect 7466 17116 7472 17128
rect 7239 17088 7472 17116
rect 7239 17085 7251 17088
rect 7193 17079 7251 17085
rect 7466 17076 7472 17088
rect 7524 17076 7530 17128
rect 8588 17125 8616 17156
rect 9398 17144 9404 17196
rect 9456 17184 9462 17196
rect 9493 17187 9551 17193
rect 9493 17184 9505 17187
rect 9456 17156 9505 17184
rect 9456 17144 9462 17156
rect 9493 17153 9505 17156
rect 9539 17153 9551 17187
rect 9493 17147 9551 17153
rect 11238 17144 11244 17196
rect 11296 17184 11302 17196
rect 13354 17184 13360 17196
rect 11296 17156 13360 17184
rect 11296 17144 11302 17156
rect 13354 17144 13360 17156
rect 13412 17144 13418 17196
rect 14366 17144 14372 17196
rect 14424 17184 14430 17196
rect 14642 17184 14648 17196
rect 14424 17156 14648 17184
rect 14424 17144 14430 17156
rect 14642 17144 14648 17156
rect 14700 17144 14706 17196
rect 8573 17119 8631 17125
rect 8573 17085 8585 17119
rect 8619 17085 8631 17119
rect 8573 17079 8631 17085
rect 8938 17076 8944 17128
rect 8996 17116 9002 17128
rect 9677 17119 9735 17125
rect 9677 17116 9689 17119
rect 8996 17088 9689 17116
rect 8996 17076 9002 17088
rect 9677 17085 9689 17088
rect 9723 17085 9735 17119
rect 10226 17116 10232 17128
rect 10187 17088 10232 17116
rect 9677 17079 9735 17085
rect 10226 17076 10232 17088
rect 10284 17076 10290 17128
rect 10502 17116 10508 17128
rect 10463 17088 10508 17116
rect 10502 17076 10508 17088
rect 10560 17076 10566 17128
rect 12434 17116 12440 17128
rect 12395 17088 12440 17116
rect 12434 17076 12440 17088
rect 12492 17076 12498 17128
rect 12570 17119 12628 17125
rect 12570 17085 12582 17119
rect 12616 17116 12628 17119
rect 14001 17119 14059 17125
rect 12616 17088 12756 17116
rect 12616 17085 12628 17088
rect 12570 17079 12628 17085
rect 1719 17020 2268 17048
rect 4801 17051 4859 17057
rect 1719 17017 1731 17020
rect 1673 17011 1731 17017
rect 4801 17017 4813 17051
rect 4847 17048 4859 17051
rect 5460 17048 5488 17076
rect 7282 17048 7288 17060
rect 4847 17020 5488 17048
rect 7243 17020 7288 17048
rect 4847 17017 4859 17020
rect 4801 17011 4859 17017
rect 7282 17008 7288 17020
rect 7340 17008 7346 17060
rect 7377 17051 7435 17057
rect 7377 17017 7389 17051
rect 7423 17048 7435 17051
rect 7650 17048 7656 17060
rect 7423 17020 7656 17048
rect 7423 17017 7435 17020
rect 7377 17011 7435 17017
rect 7650 17008 7656 17020
rect 7708 17008 7714 17060
rect 7745 17051 7803 17057
rect 7745 17017 7757 17051
rect 7791 17048 7803 17051
rect 8202 17048 8208 17060
rect 7791 17020 8208 17048
rect 7791 17017 7803 17020
rect 7745 17011 7803 17017
rect 8202 17008 8208 17020
rect 8260 17008 8266 17060
rect 8481 17051 8539 17057
rect 8481 17017 8493 17051
rect 8527 17048 8539 17051
rect 10520 17048 10548 17076
rect 8527 17020 10548 17048
rect 8527 17017 8539 17020
rect 8481 17011 8539 17017
rect 11974 17008 11980 17060
rect 12032 17048 12038 17060
rect 12253 17051 12311 17057
rect 12253 17048 12265 17051
rect 12032 17020 12265 17048
rect 12032 17008 12038 17020
rect 12253 17017 12265 17020
rect 12299 17048 12311 17051
rect 12728 17048 12756 17088
rect 14001 17085 14013 17119
rect 14047 17116 14059 17119
rect 14277 17119 14335 17125
rect 14277 17116 14289 17119
rect 14047 17088 14289 17116
rect 14047 17085 14059 17088
rect 14001 17079 14059 17085
rect 14277 17085 14289 17088
rect 14323 17085 14335 17119
rect 14277 17079 14335 17085
rect 14550 17076 14556 17128
rect 14608 17116 14614 17128
rect 14829 17119 14887 17125
rect 14829 17116 14841 17119
rect 14608 17088 14841 17116
rect 14608 17076 14614 17088
rect 14829 17085 14841 17088
rect 14875 17085 14887 17119
rect 15010 17116 15016 17128
rect 14971 17088 15016 17116
rect 14829 17079 14887 17085
rect 15010 17076 15016 17088
rect 15068 17076 15074 17128
rect 15105 17119 15163 17125
rect 15105 17085 15117 17119
rect 15151 17116 15163 17119
rect 15286 17116 15292 17128
rect 15151 17088 15292 17116
rect 15151 17085 15163 17088
rect 15105 17079 15163 17085
rect 15286 17076 15292 17088
rect 15344 17116 15350 17128
rect 15657 17119 15715 17125
rect 15657 17116 15669 17119
rect 15344 17088 15669 17116
rect 15344 17076 15350 17088
rect 15657 17085 15669 17088
rect 15703 17085 15715 17119
rect 15657 17079 15715 17085
rect 13354 17048 13360 17060
rect 12299 17020 12756 17048
rect 13267 17020 13360 17048
rect 12299 17017 12311 17020
rect 12253 17011 12311 17017
rect 13354 17008 13360 17020
rect 13412 17048 13418 17060
rect 16316 17048 16344 17215
rect 18046 17212 18052 17264
rect 18104 17252 18110 17264
rect 18414 17252 18420 17264
rect 18104 17224 18420 17252
rect 18104 17212 18110 17224
rect 18414 17212 18420 17224
rect 18472 17212 18478 17264
rect 19245 17255 19303 17261
rect 19245 17221 19257 17255
rect 19291 17221 19303 17255
rect 19245 17215 19303 17221
rect 16393 17187 16451 17193
rect 16393 17153 16405 17187
rect 16439 17184 16451 17187
rect 16439 17156 16620 17184
rect 16439 17153 16451 17156
rect 16393 17147 16451 17153
rect 16485 17119 16543 17125
rect 16485 17085 16497 17119
rect 16531 17085 16543 17119
rect 16485 17079 16543 17085
rect 13412 17020 16344 17048
rect 13412 17008 13418 17020
rect 2038 16940 2044 16992
rect 2096 16980 2102 16992
rect 3510 16980 3516 16992
rect 2096 16952 3516 16980
rect 2096 16940 2102 16952
rect 3510 16940 3516 16952
rect 3568 16940 3574 16992
rect 6638 16980 6644 16992
rect 6599 16952 6644 16980
rect 6638 16940 6644 16952
rect 6696 16940 6702 16992
rect 9766 16980 9772 16992
rect 9727 16952 9772 16980
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 11330 16980 11336 16992
rect 11291 16952 11336 16980
rect 11330 16940 11336 16952
rect 11388 16940 11394 16992
rect 11606 16980 11612 16992
rect 11567 16952 11612 16980
rect 11606 16940 11612 16952
rect 11664 16940 11670 16992
rect 13630 16980 13636 16992
rect 13591 16952 13636 16980
rect 13630 16940 13636 16952
rect 13688 16940 13694 16992
rect 14277 16983 14335 16989
rect 14277 16949 14289 16983
rect 14323 16980 14335 16983
rect 14553 16983 14611 16989
rect 14553 16980 14565 16983
rect 14323 16952 14565 16980
rect 14323 16949 14335 16952
rect 14277 16943 14335 16949
rect 14553 16949 14565 16952
rect 14599 16980 14611 16983
rect 14918 16980 14924 16992
rect 14599 16952 14924 16980
rect 14599 16949 14611 16952
rect 14553 16943 14611 16949
rect 14918 16940 14924 16952
rect 14976 16940 14982 16992
rect 15657 16983 15715 16989
rect 15657 16949 15669 16983
rect 15703 16980 15715 16983
rect 15933 16983 15991 16989
rect 15933 16980 15945 16983
rect 15703 16952 15945 16980
rect 15703 16949 15715 16952
rect 15657 16943 15715 16949
rect 15933 16949 15945 16952
rect 15979 16980 15991 16983
rect 16500 16980 16528 17079
rect 16592 17048 16620 17156
rect 16666 17144 16672 17196
rect 16724 17184 16730 17196
rect 19260 17184 19288 17215
rect 19426 17212 19432 17264
rect 19484 17252 19490 17264
rect 19886 17252 19892 17264
rect 19484 17224 19892 17252
rect 19484 17212 19490 17224
rect 19886 17212 19892 17224
rect 19944 17212 19950 17264
rect 22002 17252 22008 17264
rect 21928 17224 22008 17252
rect 16724 17156 19288 17184
rect 16724 17144 16730 17156
rect 16850 17076 16856 17128
rect 16908 17116 16914 17128
rect 17218 17116 17224 17128
rect 16908 17088 17224 17116
rect 16908 17076 16914 17088
rect 17218 17076 17224 17088
rect 17276 17076 17282 17128
rect 18049 17119 18107 17125
rect 18049 17085 18061 17119
rect 18095 17116 18107 17119
rect 18095 17088 18368 17116
rect 18095 17085 18107 17088
rect 18049 17079 18107 17085
rect 17310 17048 17316 17060
rect 16592 17020 17316 17048
rect 17310 17008 17316 17020
rect 17368 17048 17374 17060
rect 17494 17048 17500 17060
rect 17368 17020 17500 17048
rect 17368 17008 17374 17020
rect 17494 17008 17500 17020
rect 17552 17008 17558 17060
rect 18340 16992 18368 17088
rect 18690 17076 18696 17128
rect 18748 17116 18754 17128
rect 19061 17119 19119 17125
rect 19061 17116 19073 17119
rect 18748 17088 19073 17116
rect 18748 17076 18754 17088
rect 19061 17085 19073 17088
rect 19107 17085 19119 17119
rect 19061 17079 19119 17085
rect 19076 17048 19104 17079
rect 19334 17076 19340 17128
rect 19392 17116 19398 17128
rect 20073 17119 20131 17125
rect 20073 17116 20085 17119
rect 19392 17088 20085 17116
rect 19392 17076 19398 17088
rect 20073 17085 20085 17088
rect 20119 17116 20131 17119
rect 20533 17119 20591 17125
rect 20533 17116 20545 17119
rect 20119 17088 20545 17116
rect 20119 17085 20131 17088
rect 20073 17079 20131 17085
rect 20533 17085 20545 17088
rect 20579 17085 20591 17119
rect 20533 17079 20591 17085
rect 21358 17076 21364 17128
rect 21416 17116 21422 17128
rect 21928 17125 21956 17224
rect 22002 17212 22008 17224
rect 22060 17212 22066 17264
rect 22186 17212 22192 17264
rect 22244 17252 22250 17264
rect 26050 17261 26056 17264
rect 22281 17255 22339 17261
rect 22281 17252 22293 17255
rect 22244 17224 22293 17252
rect 22244 17212 22250 17224
rect 22281 17221 22293 17224
rect 22327 17221 22339 17255
rect 22281 17215 22339 17221
rect 25777 17255 25835 17261
rect 25777 17221 25789 17255
rect 25823 17252 25835 17255
rect 26007 17255 26056 17261
rect 26007 17252 26019 17255
rect 25823 17224 26019 17252
rect 25823 17221 25835 17224
rect 25777 17215 25835 17221
rect 26007 17221 26019 17224
rect 26053 17221 26056 17255
rect 26007 17215 26056 17221
rect 26050 17212 26056 17215
rect 26108 17252 26114 17264
rect 31294 17252 31300 17264
rect 26108 17224 26155 17252
rect 31128 17224 31300 17252
rect 26108 17212 26114 17224
rect 26237 17187 26295 17193
rect 26237 17184 26249 17187
rect 25332 17156 26249 17184
rect 21453 17119 21511 17125
rect 21453 17116 21465 17119
rect 21416 17088 21465 17116
rect 21416 17076 21422 17088
rect 21453 17085 21465 17088
rect 21499 17085 21511 17119
rect 21453 17079 21511 17085
rect 21913 17119 21971 17125
rect 21913 17085 21925 17119
rect 21959 17085 21971 17119
rect 21913 17079 21971 17085
rect 22281 17119 22339 17125
rect 22281 17085 22293 17119
rect 22327 17085 22339 17119
rect 22281 17079 22339 17085
rect 19521 17051 19579 17057
rect 19521 17048 19533 17051
rect 19076 17020 19533 17048
rect 19521 17017 19533 17020
rect 19567 17017 19579 17051
rect 19521 17011 19579 17017
rect 20714 17008 20720 17060
rect 20772 17048 20778 17060
rect 20993 17051 21051 17057
rect 20993 17048 21005 17051
rect 20772 17020 21005 17048
rect 20772 17008 20778 17020
rect 20993 17017 21005 17020
rect 21039 17048 21051 17051
rect 22296 17048 22324 17079
rect 23474 17076 23480 17128
rect 23532 17116 23538 17128
rect 24026 17116 24032 17128
rect 23532 17088 24032 17116
rect 23532 17076 23538 17088
rect 24026 17076 24032 17088
rect 24084 17116 24090 17128
rect 24213 17119 24271 17125
rect 24213 17116 24225 17119
rect 24084 17088 24225 17116
rect 24084 17076 24090 17088
rect 24213 17085 24225 17088
rect 24259 17085 24271 17119
rect 24213 17079 24271 17085
rect 22922 17048 22928 17060
rect 21039 17020 22928 17048
rect 21039 17017 21051 17020
rect 20993 17011 21051 17017
rect 22922 17008 22928 17020
rect 22980 17008 22986 17060
rect 17218 16980 17224 16992
rect 15979 16952 17224 16980
rect 15979 16949 15991 16952
rect 15933 16943 15991 16949
rect 17218 16940 17224 16952
rect 17276 16940 17282 16992
rect 18322 16940 18328 16992
rect 18380 16980 18386 16992
rect 18509 16983 18567 16989
rect 18509 16980 18521 16983
rect 18380 16952 18521 16980
rect 18380 16940 18386 16952
rect 18509 16949 18521 16952
rect 18555 16949 18567 16983
rect 21358 16980 21364 16992
rect 21271 16952 21364 16980
rect 18509 16943 18567 16949
rect 21358 16940 21364 16952
rect 21416 16980 21422 16992
rect 23198 16980 23204 16992
rect 21416 16952 23204 16980
rect 21416 16940 21422 16952
rect 23198 16940 23204 16952
rect 23256 16940 23262 16992
rect 24118 16980 24124 16992
rect 24079 16952 24124 16980
rect 24118 16940 24124 16952
rect 24176 16940 24182 16992
rect 24302 16940 24308 16992
rect 24360 16980 24366 16992
rect 24397 16983 24455 16989
rect 24397 16980 24409 16983
rect 24360 16952 24409 16980
rect 24360 16940 24366 16952
rect 24397 16949 24409 16952
rect 24443 16949 24455 16983
rect 24397 16943 24455 16949
rect 24857 16983 24915 16989
rect 24857 16949 24869 16983
rect 24903 16980 24915 16983
rect 24946 16980 24952 16992
rect 24903 16952 24952 16980
rect 24903 16949 24915 16952
rect 24857 16943 24915 16949
rect 24946 16940 24952 16952
rect 25004 16980 25010 16992
rect 25332 16989 25360 17156
rect 26237 17153 26249 17156
rect 26283 17184 26295 17187
rect 26786 17184 26792 17196
rect 26283 17156 26792 17184
rect 26283 17153 26295 17156
rect 26237 17147 26295 17153
rect 26786 17144 26792 17156
rect 26844 17144 26850 17196
rect 28353 17187 28411 17193
rect 28353 17153 28365 17187
rect 28399 17184 28411 17187
rect 29086 17184 29092 17196
rect 28399 17156 29092 17184
rect 28399 17153 28411 17156
rect 28353 17147 28411 17153
rect 29086 17144 29092 17156
rect 29144 17144 29150 17196
rect 30006 17184 30012 17196
rect 29967 17156 30012 17184
rect 30006 17144 30012 17156
rect 30064 17144 30070 17196
rect 31128 17193 31156 17224
rect 31294 17212 31300 17224
rect 31352 17212 31358 17264
rect 31113 17187 31171 17193
rect 31113 17153 31125 17187
rect 31159 17153 31171 17187
rect 31113 17147 31171 17153
rect 31202 17144 31208 17196
rect 31260 17184 31266 17196
rect 31260 17156 32168 17184
rect 31260 17144 31266 17156
rect 25869 17119 25927 17125
rect 25869 17085 25881 17119
rect 25915 17116 25927 17119
rect 25958 17116 25964 17128
rect 25915 17088 25964 17116
rect 25915 17085 25927 17088
rect 25869 17079 25927 17085
rect 25958 17076 25964 17088
rect 26016 17076 26022 17128
rect 27890 17116 27896 17128
rect 27803 17088 27896 17116
rect 27890 17076 27896 17088
rect 27948 17116 27954 17128
rect 29362 17116 29368 17128
rect 27948 17088 29368 17116
rect 27948 17076 27954 17088
rect 29362 17076 29368 17088
rect 29420 17116 29426 17128
rect 29549 17119 29607 17125
rect 29549 17116 29561 17119
rect 29420 17088 29561 17116
rect 29420 17076 29426 17088
rect 29549 17085 29561 17088
rect 29595 17085 29607 17119
rect 31662 17116 31668 17128
rect 31623 17088 31668 17116
rect 29549 17079 29607 17085
rect 31662 17076 31668 17088
rect 31720 17076 31726 17128
rect 32140 17125 32168 17156
rect 33318 17144 33324 17196
rect 33376 17184 33382 17196
rect 33965 17187 34023 17193
rect 33965 17184 33977 17187
rect 33376 17156 33977 17184
rect 33376 17144 33382 17156
rect 33965 17153 33977 17156
rect 34011 17184 34023 17187
rect 34609 17187 34667 17193
rect 34609 17184 34621 17187
rect 34011 17156 34621 17184
rect 34011 17153 34023 17156
rect 33965 17147 34023 17153
rect 34609 17153 34621 17156
rect 34655 17153 34667 17187
rect 34609 17147 34667 17153
rect 31941 17119 31999 17125
rect 31941 17085 31953 17119
rect 31987 17085 31999 17119
rect 31941 17079 31999 17085
rect 32125 17119 32183 17125
rect 32125 17085 32137 17119
rect 32171 17116 32183 17119
rect 32490 17116 32496 17128
rect 32171 17088 32496 17116
rect 32171 17085 32183 17088
rect 32125 17079 32183 17085
rect 27062 17008 27068 17060
rect 27120 17048 27126 17060
rect 27614 17048 27620 17060
rect 27120 17020 27620 17048
rect 27120 17008 27126 17020
rect 27614 17008 27620 17020
rect 27672 17008 27678 17060
rect 27706 17008 27712 17060
rect 27764 17048 27770 17060
rect 27985 17051 28043 17057
rect 27985 17048 27997 17051
rect 27764 17020 27997 17048
rect 27764 17008 27770 17020
rect 27985 17017 27997 17020
rect 28031 17048 28043 17051
rect 28534 17048 28540 17060
rect 28031 17020 28540 17048
rect 28031 17017 28043 17020
rect 27985 17011 28043 17017
rect 28534 17008 28540 17020
rect 28592 17008 28598 17060
rect 29089 17051 29147 17057
rect 29089 17017 29101 17051
rect 29135 17048 29147 17051
rect 29270 17048 29276 17060
rect 29135 17020 29276 17048
rect 29135 17017 29147 17020
rect 29089 17011 29147 17017
rect 29270 17008 29276 17020
rect 29328 17008 29334 17060
rect 29641 17051 29699 17057
rect 29641 17017 29653 17051
rect 29687 17048 29699 17051
rect 29730 17048 29736 17060
rect 29687 17020 29736 17048
rect 29687 17017 29699 17020
rect 29641 17011 29699 17017
rect 29730 17008 29736 17020
rect 29788 17008 29794 17060
rect 31294 17008 31300 17060
rect 31352 17048 31358 17060
rect 31754 17048 31760 17060
rect 31352 17020 31760 17048
rect 31352 17008 31358 17020
rect 31754 17008 31760 17020
rect 31812 17048 31818 17060
rect 31956 17048 31984 17079
rect 32490 17076 32496 17088
rect 32548 17076 32554 17128
rect 32858 17076 32864 17128
rect 32916 17116 32922 17128
rect 33505 17119 33563 17125
rect 33505 17116 33517 17119
rect 32916 17088 33517 17116
rect 32916 17076 32922 17088
rect 33505 17085 33517 17088
rect 33551 17085 33563 17119
rect 33778 17116 33784 17128
rect 33739 17088 33784 17116
rect 33505 17079 33563 17085
rect 33778 17076 33784 17088
rect 33836 17076 33842 17128
rect 31812 17020 31984 17048
rect 32953 17051 33011 17057
rect 31812 17008 31818 17020
rect 32953 17017 32965 17051
rect 32999 17048 33011 17051
rect 33594 17048 33600 17060
rect 32999 17020 33600 17048
rect 32999 17017 33011 17020
rect 32953 17011 33011 17017
rect 33594 17008 33600 17020
rect 33652 17008 33658 17060
rect 33796 17048 33824 17076
rect 34241 17051 34299 17057
rect 34241 17048 34253 17051
rect 33796 17020 34253 17048
rect 34241 17017 34253 17020
rect 34287 17017 34299 17051
rect 34241 17011 34299 17017
rect 25317 16983 25375 16989
rect 25317 16980 25329 16983
rect 25004 16952 25329 16980
rect 25004 16940 25010 16952
rect 25317 16949 25329 16952
rect 25363 16949 25375 16983
rect 25317 16943 25375 16949
rect 26510 16940 26516 16992
rect 26568 16980 26574 16992
rect 26881 16983 26939 16989
rect 26881 16980 26893 16983
rect 26568 16952 26893 16980
rect 26568 16940 26574 16952
rect 26881 16949 26893 16952
rect 26927 16949 26939 16983
rect 26881 16943 26939 16949
rect 27525 16983 27583 16989
rect 27525 16949 27537 16983
rect 27571 16980 27583 16983
rect 27801 16983 27859 16989
rect 27801 16980 27813 16983
rect 27571 16952 27813 16980
rect 27571 16949 27583 16952
rect 27525 16943 27583 16949
rect 27801 16949 27813 16952
rect 27847 16980 27859 16983
rect 28074 16980 28080 16992
rect 27847 16952 28080 16980
rect 27847 16949 27859 16952
rect 27801 16943 27859 16949
rect 28074 16940 28080 16952
rect 28132 16940 28138 16992
rect 29454 16980 29460 16992
rect 29415 16952 29460 16980
rect 29454 16940 29460 16952
rect 29512 16940 29518 16992
rect 1104 16890 38548 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 38548 16890
rect 1104 16816 38548 16838
rect 1394 16736 1400 16788
rect 1452 16776 1458 16788
rect 1673 16779 1731 16785
rect 1673 16776 1685 16779
rect 1452 16748 1685 16776
rect 1452 16736 1458 16748
rect 1673 16745 1685 16748
rect 1719 16776 1731 16779
rect 1854 16776 1860 16788
rect 1719 16748 1860 16776
rect 1719 16745 1731 16748
rect 1673 16739 1731 16745
rect 1854 16736 1860 16748
rect 1912 16736 1918 16788
rect 2038 16776 2044 16788
rect 1999 16748 2044 16776
rect 2038 16736 2044 16748
rect 2096 16736 2102 16788
rect 2406 16776 2412 16788
rect 2367 16748 2412 16776
rect 2406 16736 2412 16748
rect 2464 16776 2470 16788
rect 2685 16779 2743 16785
rect 2685 16776 2697 16779
rect 2464 16748 2697 16776
rect 2464 16736 2470 16748
rect 2685 16745 2697 16748
rect 2731 16745 2743 16779
rect 3142 16776 3148 16788
rect 3103 16748 3148 16776
rect 2685 16739 2743 16745
rect 3142 16736 3148 16748
rect 3200 16736 3206 16788
rect 3513 16779 3571 16785
rect 3513 16745 3525 16779
rect 3559 16776 3571 16779
rect 3970 16776 3976 16788
rect 3559 16748 3976 16776
rect 3559 16745 3571 16748
rect 3513 16739 3571 16745
rect 3970 16736 3976 16748
rect 4028 16736 4034 16788
rect 4433 16779 4491 16785
rect 4433 16745 4445 16779
rect 4479 16776 4491 16779
rect 5350 16776 5356 16788
rect 4479 16748 5356 16776
rect 4479 16745 4491 16748
rect 4433 16739 4491 16745
rect 5350 16736 5356 16748
rect 5408 16736 5414 16788
rect 6825 16779 6883 16785
rect 6825 16745 6837 16779
rect 6871 16776 6883 16779
rect 7098 16776 7104 16788
rect 6871 16748 7104 16776
rect 6871 16745 6883 16748
rect 6825 16739 6883 16745
rect 7098 16736 7104 16748
rect 7156 16736 7162 16788
rect 9306 16776 9312 16788
rect 7484 16748 9312 16776
rect 7484 16720 7512 16748
rect 9306 16736 9312 16748
rect 9364 16776 9370 16788
rect 9401 16779 9459 16785
rect 9401 16776 9413 16779
rect 9364 16748 9413 16776
rect 9364 16736 9370 16748
rect 9401 16745 9413 16748
rect 9447 16745 9459 16779
rect 9401 16739 9459 16745
rect 4062 16668 4068 16720
rect 4120 16708 4126 16720
rect 6181 16711 6239 16717
rect 4120 16680 5212 16708
rect 4120 16668 4126 16680
rect 5184 16652 5212 16680
rect 6181 16677 6193 16711
rect 6227 16708 6239 16711
rect 6549 16711 6607 16717
rect 6549 16708 6561 16711
rect 6227 16680 6561 16708
rect 6227 16677 6239 16680
rect 6181 16671 6239 16677
rect 6549 16677 6561 16680
rect 6595 16708 6607 16711
rect 7282 16708 7288 16720
rect 6595 16680 7288 16708
rect 6595 16677 6607 16680
rect 6549 16671 6607 16677
rect 7282 16668 7288 16680
rect 7340 16668 7346 16720
rect 7466 16708 7472 16720
rect 7427 16680 7472 16708
rect 7466 16668 7472 16680
rect 7524 16668 7530 16720
rect 7745 16711 7803 16717
rect 7745 16677 7757 16711
rect 7791 16708 7803 16711
rect 7834 16708 7840 16720
rect 7791 16680 7840 16708
rect 7791 16677 7803 16680
rect 7745 16671 7803 16677
rect 3881 16643 3939 16649
rect 3881 16609 3893 16643
rect 3927 16640 3939 16643
rect 4890 16640 4896 16652
rect 3927 16612 4896 16640
rect 3927 16609 3939 16612
rect 3881 16603 3939 16609
rect 4890 16600 4896 16612
rect 4948 16600 4954 16652
rect 4985 16643 5043 16649
rect 4985 16609 4997 16643
rect 5031 16609 5043 16643
rect 5166 16640 5172 16652
rect 5127 16612 5172 16640
rect 4985 16603 5043 16609
rect 5000 16516 5028 16603
rect 5166 16600 5172 16612
rect 5224 16600 5230 16652
rect 5350 16640 5356 16652
rect 5311 16612 5356 16640
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 5626 16640 5632 16652
rect 5587 16612 5632 16640
rect 5626 16600 5632 16612
rect 5684 16600 5690 16652
rect 6638 16640 6644 16652
rect 6551 16612 6644 16640
rect 6638 16600 6644 16612
rect 6696 16640 6702 16652
rect 7760 16640 7788 16671
rect 7834 16668 7840 16680
rect 7892 16668 7898 16720
rect 8018 16708 8024 16720
rect 7979 16680 8024 16708
rect 8018 16668 8024 16680
rect 8076 16668 8082 16720
rect 8113 16711 8171 16717
rect 8113 16677 8125 16711
rect 8159 16708 8171 16711
rect 8570 16708 8576 16720
rect 8159 16680 8576 16708
rect 8159 16677 8171 16680
rect 8113 16671 8171 16677
rect 7926 16640 7932 16652
rect 6696 16612 7788 16640
rect 7887 16612 7932 16640
rect 6696 16600 6702 16612
rect 7926 16600 7932 16612
rect 7984 16600 7990 16652
rect 4982 16464 4988 16516
rect 5040 16464 5046 16516
rect 3142 16396 3148 16448
rect 3200 16436 3206 16448
rect 8128 16436 8156 16671
rect 8570 16668 8576 16680
rect 8628 16668 8634 16720
rect 9416 16708 9444 16739
rect 9674 16736 9680 16788
rect 9732 16776 9738 16788
rect 9953 16779 10011 16785
rect 9953 16776 9965 16779
rect 9732 16748 9965 16776
rect 9732 16736 9738 16748
rect 9953 16745 9965 16748
rect 9999 16745 10011 16779
rect 9953 16739 10011 16745
rect 11054 16736 11060 16788
rect 11112 16776 11118 16788
rect 11793 16779 11851 16785
rect 11793 16776 11805 16779
rect 11112 16748 11805 16776
rect 11112 16736 11118 16748
rect 11793 16745 11805 16748
rect 11839 16745 11851 16779
rect 13357 16779 13415 16785
rect 13357 16776 13369 16779
rect 11793 16739 11851 16745
rect 12544 16748 13369 16776
rect 10226 16708 10232 16720
rect 9416 16680 10232 16708
rect 10226 16668 10232 16680
rect 10284 16668 10290 16720
rect 11149 16711 11207 16717
rect 11149 16677 11161 16711
rect 11195 16708 11207 16711
rect 11698 16708 11704 16720
rect 11195 16680 11704 16708
rect 11195 16677 11207 16680
rect 11149 16671 11207 16677
rect 11698 16668 11704 16680
rect 11756 16668 11762 16720
rect 11808 16708 11836 16739
rect 11808 16680 12204 16708
rect 8386 16600 8392 16652
rect 8444 16640 8450 16652
rect 8481 16643 8539 16649
rect 8481 16640 8493 16643
rect 8444 16612 8493 16640
rect 8444 16600 8450 16612
rect 8481 16609 8493 16612
rect 8527 16609 8539 16643
rect 8481 16603 8539 16609
rect 9769 16643 9827 16649
rect 9769 16609 9781 16643
rect 9815 16640 9827 16643
rect 9858 16640 9864 16652
rect 9815 16612 9864 16640
rect 9815 16609 9827 16612
rect 9769 16603 9827 16609
rect 9858 16600 9864 16612
rect 9916 16600 9922 16652
rect 10965 16643 11023 16649
rect 10965 16640 10977 16643
rect 10612 16612 10977 16640
rect 3200 16408 8156 16436
rect 3200 16396 3206 16408
rect 8938 16396 8944 16448
rect 8996 16436 9002 16448
rect 9033 16439 9091 16445
rect 9033 16436 9045 16439
rect 8996 16408 9045 16436
rect 8996 16396 9002 16408
rect 9033 16405 9045 16408
rect 9079 16405 9091 16439
rect 9033 16399 9091 16405
rect 10502 16396 10508 16448
rect 10560 16436 10566 16448
rect 10612 16445 10640 16612
rect 10965 16609 10977 16612
rect 11011 16609 11023 16643
rect 10965 16603 11023 16609
rect 11054 16600 11060 16652
rect 11112 16640 11118 16652
rect 11238 16640 11244 16652
rect 11112 16612 11244 16640
rect 11112 16600 11118 16612
rect 11238 16600 11244 16612
rect 11296 16600 11302 16652
rect 10781 16575 10839 16581
rect 10781 16541 10793 16575
rect 10827 16572 10839 16575
rect 10870 16572 10876 16584
rect 10827 16544 10876 16572
rect 10827 16541 10839 16544
rect 10781 16535 10839 16541
rect 10870 16532 10876 16544
rect 10928 16532 10934 16584
rect 11514 16572 11520 16584
rect 11475 16544 11520 16572
rect 11514 16532 11520 16544
rect 11572 16532 11578 16584
rect 12176 16504 12204 16680
rect 12544 16652 12572 16748
rect 13357 16745 13369 16748
rect 13403 16745 13415 16779
rect 14090 16776 14096 16788
rect 14051 16748 14096 16776
rect 13357 16739 13415 16745
rect 14090 16736 14096 16748
rect 14148 16736 14154 16788
rect 14734 16776 14740 16788
rect 14695 16748 14740 16776
rect 14734 16736 14740 16748
rect 14792 16736 14798 16788
rect 16022 16776 16028 16788
rect 15983 16748 16028 16776
rect 16022 16736 16028 16748
rect 16080 16736 16086 16788
rect 16485 16779 16543 16785
rect 16485 16745 16497 16779
rect 16531 16776 16543 16779
rect 16574 16776 16580 16788
rect 16531 16748 16580 16776
rect 16531 16745 16543 16748
rect 16485 16739 16543 16745
rect 16574 16736 16580 16748
rect 16632 16736 16638 16788
rect 18138 16736 18144 16788
rect 18196 16776 18202 16788
rect 18417 16779 18475 16785
rect 18417 16776 18429 16779
rect 18196 16748 18429 16776
rect 18196 16736 18202 16748
rect 18417 16745 18429 16748
rect 18463 16745 18475 16779
rect 20714 16776 20720 16788
rect 20675 16748 20720 16776
rect 18417 16739 18475 16745
rect 20714 16736 20720 16748
rect 20772 16736 20778 16788
rect 24854 16736 24860 16788
rect 24912 16776 24918 16788
rect 25409 16779 25467 16785
rect 25409 16776 25421 16779
rect 24912 16748 25421 16776
rect 24912 16736 24918 16748
rect 25409 16745 25421 16748
rect 25455 16745 25467 16779
rect 25409 16739 25467 16745
rect 26329 16779 26387 16785
rect 26329 16745 26341 16779
rect 26375 16776 26387 16779
rect 26602 16776 26608 16788
rect 26375 16748 26608 16776
rect 26375 16745 26387 16748
rect 26329 16739 26387 16745
rect 26602 16736 26608 16748
rect 26660 16776 26666 16788
rect 27709 16779 27767 16785
rect 27709 16776 27721 16779
rect 26660 16748 27721 16776
rect 26660 16736 26666 16748
rect 27709 16745 27721 16748
rect 27755 16776 27767 16779
rect 27890 16776 27896 16788
rect 27755 16748 27896 16776
rect 27755 16745 27767 16748
rect 27709 16739 27767 16745
rect 27890 16736 27896 16748
rect 27948 16736 27954 16788
rect 28534 16736 28540 16788
rect 28592 16776 28598 16788
rect 29730 16776 29736 16788
rect 28592 16748 29736 16776
rect 28592 16736 28598 16748
rect 13081 16711 13139 16717
rect 13081 16677 13093 16711
rect 13127 16708 13139 16711
rect 13170 16708 13176 16720
rect 13127 16680 13176 16708
rect 13127 16677 13139 16680
rect 13081 16671 13139 16677
rect 13170 16668 13176 16680
rect 13228 16668 13234 16720
rect 14274 16668 14280 16720
rect 14332 16708 14338 16720
rect 15010 16708 15016 16720
rect 14332 16680 15016 16708
rect 14332 16668 14338 16680
rect 15010 16668 15016 16680
rect 15068 16668 15074 16720
rect 17129 16711 17187 16717
rect 17129 16677 17141 16711
rect 17175 16708 17187 16711
rect 17218 16708 17224 16720
rect 17175 16680 17224 16708
rect 17175 16677 17187 16680
rect 17129 16671 17187 16677
rect 17218 16668 17224 16680
rect 17276 16668 17282 16720
rect 17310 16668 17316 16720
rect 17368 16708 17374 16720
rect 17368 16680 18828 16708
rect 17368 16668 17374 16680
rect 12253 16643 12311 16649
rect 12253 16609 12265 16643
rect 12299 16640 12311 16643
rect 12342 16640 12348 16652
rect 12299 16612 12348 16640
rect 12299 16609 12311 16612
rect 12253 16603 12311 16609
rect 12342 16600 12348 16612
rect 12400 16600 12406 16652
rect 12526 16640 12532 16652
rect 12487 16612 12532 16640
rect 12526 16600 12532 16612
rect 12584 16600 12590 16652
rect 12618 16600 12624 16652
rect 12676 16640 12682 16652
rect 13725 16643 13783 16649
rect 13725 16640 13737 16643
rect 12676 16612 13737 16640
rect 12676 16600 12682 16612
rect 13725 16609 13737 16612
rect 13771 16609 13783 16643
rect 13909 16643 13967 16649
rect 13909 16640 13921 16643
rect 13725 16603 13783 16609
rect 13832 16612 13921 16640
rect 13630 16532 13636 16584
rect 13688 16572 13694 16584
rect 13832 16572 13860 16612
rect 13909 16609 13921 16612
rect 13955 16640 13967 16643
rect 14182 16640 14188 16652
rect 13955 16612 14188 16640
rect 13955 16609 13967 16612
rect 13909 16603 13967 16609
rect 14182 16600 14188 16612
rect 14240 16600 14246 16652
rect 14366 16640 14372 16652
rect 14327 16612 14372 16640
rect 14366 16600 14372 16612
rect 14424 16600 14430 16652
rect 15562 16640 15568 16652
rect 15523 16612 15568 16640
rect 15562 16600 15568 16612
rect 15620 16600 15626 16652
rect 16666 16640 16672 16652
rect 16627 16612 16672 16640
rect 16666 16600 16672 16612
rect 16724 16600 16730 16652
rect 16942 16600 16948 16652
rect 17000 16640 17006 16652
rect 17405 16643 17463 16649
rect 17405 16640 17417 16643
rect 17000 16612 17417 16640
rect 17000 16600 17006 16612
rect 17405 16609 17417 16612
rect 17451 16640 17463 16643
rect 17494 16640 17500 16652
rect 17451 16612 17500 16640
rect 17451 16609 17463 16612
rect 17405 16603 17463 16609
rect 17494 16600 17500 16612
rect 17552 16600 17558 16652
rect 18601 16643 18659 16649
rect 18601 16609 18613 16643
rect 18647 16640 18659 16643
rect 18690 16640 18696 16652
rect 18647 16612 18696 16640
rect 18647 16609 18659 16612
rect 18601 16603 18659 16609
rect 18690 16600 18696 16612
rect 18748 16600 18754 16652
rect 18800 16649 18828 16680
rect 19150 16668 19156 16720
rect 19208 16708 19214 16720
rect 19429 16711 19487 16717
rect 19429 16708 19441 16711
rect 19208 16680 19441 16708
rect 19208 16668 19214 16680
rect 19429 16677 19441 16680
rect 19475 16677 19487 16711
rect 19794 16708 19800 16720
rect 19755 16680 19800 16708
rect 19429 16671 19487 16677
rect 19794 16668 19800 16680
rect 19852 16668 19858 16720
rect 20349 16711 20407 16717
rect 20349 16677 20361 16711
rect 20395 16708 20407 16711
rect 22922 16708 22928 16720
rect 20395 16680 21956 16708
rect 22883 16680 22928 16708
rect 20395 16677 20407 16680
rect 20349 16671 20407 16677
rect 21928 16652 21956 16680
rect 22922 16668 22928 16680
rect 22980 16668 22986 16720
rect 25958 16668 25964 16720
rect 26016 16708 26022 16720
rect 26513 16711 26571 16717
rect 26513 16708 26525 16711
rect 26016 16680 26525 16708
rect 26016 16668 26022 16680
rect 26513 16677 26525 16680
rect 26559 16677 26571 16711
rect 27246 16708 27252 16720
rect 27207 16680 27252 16708
rect 26513 16671 26571 16677
rect 27246 16668 27252 16680
rect 27304 16668 27310 16720
rect 29196 16717 29224 16748
rect 29730 16736 29736 16748
rect 29788 16736 29794 16788
rect 29822 16736 29828 16788
rect 29880 16776 29886 16788
rect 31294 16776 31300 16788
rect 29880 16748 29925 16776
rect 31255 16748 31300 16776
rect 29880 16736 29886 16748
rect 31294 16736 31300 16748
rect 31352 16736 31358 16788
rect 31386 16736 31392 16788
rect 31444 16776 31450 16788
rect 31573 16779 31631 16785
rect 31573 16776 31585 16779
rect 31444 16748 31585 16776
rect 31444 16736 31450 16748
rect 31573 16745 31585 16748
rect 31619 16745 31631 16779
rect 32858 16776 32864 16788
rect 32819 16748 32864 16776
rect 31573 16739 31631 16745
rect 32858 16736 32864 16748
rect 32916 16736 32922 16788
rect 33594 16736 33600 16788
rect 33652 16776 33658 16788
rect 34790 16776 34796 16788
rect 33652 16748 34796 16776
rect 33652 16736 33658 16748
rect 34790 16736 34796 16748
rect 34848 16776 34854 16788
rect 35250 16776 35256 16788
rect 34848 16748 35256 16776
rect 34848 16736 34854 16748
rect 35250 16736 35256 16748
rect 35308 16736 35314 16788
rect 29181 16711 29239 16717
rect 29181 16677 29193 16711
rect 29227 16677 29239 16711
rect 29181 16671 29239 16677
rect 29454 16668 29460 16720
rect 29512 16708 29518 16720
rect 30282 16708 30288 16720
rect 29512 16680 30288 16708
rect 29512 16668 29518 16680
rect 30282 16668 30288 16680
rect 30340 16668 30346 16720
rect 31018 16668 31024 16720
rect 31076 16708 31082 16720
rect 31662 16708 31668 16720
rect 31076 16680 31668 16708
rect 31076 16668 31082 16680
rect 31662 16668 31668 16680
rect 31720 16708 31726 16720
rect 32876 16708 32904 16736
rect 33318 16708 33324 16720
rect 31720 16680 32904 16708
rect 32968 16680 33324 16708
rect 31720 16668 31726 16680
rect 18785 16643 18843 16649
rect 18785 16609 18797 16643
rect 18831 16640 18843 16643
rect 19242 16640 19248 16652
rect 18831 16612 19248 16640
rect 18831 16609 18843 16612
rect 18785 16603 18843 16609
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 20990 16600 20996 16652
rect 21048 16640 21054 16652
rect 21545 16643 21603 16649
rect 21545 16640 21557 16643
rect 21048 16612 21557 16640
rect 21048 16600 21054 16612
rect 21545 16609 21557 16612
rect 21591 16609 21603 16643
rect 21910 16640 21916 16652
rect 21871 16612 21916 16640
rect 21545 16603 21603 16609
rect 21910 16600 21916 16612
rect 21968 16600 21974 16652
rect 22094 16600 22100 16652
rect 22152 16640 22158 16652
rect 22373 16643 22431 16649
rect 22373 16640 22385 16643
rect 22152 16612 22385 16640
rect 22152 16600 22158 16612
rect 22373 16609 22385 16612
rect 22419 16640 22431 16643
rect 22741 16643 22799 16649
rect 22741 16640 22753 16643
rect 22419 16612 22753 16640
rect 22419 16609 22431 16612
rect 22373 16603 22431 16609
rect 22741 16609 22753 16612
rect 22787 16640 22799 16643
rect 23753 16643 23811 16649
rect 23753 16640 23765 16643
rect 22787 16612 23765 16640
rect 22787 16609 22799 16612
rect 22741 16603 22799 16609
rect 23753 16609 23765 16612
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 24118 16600 24124 16652
rect 24176 16640 24182 16652
rect 24305 16643 24363 16649
rect 24305 16640 24317 16643
rect 24176 16612 24317 16640
rect 24176 16600 24182 16612
rect 24305 16609 24317 16612
rect 24351 16640 24363 16643
rect 24670 16640 24676 16652
rect 24351 16612 24676 16640
rect 24351 16609 24363 16612
rect 24305 16603 24363 16609
rect 24670 16600 24676 16612
rect 24728 16640 24734 16652
rect 24765 16643 24823 16649
rect 24765 16640 24777 16643
rect 24728 16612 24777 16640
rect 24728 16600 24734 16612
rect 24765 16609 24777 16612
rect 24811 16609 24823 16643
rect 24765 16603 24823 16609
rect 24946 16600 24952 16652
rect 25004 16600 25010 16652
rect 26050 16600 26056 16652
rect 26108 16640 26114 16652
rect 28997 16643 29055 16649
rect 28997 16640 29009 16643
rect 26108 16612 26280 16640
rect 26108 16600 26114 16612
rect 13688 16544 13860 16572
rect 16577 16575 16635 16581
rect 13688 16532 13694 16544
rect 16577 16541 16589 16575
rect 16623 16572 16635 16575
rect 17310 16572 17316 16584
rect 16623 16544 17316 16572
rect 16623 16541 16635 16544
rect 16577 16535 16635 16541
rect 17310 16532 17316 16544
rect 17368 16532 17374 16584
rect 19153 16575 19211 16581
rect 19153 16541 19165 16575
rect 19199 16572 19211 16575
rect 19334 16572 19340 16584
rect 19199 16544 19340 16572
rect 19199 16541 19211 16544
rect 19153 16535 19211 16541
rect 19334 16532 19340 16544
rect 19392 16532 19398 16584
rect 21174 16532 21180 16584
rect 21232 16572 21238 16584
rect 21358 16572 21364 16584
rect 21232 16544 21364 16572
rect 21232 16532 21238 16544
rect 21358 16532 21364 16544
rect 21416 16532 21422 16584
rect 21634 16532 21640 16584
rect 21692 16572 21698 16584
rect 21821 16575 21879 16581
rect 21821 16572 21833 16575
rect 21692 16544 21833 16572
rect 21692 16532 21698 16544
rect 21821 16541 21833 16544
rect 21867 16541 21879 16575
rect 21821 16535 21879 16541
rect 23106 16532 23112 16584
rect 23164 16572 23170 16584
rect 23477 16575 23535 16581
rect 23477 16572 23489 16575
rect 23164 16544 23489 16572
rect 23164 16532 23170 16544
rect 23477 16541 23489 16544
rect 23523 16541 23535 16575
rect 23934 16572 23940 16584
rect 23895 16544 23940 16572
rect 23477 16535 23535 16541
rect 23934 16532 23940 16544
rect 23992 16532 23998 16584
rect 24394 16532 24400 16584
rect 24452 16572 24458 16584
rect 24964 16572 24992 16600
rect 25133 16575 25191 16581
rect 25133 16572 25145 16575
rect 24452 16544 25145 16572
rect 24452 16532 24458 16544
rect 25133 16541 25145 16544
rect 25179 16541 25191 16575
rect 26252 16572 26280 16612
rect 28092 16612 29009 16640
rect 26326 16572 26332 16584
rect 26252 16544 26332 16572
rect 25133 16535 25191 16541
rect 26326 16532 26332 16544
rect 26384 16532 26390 16584
rect 26694 16532 26700 16584
rect 26752 16572 26758 16584
rect 26881 16575 26939 16581
rect 26881 16572 26893 16575
rect 26752 16544 26893 16572
rect 26752 16532 26758 16544
rect 26881 16541 26893 16544
rect 26927 16541 26939 16575
rect 26881 16535 26939 16541
rect 12345 16507 12403 16513
rect 12345 16504 12357 16507
rect 12176 16476 12357 16504
rect 12345 16473 12357 16476
rect 12391 16473 12403 16507
rect 26789 16507 26847 16513
rect 26789 16504 26801 16507
rect 12345 16467 12403 16473
rect 25884 16476 26801 16504
rect 25884 16448 25912 16476
rect 26789 16473 26801 16476
rect 26835 16473 26847 16507
rect 26789 16467 26847 16473
rect 28092 16448 28120 16612
rect 28997 16609 29009 16612
rect 29043 16609 29055 16643
rect 28997 16603 29055 16609
rect 29089 16643 29147 16649
rect 29089 16609 29101 16643
rect 29135 16640 29147 16643
rect 29362 16640 29368 16652
rect 29135 16612 29368 16640
rect 29135 16609 29147 16612
rect 29089 16603 29147 16609
rect 29362 16600 29368 16612
rect 29420 16600 29426 16652
rect 30190 16600 30196 16652
rect 30248 16640 30254 16652
rect 30561 16643 30619 16649
rect 30561 16640 30573 16643
rect 30248 16612 30573 16640
rect 30248 16600 30254 16612
rect 30561 16609 30573 16612
rect 30607 16609 30619 16643
rect 30742 16640 30748 16652
rect 30703 16612 30748 16640
rect 30561 16603 30619 16609
rect 30742 16600 30748 16612
rect 30800 16600 30806 16652
rect 32401 16643 32459 16649
rect 32401 16609 32413 16643
rect 32447 16640 32459 16643
rect 32490 16640 32496 16652
rect 32447 16612 32496 16640
rect 32447 16609 32459 16612
rect 32401 16603 32459 16609
rect 32490 16600 32496 16612
rect 32548 16640 32554 16652
rect 32968 16640 32996 16680
rect 33318 16668 33324 16680
rect 33376 16668 33382 16720
rect 34517 16711 34575 16717
rect 34517 16677 34529 16711
rect 34563 16708 34575 16711
rect 34698 16708 34704 16720
rect 34563 16680 34704 16708
rect 34563 16677 34575 16680
rect 34517 16671 34575 16677
rect 34698 16668 34704 16680
rect 34756 16668 34762 16720
rect 32548 16612 32996 16640
rect 33505 16643 33563 16649
rect 32548 16600 32554 16612
rect 33505 16609 33517 16643
rect 33551 16640 33563 16643
rect 33686 16640 33692 16652
rect 33551 16612 33692 16640
rect 33551 16609 33563 16612
rect 33505 16603 33563 16609
rect 33686 16600 33692 16612
rect 33744 16600 33750 16652
rect 33781 16643 33839 16649
rect 33781 16609 33793 16643
rect 33827 16609 33839 16643
rect 33781 16603 33839 16609
rect 28813 16575 28871 16581
rect 28813 16541 28825 16575
rect 28859 16572 28871 16575
rect 29270 16572 29276 16584
rect 28859 16544 29276 16572
rect 28859 16541 28871 16544
rect 28813 16535 28871 16541
rect 29270 16532 29276 16544
rect 29328 16532 29334 16584
rect 29549 16575 29607 16581
rect 29549 16541 29561 16575
rect 29595 16541 29607 16575
rect 29549 16535 29607 16541
rect 10597 16439 10655 16445
rect 10597 16436 10609 16439
rect 10560 16408 10609 16436
rect 10560 16396 10566 16408
rect 10597 16405 10609 16408
rect 10643 16405 10655 16439
rect 10597 16399 10655 16405
rect 15749 16439 15807 16445
rect 15749 16405 15761 16439
rect 15795 16436 15807 16439
rect 16206 16436 16212 16448
rect 15795 16408 16212 16436
rect 15795 16405 15807 16408
rect 15749 16399 15807 16405
rect 16206 16396 16212 16408
rect 16264 16396 16270 16448
rect 17770 16396 17776 16448
rect 17828 16436 17834 16448
rect 18049 16439 18107 16445
rect 18049 16436 18061 16439
rect 17828 16408 18061 16436
rect 17828 16396 17834 16408
rect 18049 16405 18061 16408
rect 18095 16436 18107 16439
rect 18322 16436 18328 16448
rect 18095 16408 18328 16436
rect 18095 16405 18107 16408
rect 18049 16399 18107 16405
rect 18322 16396 18328 16408
rect 18380 16396 18386 16448
rect 21177 16439 21235 16445
rect 21177 16405 21189 16439
rect 21223 16436 21235 16439
rect 21542 16436 21548 16448
rect 21223 16408 21548 16436
rect 21223 16405 21235 16408
rect 21177 16399 21235 16405
rect 21542 16396 21548 16408
rect 21600 16396 21606 16448
rect 24673 16439 24731 16445
rect 24673 16405 24685 16439
rect 24719 16436 24731 16439
rect 24854 16436 24860 16448
rect 24719 16408 24860 16436
rect 24719 16405 24731 16408
rect 24673 16399 24731 16405
rect 24854 16396 24860 16408
rect 24912 16445 24918 16448
rect 24912 16439 24961 16445
rect 24912 16405 24915 16439
rect 24949 16405 24961 16439
rect 25038 16436 25044 16448
rect 24999 16408 25044 16436
rect 24912 16399 24961 16405
rect 24912 16396 24918 16399
rect 25038 16396 25044 16408
rect 25096 16436 25102 16448
rect 25866 16436 25872 16448
rect 25096 16408 25872 16436
rect 25096 16396 25102 16408
rect 25866 16396 25872 16408
rect 25924 16396 25930 16448
rect 26602 16396 26608 16448
rect 26660 16445 26666 16448
rect 26660 16439 26709 16445
rect 26660 16405 26663 16439
rect 26697 16405 26709 16439
rect 28074 16436 28080 16448
rect 28035 16408 28080 16436
rect 26660 16399 26709 16405
rect 26660 16396 26666 16399
rect 28074 16396 28080 16408
rect 28132 16396 28138 16448
rect 28534 16396 28540 16448
rect 28592 16436 28598 16448
rect 28629 16439 28687 16445
rect 28629 16436 28641 16439
rect 28592 16408 28641 16436
rect 28592 16396 28598 16408
rect 28629 16405 28641 16408
rect 28675 16405 28687 16439
rect 28629 16399 28687 16405
rect 28810 16396 28816 16448
rect 28868 16436 28874 16448
rect 29564 16436 29592 16535
rect 32858 16532 32864 16584
rect 32916 16572 32922 16584
rect 33042 16572 33048 16584
rect 32916 16544 33048 16572
rect 32916 16532 32922 16544
rect 33042 16532 33048 16544
rect 33100 16532 33106 16584
rect 33796 16572 33824 16603
rect 33870 16572 33876 16584
rect 33704 16544 33876 16572
rect 32214 16464 32220 16516
rect 32272 16504 32278 16516
rect 33704 16504 33732 16544
rect 33870 16532 33876 16544
rect 33928 16532 33934 16584
rect 34054 16572 34060 16584
rect 34015 16544 34060 16572
rect 34054 16532 34060 16544
rect 34112 16532 34118 16584
rect 32272 16476 33732 16504
rect 32272 16464 32278 16476
rect 30926 16436 30932 16448
rect 28868 16408 29592 16436
rect 30887 16408 30932 16436
rect 28868 16396 28874 16408
rect 30926 16396 30932 16408
rect 30984 16396 30990 16448
rect 1104 16346 38548 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 38548 16346
rect 1104 16272 38548 16294
rect 3513 16235 3571 16241
rect 3513 16201 3525 16235
rect 3559 16232 3571 16235
rect 4062 16232 4068 16244
rect 3559 16204 4068 16232
rect 3559 16201 3571 16204
rect 3513 16195 3571 16201
rect 4062 16192 4068 16204
rect 4120 16192 4126 16244
rect 4798 16232 4804 16244
rect 4711 16204 4804 16232
rect 4798 16192 4804 16204
rect 4856 16232 4862 16244
rect 5350 16232 5356 16244
rect 4856 16204 5356 16232
rect 4856 16192 4862 16204
rect 5350 16192 5356 16204
rect 5408 16192 5414 16244
rect 6273 16235 6331 16241
rect 6273 16201 6285 16235
rect 6319 16232 6331 16235
rect 6638 16232 6644 16244
rect 6319 16204 6644 16232
rect 6319 16201 6331 16204
rect 6273 16195 6331 16201
rect 6638 16192 6644 16204
rect 6696 16192 6702 16244
rect 7834 16192 7840 16244
rect 7892 16232 7898 16244
rect 8297 16235 8355 16241
rect 8297 16232 8309 16235
rect 7892 16204 8309 16232
rect 7892 16192 7898 16204
rect 8297 16201 8309 16204
rect 8343 16232 8355 16235
rect 10870 16232 10876 16244
rect 8343 16204 10876 16232
rect 8343 16201 8355 16204
rect 8297 16195 8355 16201
rect 10870 16192 10876 16204
rect 10928 16232 10934 16244
rect 10965 16235 11023 16241
rect 10965 16232 10977 16235
rect 10928 16204 10977 16232
rect 10928 16192 10934 16204
rect 10965 16201 10977 16204
rect 11011 16232 11023 16235
rect 11241 16235 11299 16241
rect 11241 16232 11253 16235
rect 11011 16204 11253 16232
rect 11011 16201 11023 16204
rect 10965 16195 11023 16201
rect 11241 16201 11253 16204
rect 11287 16201 11299 16235
rect 11241 16195 11299 16201
rect 13446 16192 13452 16244
rect 13504 16232 13510 16244
rect 14277 16235 14335 16241
rect 14277 16232 14289 16235
rect 13504 16204 14289 16232
rect 13504 16192 13510 16204
rect 14277 16201 14289 16204
rect 14323 16201 14335 16235
rect 16666 16232 16672 16244
rect 16627 16204 16672 16232
rect 14277 16195 14335 16201
rect 16666 16192 16672 16204
rect 16724 16192 16730 16244
rect 17037 16235 17095 16241
rect 17037 16201 17049 16235
rect 17083 16232 17095 16235
rect 17310 16232 17316 16244
rect 17083 16204 17316 16232
rect 17083 16201 17095 16204
rect 17037 16195 17095 16201
rect 4614 16164 4620 16176
rect 4527 16136 4620 16164
rect 4614 16124 4620 16136
rect 4672 16164 4678 16176
rect 5074 16164 5080 16176
rect 4672 16136 5080 16164
rect 4672 16124 4678 16136
rect 5074 16124 5080 16136
rect 5132 16164 5138 16176
rect 5718 16164 5724 16176
rect 5132 16136 5724 16164
rect 5132 16124 5138 16136
rect 5718 16124 5724 16136
rect 5776 16124 5782 16176
rect 7929 16167 7987 16173
rect 7929 16133 7941 16167
rect 7975 16164 7987 16167
rect 8018 16164 8024 16176
rect 7975 16136 8024 16164
rect 7975 16133 7987 16136
rect 7929 16127 7987 16133
rect 8018 16124 8024 16136
rect 8076 16124 8082 16176
rect 9306 16124 9312 16176
rect 9364 16164 9370 16176
rect 9950 16164 9956 16176
rect 9364 16136 9956 16164
rect 9364 16124 9370 16136
rect 9950 16124 9956 16136
rect 10008 16124 10014 16176
rect 13541 16167 13599 16173
rect 13541 16133 13553 16167
rect 13587 16164 13599 16167
rect 13630 16164 13636 16176
rect 13587 16136 13636 16164
rect 13587 16133 13599 16136
rect 13541 16127 13599 16133
rect 1394 16096 1400 16108
rect 1355 16068 1400 16096
rect 1394 16056 1400 16068
rect 1452 16056 1458 16108
rect 1670 16096 1676 16108
rect 1631 16068 1676 16096
rect 1670 16056 1676 16068
rect 1728 16056 1734 16108
rect 3881 16099 3939 16105
rect 3881 16065 3893 16099
rect 3927 16096 3939 16099
rect 4706 16096 4712 16108
rect 3927 16068 4712 16096
rect 3927 16065 3939 16068
rect 3881 16059 3939 16065
rect 4706 16056 4712 16068
rect 4764 16096 4770 16108
rect 5258 16096 5264 16108
rect 4764 16068 5264 16096
rect 4764 16056 4770 16068
rect 5258 16056 5264 16068
rect 5316 16056 5322 16108
rect 7561 16099 7619 16105
rect 7561 16096 7573 16099
rect 5368 16068 7573 16096
rect 5368 16040 5396 16068
rect 7561 16065 7573 16068
rect 7607 16065 7619 16099
rect 10226 16096 10232 16108
rect 10187 16068 10232 16096
rect 7561 16059 7619 16065
rect 10226 16056 10232 16068
rect 10284 16056 10290 16108
rect 5350 16028 5356 16040
rect 5263 16000 5356 16028
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 5718 16028 5724 16040
rect 5679 16000 5724 16028
rect 5718 15988 5724 16000
rect 5776 15988 5782 16040
rect 5905 16031 5963 16037
rect 5905 15997 5917 16031
rect 5951 16028 5963 16031
rect 6270 16028 6276 16040
rect 5951 16000 6276 16028
rect 5951 15997 5963 16000
rect 5905 15991 5963 15997
rect 6270 15988 6276 16000
rect 6328 15988 6334 16040
rect 6638 15988 6644 16040
rect 6696 16028 6702 16040
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 6696 16000 6837 16028
rect 6696 15988 6702 16000
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 6825 15991 6883 15997
rect 6914 15988 6920 16040
rect 6972 16028 6978 16040
rect 7101 16031 7159 16037
rect 7101 16028 7113 16031
rect 6972 16000 7113 16028
rect 6972 15988 6978 16000
rect 7101 15997 7113 16000
rect 7147 15997 7159 16031
rect 7101 15991 7159 15997
rect 8665 16031 8723 16037
rect 8665 15997 8677 16031
rect 8711 16028 8723 16031
rect 8846 16028 8852 16040
rect 8711 16000 8852 16028
rect 8711 15997 8723 16000
rect 8665 15991 8723 15997
rect 8846 15988 8852 16000
rect 8904 15988 8910 16040
rect 9214 16028 9220 16040
rect 9175 16000 9220 16028
rect 9214 15988 9220 16000
rect 9272 15988 9278 16040
rect 9769 16031 9827 16037
rect 9769 15997 9781 16031
rect 9815 16028 9827 16031
rect 9950 16028 9956 16040
rect 9815 16000 9956 16028
rect 9815 15997 9827 16000
rect 9769 15991 9827 15997
rect 9950 15988 9956 16000
rect 10008 15988 10014 16040
rect 10137 16031 10195 16037
rect 10137 15997 10149 16031
rect 10183 16028 10195 16031
rect 10686 16028 10692 16040
rect 10183 16000 10692 16028
rect 10183 15997 10195 16000
rect 10137 15991 10195 15997
rect 10686 15988 10692 16000
rect 10744 15988 10750 16040
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 16028 11115 16031
rect 11333 16031 11391 16037
rect 11333 16028 11345 16031
rect 11103 16000 11345 16028
rect 11103 15997 11115 16000
rect 11057 15991 11115 15997
rect 11333 15997 11345 16000
rect 11379 15997 11391 16031
rect 12621 16031 12679 16037
rect 12621 16028 12633 16031
rect 11333 15991 11391 15997
rect 12176 16000 12633 16028
rect 3053 15963 3111 15969
rect 3053 15929 3065 15963
rect 3099 15960 3111 15963
rect 3878 15960 3884 15972
rect 3099 15932 3884 15960
rect 3099 15929 3111 15932
rect 3053 15923 3111 15929
rect 3878 15920 3884 15932
rect 3936 15920 3942 15972
rect 4249 15963 4307 15969
rect 4249 15929 4261 15963
rect 4295 15960 4307 15963
rect 5626 15960 5632 15972
rect 4295 15932 5632 15960
rect 4295 15929 4307 15932
rect 4249 15923 4307 15929
rect 5626 15920 5632 15932
rect 5684 15920 5690 15972
rect 7190 15960 7196 15972
rect 6932 15932 7196 15960
rect 6822 15852 6828 15904
rect 6880 15892 6886 15904
rect 6932 15892 6960 15932
rect 7190 15920 7196 15932
rect 7248 15920 7254 15972
rect 11146 15920 11152 15972
rect 11204 15960 11210 15972
rect 12176 15969 12204 16000
rect 12621 15997 12633 16000
rect 12667 16028 12679 16031
rect 13354 16028 13360 16040
rect 12667 16000 13360 16028
rect 12667 15997 12679 16000
rect 12621 15991 12679 15997
rect 13354 15988 13360 16000
rect 13412 16028 13418 16040
rect 13556 16028 13584 16127
rect 13630 16124 13636 16136
rect 13688 16124 13694 16176
rect 14550 16124 14556 16176
rect 14608 16164 14614 16176
rect 15102 16164 15108 16176
rect 14608 16136 15108 16164
rect 14608 16124 14614 16136
rect 15102 16124 15108 16136
rect 15160 16124 15166 16176
rect 15194 16124 15200 16176
rect 15252 16164 15258 16176
rect 16209 16167 16267 16173
rect 16209 16164 16221 16167
rect 15252 16136 16221 16164
rect 15252 16124 15258 16136
rect 16209 16133 16221 16136
rect 16255 16133 16267 16167
rect 16209 16127 16267 16133
rect 15562 16096 15568 16108
rect 14016 16068 15568 16096
rect 13906 16028 13912 16040
rect 13412 16000 13584 16028
rect 13819 16000 13912 16028
rect 13412 15988 13418 16000
rect 13906 15988 13912 16000
rect 13964 16028 13970 16040
rect 14016 16037 14044 16068
rect 15562 16056 15568 16068
rect 15620 16056 15626 16108
rect 14001 16031 14059 16037
rect 14001 16028 14013 16031
rect 13964 16000 14013 16028
rect 13964 15988 13970 16000
rect 14001 15997 14013 16000
rect 14047 15997 14059 16031
rect 14001 15991 14059 15997
rect 14185 16031 14243 16037
rect 14185 15997 14197 16031
rect 14231 15997 14243 16031
rect 14185 15991 14243 15997
rect 16025 16031 16083 16037
rect 16025 15997 16037 16031
rect 16071 16028 16083 16031
rect 16114 16028 16120 16040
rect 16071 16000 16120 16028
rect 16071 15997 16083 16000
rect 16025 15991 16083 15997
rect 12161 15963 12219 15969
rect 12161 15960 12173 15963
rect 11204 15932 12173 15960
rect 11204 15920 11210 15932
rect 12161 15929 12173 15932
rect 12207 15929 12219 15963
rect 12434 15960 12440 15972
rect 12161 15923 12219 15929
rect 12268 15932 12440 15960
rect 6880 15864 6960 15892
rect 7009 15895 7067 15901
rect 6880 15852 6886 15864
rect 7009 15861 7021 15895
rect 7055 15892 7067 15895
rect 7282 15892 7288 15904
rect 7055 15864 7288 15892
rect 7055 15861 7067 15864
rect 7009 15855 7067 15861
rect 7282 15852 7288 15864
rect 7340 15852 7346 15904
rect 9858 15852 9864 15904
rect 9916 15892 9922 15904
rect 10597 15895 10655 15901
rect 10597 15892 10609 15895
rect 9916 15864 10609 15892
rect 9916 15852 9922 15864
rect 10597 15861 10609 15864
rect 10643 15892 10655 15895
rect 11238 15892 11244 15904
rect 10643 15864 11244 15892
rect 10643 15861 10655 15864
rect 10597 15855 10655 15861
rect 11238 15852 11244 15864
rect 11296 15852 11302 15904
rect 11333 15895 11391 15901
rect 11333 15861 11345 15895
rect 11379 15892 11391 15895
rect 11606 15892 11612 15904
rect 11379 15864 11612 15892
rect 11379 15861 11391 15864
rect 11333 15855 11391 15861
rect 11606 15852 11612 15864
rect 11664 15892 11670 15904
rect 12268 15892 12296 15932
rect 12434 15920 12440 15932
rect 12492 15960 12498 15972
rect 12802 15960 12808 15972
rect 12492 15932 12537 15960
rect 12763 15932 12808 15960
rect 12492 15920 12498 15932
rect 12802 15920 12808 15932
rect 12860 15920 12866 15972
rect 13170 15960 13176 15972
rect 13131 15932 13176 15960
rect 13170 15920 13176 15932
rect 13228 15920 13234 15972
rect 14200 15904 14228 15991
rect 16114 15988 16120 16000
rect 16172 16028 16178 16040
rect 17052 16028 17080 16195
rect 17310 16192 17316 16204
rect 17368 16192 17374 16244
rect 19150 16192 19156 16244
rect 19208 16232 19214 16244
rect 19889 16235 19947 16241
rect 19889 16232 19901 16235
rect 19208 16204 19901 16232
rect 19208 16192 19214 16204
rect 19889 16201 19901 16204
rect 19935 16201 19947 16235
rect 19889 16195 19947 16201
rect 21174 16192 21180 16244
rect 21232 16232 21238 16244
rect 21361 16235 21419 16241
rect 21361 16232 21373 16235
rect 21232 16204 21373 16232
rect 21232 16192 21238 16204
rect 21361 16201 21373 16204
rect 21407 16232 21419 16235
rect 21634 16232 21640 16244
rect 21407 16204 21640 16232
rect 21407 16201 21419 16204
rect 21361 16195 21419 16201
rect 21634 16192 21640 16204
rect 21692 16192 21698 16244
rect 23017 16235 23075 16241
rect 23017 16201 23029 16235
rect 23063 16232 23075 16235
rect 23934 16232 23940 16244
rect 23063 16204 23940 16232
rect 23063 16201 23075 16204
rect 23017 16195 23075 16201
rect 23934 16192 23940 16204
rect 23992 16192 23998 16244
rect 25222 16232 25228 16244
rect 25183 16204 25228 16232
rect 25222 16192 25228 16204
rect 25280 16192 25286 16244
rect 26234 16192 26240 16244
rect 26292 16232 26298 16244
rect 26605 16235 26663 16241
rect 26605 16232 26617 16235
rect 26292 16204 26617 16232
rect 26292 16192 26298 16204
rect 26605 16201 26617 16204
rect 26651 16201 26663 16235
rect 26605 16195 26663 16201
rect 27798 16192 27804 16244
rect 27856 16232 27862 16244
rect 28629 16235 28687 16241
rect 28629 16232 28641 16235
rect 27856 16204 28641 16232
rect 27856 16192 27862 16204
rect 17218 16124 17224 16176
rect 17276 16164 17282 16176
rect 17405 16167 17463 16173
rect 17405 16164 17417 16167
rect 17276 16136 17417 16164
rect 17276 16124 17282 16136
rect 17405 16133 17417 16136
rect 17451 16133 17463 16167
rect 22370 16164 22376 16176
rect 22331 16136 22376 16164
rect 17405 16127 17463 16133
rect 22370 16124 22376 16136
rect 22428 16124 22434 16176
rect 25038 16164 25044 16176
rect 24999 16136 25044 16164
rect 25038 16124 25044 16136
rect 25096 16124 25102 16176
rect 26050 16124 26056 16176
rect 26108 16164 26114 16176
rect 26510 16173 26516 16176
rect 26494 16167 26516 16173
rect 26494 16164 26506 16167
rect 26108 16136 26506 16164
rect 26108 16124 26114 16136
rect 26494 16133 26506 16136
rect 26494 16127 26516 16133
rect 26510 16124 26516 16127
rect 26568 16124 26574 16176
rect 26789 16167 26847 16173
rect 26789 16164 26801 16167
rect 26620 16136 26801 16164
rect 18782 16096 18788 16108
rect 18432 16068 18788 16096
rect 16172 16000 17080 16028
rect 16172 15988 16178 16000
rect 17770 15988 17776 16040
rect 17828 16028 17834 16040
rect 18325 16031 18383 16037
rect 18325 16028 18337 16031
rect 17828 16000 18337 16028
rect 17828 15988 17834 16000
rect 18325 15997 18337 16000
rect 18371 15997 18383 16031
rect 18325 15991 18383 15997
rect 15562 15920 15568 15972
rect 15620 15960 15626 15972
rect 18432 15969 18460 16068
rect 18782 16056 18788 16068
rect 18840 16056 18846 16108
rect 20993 16099 21051 16105
rect 20993 16065 21005 16099
rect 21039 16096 21051 16099
rect 21358 16096 21364 16108
rect 21039 16068 21364 16096
rect 21039 16065 21051 16068
rect 20993 16059 21051 16065
rect 21358 16056 21364 16068
rect 21416 16056 21422 16108
rect 21729 16099 21787 16105
rect 21729 16065 21741 16099
rect 21775 16096 21787 16099
rect 22094 16096 22100 16108
rect 21775 16068 22100 16096
rect 21775 16065 21787 16068
rect 21729 16059 21787 16065
rect 22094 16056 22100 16068
rect 22152 16056 22158 16108
rect 24673 16099 24731 16105
rect 24673 16065 24685 16099
rect 24719 16096 24731 16099
rect 25133 16099 25191 16105
rect 25133 16096 25145 16099
rect 24719 16068 25145 16096
rect 24719 16065 24731 16068
rect 24673 16059 24731 16065
rect 25133 16065 25145 16068
rect 25179 16096 25191 16099
rect 25777 16099 25835 16105
rect 25777 16096 25789 16099
rect 25179 16068 25789 16096
rect 25179 16065 25191 16068
rect 25133 16059 25191 16065
rect 25777 16065 25789 16068
rect 25823 16065 25835 16099
rect 25777 16059 25835 16065
rect 18506 15988 18512 16040
rect 18564 16028 18570 16040
rect 18966 16028 18972 16040
rect 18564 16000 18972 16028
rect 18564 15988 18570 16000
rect 18966 15988 18972 16000
rect 19024 15988 19030 16040
rect 19242 15988 19248 16040
rect 19300 16028 19306 16040
rect 19613 16031 19671 16037
rect 19613 16028 19625 16031
rect 19300 16000 19625 16028
rect 19300 15988 19306 16000
rect 19613 15997 19625 16000
rect 19659 15997 19671 16031
rect 19613 15991 19671 15997
rect 19705 16031 19763 16037
rect 19705 15997 19717 16031
rect 19751 16028 19763 16031
rect 19978 16028 19984 16040
rect 19751 16000 19984 16028
rect 19751 15997 19763 16000
rect 19705 15991 19763 15997
rect 15657 15963 15715 15969
rect 15657 15960 15669 15963
rect 15620 15932 15669 15960
rect 15620 15920 15626 15932
rect 15657 15929 15669 15932
rect 15703 15960 15715 15963
rect 18049 15963 18107 15969
rect 15703 15932 17724 15960
rect 15703 15929 15715 15932
rect 15657 15923 15715 15929
rect 17696 15904 17724 15932
rect 18049 15929 18061 15963
rect 18095 15929 18107 15963
rect 18417 15963 18475 15969
rect 18417 15960 18429 15963
rect 18049 15923 18107 15929
rect 18340 15932 18429 15960
rect 11664 15864 12296 15892
rect 11664 15852 11670 15864
rect 12342 15852 12348 15904
rect 12400 15892 12406 15904
rect 12526 15892 12532 15904
rect 12400 15864 12532 15892
rect 12400 15852 12406 15864
rect 12526 15852 12532 15864
rect 12584 15892 12590 15904
rect 12713 15895 12771 15901
rect 12713 15892 12725 15895
rect 12584 15864 12725 15892
rect 12584 15852 12590 15864
rect 12713 15861 12725 15864
rect 12759 15861 12771 15895
rect 12713 15855 12771 15861
rect 14182 15852 14188 15904
rect 14240 15892 14246 15904
rect 14829 15895 14887 15901
rect 14829 15892 14841 15895
rect 14240 15864 14841 15892
rect 14240 15852 14246 15864
rect 14829 15861 14841 15864
rect 14875 15861 14887 15895
rect 15194 15892 15200 15904
rect 15155 15864 15200 15892
rect 14829 15855 14887 15861
rect 15194 15852 15200 15864
rect 15252 15852 15258 15904
rect 17678 15852 17684 15904
rect 17736 15892 17742 15904
rect 17773 15895 17831 15901
rect 17773 15892 17785 15895
rect 17736 15864 17785 15892
rect 17736 15852 17742 15864
rect 17773 15861 17785 15864
rect 17819 15892 17831 15895
rect 18064 15892 18092 15923
rect 18340 15904 18368 15932
rect 18417 15929 18429 15932
rect 18463 15929 18475 15963
rect 18782 15960 18788 15972
rect 18743 15932 18788 15960
rect 18417 15923 18475 15929
rect 18782 15920 18788 15932
rect 18840 15920 18846 15972
rect 17819 15864 18092 15892
rect 17819 15861 17831 15864
rect 17773 15855 17831 15861
rect 18138 15852 18144 15904
rect 18196 15892 18202 15904
rect 18233 15895 18291 15901
rect 18233 15892 18245 15895
rect 18196 15864 18245 15892
rect 18196 15852 18202 15864
rect 18233 15861 18245 15864
rect 18279 15861 18291 15895
rect 18233 15855 18291 15861
rect 18322 15852 18328 15904
rect 18380 15852 18386 15904
rect 18690 15852 18696 15904
rect 18748 15892 18754 15904
rect 19061 15895 19119 15901
rect 19061 15892 19073 15895
rect 18748 15864 19073 15892
rect 18748 15852 18754 15864
rect 19061 15861 19073 15864
rect 19107 15861 19119 15895
rect 19061 15855 19119 15861
rect 19521 15895 19579 15901
rect 19521 15861 19533 15895
rect 19567 15892 19579 15895
rect 19628 15892 19656 15991
rect 19978 15988 19984 16000
rect 20036 15988 20042 16040
rect 21818 15988 21824 16040
rect 21876 16028 21882 16040
rect 21913 16031 21971 16037
rect 21913 16028 21925 16031
rect 21876 16000 21925 16028
rect 21876 15988 21882 16000
rect 21913 15997 21925 16000
rect 21959 15997 21971 16031
rect 21913 15991 21971 15997
rect 22465 16031 22523 16037
rect 22465 15997 22477 16031
rect 22511 16028 22523 16031
rect 22922 16028 22928 16040
rect 22511 16000 22928 16028
rect 22511 15997 22523 16000
rect 22465 15991 22523 15997
rect 22922 15988 22928 16000
rect 22980 15988 22986 16040
rect 23661 16031 23719 16037
rect 23661 15997 23673 16031
rect 23707 16028 23719 16031
rect 23750 16028 23756 16040
rect 23707 16000 23756 16028
rect 23707 15997 23719 16000
rect 23661 15991 23719 15997
rect 23750 15988 23756 16000
rect 23808 15988 23814 16040
rect 24854 16028 24860 16040
rect 23860 16000 24860 16028
rect 20254 15892 20260 15904
rect 19567 15864 20260 15892
rect 19567 15861 19579 15864
rect 19521 15855 19579 15861
rect 20254 15852 20260 15864
rect 20312 15892 20318 15904
rect 20441 15895 20499 15901
rect 20441 15892 20453 15895
rect 20312 15864 20453 15892
rect 20312 15852 20318 15864
rect 20441 15861 20453 15864
rect 20487 15861 20499 15895
rect 23474 15892 23480 15904
rect 23435 15864 23480 15892
rect 20441 15855 20499 15861
rect 23474 15852 23480 15864
rect 23532 15852 23538 15904
rect 23860 15901 23888 16000
rect 24854 15988 24860 16000
rect 24912 16037 24918 16040
rect 24912 16031 24970 16037
rect 24912 15997 24924 16031
rect 24958 16028 24970 16031
rect 25314 16028 25320 16040
rect 24958 16000 25320 16028
rect 24958 15997 24970 16000
rect 24912 15991 24970 15997
rect 24912 15988 24918 15991
rect 25314 15988 25320 16000
rect 25372 15988 25378 16040
rect 25792 16028 25820 16059
rect 26142 16056 26148 16108
rect 26200 16096 26206 16108
rect 26620 16096 26648 16136
rect 26789 16133 26801 16136
rect 26835 16133 26847 16167
rect 26789 16127 26847 16133
rect 26200 16068 26648 16096
rect 26200 16056 26206 16068
rect 26694 16056 26700 16108
rect 26752 16096 26758 16108
rect 26752 16068 26845 16096
rect 26752 16056 26758 16068
rect 26712 16028 26740 16056
rect 28184 16037 28212 16204
rect 28629 16201 28641 16204
rect 28675 16232 28687 16235
rect 28810 16232 28816 16244
rect 28675 16204 28816 16232
rect 28675 16201 28687 16204
rect 28629 16195 28687 16201
rect 28810 16192 28816 16204
rect 28868 16192 28874 16244
rect 29089 16235 29147 16241
rect 29089 16201 29101 16235
rect 29135 16232 29147 16235
rect 29270 16232 29276 16244
rect 29135 16204 29276 16232
rect 29135 16201 29147 16204
rect 29089 16195 29147 16201
rect 29270 16192 29276 16204
rect 29328 16192 29334 16244
rect 30742 16192 30748 16244
rect 30800 16232 30806 16244
rect 30837 16235 30895 16241
rect 30837 16232 30849 16235
rect 30800 16204 30849 16232
rect 30800 16192 30806 16204
rect 30837 16201 30849 16204
rect 30883 16201 30895 16235
rect 30837 16195 30895 16201
rect 33870 16192 33876 16244
rect 33928 16232 33934 16244
rect 33965 16235 34023 16241
rect 33965 16232 33977 16235
rect 33928 16204 33977 16232
rect 33928 16192 33934 16204
rect 33965 16201 33977 16204
rect 34011 16201 34023 16235
rect 33965 16195 34023 16201
rect 30561 16167 30619 16173
rect 30561 16133 30573 16167
rect 30607 16164 30619 16167
rect 31018 16164 31024 16176
rect 30607 16136 31024 16164
rect 30607 16133 30619 16136
rect 30561 16127 30619 16133
rect 31018 16124 31024 16136
rect 31076 16124 31082 16176
rect 30190 16096 30196 16108
rect 30151 16068 30196 16096
rect 30190 16056 30196 16068
rect 30248 16056 30254 16108
rect 30926 16056 30932 16108
rect 30984 16096 30990 16108
rect 32217 16099 32275 16105
rect 32217 16096 32229 16099
rect 30984 16068 32229 16096
rect 30984 16056 30990 16068
rect 32217 16065 32229 16068
rect 32263 16096 32275 16099
rect 32263 16068 33180 16096
rect 32263 16065 32275 16068
rect 32217 16059 32275 16065
rect 27341 16031 27399 16037
rect 27341 16028 27353 16031
rect 25792 16000 27353 16028
rect 27341 15997 27353 16000
rect 27387 15997 27399 16031
rect 27341 15991 27399 15997
rect 28169 16031 28227 16037
rect 28169 15997 28181 16031
rect 28215 15997 28227 16031
rect 28169 15991 28227 15997
rect 29733 16031 29791 16037
rect 29733 15997 29745 16031
rect 29779 15997 29791 16031
rect 29733 15991 29791 15997
rect 24670 15920 24676 15972
rect 24728 15960 24734 15972
rect 24765 15963 24823 15969
rect 24765 15960 24777 15963
rect 24728 15932 24777 15960
rect 24728 15920 24734 15932
rect 24765 15929 24777 15932
rect 24811 15960 24823 15963
rect 26329 15963 26387 15969
rect 26329 15960 26341 15963
rect 24811 15932 26341 15960
rect 24811 15929 24823 15932
rect 24765 15923 24823 15929
rect 26329 15929 26341 15932
rect 26375 15960 26387 15963
rect 27890 15960 27896 15972
rect 26375 15932 27896 15960
rect 26375 15929 26387 15932
rect 26329 15923 26387 15929
rect 27890 15920 27896 15932
rect 27948 15920 27954 15972
rect 29086 15920 29092 15972
rect 29144 15960 29150 15972
rect 29748 15960 29776 15991
rect 29822 15988 29828 16040
rect 29880 16028 29886 16040
rect 30285 16031 30343 16037
rect 30285 16028 30297 16031
rect 29880 16000 30297 16028
rect 29880 15988 29886 16000
rect 30285 15997 30297 16000
rect 30331 15997 30343 16031
rect 31846 16028 31852 16040
rect 31759 16000 31852 16028
rect 30285 15991 30343 15997
rect 31846 15988 31852 16000
rect 31904 16028 31910 16040
rect 33152 16037 33180 16068
rect 32861 16031 32919 16037
rect 32861 16028 32873 16031
rect 31904 16000 32873 16028
rect 31904 15988 31910 16000
rect 32861 15997 32873 16000
rect 32907 15997 32919 16031
rect 32861 15991 32919 15997
rect 33137 16031 33195 16037
rect 33137 15997 33149 16031
rect 33183 15997 33195 16031
rect 33318 16028 33324 16040
rect 33231 16000 33324 16028
rect 33137 15991 33195 15997
rect 33318 15988 33324 16000
rect 33376 16028 33382 16040
rect 33502 16028 33508 16040
rect 33376 16000 33508 16028
rect 33376 15988 33382 16000
rect 33502 15988 33508 16000
rect 33560 15988 33566 16040
rect 34882 16028 34888 16040
rect 34843 16000 34888 16028
rect 34882 15988 34888 16000
rect 34940 16028 34946 16040
rect 35345 16031 35403 16037
rect 35345 16028 35357 16031
rect 34940 16000 35357 16028
rect 34940 15988 34946 16000
rect 35345 15997 35357 16000
rect 35391 15997 35403 16031
rect 35345 15991 35403 15997
rect 31205 15963 31263 15969
rect 31205 15960 31217 15963
rect 29144 15932 31217 15960
rect 29144 15920 29150 15932
rect 31205 15929 31217 15932
rect 31251 15929 31263 15963
rect 31205 15923 31263 15929
rect 32214 15920 32220 15972
rect 32272 15960 32278 15972
rect 32309 15963 32367 15969
rect 32309 15960 32321 15963
rect 32272 15932 32321 15960
rect 32272 15920 32278 15932
rect 32309 15929 32321 15932
rect 32355 15929 32367 15963
rect 33597 15963 33655 15969
rect 33597 15960 33609 15963
rect 32309 15923 32367 15929
rect 32876 15932 33609 15960
rect 32876 15904 32904 15932
rect 33597 15929 33609 15932
rect 33643 15929 33655 15963
rect 33597 15923 33655 15929
rect 23845 15895 23903 15901
rect 23845 15861 23857 15895
rect 23891 15892 23903 15895
rect 23934 15892 23940 15904
rect 23891 15864 23940 15892
rect 23891 15861 23903 15864
rect 23845 15855 23903 15861
rect 23934 15852 23940 15864
rect 23992 15852 23998 15904
rect 24302 15892 24308 15904
rect 24263 15864 24308 15892
rect 24302 15852 24308 15864
rect 24360 15852 24366 15904
rect 26234 15892 26240 15904
rect 26195 15864 26240 15892
rect 26234 15852 26240 15864
rect 26292 15852 26298 15904
rect 28074 15892 28080 15904
rect 28035 15864 28080 15892
rect 28074 15852 28080 15864
rect 28132 15852 28138 15904
rect 28353 15895 28411 15901
rect 28353 15861 28365 15895
rect 28399 15892 28411 15895
rect 28534 15892 28540 15904
rect 28399 15864 28540 15892
rect 28399 15861 28411 15864
rect 28353 15855 28411 15861
rect 28534 15852 28540 15864
rect 28592 15852 28598 15904
rect 32858 15852 32864 15904
rect 32916 15852 32922 15904
rect 33502 15852 33508 15904
rect 33560 15892 33566 15904
rect 35069 15895 35127 15901
rect 35069 15892 35081 15895
rect 33560 15864 35081 15892
rect 33560 15852 33566 15864
rect 35069 15861 35081 15864
rect 35115 15861 35127 15895
rect 35069 15855 35127 15861
rect 1104 15802 38548 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 38548 15802
rect 1104 15728 38548 15750
rect 1670 15688 1676 15700
rect 1631 15660 1676 15688
rect 1670 15648 1676 15660
rect 1728 15648 1734 15700
rect 4433 15691 4491 15697
rect 4433 15657 4445 15691
rect 4479 15688 4491 15691
rect 4798 15688 4804 15700
rect 4479 15660 4804 15688
rect 4479 15657 4491 15660
rect 4433 15651 4491 15657
rect 4798 15648 4804 15660
rect 4856 15648 4862 15700
rect 5350 15648 5356 15700
rect 5408 15688 5414 15700
rect 5445 15691 5503 15697
rect 5445 15688 5457 15691
rect 5408 15660 5457 15688
rect 5408 15648 5414 15660
rect 5445 15657 5457 15660
rect 5491 15657 5503 15691
rect 5445 15651 5503 15657
rect 6914 15648 6920 15700
rect 6972 15688 6978 15700
rect 7377 15691 7435 15697
rect 7377 15688 7389 15691
rect 6972 15660 7389 15688
rect 6972 15648 6978 15660
rect 7377 15657 7389 15660
rect 7423 15657 7435 15691
rect 7377 15651 7435 15657
rect 7837 15691 7895 15697
rect 7837 15657 7849 15691
rect 7883 15688 7895 15691
rect 7926 15688 7932 15700
rect 7883 15660 7932 15688
rect 7883 15657 7895 15660
rect 7837 15651 7895 15657
rect 7926 15648 7932 15660
rect 7984 15648 7990 15700
rect 8294 15648 8300 15700
rect 8352 15688 8358 15700
rect 8573 15691 8631 15697
rect 8573 15688 8585 15691
rect 8352 15660 8585 15688
rect 8352 15648 8358 15660
rect 8573 15657 8585 15660
rect 8619 15657 8631 15691
rect 8573 15651 8631 15657
rect 10781 15691 10839 15697
rect 10781 15657 10793 15691
rect 10827 15688 10839 15691
rect 10870 15688 10876 15700
rect 10827 15660 10876 15688
rect 10827 15657 10839 15660
rect 10781 15651 10839 15657
rect 10870 15648 10876 15660
rect 10928 15688 10934 15700
rect 11330 15688 11336 15700
rect 10928 15660 11336 15688
rect 10928 15648 10934 15660
rect 11330 15648 11336 15660
rect 11388 15648 11394 15700
rect 12986 15688 12992 15700
rect 12947 15660 12992 15688
rect 12986 15648 12992 15660
rect 13044 15648 13050 15700
rect 16114 15688 16120 15700
rect 16075 15660 16120 15688
rect 16114 15648 16120 15660
rect 16172 15648 16178 15700
rect 16669 15691 16727 15697
rect 16669 15657 16681 15691
rect 16715 15688 16727 15691
rect 17126 15688 17132 15700
rect 16715 15660 17132 15688
rect 16715 15657 16727 15660
rect 16669 15651 16727 15657
rect 17126 15648 17132 15660
rect 17184 15648 17190 15700
rect 17770 15648 17776 15700
rect 17828 15688 17834 15700
rect 18693 15691 18751 15697
rect 18693 15688 18705 15691
rect 17828 15660 18705 15688
rect 17828 15648 17834 15660
rect 18693 15657 18705 15660
rect 18739 15688 18751 15691
rect 19150 15688 19156 15700
rect 18739 15660 19156 15688
rect 18739 15657 18751 15660
rect 18693 15651 18751 15657
rect 19150 15648 19156 15660
rect 19208 15648 19214 15700
rect 20349 15691 20407 15697
rect 20349 15657 20361 15691
rect 20395 15688 20407 15691
rect 20622 15688 20628 15700
rect 20395 15660 20628 15688
rect 20395 15657 20407 15660
rect 20349 15651 20407 15657
rect 20622 15648 20628 15660
rect 20680 15648 20686 15700
rect 20717 15691 20775 15697
rect 20717 15657 20729 15691
rect 20763 15688 20775 15691
rect 21818 15688 21824 15700
rect 20763 15660 21824 15688
rect 20763 15657 20775 15660
rect 20717 15651 20775 15657
rect 21818 15648 21824 15660
rect 21876 15648 21882 15700
rect 22005 15691 22063 15697
rect 22005 15657 22017 15691
rect 22051 15657 22063 15691
rect 22005 15651 22063 15657
rect 5534 15580 5540 15632
rect 5592 15620 5598 15632
rect 5629 15623 5687 15629
rect 5629 15620 5641 15623
rect 5592 15592 5641 15620
rect 5592 15580 5598 15592
rect 5629 15589 5641 15592
rect 5675 15589 5687 15623
rect 5629 15583 5687 15589
rect 5902 15580 5908 15632
rect 5960 15620 5966 15632
rect 11241 15623 11299 15629
rect 5960 15592 6500 15620
rect 5960 15580 5966 15592
rect 4617 15555 4675 15561
rect 4617 15521 4629 15555
rect 4663 15552 4675 15555
rect 4890 15552 4896 15564
rect 4663 15524 4896 15552
rect 4663 15521 4675 15524
rect 4617 15515 4675 15521
rect 4890 15512 4896 15524
rect 4948 15512 4954 15564
rect 5810 15512 5816 15564
rect 5868 15552 5874 15564
rect 6089 15555 6147 15561
rect 6089 15552 6101 15555
rect 5868 15524 6101 15552
rect 5868 15512 5874 15524
rect 6089 15521 6101 15524
rect 6135 15521 6147 15555
rect 6089 15515 6147 15521
rect 6178 15512 6184 15564
rect 6236 15552 6242 15564
rect 6472 15561 6500 15592
rect 11241 15589 11253 15623
rect 11287 15620 11299 15623
rect 11606 15620 11612 15632
rect 11287 15592 11376 15620
rect 11567 15592 11612 15620
rect 11287 15589 11299 15592
rect 11241 15583 11299 15589
rect 6273 15555 6331 15561
rect 6273 15552 6285 15555
rect 6236 15524 6285 15552
rect 6236 15512 6242 15524
rect 6273 15521 6285 15524
rect 6319 15521 6331 15555
rect 6273 15515 6331 15521
rect 6457 15555 6515 15561
rect 6457 15521 6469 15555
rect 6503 15521 6515 15555
rect 7098 15552 7104 15564
rect 7059 15524 7104 15552
rect 6457 15515 6515 15521
rect 7098 15512 7104 15524
rect 7156 15512 7162 15564
rect 7834 15512 7840 15564
rect 7892 15552 7898 15564
rect 7929 15555 7987 15561
rect 7929 15552 7941 15555
rect 7892 15524 7941 15552
rect 7892 15512 7898 15524
rect 7929 15521 7941 15524
rect 7975 15521 7987 15555
rect 7929 15515 7987 15521
rect 9674 15512 9680 15564
rect 9732 15552 9738 15564
rect 9732 15524 9777 15552
rect 9732 15512 9738 15524
rect 10502 15512 10508 15564
rect 10560 15552 10566 15564
rect 10686 15552 10692 15564
rect 10560 15524 10692 15552
rect 10560 15512 10566 15524
rect 10686 15512 10692 15524
rect 10744 15552 10750 15564
rect 11057 15555 11115 15561
rect 11057 15552 11069 15555
rect 10744 15524 11069 15552
rect 10744 15512 10750 15524
rect 11057 15521 11069 15524
rect 11103 15521 11115 15555
rect 11057 15515 11115 15521
rect 11146 15512 11152 15564
rect 11204 15552 11210 15564
rect 11348 15552 11376 15592
rect 11606 15580 11612 15592
rect 11664 15580 11670 15632
rect 12434 15580 12440 15632
rect 12492 15620 12498 15632
rect 12529 15623 12587 15629
rect 12529 15620 12541 15623
rect 12492 15592 12541 15620
rect 12492 15580 12498 15592
rect 12529 15589 12541 15592
rect 12575 15620 12587 15623
rect 13078 15620 13084 15632
rect 12575 15592 13084 15620
rect 12575 15589 12587 15592
rect 12529 15583 12587 15589
rect 13078 15580 13084 15592
rect 13136 15620 13142 15632
rect 16206 15620 16212 15632
rect 13136 15592 16212 15620
rect 13136 15580 13142 15592
rect 16206 15580 16212 15592
rect 16264 15620 16270 15632
rect 16485 15623 16543 15629
rect 16485 15620 16497 15623
rect 16264 15592 16497 15620
rect 16264 15580 16270 15592
rect 16485 15589 16497 15592
rect 16531 15589 16543 15623
rect 16485 15583 16543 15589
rect 16853 15623 16911 15629
rect 16853 15589 16865 15623
rect 16899 15620 16911 15623
rect 17218 15620 17224 15632
rect 16899 15592 17224 15620
rect 16899 15589 16911 15592
rect 16853 15583 16911 15589
rect 17218 15580 17224 15592
rect 17276 15620 17282 15632
rect 18138 15620 18144 15632
rect 17276 15592 18144 15620
rect 17276 15580 17282 15592
rect 18138 15580 18144 15592
rect 18196 15580 18202 15632
rect 18966 15580 18972 15632
rect 19024 15620 19030 15632
rect 19245 15623 19303 15629
rect 19245 15620 19257 15623
rect 19024 15592 19257 15620
rect 19024 15580 19030 15592
rect 19245 15589 19257 15592
rect 19291 15620 19303 15623
rect 19426 15620 19432 15632
rect 19291 15592 19432 15620
rect 19291 15589 19303 15592
rect 19245 15583 19303 15589
rect 19426 15580 19432 15592
rect 19484 15580 19490 15632
rect 20990 15580 20996 15632
rect 21048 15620 21054 15632
rect 21085 15623 21143 15629
rect 21085 15620 21097 15623
rect 21048 15592 21097 15620
rect 21048 15580 21054 15592
rect 21085 15589 21097 15592
rect 21131 15620 21143 15623
rect 21542 15620 21548 15632
rect 21131 15592 21548 15620
rect 21131 15589 21143 15592
rect 21085 15583 21143 15589
rect 21542 15580 21548 15592
rect 21600 15580 21606 15632
rect 21726 15580 21732 15632
rect 21784 15620 21790 15632
rect 22020 15620 22048 15651
rect 22278 15648 22284 15700
rect 22336 15688 22342 15700
rect 22373 15691 22431 15697
rect 22373 15688 22385 15691
rect 22336 15660 22385 15688
rect 22336 15648 22342 15660
rect 22373 15657 22385 15660
rect 22419 15688 22431 15691
rect 22738 15688 22744 15700
rect 22419 15660 22744 15688
rect 22419 15657 22431 15660
rect 22373 15651 22431 15657
rect 22738 15648 22744 15660
rect 22796 15648 22802 15700
rect 23017 15691 23075 15697
rect 23017 15657 23029 15691
rect 23063 15688 23075 15691
rect 23290 15688 23296 15700
rect 23063 15660 23296 15688
rect 23063 15657 23075 15660
rect 23017 15651 23075 15657
rect 23290 15648 23296 15660
rect 23348 15648 23354 15700
rect 24302 15648 24308 15700
rect 24360 15688 24366 15700
rect 24857 15691 24915 15697
rect 24857 15688 24869 15691
rect 24360 15660 24869 15688
rect 24360 15648 24366 15660
rect 24857 15657 24869 15660
rect 24903 15688 24915 15691
rect 25038 15688 25044 15700
rect 24903 15660 25044 15688
rect 24903 15657 24915 15660
rect 24857 15651 24915 15657
rect 25038 15648 25044 15660
rect 25096 15688 25102 15700
rect 26237 15691 26295 15697
rect 26237 15688 26249 15691
rect 25096 15660 26249 15688
rect 25096 15648 25102 15660
rect 26237 15657 26249 15660
rect 26283 15657 26295 15691
rect 26237 15651 26295 15657
rect 26970 15648 26976 15700
rect 27028 15688 27034 15700
rect 27157 15691 27215 15697
rect 27157 15688 27169 15691
rect 27028 15660 27169 15688
rect 27028 15648 27034 15660
rect 27157 15657 27169 15660
rect 27203 15657 27215 15691
rect 27890 15688 27896 15700
rect 27851 15660 27896 15688
rect 27157 15651 27215 15657
rect 27890 15648 27896 15660
rect 27948 15648 27954 15700
rect 28442 15648 28448 15700
rect 28500 15688 28506 15700
rect 28537 15691 28595 15697
rect 28537 15688 28549 15691
rect 28500 15660 28549 15688
rect 28500 15648 28506 15660
rect 28537 15657 28549 15660
rect 28583 15657 28595 15691
rect 28537 15651 28595 15657
rect 28644 15660 30236 15688
rect 28644 15632 28672 15660
rect 21784 15592 22048 15620
rect 22649 15623 22707 15629
rect 21784 15580 21790 15592
rect 22649 15589 22661 15623
rect 22695 15620 22707 15623
rect 23106 15620 23112 15632
rect 22695 15592 23112 15620
rect 22695 15589 22707 15592
rect 22649 15583 22707 15589
rect 23106 15580 23112 15592
rect 23164 15580 23170 15632
rect 23385 15623 23443 15629
rect 23385 15589 23397 15623
rect 23431 15620 23443 15623
rect 23474 15620 23480 15632
rect 23431 15592 23480 15620
rect 23431 15589 23443 15592
rect 23385 15583 23443 15589
rect 23474 15580 23480 15592
rect 23532 15620 23538 15632
rect 23845 15623 23903 15629
rect 23845 15620 23857 15623
rect 23532 15592 23857 15620
rect 23532 15580 23538 15592
rect 23845 15589 23857 15592
rect 23891 15620 23903 15623
rect 24670 15620 24676 15632
rect 23891 15592 24676 15620
rect 23891 15589 23903 15592
rect 23845 15583 23903 15589
rect 24670 15580 24676 15592
rect 24728 15580 24734 15632
rect 25958 15620 25964 15632
rect 25919 15592 25964 15620
rect 25958 15580 25964 15592
rect 26016 15620 26022 15632
rect 26513 15623 26571 15629
rect 26513 15620 26525 15623
rect 26016 15592 26525 15620
rect 26016 15580 26022 15592
rect 26513 15589 26525 15592
rect 26559 15589 26571 15623
rect 28626 15620 28632 15632
rect 28539 15592 28632 15620
rect 26513 15583 26571 15589
rect 28626 15580 28632 15592
rect 28684 15580 28690 15632
rect 28997 15623 29055 15629
rect 28997 15589 29009 15623
rect 29043 15620 29055 15623
rect 29086 15620 29092 15632
rect 29043 15592 29092 15620
rect 29043 15589 29055 15592
rect 28997 15583 29055 15589
rect 29086 15580 29092 15592
rect 29144 15580 29150 15632
rect 29362 15620 29368 15632
rect 29323 15592 29368 15620
rect 29362 15580 29368 15592
rect 29420 15580 29426 15632
rect 30208 15629 30236 15660
rect 30466 15648 30472 15700
rect 30524 15688 30530 15700
rect 31205 15691 31263 15697
rect 31205 15688 31217 15691
rect 30524 15660 31217 15688
rect 30524 15648 30530 15660
rect 31205 15657 31217 15660
rect 31251 15657 31263 15691
rect 31205 15651 31263 15657
rect 31754 15648 31760 15700
rect 31812 15688 31818 15700
rect 32217 15691 32275 15697
rect 32217 15688 32229 15691
rect 31812 15660 32229 15688
rect 31812 15648 31818 15660
rect 32217 15657 32229 15660
rect 32263 15657 32275 15691
rect 32217 15651 32275 15657
rect 33229 15691 33287 15697
rect 33229 15657 33241 15691
rect 33275 15688 33287 15691
rect 33686 15688 33692 15700
rect 33275 15660 33692 15688
rect 33275 15657 33287 15660
rect 33229 15651 33287 15657
rect 33686 15648 33692 15660
rect 33744 15648 33750 15700
rect 30193 15623 30251 15629
rect 30193 15589 30205 15623
rect 30239 15620 30251 15623
rect 30282 15620 30288 15632
rect 30239 15592 30288 15620
rect 30239 15589 30251 15592
rect 30193 15583 30251 15589
rect 30282 15580 30288 15592
rect 30340 15580 30346 15632
rect 11790 15552 11796 15564
rect 11204 15524 11249 15552
rect 11348 15524 11796 15552
rect 11204 15512 11210 15524
rect 11790 15512 11796 15524
rect 11848 15552 11854 15564
rect 12250 15552 12256 15564
rect 11848 15524 12256 15552
rect 11848 15512 11854 15524
rect 12250 15512 12256 15524
rect 12308 15512 12314 15564
rect 13170 15552 13176 15564
rect 13131 15524 13176 15552
rect 13170 15512 13176 15524
rect 13228 15512 13234 15564
rect 13630 15552 13636 15564
rect 13591 15524 13636 15552
rect 13630 15512 13636 15524
rect 13688 15512 13694 15564
rect 13725 15555 13783 15561
rect 13725 15521 13737 15555
rect 13771 15521 13783 15555
rect 13725 15515 13783 15521
rect 14277 15555 14335 15561
rect 14277 15521 14289 15555
rect 14323 15552 14335 15555
rect 14734 15552 14740 15564
rect 14323 15524 14740 15552
rect 14323 15521 14335 15524
rect 14277 15515 14335 15521
rect 3234 15444 3240 15496
rect 3292 15484 3298 15496
rect 3513 15487 3571 15493
rect 3513 15484 3525 15487
rect 3292 15456 3525 15484
rect 3292 15444 3298 15456
rect 3513 15453 3525 15456
rect 3559 15484 3571 15487
rect 5074 15484 5080 15496
rect 3559 15456 5080 15484
rect 3559 15453 3571 15456
rect 3513 15447 3571 15453
rect 5074 15444 5080 15456
rect 5132 15444 5138 15496
rect 5718 15444 5724 15496
rect 5776 15484 5782 15496
rect 6733 15487 6791 15493
rect 6733 15484 6745 15487
rect 5776 15456 6745 15484
rect 5776 15444 5782 15456
rect 6733 15453 6745 15456
rect 6779 15453 6791 15487
rect 8294 15484 8300 15496
rect 8255 15456 8300 15484
rect 6733 15447 6791 15453
rect 8294 15444 8300 15456
rect 8352 15444 8358 15496
rect 10870 15484 10876 15496
rect 10831 15456 10876 15484
rect 10870 15444 10876 15456
rect 10928 15444 10934 15496
rect 13740 15484 13768 15515
rect 14734 15512 14740 15524
rect 14792 15512 14798 15564
rect 15286 15552 15292 15564
rect 15247 15524 15292 15552
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 16758 15512 16764 15564
rect 16816 15552 16822 15564
rect 16816 15524 16861 15552
rect 16816 15512 16822 15524
rect 18046 15512 18052 15564
rect 18104 15552 18110 15564
rect 19061 15555 19119 15561
rect 19061 15552 19073 15555
rect 18104 15524 19073 15552
rect 18104 15512 18110 15524
rect 19061 15521 19073 15524
rect 19107 15521 19119 15555
rect 21818 15552 21824 15564
rect 21779 15524 21824 15552
rect 19061 15515 19119 15521
rect 21818 15512 21824 15524
rect 21876 15512 21882 15564
rect 22833 15555 22891 15561
rect 22833 15521 22845 15555
rect 22879 15521 22891 15555
rect 22833 15515 22891 15521
rect 12912 15456 13768 15484
rect 3145 15419 3203 15425
rect 3145 15385 3157 15419
rect 3191 15416 3203 15419
rect 4706 15416 4712 15428
rect 3191 15388 4712 15416
rect 3191 15385 3203 15388
rect 3145 15379 3203 15385
rect 4706 15376 4712 15388
rect 4764 15376 4770 15428
rect 4801 15419 4859 15425
rect 4801 15385 4813 15419
rect 4847 15416 4859 15419
rect 5442 15416 5448 15428
rect 4847 15388 5448 15416
rect 4847 15385 4859 15388
rect 4801 15379 4859 15385
rect 5442 15376 5448 15388
rect 5500 15376 5506 15428
rect 6822 15376 6828 15428
rect 6880 15416 6886 15428
rect 8205 15419 8263 15425
rect 8205 15416 8217 15419
rect 6880 15388 8217 15416
rect 6880 15376 6886 15388
rect 8205 15385 8217 15388
rect 8251 15385 8263 15419
rect 9861 15419 9919 15425
rect 9861 15416 9873 15419
rect 8205 15379 8263 15385
rect 8956 15388 9873 15416
rect 8956 15360 8984 15388
rect 9861 15385 9873 15388
rect 9907 15385 9919 15419
rect 9861 15379 9919 15385
rect 12912 15360 12940 15456
rect 16666 15444 16672 15496
rect 16724 15484 16730 15496
rect 17221 15487 17279 15493
rect 17221 15484 17233 15487
rect 16724 15456 17233 15484
rect 16724 15444 16730 15456
rect 17221 15453 17233 15456
rect 17267 15453 17279 15487
rect 17221 15447 17279 15453
rect 18598 15444 18604 15496
rect 18656 15484 18662 15496
rect 18877 15487 18935 15493
rect 18877 15484 18889 15487
rect 18656 15456 18889 15484
rect 18656 15444 18662 15456
rect 18877 15453 18889 15456
rect 18923 15453 18935 15487
rect 18877 15447 18935 15453
rect 19334 15444 19340 15496
rect 19392 15484 19398 15496
rect 19613 15487 19671 15493
rect 19613 15484 19625 15487
rect 19392 15456 19625 15484
rect 19392 15444 19398 15456
rect 19613 15453 19625 15456
rect 19659 15453 19671 15487
rect 19613 15447 19671 15453
rect 15194 15376 15200 15428
rect 15252 15416 15258 15428
rect 15473 15419 15531 15425
rect 15473 15416 15485 15419
rect 15252 15388 15485 15416
rect 15252 15376 15258 15388
rect 15473 15385 15485 15388
rect 15519 15385 15531 15419
rect 15473 15379 15531 15385
rect 17773 15419 17831 15425
rect 17773 15385 17785 15419
rect 17819 15416 17831 15419
rect 17954 15416 17960 15428
rect 17819 15388 17960 15416
rect 17819 15385 17831 15388
rect 17773 15379 17831 15385
rect 17954 15376 17960 15388
rect 18012 15376 18018 15428
rect 21729 15419 21787 15425
rect 21729 15385 21741 15419
rect 21775 15416 21787 15419
rect 22554 15416 22560 15428
rect 21775 15388 22560 15416
rect 21775 15385 21787 15388
rect 21729 15379 21787 15385
rect 22554 15376 22560 15388
rect 22612 15376 22618 15428
rect 22738 15376 22744 15428
rect 22796 15416 22802 15428
rect 22848 15416 22876 15515
rect 23934 15512 23940 15564
rect 23992 15561 23998 15564
rect 23992 15555 24050 15561
rect 23992 15521 24004 15555
rect 24038 15521 24050 15555
rect 23992 15515 24050 15521
rect 25409 15555 25467 15561
rect 25409 15521 25421 15555
rect 25455 15552 25467 15555
rect 25498 15552 25504 15564
rect 25455 15524 25504 15552
rect 25455 15521 25467 15524
rect 25409 15515 25467 15521
rect 23992 15512 23998 15515
rect 25498 15512 25504 15524
rect 25556 15512 25562 15564
rect 26326 15512 26332 15564
rect 26384 15552 26390 15564
rect 26660 15555 26718 15561
rect 26660 15552 26672 15555
rect 26384 15524 26672 15552
rect 26384 15512 26390 15524
rect 26660 15521 26672 15524
rect 26706 15521 26718 15555
rect 26660 15515 26718 15521
rect 28350 15512 28356 15564
rect 28408 15552 28414 15564
rect 28445 15555 28503 15561
rect 28445 15552 28457 15555
rect 28408 15524 28457 15552
rect 28408 15512 28414 15524
rect 28445 15521 28457 15524
rect 28491 15552 28503 15555
rect 29454 15552 29460 15564
rect 28491 15524 29460 15552
rect 28491 15521 28503 15524
rect 28445 15515 28503 15521
rect 29454 15512 29460 15524
rect 29512 15512 29518 15564
rect 30006 15552 30012 15564
rect 29967 15524 30012 15552
rect 30006 15512 30012 15524
rect 30064 15512 30070 15564
rect 30101 15555 30159 15561
rect 30101 15521 30113 15555
rect 30147 15521 30159 15555
rect 30101 15515 30159 15521
rect 23290 15444 23296 15496
rect 23348 15484 23354 15496
rect 23952 15484 23980 15512
rect 23348 15456 23980 15484
rect 24213 15487 24271 15493
rect 23348 15444 23354 15456
rect 24213 15453 24225 15487
rect 24259 15484 24271 15487
rect 24394 15484 24400 15496
rect 24259 15456 24400 15484
rect 24259 15453 24271 15456
rect 24213 15447 24271 15453
rect 24394 15444 24400 15456
rect 24452 15444 24458 15496
rect 25314 15484 25320 15496
rect 25227 15456 25320 15484
rect 25314 15444 25320 15456
rect 25372 15484 25378 15496
rect 26050 15484 26056 15496
rect 25372 15456 26056 15484
rect 25372 15444 25378 15456
rect 26050 15444 26056 15456
rect 26108 15444 26114 15496
rect 26786 15444 26792 15496
rect 26844 15484 26850 15496
rect 26881 15487 26939 15493
rect 26881 15484 26893 15487
rect 26844 15456 26893 15484
rect 26844 15444 26850 15456
rect 26881 15453 26893 15456
rect 26927 15484 26939 15487
rect 27338 15484 27344 15496
rect 26927 15456 27344 15484
rect 26927 15453 26939 15456
rect 26881 15447 26939 15453
rect 27338 15444 27344 15456
rect 27396 15444 27402 15496
rect 27614 15444 27620 15496
rect 27672 15444 27678 15496
rect 28261 15487 28319 15493
rect 28261 15453 28273 15487
rect 28307 15453 28319 15487
rect 28261 15447 28319 15453
rect 24305 15419 24363 15425
rect 24305 15416 24317 15419
rect 22796 15388 24317 15416
rect 22796 15376 22802 15388
rect 24305 15385 24317 15388
rect 24351 15385 24363 15419
rect 24305 15379 24363 15385
rect 25593 15419 25651 15425
rect 25593 15385 25605 15419
rect 25639 15416 25651 15419
rect 27632 15416 27660 15444
rect 27890 15416 27896 15428
rect 25639 15388 27896 15416
rect 25639 15385 25651 15388
rect 25593 15379 25651 15385
rect 27890 15376 27896 15388
rect 27948 15416 27954 15428
rect 28276 15416 28304 15447
rect 29270 15444 29276 15496
rect 29328 15484 29334 15496
rect 29825 15487 29883 15493
rect 29825 15484 29837 15487
rect 29328 15456 29837 15484
rect 29328 15444 29334 15456
rect 29825 15453 29837 15456
rect 29871 15453 29883 15487
rect 30116 15484 30144 15515
rect 31938 15512 31944 15564
rect 31996 15552 32002 15564
rect 32125 15555 32183 15561
rect 32125 15552 32137 15555
rect 31996 15524 32137 15552
rect 31996 15512 32002 15524
rect 32125 15521 32137 15524
rect 32171 15521 32183 15555
rect 32125 15515 32183 15521
rect 32214 15512 32220 15564
rect 32272 15552 32278 15564
rect 32398 15552 32404 15564
rect 32272 15524 32404 15552
rect 32272 15512 32278 15524
rect 32398 15512 32404 15524
rect 32456 15512 32462 15564
rect 32490 15512 32496 15564
rect 32548 15552 32554 15564
rect 32585 15555 32643 15561
rect 32585 15552 32597 15555
rect 32548 15524 32597 15552
rect 32548 15512 32554 15524
rect 32585 15521 32597 15524
rect 32631 15552 32643 15555
rect 33134 15552 33140 15564
rect 32631 15524 33140 15552
rect 32631 15521 32643 15524
rect 32585 15515 32643 15521
rect 33134 15512 33140 15524
rect 33192 15512 33198 15564
rect 34422 15552 34428 15564
rect 34383 15524 34428 15552
rect 34422 15512 34428 15524
rect 34480 15512 34486 15564
rect 34790 15552 34796 15564
rect 34751 15524 34796 15552
rect 34790 15512 34796 15524
rect 34848 15512 34854 15564
rect 30558 15484 30564 15496
rect 29825 15447 29883 15453
rect 30024 15456 30144 15484
rect 30471 15456 30564 15484
rect 27948 15388 28304 15416
rect 27948 15376 27954 15388
rect 28442 15376 28448 15428
rect 28500 15416 28506 15428
rect 29914 15416 29920 15428
rect 28500 15388 29920 15416
rect 28500 15376 28506 15388
rect 29914 15376 29920 15388
rect 29972 15416 29978 15428
rect 30024 15416 30052 15456
rect 30558 15444 30564 15456
rect 30616 15484 30622 15496
rect 30837 15487 30895 15493
rect 30837 15484 30849 15487
rect 30616 15456 30849 15484
rect 30616 15444 30622 15456
rect 30837 15453 30849 15456
rect 30883 15453 30895 15487
rect 30837 15447 30895 15453
rect 34149 15487 34207 15493
rect 34149 15453 34161 15487
rect 34195 15484 34207 15487
rect 34330 15484 34336 15496
rect 34195 15456 34336 15484
rect 34195 15453 34207 15456
rect 34149 15447 34207 15453
rect 34330 15444 34336 15456
rect 34388 15444 34394 15496
rect 34790 15416 34796 15428
rect 29972 15388 30052 15416
rect 34751 15388 34796 15416
rect 29972 15376 29978 15388
rect 34790 15376 34796 15388
rect 34848 15376 34854 15428
rect 3881 15351 3939 15357
rect 3881 15317 3893 15351
rect 3927 15348 3939 15351
rect 4982 15348 4988 15360
rect 3927 15320 4988 15348
rect 3927 15317 3939 15320
rect 3881 15311 3939 15317
rect 4982 15308 4988 15320
rect 5040 15308 5046 15360
rect 5169 15351 5227 15357
rect 5169 15317 5181 15351
rect 5215 15348 5227 15351
rect 6270 15348 6276 15360
rect 5215 15320 6276 15348
rect 5215 15317 5227 15320
rect 5169 15311 5227 15317
rect 6270 15308 6276 15320
rect 6328 15308 6334 15360
rect 8018 15308 8024 15360
rect 8076 15357 8082 15360
rect 8076 15351 8125 15357
rect 8076 15317 8079 15351
rect 8113 15317 8125 15351
rect 8938 15348 8944 15360
rect 8899 15320 8944 15348
rect 8076 15311 8125 15317
rect 8076 15308 8082 15311
rect 8938 15308 8944 15320
rect 8996 15308 9002 15360
rect 9214 15308 9220 15360
rect 9272 15348 9278 15360
rect 9309 15351 9367 15357
rect 9309 15348 9321 15351
rect 9272 15320 9321 15348
rect 9272 15308 9278 15320
rect 9309 15317 9321 15320
rect 9355 15317 9367 15351
rect 9309 15311 9367 15317
rect 9950 15308 9956 15360
rect 10008 15348 10014 15360
rect 10229 15351 10287 15357
rect 10229 15348 10241 15351
rect 10008 15320 10241 15348
rect 10008 15308 10014 15320
rect 10229 15317 10241 15320
rect 10275 15348 10287 15351
rect 10502 15348 10508 15360
rect 10275 15320 10508 15348
rect 10275 15317 10287 15320
rect 10229 15311 10287 15317
rect 10502 15308 10508 15320
rect 10560 15308 10566 15360
rect 12161 15351 12219 15357
rect 12161 15317 12173 15351
rect 12207 15348 12219 15351
rect 12894 15348 12900 15360
rect 12207 15320 12900 15348
rect 12207 15317 12219 15320
rect 12161 15311 12219 15317
rect 12894 15308 12900 15320
rect 12952 15308 12958 15360
rect 14734 15348 14740 15360
rect 14695 15320 14740 15348
rect 14734 15308 14740 15320
rect 14792 15308 14798 15360
rect 15102 15348 15108 15360
rect 15063 15320 15108 15348
rect 15102 15308 15108 15320
rect 15160 15308 15166 15360
rect 18046 15348 18052 15360
rect 18007 15320 18052 15348
rect 18046 15308 18052 15320
rect 18104 15308 18110 15360
rect 19150 15308 19156 15360
rect 19208 15348 19214 15360
rect 19889 15351 19947 15357
rect 19889 15348 19901 15351
rect 19208 15320 19901 15348
rect 19208 15308 19214 15320
rect 19889 15317 19901 15320
rect 19935 15317 19947 15351
rect 19889 15311 19947 15317
rect 23753 15351 23811 15357
rect 23753 15317 23765 15351
rect 23799 15348 23811 15351
rect 23842 15348 23848 15360
rect 23799 15320 23848 15348
rect 23799 15317 23811 15320
rect 23753 15311 23811 15317
rect 23842 15308 23848 15320
rect 23900 15308 23906 15360
rect 24121 15351 24179 15357
rect 24121 15317 24133 15351
rect 24167 15348 24179 15351
rect 24210 15348 24216 15360
rect 24167 15320 24216 15348
rect 24167 15317 24179 15320
rect 24121 15311 24179 15317
rect 24210 15308 24216 15320
rect 24268 15308 24274 15360
rect 26786 15348 26792 15360
rect 26747 15320 26792 15348
rect 26786 15308 26792 15320
rect 26844 15308 26850 15360
rect 27430 15308 27436 15360
rect 27488 15348 27494 15360
rect 27617 15351 27675 15357
rect 27617 15348 27629 15351
rect 27488 15320 27629 15348
rect 27488 15308 27494 15320
rect 27617 15317 27629 15320
rect 27663 15317 27675 15351
rect 27617 15311 27675 15317
rect 29733 15351 29791 15357
rect 29733 15317 29745 15351
rect 29779 15348 29791 15351
rect 30190 15348 30196 15360
rect 29779 15320 30196 15348
rect 29779 15317 29791 15320
rect 29733 15311 29791 15317
rect 30190 15308 30196 15320
rect 30248 15308 30254 15360
rect 1104 15258 38548 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 38548 15258
rect 1104 15184 38548 15206
rect 2866 15104 2872 15156
rect 2924 15144 2930 15156
rect 2961 15147 3019 15153
rect 2961 15144 2973 15147
rect 2924 15116 2973 15144
rect 2924 15104 2930 15116
rect 2961 15113 2973 15116
rect 3007 15113 3019 15147
rect 2961 15107 3019 15113
rect 5721 15147 5779 15153
rect 5721 15113 5733 15147
rect 5767 15144 5779 15147
rect 5810 15144 5816 15156
rect 5767 15116 5816 15144
rect 5767 15113 5779 15116
rect 5721 15107 5779 15113
rect 5810 15104 5816 15116
rect 5868 15104 5874 15156
rect 8478 15144 8484 15156
rect 8439 15116 8484 15144
rect 8478 15104 8484 15116
rect 8536 15104 8542 15156
rect 10962 15153 10968 15156
rect 10946 15147 10968 15153
rect 10946 15113 10958 15147
rect 10946 15107 10968 15113
rect 10962 15104 10968 15107
rect 11020 15104 11026 15156
rect 11054 15104 11060 15156
rect 11112 15144 11118 15156
rect 11112 15116 11157 15144
rect 11112 15104 11118 15116
rect 11330 15104 11336 15156
rect 11388 15144 11394 15156
rect 11793 15147 11851 15153
rect 11793 15144 11805 15147
rect 11388 15116 11805 15144
rect 11388 15104 11394 15116
rect 11793 15113 11805 15116
rect 11839 15113 11851 15147
rect 11793 15107 11851 15113
rect 7650 15076 7656 15088
rect 7611 15048 7656 15076
rect 7650 15036 7656 15048
rect 7708 15076 7714 15088
rect 8386 15076 8392 15088
rect 7708 15048 8392 15076
rect 7708 15036 7714 15048
rect 8386 15036 8392 15048
rect 8444 15036 8450 15088
rect 9674 15036 9680 15088
rect 9732 15076 9738 15088
rect 9953 15079 10011 15085
rect 9953 15076 9965 15079
rect 9732 15048 9965 15076
rect 9732 15036 9738 15048
rect 9953 15045 9965 15048
rect 9999 15045 10011 15079
rect 11238 15076 11244 15088
rect 11199 15048 11244 15076
rect 9953 15039 10011 15045
rect 1394 15008 1400 15020
rect 1355 14980 1400 15008
rect 1394 14968 1400 14980
rect 1452 14968 1458 15020
rect 1578 14968 1584 15020
rect 1636 15008 1642 15020
rect 1673 15011 1731 15017
rect 1673 15008 1685 15011
rect 1636 14980 1685 15008
rect 1636 14968 1642 14980
rect 1673 14977 1685 14980
rect 1719 14977 1731 15011
rect 1673 14971 1731 14977
rect 2866 14968 2872 15020
rect 2924 15008 2930 15020
rect 3418 15008 3424 15020
rect 2924 14980 3424 15008
rect 2924 14968 2930 14980
rect 3418 14968 3424 14980
rect 3476 14968 3482 15020
rect 4706 14968 4712 15020
rect 4764 15008 4770 15020
rect 4764 14980 4936 15008
rect 4764 14968 4770 14980
rect 3789 14943 3847 14949
rect 3789 14909 3801 14943
rect 3835 14940 3847 14943
rect 4338 14940 4344 14952
rect 3835 14912 4344 14940
rect 3835 14909 3847 14912
rect 3789 14903 3847 14909
rect 4338 14900 4344 14912
rect 4396 14900 4402 14952
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14940 4583 14943
rect 4798 14940 4804 14952
rect 4571 14912 4804 14940
rect 4571 14909 4583 14912
rect 4525 14903 4583 14909
rect 4798 14900 4804 14912
rect 4856 14900 4862 14952
rect 4908 14949 4936 14980
rect 7190 14968 7196 15020
rect 7248 15008 7254 15020
rect 7745 15011 7803 15017
rect 7745 15008 7757 15011
rect 7248 14980 7757 15008
rect 7248 14968 7254 14980
rect 7745 14977 7757 14980
rect 7791 14977 7803 15011
rect 7745 14971 7803 14977
rect 7834 14968 7840 15020
rect 7892 15008 7898 15020
rect 8849 15011 8907 15017
rect 7892 14980 7937 15008
rect 7892 14968 7898 14980
rect 8849 14977 8861 15011
rect 8895 15008 8907 15011
rect 9398 15008 9404 15020
rect 8895 14980 9404 15008
rect 8895 14977 8907 14980
rect 8849 14971 8907 14977
rect 9398 14968 9404 14980
rect 9456 14968 9462 15020
rect 9968 15008 9996 15039
rect 11238 15036 11244 15048
rect 11296 15036 11302 15088
rect 11149 15011 11207 15017
rect 9968 14980 11100 15008
rect 4893 14943 4951 14949
rect 4893 14909 4905 14943
rect 4939 14909 4951 14943
rect 5074 14940 5080 14952
rect 4987 14912 5080 14940
rect 4893 14903 4951 14909
rect 5074 14900 5080 14912
rect 5132 14940 5138 14952
rect 7098 14940 7104 14952
rect 5132 14912 7104 14940
rect 5132 14900 5138 14912
rect 7098 14900 7104 14912
rect 7156 14900 7162 14952
rect 7466 14900 7472 14952
rect 7524 14949 7530 14952
rect 7524 14943 7582 14949
rect 7524 14909 7536 14943
rect 7570 14940 7582 14943
rect 9677 14943 9735 14949
rect 9677 14940 9689 14943
rect 7570 14912 9689 14940
rect 7570 14909 7582 14912
rect 7524 14903 7582 14909
rect 9677 14909 9689 14912
rect 9723 14909 9735 14943
rect 10778 14940 10784 14952
rect 10739 14912 10784 14940
rect 9677 14903 9735 14909
rect 7524 14900 7530 14903
rect 10778 14900 10784 14912
rect 10836 14900 10842 14952
rect 11072 14940 11100 14980
rect 11149 14977 11161 15011
rect 11195 15008 11207 15011
rect 11514 15008 11520 15020
rect 11195 14980 11520 15008
rect 11195 14977 11207 14980
rect 11149 14971 11207 14977
rect 11514 14968 11520 14980
rect 11572 14968 11578 15020
rect 11808 14952 11836 15107
rect 13170 15104 13176 15156
rect 13228 15144 13234 15156
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 13228 15116 13461 15144
rect 13228 15104 13234 15116
rect 13449 15113 13461 15116
rect 13495 15113 13507 15147
rect 13449 15107 13507 15113
rect 13630 15104 13636 15156
rect 13688 15144 13694 15156
rect 13817 15147 13875 15153
rect 13817 15144 13829 15147
rect 13688 15116 13829 15144
rect 13688 15104 13694 15116
rect 13817 15113 13829 15116
rect 13863 15113 13875 15147
rect 13817 15107 13875 15113
rect 14369 15147 14427 15153
rect 14369 15113 14381 15147
rect 14415 15144 14427 15147
rect 15286 15144 15292 15156
rect 14415 15116 15292 15144
rect 14415 15113 14427 15116
rect 14369 15107 14427 15113
rect 15286 15104 15292 15116
rect 15344 15104 15350 15156
rect 16206 15104 16212 15156
rect 16264 15144 16270 15156
rect 16577 15147 16635 15153
rect 16577 15144 16589 15147
rect 16264 15116 16589 15144
rect 16264 15104 16270 15116
rect 16577 15113 16589 15116
rect 16623 15113 16635 15147
rect 16577 15107 16635 15113
rect 16758 15104 16764 15156
rect 16816 15144 16822 15156
rect 17589 15147 17647 15153
rect 17589 15144 17601 15147
rect 16816 15116 17601 15144
rect 16816 15104 16822 15116
rect 17589 15113 17601 15116
rect 17635 15144 17647 15147
rect 17770 15144 17776 15156
rect 17635 15116 17776 15144
rect 17635 15113 17647 15116
rect 17589 15107 17647 15113
rect 17770 15104 17776 15116
rect 17828 15104 17834 15156
rect 17954 15104 17960 15156
rect 18012 15144 18018 15156
rect 18601 15147 18659 15153
rect 18601 15144 18613 15147
rect 18012 15116 18613 15144
rect 18012 15104 18018 15116
rect 18601 15113 18613 15116
rect 18647 15144 18659 15147
rect 19242 15144 19248 15156
rect 18647 15116 19248 15144
rect 18647 15113 18659 15116
rect 18601 15107 18659 15113
rect 19242 15104 19248 15116
rect 19300 15104 19306 15156
rect 21177 15147 21235 15153
rect 21177 15113 21189 15147
rect 21223 15144 21235 15147
rect 21818 15144 21824 15156
rect 21223 15116 21824 15144
rect 21223 15113 21235 15116
rect 21177 15107 21235 15113
rect 21818 15104 21824 15116
rect 21876 15104 21882 15156
rect 23109 15147 23167 15153
rect 23109 15113 23121 15147
rect 23155 15144 23167 15147
rect 23290 15144 23296 15156
rect 23155 15116 23296 15144
rect 23155 15113 23167 15116
rect 23109 15107 23167 15113
rect 23290 15104 23296 15116
rect 23348 15104 23354 15156
rect 23477 15147 23535 15153
rect 23477 15113 23489 15147
rect 23523 15144 23535 15147
rect 24302 15144 24308 15156
rect 23523 15116 24308 15144
rect 23523 15113 23535 15116
rect 23477 15107 23535 15113
rect 24302 15104 24308 15116
rect 24360 15104 24366 15156
rect 24486 15144 24492 15156
rect 24447 15116 24492 15144
rect 24486 15104 24492 15116
rect 24544 15104 24550 15156
rect 26050 15104 26056 15156
rect 26108 15153 26114 15156
rect 26108 15147 26157 15153
rect 26108 15113 26111 15147
rect 26145 15113 26157 15147
rect 26108 15107 26157 15113
rect 26108 15104 26114 15107
rect 26326 15104 26332 15156
rect 26384 15144 26390 15156
rect 27062 15144 27068 15156
rect 26384 15116 27068 15144
rect 26384 15104 26390 15116
rect 27062 15104 27068 15116
rect 27120 15144 27126 15156
rect 27341 15147 27399 15153
rect 27341 15144 27353 15147
rect 27120 15116 27353 15144
rect 27120 15104 27126 15116
rect 27341 15113 27353 15116
rect 27387 15144 27399 15147
rect 28261 15147 28319 15153
rect 28261 15144 28273 15147
rect 27387 15116 28273 15144
rect 27387 15113 27399 15116
rect 27341 15107 27399 15113
rect 28261 15113 28273 15116
rect 28307 15144 28319 15147
rect 28442 15144 28448 15156
rect 28307 15116 28448 15144
rect 28307 15113 28319 15116
rect 28261 15107 28319 15113
rect 28442 15104 28448 15116
rect 28500 15104 28506 15156
rect 28626 15144 28632 15156
rect 28587 15116 28632 15144
rect 28626 15104 28632 15116
rect 28684 15104 28690 15156
rect 29270 15104 29276 15156
rect 29328 15144 29334 15156
rect 29457 15147 29515 15153
rect 29457 15144 29469 15147
rect 29328 15116 29469 15144
rect 29328 15104 29334 15116
rect 29457 15113 29469 15116
rect 29503 15113 29515 15147
rect 29457 15107 29515 15113
rect 30745 15147 30803 15153
rect 30745 15113 30757 15147
rect 30791 15144 30803 15147
rect 31846 15144 31852 15156
rect 30791 15116 31852 15144
rect 30791 15113 30803 15116
rect 30745 15107 30803 15113
rect 31846 15104 31852 15116
rect 31904 15104 31910 15156
rect 31938 15104 31944 15156
rect 31996 15144 32002 15156
rect 32401 15147 32459 15153
rect 31996 15116 32041 15144
rect 31996 15104 32002 15116
rect 32401 15113 32413 15147
rect 32447 15144 32459 15147
rect 32582 15144 32588 15156
rect 32447 15116 32588 15144
rect 32447 15113 32459 15116
rect 32401 15107 32459 15113
rect 32582 15104 32588 15116
rect 32640 15104 32646 15156
rect 33134 15104 33140 15156
rect 33192 15144 33198 15156
rect 33781 15147 33839 15153
rect 33781 15144 33793 15147
rect 33192 15116 33793 15144
rect 33192 15104 33198 15116
rect 33781 15113 33793 15116
rect 33827 15113 33839 15147
rect 33781 15107 33839 15113
rect 34241 15147 34299 15153
rect 34241 15113 34253 15147
rect 34287 15144 34299 15147
rect 34330 15144 34336 15156
rect 34287 15116 34336 15144
rect 34287 15113 34299 15116
rect 34241 15107 34299 15113
rect 34330 15104 34336 15116
rect 34388 15104 34394 15156
rect 34609 15147 34667 15153
rect 34609 15113 34621 15147
rect 34655 15144 34667 15147
rect 34698 15144 34704 15156
rect 34655 15116 34704 15144
rect 34655 15113 34667 15116
rect 34609 15107 34667 15113
rect 34698 15104 34704 15116
rect 34756 15104 34762 15156
rect 12342 15036 12348 15088
rect 12400 15076 12406 15088
rect 16022 15076 16028 15088
rect 12400 15048 16028 15076
rect 12400 15036 12406 15048
rect 16022 15036 16028 15048
rect 16080 15076 16086 15088
rect 18322 15076 18328 15088
rect 16080 15048 18328 15076
rect 16080 15036 16086 15048
rect 18322 15036 18328 15048
rect 18380 15036 18386 15088
rect 19886 15076 19892 15088
rect 18616 15048 19892 15076
rect 12069 15011 12127 15017
rect 12069 14977 12081 15011
rect 12115 15008 12127 15011
rect 12437 15011 12495 15017
rect 12437 15008 12449 15011
rect 12115 14980 12449 15008
rect 12115 14977 12127 14980
rect 12069 14971 12127 14977
rect 12437 14977 12449 14980
rect 12483 14977 12495 15011
rect 12437 14971 12495 14977
rect 12894 14968 12900 15020
rect 12952 15008 12958 15020
rect 13173 15011 13231 15017
rect 13173 15008 13185 15011
rect 12952 14980 13185 15008
rect 12952 14968 12958 14980
rect 13173 14977 13185 14980
rect 13219 14977 13231 15011
rect 13173 14971 13231 14977
rect 14553 15011 14611 15017
rect 14553 14977 14565 15011
rect 14599 14977 14611 15011
rect 16574 15008 16580 15020
rect 14553 14971 14611 14977
rect 15212 14980 16580 15008
rect 11609 14943 11667 14949
rect 11609 14940 11621 14943
rect 11072 14912 11621 14940
rect 11609 14909 11621 14912
rect 11655 14909 11667 14943
rect 11790 14940 11796 14952
rect 11703 14912 11796 14940
rect 11609 14903 11667 14909
rect 11790 14900 11796 14912
rect 11848 14940 11854 14952
rect 12713 14943 12771 14949
rect 12713 14940 12725 14943
rect 11848 14912 12725 14940
rect 11848 14900 11854 14912
rect 12713 14909 12725 14912
rect 12759 14909 12771 14943
rect 12713 14903 12771 14909
rect 13998 14900 14004 14952
rect 14056 14940 14062 14952
rect 14461 14943 14519 14949
rect 14461 14940 14473 14943
rect 14056 14912 14473 14940
rect 14056 14900 14062 14912
rect 14461 14909 14473 14912
rect 14507 14909 14519 14943
rect 14461 14903 14519 14909
rect 7374 14872 7380 14884
rect 7335 14844 7380 14872
rect 7374 14832 7380 14844
rect 7432 14832 7438 14884
rect 7926 14832 7932 14884
rect 7984 14872 7990 14884
rect 8938 14872 8944 14884
rect 7984 14844 8944 14872
rect 7984 14832 7990 14844
rect 8938 14832 8944 14844
rect 8996 14832 9002 14884
rect 9309 14875 9367 14881
rect 9309 14841 9321 14875
rect 9355 14872 9367 14875
rect 9582 14872 9588 14884
rect 9355 14844 9588 14872
rect 9355 14841 9367 14844
rect 9309 14835 9367 14841
rect 9582 14832 9588 14844
rect 9640 14872 9646 14884
rect 9858 14872 9864 14884
rect 9640 14844 9864 14872
rect 9640 14832 9646 14844
rect 9858 14832 9864 14844
rect 9916 14832 9922 14884
rect 12802 14872 12808 14884
rect 12763 14844 12808 14872
rect 12802 14832 12808 14844
rect 12860 14832 12866 14884
rect 3418 14804 3424 14816
rect 3379 14776 3424 14804
rect 3418 14764 3424 14776
rect 3476 14764 3482 14816
rect 3970 14804 3976 14816
rect 3931 14776 3976 14804
rect 3970 14764 3976 14776
rect 4028 14764 4034 14816
rect 5902 14764 5908 14816
rect 5960 14804 5966 14816
rect 5997 14807 6055 14813
rect 5997 14804 6009 14807
rect 5960 14776 6009 14804
rect 5960 14764 5966 14776
rect 5997 14773 6009 14776
rect 6043 14773 6055 14807
rect 5997 14767 6055 14773
rect 6178 14764 6184 14816
rect 6236 14804 6242 14816
rect 6457 14807 6515 14813
rect 6457 14804 6469 14807
rect 6236 14776 6469 14804
rect 6236 14764 6242 14776
rect 6457 14773 6469 14776
rect 6503 14804 6515 14807
rect 7006 14804 7012 14816
rect 6503 14776 7012 14804
rect 6503 14773 6515 14776
rect 6457 14767 6515 14773
rect 7006 14764 7012 14776
rect 7064 14764 7070 14816
rect 7190 14804 7196 14816
rect 7151 14776 7196 14804
rect 7190 14764 7196 14776
rect 7248 14764 7254 14816
rect 9122 14804 9128 14816
rect 9083 14776 9128 14804
rect 9122 14764 9128 14776
rect 9180 14764 9186 14816
rect 9217 14807 9275 14813
rect 9217 14773 9229 14807
rect 9263 14804 9275 14807
rect 9398 14804 9404 14816
rect 9263 14776 9404 14804
rect 9263 14773 9275 14776
rect 9217 14767 9275 14773
rect 9398 14764 9404 14776
rect 9456 14764 9462 14816
rect 10689 14807 10747 14813
rect 10689 14773 10701 14807
rect 10735 14804 10747 14807
rect 11146 14804 11152 14816
rect 10735 14776 11152 14804
rect 10735 14773 10747 14776
rect 10689 14767 10747 14773
rect 11146 14764 11152 14776
rect 11204 14764 11210 14816
rect 11609 14807 11667 14813
rect 11609 14773 11621 14807
rect 11655 14804 11667 14807
rect 12069 14807 12127 14813
rect 12069 14804 12081 14807
rect 11655 14776 12081 14804
rect 11655 14773 11667 14776
rect 11609 14767 11667 14773
rect 12069 14773 12081 14776
rect 12115 14804 12127 14807
rect 12161 14807 12219 14813
rect 12161 14804 12173 14807
rect 12115 14776 12173 14804
rect 12115 14773 12127 14776
rect 12069 14767 12127 14773
rect 12161 14773 12173 14776
rect 12207 14773 12219 14807
rect 12161 14767 12219 14773
rect 12526 14764 12532 14816
rect 12584 14804 12590 14816
rect 12621 14807 12679 14813
rect 12621 14804 12633 14807
rect 12584 14776 12633 14804
rect 12584 14764 12590 14776
rect 12621 14773 12633 14776
rect 12667 14773 12679 14807
rect 12621 14767 12679 14773
rect 13814 14764 13820 14816
rect 13872 14804 13878 14816
rect 14568 14804 14596 14971
rect 15212 14949 15240 14980
rect 16574 14968 16580 14980
rect 16632 14968 16638 15020
rect 17494 14968 17500 15020
rect 17552 15008 17558 15020
rect 18472 15011 18530 15017
rect 18472 15008 18484 15011
rect 17552 14980 18484 15008
rect 17552 14968 17558 14980
rect 18472 14977 18484 14980
rect 18518 15008 18530 15011
rect 18616 15008 18644 15048
rect 19886 15036 19892 15048
rect 19944 15036 19950 15088
rect 22462 15076 22468 15088
rect 22423 15048 22468 15076
rect 22462 15036 22468 15048
rect 22520 15036 22526 15088
rect 25866 15036 25872 15088
rect 25924 15076 25930 15088
rect 26237 15079 26295 15085
rect 26237 15076 26249 15079
rect 25924 15048 26249 15076
rect 25924 15036 25930 15048
rect 26237 15045 26249 15048
rect 26283 15076 26295 15079
rect 26786 15076 26792 15088
rect 26283 15048 26792 15076
rect 26283 15045 26295 15048
rect 26237 15039 26295 15045
rect 26786 15036 26792 15048
rect 26844 15076 26850 15088
rect 26973 15079 27031 15085
rect 26973 15076 26985 15079
rect 26844 15048 26985 15076
rect 26844 15036 26850 15048
rect 26973 15045 26985 15048
rect 27019 15045 27031 15079
rect 27706 15076 27712 15088
rect 27667 15048 27712 15076
rect 26973 15039 27031 15045
rect 27706 15036 27712 15048
rect 27764 15036 27770 15088
rect 18518 14980 18644 15008
rect 18693 15011 18751 15017
rect 18518 14977 18530 14980
rect 18472 14971 18530 14977
rect 18693 14977 18705 15011
rect 18739 15008 18751 15011
rect 18782 15008 18788 15020
rect 18739 14980 18788 15008
rect 18739 14977 18751 14980
rect 18693 14971 18751 14977
rect 18782 14968 18788 14980
rect 18840 14968 18846 15020
rect 19061 15011 19119 15017
rect 19061 14977 19073 15011
rect 19107 15008 19119 15011
rect 19242 15008 19248 15020
rect 19107 14980 19248 15008
rect 19107 14977 19119 14980
rect 19061 14971 19119 14977
rect 19242 14968 19248 14980
rect 19300 14968 19306 15020
rect 23842 14968 23848 15020
rect 23900 15008 23906 15020
rect 24394 15008 24400 15020
rect 23900 14980 24400 15008
rect 23900 14968 23906 14980
rect 24394 14968 24400 14980
rect 24452 14968 24458 15020
rect 26326 15008 26332 15020
rect 26239 14980 26332 15008
rect 26326 14968 26332 14980
rect 26384 15008 26390 15020
rect 26694 15008 26700 15020
rect 26384 14980 26700 15008
rect 26384 14968 26390 14980
rect 26694 14968 26700 14980
rect 26752 14968 26758 15020
rect 29822 14968 29828 15020
rect 29880 15008 29886 15020
rect 30558 15008 30564 15020
rect 29880 14980 30420 15008
rect 30519 14980 30564 15008
rect 29880 14968 29886 14980
rect 15197 14943 15255 14949
rect 15197 14909 15209 14943
rect 15243 14909 15255 14943
rect 15197 14903 15255 14909
rect 15289 14943 15347 14949
rect 15289 14909 15301 14943
rect 15335 14909 15347 14943
rect 15289 14903 15347 14909
rect 15304 14872 15332 14903
rect 15378 14900 15384 14952
rect 15436 14940 15442 14952
rect 15654 14940 15660 14952
rect 15436 14912 15660 14940
rect 15436 14900 15442 14912
rect 15654 14900 15660 14912
rect 15712 14900 15718 14952
rect 16298 14900 16304 14952
rect 16356 14940 16362 14952
rect 16761 14943 16819 14949
rect 16761 14940 16773 14943
rect 16356 14912 16773 14940
rect 16356 14900 16362 14912
rect 16761 14909 16773 14912
rect 16807 14940 16819 14943
rect 17221 14943 17279 14949
rect 17221 14940 17233 14943
rect 16807 14912 17233 14940
rect 16807 14909 16819 14912
rect 16761 14903 16819 14909
rect 17221 14909 17233 14912
rect 17267 14940 17279 14943
rect 18046 14940 18052 14952
rect 17267 14912 18052 14940
rect 17267 14909 17279 14912
rect 17221 14903 17279 14909
rect 18046 14900 18052 14912
rect 18104 14900 18110 14952
rect 18322 14940 18328 14952
rect 18235 14912 18328 14940
rect 18322 14900 18328 14912
rect 18380 14940 18386 14952
rect 19150 14940 19156 14952
rect 18380 14912 19156 14940
rect 18380 14900 18386 14912
rect 19150 14900 19156 14912
rect 19208 14900 19214 14952
rect 19334 14900 19340 14952
rect 19392 14940 19398 14952
rect 19705 14943 19763 14949
rect 19705 14940 19717 14943
rect 19392 14912 19717 14940
rect 19392 14900 19398 14912
rect 19705 14909 19717 14912
rect 19751 14909 19763 14943
rect 20162 14940 20168 14952
rect 20123 14912 20168 14940
rect 19705 14903 19763 14909
rect 20162 14900 20168 14912
rect 20220 14900 20226 14952
rect 21637 14943 21695 14949
rect 21637 14909 21649 14943
rect 21683 14909 21695 14943
rect 21637 14903 21695 14909
rect 22189 14943 22247 14949
rect 22189 14909 22201 14943
rect 22235 14940 22247 14943
rect 22278 14940 22284 14952
rect 22235 14912 22284 14940
rect 22235 14909 22247 14912
rect 22189 14903 22247 14909
rect 15562 14872 15568 14884
rect 15304 14844 15568 14872
rect 15562 14832 15568 14844
rect 15620 14832 15626 14884
rect 19242 14832 19248 14884
rect 19300 14872 19306 14884
rect 19889 14875 19947 14881
rect 19889 14872 19901 14875
rect 19300 14844 19901 14872
rect 19300 14832 19306 14844
rect 19889 14841 19901 14844
rect 19935 14841 19947 14875
rect 19889 14835 19947 14841
rect 13872 14776 14596 14804
rect 16945 14807 17003 14813
rect 13872 14764 13878 14776
rect 16945 14773 16957 14807
rect 16991 14804 17003 14807
rect 17126 14804 17132 14816
rect 16991 14776 17132 14804
rect 16991 14773 17003 14776
rect 16945 14767 17003 14773
rect 17126 14764 17132 14776
rect 17184 14764 17190 14816
rect 18598 14764 18604 14816
rect 18656 14804 18662 14816
rect 19150 14804 19156 14816
rect 18656 14776 19156 14804
rect 18656 14764 18662 14776
rect 19150 14764 19156 14776
rect 19208 14804 19214 14816
rect 19337 14807 19395 14813
rect 19337 14804 19349 14807
rect 19208 14776 19349 14804
rect 19208 14764 19214 14776
rect 19337 14773 19349 14776
rect 19383 14773 19395 14807
rect 19337 14767 19395 14773
rect 21545 14807 21603 14813
rect 21545 14773 21557 14807
rect 21591 14804 21603 14807
rect 21652 14804 21680 14903
rect 22278 14900 22284 14912
rect 22336 14900 22342 14952
rect 22554 14940 22560 14952
rect 22515 14912 22560 14940
rect 22554 14900 22560 14912
rect 22612 14900 22618 14952
rect 23474 14900 23480 14952
rect 23532 14940 23538 14952
rect 24029 14943 24087 14949
rect 24029 14940 24041 14943
rect 23532 14912 24041 14940
rect 23532 14900 23538 14912
rect 24029 14909 24041 14912
rect 24075 14909 24087 14943
rect 24029 14903 24087 14909
rect 24118 14900 24124 14952
rect 24176 14949 24182 14952
rect 24176 14943 24234 14949
rect 24176 14909 24188 14943
rect 24222 14909 24234 14943
rect 24176 14903 24234 14909
rect 25133 14943 25191 14949
rect 25133 14909 25145 14943
rect 25179 14940 25191 14943
rect 25958 14940 25964 14952
rect 25179 14912 25964 14940
rect 25179 14909 25191 14912
rect 25133 14903 25191 14909
rect 24176 14900 24182 14903
rect 25958 14900 25964 14912
rect 26016 14900 26022 14952
rect 26602 14900 26608 14952
rect 26660 14940 26666 14952
rect 27430 14940 27436 14952
rect 26660 14912 27436 14940
rect 26660 14900 26666 14912
rect 27430 14900 27436 14912
rect 27488 14940 27494 14952
rect 27525 14943 27583 14949
rect 27525 14940 27537 14943
rect 27488 14912 27537 14940
rect 27488 14900 27494 14912
rect 27525 14909 27537 14912
rect 27571 14909 27583 14943
rect 27525 14903 27583 14909
rect 29917 14943 29975 14949
rect 29917 14909 29929 14943
rect 29963 14940 29975 14943
rect 30190 14940 30196 14952
rect 29963 14912 30196 14940
rect 29963 14909 29975 14912
rect 29917 14903 29975 14909
rect 30190 14900 30196 14912
rect 30248 14900 30254 14952
rect 30392 14940 30420 14980
rect 30558 14968 30564 14980
rect 30616 14968 30622 15020
rect 31864 15008 31892 15104
rect 34422 15036 34428 15088
rect 34480 15076 34486 15088
rect 35069 15079 35127 15085
rect 35069 15076 35081 15079
rect 34480 15048 35081 15076
rect 34480 15036 34486 15048
rect 35069 15045 35081 15048
rect 35115 15045 35127 15079
rect 35069 15039 35127 15045
rect 33042 15008 33048 15020
rect 31864 14980 33048 15008
rect 33042 14968 33048 14980
rect 33100 14968 33106 15020
rect 30469 14943 30527 14949
rect 30469 14940 30481 14943
rect 30392 14912 30481 14940
rect 30469 14909 30481 14912
rect 30515 14940 30527 14943
rect 31021 14943 31079 14949
rect 31021 14940 31033 14943
rect 30515 14912 31033 14940
rect 30515 14909 30527 14912
rect 30469 14903 30527 14909
rect 31021 14909 31033 14912
rect 31067 14909 31079 14943
rect 31021 14903 31079 14909
rect 32582 14900 32588 14952
rect 32640 14940 32646 14952
rect 33321 14943 33379 14949
rect 33321 14940 33333 14943
rect 32640 14912 33333 14940
rect 32640 14900 32646 14912
rect 33321 14909 33333 14912
rect 33367 14909 33379 14943
rect 33502 14940 33508 14952
rect 33463 14912 33508 14940
rect 33321 14903 33379 14909
rect 33502 14900 33508 14912
rect 33560 14900 33566 14952
rect 26694 14872 26700 14884
rect 26655 14844 26700 14872
rect 26694 14832 26700 14844
rect 26752 14832 26758 14884
rect 30006 14872 30012 14884
rect 29012 14844 30012 14872
rect 21818 14804 21824 14816
rect 21591 14776 21824 14804
rect 21591 14773 21603 14776
rect 21545 14767 21603 14773
rect 21818 14764 21824 14776
rect 21876 14764 21882 14816
rect 23937 14807 23995 14813
rect 23937 14773 23949 14807
rect 23983 14804 23995 14807
rect 24210 14804 24216 14816
rect 23983 14776 24216 14804
rect 23983 14773 23995 14776
rect 23937 14767 23995 14773
rect 24210 14764 24216 14776
rect 24268 14764 24274 14816
rect 25498 14804 25504 14816
rect 25459 14776 25504 14804
rect 25498 14764 25504 14776
rect 25556 14764 25562 14816
rect 25866 14804 25872 14816
rect 25827 14776 25872 14804
rect 25866 14764 25872 14776
rect 25924 14764 25930 14816
rect 28074 14764 28080 14816
rect 28132 14804 28138 14816
rect 29012 14813 29040 14844
rect 30006 14832 30012 14844
rect 30064 14832 30070 14884
rect 30374 14832 30380 14884
rect 30432 14872 30438 14884
rect 31389 14875 31447 14881
rect 31389 14872 31401 14875
rect 30432 14844 31401 14872
rect 30432 14832 30438 14844
rect 31389 14841 31401 14844
rect 31435 14841 31447 14875
rect 31389 14835 31447 14841
rect 32493 14875 32551 14881
rect 32493 14841 32505 14875
rect 32539 14872 32551 14875
rect 33594 14872 33600 14884
rect 32539 14844 33600 14872
rect 32539 14841 32551 14844
rect 32493 14835 32551 14841
rect 33594 14832 33600 14844
rect 33652 14832 33658 14884
rect 28997 14807 29055 14813
rect 28997 14804 29009 14807
rect 28132 14776 29009 14804
rect 28132 14764 28138 14776
rect 28997 14773 29009 14776
rect 29043 14773 29055 14807
rect 28997 14767 29055 14773
rect 1104 14714 38548 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 38548 14714
rect 1104 14640 38548 14662
rect 1394 14560 1400 14612
rect 1452 14600 1458 14612
rect 1949 14603 2007 14609
rect 1949 14600 1961 14603
rect 1452 14572 1961 14600
rect 1452 14560 1458 14572
rect 1949 14569 1961 14572
rect 1995 14600 2007 14603
rect 2682 14600 2688 14612
rect 1995 14572 2688 14600
rect 1995 14569 2007 14572
rect 1949 14563 2007 14569
rect 2682 14560 2688 14572
rect 2740 14560 2746 14612
rect 3510 14600 3516 14612
rect 3471 14572 3516 14600
rect 3510 14560 3516 14572
rect 3568 14560 3574 14612
rect 3878 14600 3884 14612
rect 3839 14572 3884 14600
rect 3878 14560 3884 14572
rect 3936 14560 3942 14612
rect 4338 14600 4344 14612
rect 4299 14572 4344 14600
rect 4338 14560 4344 14572
rect 4396 14560 4402 14612
rect 5350 14600 5356 14612
rect 5311 14572 5356 14600
rect 5350 14560 5356 14572
rect 5408 14560 5414 14612
rect 6086 14600 6092 14612
rect 6047 14572 6092 14600
rect 6086 14560 6092 14572
rect 6144 14560 6150 14612
rect 7469 14603 7527 14609
rect 7469 14569 7481 14603
rect 7515 14600 7527 14603
rect 8110 14600 8116 14612
rect 7515 14572 8116 14600
rect 7515 14569 7527 14572
rect 7469 14563 7527 14569
rect 8110 14560 8116 14572
rect 8168 14560 8174 14612
rect 8202 14560 8208 14612
rect 8260 14560 8266 14612
rect 10870 14600 10876 14612
rect 9968 14572 10876 14600
rect 2498 14492 2504 14544
rect 2556 14532 2562 14544
rect 3145 14535 3203 14541
rect 3145 14532 3157 14535
rect 2556 14504 3157 14532
rect 2556 14492 2562 14504
rect 3145 14501 3157 14504
rect 3191 14532 3203 14535
rect 4798 14532 4804 14544
rect 3191 14504 4804 14532
rect 3191 14501 3203 14504
rect 3145 14495 3203 14501
rect 4798 14492 4804 14504
rect 4856 14492 4862 14544
rect 7101 14535 7159 14541
rect 7101 14501 7113 14535
rect 7147 14532 7159 14535
rect 8220 14532 8248 14560
rect 7147 14504 8248 14532
rect 8297 14535 8355 14541
rect 7147 14501 7159 14504
rect 7101 14495 7159 14501
rect 8297 14501 8309 14535
rect 8343 14532 8355 14535
rect 8478 14532 8484 14544
rect 8343 14504 8484 14532
rect 8343 14501 8355 14504
rect 8297 14495 8355 14501
rect 8478 14492 8484 14504
rect 8536 14492 8542 14544
rect 9858 14492 9864 14544
rect 9916 14532 9922 14544
rect 9968 14541 9996 14572
rect 10870 14560 10876 14572
rect 10928 14600 10934 14612
rect 10965 14603 11023 14609
rect 10965 14600 10977 14603
rect 10928 14572 10977 14600
rect 10928 14560 10934 14572
rect 10965 14569 10977 14572
rect 11011 14569 11023 14603
rect 10965 14563 11023 14569
rect 11514 14560 11520 14612
rect 11572 14600 11578 14612
rect 11701 14603 11759 14609
rect 11701 14600 11713 14603
rect 11572 14572 11713 14600
rect 11572 14560 11578 14572
rect 11701 14569 11713 14572
rect 11747 14569 11759 14603
rect 13354 14600 13360 14612
rect 13315 14572 13360 14600
rect 11701 14563 11759 14569
rect 13354 14560 13360 14572
rect 13412 14560 13418 14612
rect 14090 14560 14096 14612
rect 14148 14600 14154 14612
rect 14185 14603 14243 14609
rect 14185 14600 14197 14603
rect 14148 14572 14197 14600
rect 14148 14560 14154 14572
rect 14185 14569 14197 14572
rect 14231 14600 14243 14603
rect 14918 14600 14924 14612
rect 14231 14572 14924 14600
rect 14231 14569 14243 14572
rect 14185 14563 14243 14569
rect 14918 14560 14924 14572
rect 14976 14560 14982 14612
rect 15194 14560 15200 14612
rect 15252 14600 15258 14612
rect 16206 14600 16212 14612
rect 15252 14572 16212 14600
rect 15252 14560 15258 14572
rect 16206 14560 16212 14572
rect 16264 14600 16270 14612
rect 17494 14600 17500 14612
rect 16264 14572 16712 14600
rect 17455 14572 17500 14600
rect 16264 14560 16270 14572
rect 9953 14535 10011 14541
rect 9953 14532 9965 14535
rect 9916 14504 9965 14532
rect 9916 14492 9922 14504
rect 9953 14501 9965 14504
rect 9999 14501 10011 14535
rect 9953 14495 10011 14501
rect 10321 14535 10379 14541
rect 10321 14501 10333 14535
rect 10367 14532 10379 14535
rect 10689 14535 10747 14541
rect 10367 14504 10456 14532
rect 10367 14501 10379 14504
rect 10321 14495 10379 14501
rect 4062 14424 4068 14476
rect 4120 14464 4126 14476
rect 4157 14467 4215 14473
rect 4157 14464 4169 14467
rect 4120 14436 4169 14464
rect 4120 14424 4126 14436
rect 4157 14433 4169 14436
rect 4203 14433 4215 14467
rect 6454 14464 6460 14476
rect 6415 14436 6460 14464
rect 4157 14427 4215 14433
rect 6454 14424 6460 14436
rect 6512 14424 6518 14476
rect 7837 14467 7895 14473
rect 7837 14433 7849 14467
rect 7883 14464 7895 14467
rect 7926 14464 7932 14476
rect 7883 14436 7932 14464
rect 7883 14433 7895 14436
rect 7837 14427 7895 14433
rect 7926 14424 7932 14436
rect 7984 14424 7990 14476
rect 8110 14464 8116 14476
rect 8071 14436 8116 14464
rect 8110 14424 8116 14436
rect 8168 14424 8174 14476
rect 8202 14424 8208 14476
rect 8260 14464 8266 14476
rect 8260 14436 8305 14464
rect 8260 14424 8266 14436
rect 9490 14424 9496 14476
rect 9548 14464 9554 14476
rect 10137 14467 10195 14473
rect 10137 14464 10149 14467
rect 9548 14436 10149 14464
rect 9548 14424 9554 14436
rect 8665 14399 8723 14405
rect 8665 14396 8677 14399
rect 8036 14368 8677 14396
rect 4709 14331 4767 14337
rect 4709 14297 4721 14331
rect 4755 14328 4767 14331
rect 4890 14328 4896 14340
rect 4755 14300 4896 14328
rect 4755 14297 4767 14300
rect 4709 14291 4767 14297
rect 4890 14288 4896 14300
rect 4948 14288 4954 14340
rect 5534 14288 5540 14340
rect 5592 14328 5598 14340
rect 6641 14331 6699 14337
rect 6641 14328 6653 14331
rect 5592 14300 6653 14328
rect 5592 14288 5598 14300
rect 6641 14297 6653 14300
rect 6687 14328 6699 14331
rect 7190 14328 7196 14340
rect 6687 14300 7196 14328
rect 6687 14297 6699 14300
rect 6641 14291 6699 14297
rect 7190 14288 7196 14300
rect 7248 14288 7254 14340
rect 7374 14288 7380 14340
rect 7432 14328 7438 14340
rect 8036 14328 8064 14368
rect 8665 14365 8677 14368
rect 8711 14365 8723 14399
rect 8665 14359 8723 14365
rect 7432 14300 8064 14328
rect 7432 14288 7438 14300
rect 8570 14288 8576 14340
rect 8628 14328 8634 14340
rect 9309 14331 9367 14337
rect 9309 14328 9321 14331
rect 8628 14300 9321 14328
rect 8628 14288 8634 14300
rect 9309 14297 9321 14300
rect 9355 14328 9367 14331
rect 9858 14328 9864 14340
rect 9355 14300 9864 14328
rect 9355 14297 9367 14300
rect 9309 14291 9367 14297
rect 9858 14288 9864 14300
rect 9916 14288 9922 14340
rect 1578 14260 1584 14272
rect 1539 14232 1584 14260
rect 1578 14220 1584 14232
rect 1636 14220 1642 14272
rect 5718 14260 5724 14272
rect 5679 14232 5724 14260
rect 5718 14220 5724 14232
rect 5776 14220 5782 14272
rect 7926 14220 7932 14272
rect 7984 14260 7990 14272
rect 8202 14260 8208 14272
rect 7984 14232 8208 14260
rect 7984 14220 7990 14232
rect 8202 14220 8208 14232
rect 8260 14220 8266 14272
rect 8662 14220 8668 14272
rect 8720 14260 8726 14272
rect 8941 14263 8999 14269
rect 8941 14260 8953 14263
rect 8720 14232 8953 14260
rect 8720 14220 8726 14232
rect 8941 14229 8953 14232
rect 8987 14260 8999 14263
rect 9122 14260 9128 14272
rect 8987 14232 9128 14260
rect 8987 14229 8999 14232
rect 8941 14223 8999 14229
rect 9122 14220 9128 14232
rect 9180 14220 9186 14272
rect 10060 14260 10088 14436
rect 10137 14433 10149 14436
rect 10183 14433 10195 14467
rect 10137 14427 10195 14433
rect 10226 14424 10232 14476
rect 10284 14464 10290 14476
rect 10284 14436 10329 14464
rect 10284 14424 10290 14436
rect 10428 14396 10456 14504
rect 10689 14501 10701 14535
rect 10735 14532 10747 14535
rect 10778 14532 10784 14544
rect 10735 14504 10784 14532
rect 10735 14501 10747 14504
rect 10689 14495 10747 14501
rect 10778 14492 10784 14504
rect 10836 14492 10842 14544
rect 12250 14492 12256 14544
rect 12308 14532 12314 14544
rect 12986 14532 12992 14544
rect 12308 14504 12992 14532
rect 12308 14492 12314 14504
rect 12986 14492 12992 14504
rect 13044 14532 13050 14544
rect 13449 14535 13507 14541
rect 13449 14532 13461 14535
rect 13044 14504 13461 14532
rect 13044 14492 13050 14504
rect 13449 14501 13461 14504
rect 13495 14501 13507 14535
rect 13449 14495 13507 14501
rect 13630 14492 13636 14544
rect 13688 14532 13694 14544
rect 13817 14535 13875 14541
rect 13817 14532 13829 14535
rect 13688 14504 13829 14532
rect 13688 14492 13694 14504
rect 13817 14501 13829 14504
rect 13863 14501 13875 14535
rect 13817 14495 13875 14501
rect 15565 14535 15623 14541
rect 15565 14501 15577 14535
rect 15611 14532 15623 14535
rect 15654 14532 15660 14544
rect 15611 14504 15660 14532
rect 15611 14501 15623 14504
rect 15565 14495 15623 14501
rect 15654 14492 15660 14504
rect 15712 14492 15718 14544
rect 15930 14492 15936 14544
rect 15988 14532 15994 14544
rect 16301 14535 16359 14541
rect 15988 14504 16252 14532
rect 15988 14492 15994 14504
rect 11885 14467 11943 14473
rect 11885 14433 11897 14467
rect 11931 14464 11943 14467
rect 12066 14464 12072 14476
rect 11931 14436 12072 14464
rect 11931 14433 11943 14436
rect 11885 14427 11943 14433
rect 12066 14424 12072 14436
rect 12124 14424 12130 14476
rect 12897 14467 12955 14473
rect 12897 14433 12909 14467
rect 12943 14464 12955 14467
rect 13262 14464 13268 14476
rect 12943 14436 13268 14464
rect 12943 14433 12955 14436
rect 12897 14427 12955 14433
rect 13262 14424 13268 14436
rect 13320 14424 13326 14476
rect 15105 14467 15163 14473
rect 15105 14433 15117 14467
rect 15151 14464 15163 14467
rect 15194 14464 15200 14476
rect 15151 14436 15200 14464
rect 15151 14433 15163 14436
rect 15105 14427 15163 14433
rect 15194 14424 15200 14436
rect 15252 14464 15258 14476
rect 16224 14473 16252 14504
rect 16301 14501 16313 14535
rect 16347 14532 16359 14535
rect 16574 14532 16580 14544
rect 16347 14504 16580 14532
rect 16347 14501 16359 14504
rect 16301 14495 16359 14501
rect 16574 14492 16580 14504
rect 16632 14492 16638 14544
rect 16684 14541 16712 14572
rect 17494 14560 17500 14572
rect 17552 14560 17558 14612
rect 17770 14600 17776 14612
rect 17731 14572 17776 14600
rect 17770 14560 17776 14572
rect 17828 14560 17834 14612
rect 18693 14603 18751 14609
rect 17880 14572 18552 14600
rect 17880 14541 17908 14572
rect 16669 14535 16727 14541
rect 16669 14501 16681 14535
rect 16715 14501 16727 14535
rect 17865 14535 17923 14541
rect 17865 14532 17877 14535
rect 16669 14495 16727 14501
rect 17512 14504 17877 14532
rect 17512 14476 17540 14504
rect 17865 14501 17877 14504
rect 17911 14501 17923 14535
rect 17865 14495 17923 14501
rect 17957 14535 18015 14541
rect 17957 14501 17969 14535
rect 18003 14532 18015 14535
rect 18138 14532 18144 14544
rect 18003 14504 18144 14532
rect 18003 14501 18015 14504
rect 17957 14495 18015 14501
rect 18138 14492 18144 14504
rect 18196 14492 18202 14544
rect 18322 14532 18328 14544
rect 18283 14504 18328 14532
rect 18322 14492 18328 14504
rect 18380 14492 18386 14544
rect 18524 14532 18552 14572
rect 18693 14569 18705 14603
rect 18739 14600 18751 14603
rect 18782 14600 18788 14612
rect 18739 14572 18788 14600
rect 18739 14569 18751 14572
rect 18693 14563 18751 14569
rect 18782 14560 18788 14572
rect 18840 14560 18846 14612
rect 19058 14600 19064 14612
rect 18971 14572 19064 14600
rect 19058 14560 19064 14572
rect 19116 14600 19122 14612
rect 19242 14600 19248 14612
rect 19116 14572 19248 14600
rect 19116 14560 19122 14572
rect 19242 14560 19248 14572
rect 19300 14560 19306 14612
rect 19426 14560 19432 14612
rect 19484 14600 19490 14612
rect 20533 14603 20591 14609
rect 20533 14600 20545 14603
rect 19484 14572 20545 14600
rect 19484 14560 19490 14572
rect 20533 14569 20545 14572
rect 20579 14569 20591 14603
rect 20533 14563 20591 14569
rect 21637 14603 21695 14609
rect 21637 14569 21649 14603
rect 21683 14600 21695 14603
rect 21726 14600 21732 14612
rect 21683 14572 21732 14600
rect 21683 14569 21695 14572
rect 21637 14563 21695 14569
rect 21726 14560 21732 14572
rect 21784 14560 21790 14612
rect 22097 14603 22155 14609
rect 22097 14569 22109 14603
rect 22143 14569 22155 14603
rect 22738 14600 22744 14612
rect 22699 14572 22744 14600
rect 22097 14563 22155 14569
rect 18524 14504 19472 14532
rect 16117 14467 16175 14473
rect 16117 14464 16129 14467
rect 15252 14436 16129 14464
rect 15252 14424 15258 14436
rect 16117 14433 16129 14436
rect 16163 14433 16175 14467
rect 16117 14427 16175 14433
rect 16209 14467 16267 14473
rect 16209 14433 16221 14467
rect 16255 14433 16267 14467
rect 16209 14427 16267 14433
rect 12342 14396 12348 14408
rect 10152 14368 12348 14396
rect 10152 14340 10180 14368
rect 12342 14356 12348 14368
rect 12400 14356 12406 14408
rect 13078 14396 13084 14408
rect 13039 14368 13084 14396
rect 13078 14356 13084 14368
rect 13136 14396 13142 14408
rect 13906 14396 13912 14408
rect 13136 14368 13912 14396
rect 13136 14356 13142 14368
rect 13906 14356 13912 14368
rect 13964 14356 13970 14408
rect 15470 14356 15476 14408
rect 15528 14396 15534 14408
rect 15933 14399 15991 14405
rect 15933 14396 15945 14399
rect 15528 14368 15945 14396
rect 15528 14356 15534 14368
rect 15933 14365 15945 14368
rect 15979 14365 15991 14399
rect 16132 14396 16160 14427
rect 17494 14424 17500 14476
rect 17552 14424 17558 14476
rect 18046 14424 18052 14476
rect 18104 14464 18110 14476
rect 19334 14464 19340 14476
rect 18104 14436 19340 14464
rect 18104 14424 18110 14436
rect 19334 14424 19340 14436
rect 19392 14424 19398 14476
rect 19444 14473 19472 14504
rect 19518 14492 19524 14544
rect 19576 14532 19582 14544
rect 19886 14532 19892 14544
rect 19576 14504 19621 14532
rect 19847 14504 19892 14532
rect 19576 14492 19582 14504
rect 19886 14492 19892 14504
rect 19944 14492 19950 14544
rect 22112 14532 22140 14563
rect 22738 14560 22744 14572
rect 22796 14560 22802 14612
rect 25958 14560 25964 14612
rect 26016 14600 26022 14612
rect 26973 14603 27031 14609
rect 26973 14600 26985 14603
rect 26016 14572 26985 14600
rect 26016 14560 26022 14572
rect 26973 14569 26985 14572
rect 27019 14569 27031 14603
rect 27338 14600 27344 14612
rect 27299 14572 27344 14600
rect 26973 14563 27031 14569
rect 27338 14560 27344 14572
rect 27396 14560 27402 14612
rect 27890 14600 27896 14612
rect 27851 14572 27896 14600
rect 27890 14560 27896 14572
rect 27948 14560 27954 14612
rect 29914 14600 29920 14612
rect 29875 14572 29920 14600
rect 29914 14560 29920 14572
rect 29972 14560 29978 14612
rect 30377 14603 30435 14609
rect 30377 14569 30389 14603
rect 30423 14600 30435 14603
rect 30466 14600 30472 14612
rect 30423 14572 30472 14600
rect 30423 14569 30435 14572
rect 30377 14563 30435 14569
rect 30466 14560 30472 14572
rect 30524 14560 30530 14612
rect 32309 14603 32367 14609
rect 32309 14569 32321 14603
rect 32355 14600 32367 14603
rect 32582 14600 32588 14612
rect 32355 14572 32588 14600
rect 32355 14569 32367 14572
rect 32309 14563 32367 14569
rect 32582 14560 32588 14572
rect 32640 14560 32646 14612
rect 33042 14600 33048 14612
rect 33003 14572 33048 14600
rect 33042 14560 33048 14572
rect 33100 14560 33106 14612
rect 23474 14532 23480 14544
rect 22112 14504 23480 14532
rect 23474 14492 23480 14504
rect 23532 14492 23538 14544
rect 26053 14535 26111 14541
rect 26053 14501 26065 14535
rect 26099 14532 26111 14535
rect 26326 14532 26332 14544
rect 26099 14504 26332 14532
rect 26099 14501 26111 14504
rect 26053 14495 26111 14501
rect 26326 14492 26332 14504
rect 26384 14492 26390 14544
rect 28258 14492 28264 14544
rect 28316 14532 28322 14544
rect 28316 14504 28764 14532
rect 28316 14492 28322 14504
rect 19429 14467 19487 14473
rect 19429 14433 19441 14467
rect 19475 14464 19487 14467
rect 20162 14464 20168 14476
rect 19475 14436 20168 14464
rect 19475 14433 19487 14436
rect 19429 14427 19487 14433
rect 20162 14424 20168 14436
rect 20220 14424 20226 14476
rect 20901 14467 20959 14473
rect 20901 14433 20913 14467
rect 20947 14464 20959 14467
rect 20990 14464 20996 14476
rect 20947 14436 20996 14464
rect 20947 14433 20959 14436
rect 20901 14427 20959 14433
rect 20990 14424 20996 14436
rect 21048 14424 21054 14476
rect 21910 14464 21916 14476
rect 21871 14436 21916 14464
rect 21910 14424 21916 14436
rect 21968 14424 21974 14476
rect 22925 14467 22983 14473
rect 22925 14433 22937 14467
rect 22971 14433 22983 14467
rect 23934 14464 23940 14476
rect 23895 14436 23940 14464
rect 22925 14427 22983 14433
rect 17589 14399 17647 14405
rect 16132 14368 17080 14396
rect 15933 14359 15991 14365
rect 10134 14288 10140 14340
rect 10192 14288 10198 14340
rect 13998 14288 14004 14340
rect 14056 14328 14062 14340
rect 14461 14331 14519 14337
rect 14461 14328 14473 14331
rect 14056 14300 14473 14328
rect 14056 14288 14062 14300
rect 14461 14297 14473 14300
rect 14507 14297 14519 14331
rect 14461 14291 14519 14297
rect 10686 14260 10692 14272
rect 10060 14232 10692 14260
rect 10686 14220 10692 14232
rect 10744 14260 10750 14272
rect 11330 14260 11336 14272
rect 10744 14232 11336 14260
rect 10744 14220 10750 14232
rect 11330 14220 11336 14232
rect 11388 14220 11394 14272
rect 11422 14220 11428 14272
rect 11480 14260 11486 14272
rect 12066 14260 12072 14272
rect 11480 14232 12072 14260
rect 11480 14220 11486 14232
rect 12066 14220 12072 14232
rect 12124 14220 12130 14272
rect 12526 14260 12532 14272
rect 12439 14232 12532 14260
rect 12526 14220 12532 14232
rect 12584 14260 12590 14272
rect 12894 14260 12900 14272
rect 12584 14232 12900 14260
rect 12584 14220 12590 14232
rect 12894 14220 12900 14232
rect 12952 14220 12958 14272
rect 17052 14269 17080 14368
rect 17589 14365 17601 14399
rect 17635 14365 17647 14399
rect 19150 14396 19156 14408
rect 19111 14368 19156 14396
rect 17589 14359 17647 14365
rect 17604 14328 17632 14359
rect 19150 14356 19156 14368
rect 19208 14356 19214 14408
rect 17770 14328 17776 14340
rect 17604 14300 17776 14328
rect 17770 14288 17776 14300
rect 17828 14288 17834 14340
rect 18138 14288 18144 14340
rect 18196 14328 18202 14340
rect 20165 14331 20223 14337
rect 20165 14328 20177 14331
rect 18196 14300 20177 14328
rect 18196 14288 18202 14300
rect 20165 14297 20177 14300
rect 20211 14297 20223 14331
rect 20165 14291 20223 14297
rect 20254 14288 20260 14340
rect 20312 14328 20318 14340
rect 21085 14331 21143 14337
rect 21085 14328 21097 14331
rect 20312 14300 21097 14328
rect 20312 14288 20318 14300
rect 21085 14297 21097 14300
rect 21131 14297 21143 14331
rect 21085 14291 21143 14297
rect 22465 14331 22523 14337
rect 22465 14297 22477 14331
rect 22511 14328 22523 14331
rect 22940 14328 22968 14427
rect 23934 14424 23940 14436
rect 23992 14424 23998 14476
rect 24118 14473 24124 14476
rect 24084 14467 24124 14473
rect 24084 14433 24096 14467
rect 24176 14464 24182 14476
rect 26513 14467 26571 14473
rect 24176 14436 25360 14464
rect 24084 14427 24124 14433
rect 24099 14424 24124 14427
rect 24176 14424 24182 14436
rect 23106 14356 23112 14408
rect 23164 14396 23170 14408
rect 23477 14399 23535 14405
rect 23477 14396 23489 14399
rect 23164 14368 23489 14396
rect 23164 14356 23170 14368
rect 23477 14365 23489 14368
rect 23523 14396 23535 14399
rect 24099 14396 24127 14424
rect 24302 14396 24308 14408
rect 23523 14368 24127 14396
rect 24215 14368 24308 14396
rect 23523 14365 23535 14368
rect 23477 14359 23535 14365
rect 24302 14356 24308 14368
rect 24360 14396 24366 14408
rect 25222 14396 25228 14408
rect 24360 14368 25228 14396
rect 24360 14356 24366 14368
rect 25222 14356 25228 14368
rect 25280 14356 25286 14408
rect 24397 14331 24455 14337
rect 24397 14328 24409 14331
rect 22511 14300 24409 14328
rect 22511 14297 22523 14300
rect 22465 14291 22523 14297
rect 24397 14297 24409 14300
rect 24443 14297 24455 14331
rect 24397 14291 24455 14297
rect 17037 14263 17095 14269
rect 17037 14229 17049 14263
rect 17083 14260 17095 14263
rect 17126 14260 17132 14272
rect 17083 14232 17132 14260
rect 17083 14229 17095 14232
rect 17037 14223 17095 14229
rect 17126 14220 17132 14232
rect 17184 14220 17190 14272
rect 22278 14220 22284 14272
rect 22336 14260 22342 14272
rect 23109 14263 23167 14269
rect 23109 14260 23121 14263
rect 22336 14232 23121 14260
rect 22336 14220 22342 14232
rect 23109 14229 23121 14232
rect 23155 14229 23167 14263
rect 23842 14260 23848 14272
rect 23803 14232 23848 14260
rect 23109 14223 23167 14229
rect 23842 14220 23848 14232
rect 23900 14220 23906 14272
rect 24210 14260 24216 14272
rect 24171 14232 24216 14260
rect 24210 14220 24216 14232
rect 24268 14220 24274 14272
rect 25332 14269 25360 14436
rect 26513 14433 26525 14467
rect 26559 14464 26571 14467
rect 26786 14464 26792 14476
rect 26559 14436 26792 14464
rect 26559 14433 26571 14436
rect 26513 14427 26571 14433
rect 26786 14424 26792 14436
rect 26844 14424 26850 14476
rect 28736 14473 28764 14504
rect 31386 14492 31392 14544
rect 31444 14532 31450 14544
rect 31481 14535 31539 14541
rect 31481 14532 31493 14535
rect 31444 14504 31493 14532
rect 31444 14492 31450 14504
rect 31481 14501 31493 14504
rect 31527 14501 31539 14535
rect 31481 14495 31539 14501
rect 33594 14492 33600 14544
rect 33652 14532 33658 14544
rect 33652 14504 34284 14532
rect 33652 14492 33658 14504
rect 28629 14467 28687 14473
rect 28629 14464 28641 14467
rect 28276 14436 28641 14464
rect 25685 14399 25743 14405
rect 25685 14365 25697 14399
rect 25731 14396 25743 14399
rect 26050 14396 26056 14408
rect 25731 14368 26056 14396
rect 25731 14365 25743 14368
rect 25685 14359 25743 14365
rect 26050 14356 26056 14368
rect 26108 14356 26114 14408
rect 26510 14288 26516 14340
rect 26568 14328 26574 14340
rect 28276 14337 28304 14436
rect 28629 14433 28641 14436
rect 28675 14433 28687 14467
rect 28629 14427 28687 14433
rect 28721 14467 28779 14473
rect 28721 14433 28733 14467
rect 28767 14433 28779 14467
rect 28721 14427 28779 14433
rect 29822 14424 29828 14476
rect 29880 14464 29886 14476
rect 30101 14467 30159 14473
rect 30101 14464 30113 14467
rect 29880 14436 30113 14464
rect 29880 14424 29886 14436
rect 30101 14433 30113 14436
rect 30147 14433 30159 14467
rect 30101 14427 30159 14433
rect 30374 14424 30380 14476
rect 30432 14464 30438 14476
rect 30929 14467 30987 14473
rect 30929 14464 30941 14467
rect 30432 14436 30941 14464
rect 30432 14424 30438 14436
rect 30929 14433 30941 14436
rect 30975 14433 30987 14467
rect 30929 14427 30987 14433
rect 31018 14424 31024 14476
rect 31076 14464 31082 14476
rect 31113 14467 31171 14473
rect 31113 14464 31125 14467
rect 31076 14436 31125 14464
rect 31076 14424 31082 14436
rect 31113 14433 31125 14436
rect 31159 14464 31171 14467
rect 31662 14464 31668 14476
rect 31159 14436 31668 14464
rect 31159 14433 31171 14436
rect 31113 14427 31171 14433
rect 31662 14424 31668 14436
rect 31720 14424 31726 14476
rect 32122 14464 32128 14476
rect 32083 14436 32128 14464
rect 32122 14424 32128 14436
rect 32180 14424 32186 14476
rect 33781 14467 33839 14473
rect 33781 14464 33793 14467
rect 32232 14436 33793 14464
rect 29181 14399 29239 14405
rect 29181 14365 29193 14399
rect 29227 14396 29239 14399
rect 30190 14396 30196 14408
rect 29227 14368 30196 14396
rect 29227 14365 29239 14368
rect 29181 14359 29239 14365
rect 30190 14356 30196 14368
rect 30248 14356 30254 14408
rect 31386 14356 31392 14408
rect 31444 14396 31450 14408
rect 32232 14396 32260 14436
rect 33781 14433 33793 14436
rect 33827 14464 33839 14467
rect 34146 14464 34152 14476
rect 33827 14436 34152 14464
rect 33827 14433 33839 14436
rect 33781 14427 33839 14433
rect 34146 14424 34152 14436
rect 34204 14424 34210 14476
rect 34256 14473 34284 14504
rect 34241 14467 34299 14473
rect 34241 14433 34253 14467
rect 34287 14433 34299 14467
rect 34241 14427 34299 14433
rect 31444 14368 32260 14396
rect 33597 14399 33655 14405
rect 31444 14356 31450 14368
rect 33597 14365 33609 14399
rect 33643 14396 33655 14399
rect 33870 14396 33876 14408
rect 33643 14368 33876 14396
rect 33643 14365 33655 14368
rect 33597 14359 33655 14365
rect 33870 14356 33876 14368
rect 33928 14396 33934 14408
rect 34330 14396 34336 14408
rect 33928 14368 34336 14396
rect 33928 14356 33934 14368
rect 34330 14356 34336 14368
rect 34388 14356 34394 14408
rect 28261 14331 28319 14337
rect 28261 14328 28273 14331
rect 26568 14300 28273 14328
rect 26568 14288 26574 14300
rect 28261 14297 28273 14300
rect 28307 14328 28319 14331
rect 29454 14328 29460 14340
rect 28307 14300 29460 14328
rect 28307 14297 28319 14300
rect 28261 14291 28319 14297
rect 29454 14288 29460 14300
rect 29512 14288 29518 14340
rect 34238 14328 34244 14340
rect 34199 14300 34244 14328
rect 34238 14288 34244 14300
rect 34296 14288 34302 14340
rect 25317 14263 25375 14269
rect 25317 14229 25329 14263
rect 25363 14260 25375 14263
rect 26142 14260 26148 14272
rect 25363 14232 26148 14260
rect 25363 14229 25375 14232
rect 25317 14223 25375 14229
rect 26142 14220 26148 14232
rect 26200 14260 26206 14272
rect 26697 14263 26755 14269
rect 26697 14260 26709 14263
rect 26200 14232 26709 14260
rect 26200 14220 26206 14232
rect 26697 14229 26709 14232
rect 26743 14229 26755 14263
rect 28442 14260 28448 14272
rect 28403 14232 28448 14260
rect 26697 14223 26755 14229
rect 28442 14220 28448 14232
rect 28500 14220 28506 14272
rect 31938 14260 31944 14272
rect 31899 14232 31944 14260
rect 31938 14220 31944 14232
rect 31996 14220 32002 14272
rect 32582 14260 32588 14272
rect 32543 14232 32588 14260
rect 32582 14220 32588 14232
rect 32640 14260 32646 14272
rect 33502 14260 33508 14272
rect 32640 14232 33508 14260
rect 32640 14220 32646 14232
rect 33502 14220 33508 14232
rect 33560 14220 33566 14272
rect 1104 14170 38548 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 38548 14170
rect 1104 14096 38548 14118
rect 2682 14056 2688 14068
rect 2643 14028 2688 14056
rect 2682 14016 2688 14028
rect 2740 14016 2746 14068
rect 4617 14059 4675 14065
rect 4617 14025 4629 14059
rect 4663 14056 4675 14059
rect 4706 14056 4712 14068
rect 4663 14028 4712 14056
rect 4663 14025 4675 14028
rect 4617 14019 4675 14025
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 5261 14059 5319 14065
rect 5261 14025 5273 14059
rect 5307 14056 5319 14059
rect 5442 14056 5448 14068
rect 5307 14028 5448 14056
rect 5307 14025 5319 14028
rect 5261 14019 5319 14025
rect 5442 14016 5448 14028
rect 5500 14016 5506 14068
rect 5629 14059 5687 14065
rect 5629 14025 5641 14059
rect 5675 14056 5687 14059
rect 6454 14056 6460 14068
rect 5675 14028 6460 14056
rect 5675 14025 5687 14028
rect 5629 14019 5687 14025
rect 6454 14016 6460 14028
rect 6512 14056 6518 14068
rect 7101 14059 7159 14065
rect 7101 14056 7113 14059
rect 6512 14028 7113 14056
rect 6512 14016 6518 14028
rect 7101 14025 7113 14028
rect 7147 14025 7159 14059
rect 7101 14019 7159 14025
rect 7745 14059 7803 14065
rect 7745 14025 7757 14059
rect 7791 14056 7803 14059
rect 9398 14056 9404 14068
rect 7791 14028 9404 14056
rect 7791 14025 7803 14028
rect 7745 14019 7803 14025
rect 5905 13991 5963 13997
rect 5905 13957 5917 13991
rect 5951 13988 5963 13991
rect 6914 13988 6920 14000
rect 5951 13960 6920 13988
rect 5951 13957 5963 13960
rect 5905 13951 5963 13957
rect 6914 13948 6920 13960
rect 6972 13948 6978 14000
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13920 3203 13923
rect 3191 13892 3556 13920
rect 3191 13889 3203 13892
rect 3145 13883 3203 13889
rect 2682 13812 2688 13864
rect 2740 13852 2746 13864
rect 3528 13861 3556 13892
rect 3237 13855 3295 13861
rect 3237 13852 3249 13855
rect 2740 13824 3249 13852
rect 2740 13812 2746 13824
rect 3237 13821 3249 13824
rect 3283 13821 3295 13855
rect 3237 13815 3295 13821
rect 3513 13855 3571 13861
rect 3513 13821 3525 13855
rect 3559 13852 3571 13855
rect 3970 13852 3976 13864
rect 3559 13824 3976 13852
rect 3559 13821 3571 13824
rect 3513 13815 3571 13821
rect 3970 13812 3976 13824
rect 4028 13812 4034 13864
rect 5721 13855 5779 13861
rect 5721 13821 5733 13855
rect 5767 13852 5779 13855
rect 6273 13855 6331 13861
rect 6273 13852 6285 13855
rect 5767 13824 6285 13852
rect 5767 13821 5779 13824
rect 5721 13815 5779 13821
rect 6273 13821 6285 13824
rect 6319 13852 6331 13855
rect 6641 13855 6699 13861
rect 6641 13852 6653 13855
rect 6319 13824 6653 13852
rect 6319 13821 6331 13824
rect 6273 13815 6331 13821
rect 6641 13821 6653 13824
rect 6687 13852 6699 13855
rect 6822 13852 6828 13864
rect 6687 13824 6828 13852
rect 6687 13821 6699 13824
rect 6641 13815 6699 13821
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 6917 13855 6975 13861
rect 6917 13821 6929 13855
rect 6963 13852 6975 13855
rect 7006 13852 7012 13864
rect 6963 13824 7012 13852
rect 6963 13821 6975 13824
rect 6917 13815 6975 13821
rect 7006 13812 7012 13824
rect 7064 13852 7070 13864
rect 7760 13852 7788 14019
rect 9398 14016 9404 14028
rect 9456 14016 9462 14068
rect 9585 14059 9643 14065
rect 9585 14025 9597 14059
rect 9631 14056 9643 14059
rect 10226 14056 10232 14068
rect 9631 14028 10232 14056
rect 9631 14025 9643 14028
rect 9585 14019 9643 14025
rect 9214 13920 9220 13932
rect 9175 13892 9220 13920
rect 9214 13880 9220 13892
rect 9272 13880 9278 13932
rect 7064 13824 7788 13852
rect 8389 13855 8447 13861
rect 7064 13812 7070 13824
rect 8389 13821 8401 13855
rect 8435 13852 8447 13855
rect 8757 13855 8815 13861
rect 8757 13852 8769 13855
rect 8435 13824 8769 13852
rect 8435 13821 8447 13824
rect 8389 13815 8447 13821
rect 8757 13821 8769 13824
rect 8803 13852 8815 13855
rect 9600 13852 9628 14019
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 10318 14016 10324 14068
rect 10376 14056 10382 14068
rect 10870 14056 10876 14068
rect 10376 14028 10876 14056
rect 10376 14016 10382 14028
rect 10870 14016 10876 14028
rect 10928 14016 10934 14068
rect 12253 14059 12311 14065
rect 12253 14025 12265 14059
rect 12299 14056 12311 14059
rect 13354 14056 13360 14068
rect 12299 14028 13360 14056
rect 12299 14025 12311 14028
rect 12253 14019 12311 14025
rect 13354 14016 13360 14028
rect 13412 14016 13418 14068
rect 15378 14056 15384 14068
rect 15339 14028 15384 14056
rect 15378 14016 15384 14028
rect 15436 14016 15442 14068
rect 15930 14056 15936 14068
rect 15891 14028 15936 14056
rect 15930 14016 15936 14028
rect 15988 14016 15994 14068
rect 16574 14065 16580 14068
rect 16558 14059 16580 14065
rect 16558 14025 16570 14059
rect 16558 14019 16580 14025
rect 16574 14016 16580 14019
rect 16632 14016 16638 14068
rect 18046 14016 18052 14068
rect 18104 14056 18110 14068
rect 18417 14059 18475 14065
rect 18417 14056 18429 14059
rect 18104 14028 18429 14056
rect 18104 14016 18110 14028
rect 18417 14025 18429 14028
rect 18463 14025 18475 14059
rect 18417 14019 18475 14025
rect 18690 14016 18696 14068
rect 18748 14056 18754 14068
rect 18877 14059 18935 14065
rect 18877 14056 18889 14059
rect 18748 14028 18889 14056
rect 18748 14016 18754 14028
rect 18877 14025 18889 14028
rect 18923 14056 18935 14059
rect 19245 14059 19303 14065
rect 19245 14056 19257 14059
rect 18923 14028 19257 14056
rect 18923 14025 18935 14028
rect 18877 14019 18935 14025
rect 19245 14025 19257 14028
rect 19291 14025 19303 14059
rect 19245 14019 19303 14025
rect 19334 14016 19340 14068
rect 19392 14056 19398 14068
rect 19981 14059 20039 14065
rect 19981 14056 19993 14059
rect 19392 14028 19993 14056
rect 19392 14016 19398 14028
rect 19981 14025 19993 14028
rect 20027 14025 20039 14059
rect 19981 14019 20039 14025
rect 20162 14016 20168 14068
rect 20220 14056 20226 14068
rect 20349 14059 20407 14065
rect 20349 14056 20361 14059
rect 20220 14028 20361 14056
rect 20220 14016 20226 14028
rect 20349 14025 20361 14028
rect 20395 14025 20407 14059
rect 20990 14056 20996 14068
rect 20951 14028 20996 14056
rect 20349 14019 20407 14025
rect 20990 14016 20996 14028
rect 21048 14016 21054 14068
rect 23106 14056 23112 14068
rect 23067 14028 23112 14056
rect 23106 14016 23112 14028
rect 23164 14016 23170 14068
rect 24029 14059 24087 14065
rect 24029 14025 24041 14059
rect 24075 14056 24087 14059
rect 24302 14056 24308 14068
rect 24075 14028 24308 14056
rect 24075 14025 24087 14028
rect 24029 14019 24087 14025
rect 24302 14016 24308 14028
rect 24360 14016 24366 14068
rect 25501 14059 25559 14065
rect 25501 14025 25513 14059
rect 25547 14056 25559 14059
rect 25958 14056 25964 14068
rect 25547 14028 25964 14056
rect 25547 14025 25559 14028
rect 25501 14019 25559 14025
rect 25958 14016 25964 14028
rect 26016 14016 26022 14068
rect 26142 14065 26148 14068
rect 26126 14059 26148 14065
rect 26126 14025 26138 14059
rect 26126 14019 26148 14025
rect 26142 14016 26148 14019
rect 26200 14016 26206 14068
rect 26602 14056 26608 14068
rect 26563 14028 26608 14056
rect 26602 14016 26608 14028
rect 26660 14016 26666 14068
rect 26786 14016 26792 14068
rect 26844 14056 26850 14068
rect 26973 14059 27031 14065
rect 26973 14056 26985 14059
rect 26844 14028 26985 14056
rect 26844 14016 26850 14028
rect 26973 14025 26985 14028
rect 27019 14025 27031 14059
rect 26973 14019 27031 14025
rect 27709 14059 27767 14065
rect 27709 14025 27721 14059
rect 27755 14056 27767 14059
rect 27798 14056 27804 14068
rect 27755 14028 27804 14056
rect 27755 14025 27767 14028
rect 27709 14019 27767 14025
rect 27798 14016 27804 14028
rect 27856 14016 27862 14068
rect 28258 14016 28264 14068
rect 28316 14056 28322 14068
rect 28445 14059 28503 14065
rect 28445 14056 28457 14059
rect 28316 14028 28457 14056
rect 28316 14016 28322 14028
rect 28445 14025 28457 14028
rect 28491 14025 28503 14059
rect 28445 14019 28503 14025
rect 29822 14016 29828 14068
rect 29880 14056 29886 14068
rect 30466 14056 30472 14068
rect 29880 14028 30472 14056
rect 29880 14016 29886 14028
rect 30466 14016 30472 14028
rect 30524 14056 30530 14068
rect 30653 14059 30711 14065
rect 30653 14056 30665 14059
rect 30524 14028 30665 14056
rect 30524 14016 30530 14028
rect 30653 14025 30665 14028
rect 30699 14056 30711 14059
rect 31754 14056 31760 14068
rect 30699 14028 31760 14056
rect 30699 14025 30711 14028
rect 30653 14019 30711 14025
rect 31754 14016 31760 14028
rect 31812 14016 31818 14068
rect 32122 14016 32128 14068
rect 32180 14056 32186 14068
rect 32217 14059 32275 14065
rect 32217 14056 32229 14059
rect 32180 14028 32229 14056
rect 32180 14016 32186 14028
rect 32217 14025 32229 14028
rect 32263 14025 32275 14059
rect 32217 14019 32275 14025
rect 34146 14016 34152 14068
rect 34204 14056 34210 14068
rect 34517 14059 34575 14065
rect 34517 14056 34529 14059
rect 34204 14028 34529 14056
rect 34204 14016 34210 14028
rect 34517 14025 34529 14028
rect 34563 14025 34575 14059
rect 34517 14019 34575 14025
rect 12066 13948 12072 14000
rect 12124 13988 12130 14000
rect 13265 13991 13323 13997
rect 13265 13988 13277 13991
rect 12124 13960 13277 13988
rect 12124 13948 12130 13960
rect 13265 13957 13277 13960
rect 13311 13957 13323 13991
rect 13265 13951 13323 13957
rect 15102 13948 15108 14000
rect 15160 13988 15166 14000
rect 16666 13988 16672 14000
rect 15160 13960 16344 13988
rect 16627 13960 16672 13988
rect 15160 13948 15166 13960
rect 10781 13923 10839 13929
rect 10781 13889 10793 13923
rect 10827 13920 10839 13923
rect 11054 13920 11060 13932
rect 10827 13892 11060 13920
rect 10827 13889 10839 13892
rect 10781 13883 10839 13889
rect 11054 13880 11060 13892
rect 11112 13880 11118 13932
rect 11422 13880 11428 13932
rect 11480 13920 11486 13932
rect 11698 13920 11704 13932
rect 11480 13892 11704 13920
rect 11480 13880 11486 13892
rect 11698 13880 11704 13892
rect 11756 13880 11762 13932
rect 13173 13923 13231 13929
rect 13173 13889 13185 13923
rect 13219 13920 13231 13923
rect 13633 13923 13691 13929
rect 13633 13920 13645 13923
rect 13219 13892 13645 13920
rect 13219 13889 13231 13892
rect 13173 13883 13231 13889
rect 13633 13889 13645 13892
rect 13679 13920 13691 13923
rect 13722 13920 13728 13932
rect 13679 13892 13728 13920
rect 13679 13889 13691 13892
rect 13633 13883 13691 13889
rect 13722 13880 13728 13892
rect 13780 13880 13786 13932
rect 14737 13923 14795 13929
rect 14737 13889 14749 13923
rect 14783 13920 14795 13923
rect 16316 13920 16344 13960
rect 16666 13948 16672 13960
rect 16724 13948 16730 14000
rect 19134 13991 19192 13997
rect 16776 13960 17816 13988
rect 16776 13929 16804 13960
rect 16761 13923 16819 13929
rect 16761 13920 16773 13923
rect 14783 13892 15240 13920
rect 16316 13892 16773 13920
rect 14783 13889 14795 13892
rect 14737 13883 14795 13889
rect 15212 13864 15240 13892
rect 16761 13889 16773 13892
rect 16807 13889 16819 13923
rect 16761 13883 16819 13889
rect 16850 13880 16856 13932
rect 16908 13920 16914 13932
rect 16908 13892 16953 13920
rect 16908 13880 16914 13892
rect 10962 13852 10968 13864
rect 8803 13824 9628 13852
rect 10875 13824 10968 13852
rect 8803 13821 8815 13824
rect 8757 13815 8815 13821
rect 10962 13812 10968 13824
rect 11020 13852 11026 13864
rect 11793 13855 11851 13861
rect 11793 13852 11805 13855
rect 11020 13824 11805 13852
rect 11020 13812 11026 13824
rect 11793 13821 11805 13824
rect 11839 13821 11851 13855
rect 11793 13815 11851 13821
rect 12526 13812 12532 13864
rect 12584 13852 12590 13864
rect 12621 13855 12679 13861
rect 12621 13852 12633 13855
rect 12584 13824 12633 13852
rect 12584 13812 12590 13824
rect 12621 13821 12633 13824
rect 12667 13852 12679 13855
rect 13909 13855 13967 13861
rect 12667 13824 13216 13852
rect 12667 13821 12679 13824
rect 12621 13815 12679 13821
rect 8018 13744 8024 13796
rect 8076 13784 8082 13796
rect 8481 13787 8539 13793
rect 8481 13784 8493 13787
rect 8076 13756 8493 13784
rect 8076 13744 8082 13756
rect 8481 13753 8493 13756
rect 8527 13784 8539 13787
rect 8570 13784 8576 13796
rect 8527 13756 8576 13784
rect 8527 13753 8539 13756
rect 8481 13747 8539 13753
rect 8570 13744 8576 13756
rect 8628 13744 8634 13796
rect 8849 13787 8907 13793
rect 8849 13753 8861 13787
rect 8895 13784 8907 13787
rect 9306 13784 9312 13796
rect 8895 13756 9312 13784
rect 8895 13753 8907 13756
rect 8849 13747 8907 13753
rect 9306 13744 9312 13756
rect 9364 13744 9370 13796
rect 10045 13787 10103 13793
rect 10045 13753 10057 13787
rect 10091 13753 10103 13787
rect 10045 13747 10103 13753
rect 10413 13787 10471 13793
rect 10413 13753 10425 13787
rect 10459 13784 10471 13787
rect 10980 13784 11008 13812
rect 10459 13756 11008 13784
rect 10459 13753 10471 13756
rect 10413 13747 10471 13753
rect 8662 13716 8668 13728
rect 8623 13688 8668 13716
rect 8662 13676 8668 13688
rect 8720 13676 8726 13728
rect 9858 13716 9864 13728
rect 9819 13688 9864 13716
rect 9858 13676 9864 13688
rect 9916 13716 9922 13728
rect 10060 13716 10088 13747
rect 10226 13716 10232 13728
rect 9916 13688 10088 13716
rect 10187 13688 10232 13716
rect 9916 13676 9922 13688
rect 10226 13676 10232 13688
rect 10284 13676 10290 13728
rect 10321 13719 10379 13725
rect 10321 13685 10333 13719
rect 10367 13716 10379 13719
rect 11146 13716 11152 13728
rect 10367 13688 11152 13716
rect 10367 13685 10379 13688
rect 10321 13679 10379 13685
rect 11146 13676 11152 13688
rect 11204 13676 11210 13728
rect 11330 13676 11336 13728
rect 11388 13716 11394 13728
rect 11517 13719 11575 13725
rect 11517 13716 11529 13719
rect 11388 13688 11529 13716
rect 11388 13676 11394 13688
rect 11517 13685 11529 13688
rect 11563 13716 11575 13719
rect 11698 13716 11704 13728
rect 11563 13688 11704 13716
rect 11563 13685 11575 13688
rect 11517 13679 11575 13685
rect 11698 13676 11704 13688
rect 11756 13676 11762 13728
rect 12805 13719 12863 13725
rect 12805 13685 12817 13719
rect 12851 13716 12863 13719
rect 12894 13716 12900 13728
rect 12851 13688 12900 13716
rect 12851 13685 12863 13688
rect 12805 13679 12863 13685
rect 12894 13676 12900 13688
rect 12952 13676 12958 13728
rect 13188 13716 13216 13824
rect 13909 13821 13921 13855
rect 13955 13852 13967 13855
rect 14090 13852 14096 13864
rect 13955 13824 14096 13852
rect 13955 13821 13967 13824
rect 13909 13815 13967 13821
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 15194 13852 15200 13864
rect 15155 13824 15200 13852
rect 15194 13812 15200 13824
rect 15252 13812 15258 13864
rect 16206 13812 16212 13864
rect 16264 13852 16270 13864
rect 16393 13855 16451 13861
rect 16393 13852 16405 13855
rect 16264 13824 16405 13852
rect 16264 13812 16270 13824
rect 16393 13821 16405 13824
rect 16439 13821 16451 13855
rect 16393 13815 16451 13821
rect 17678 13812 17684 13864
rect 17736 13812 17742 13864
rect 17788 13852 17816 13960
rect 19134 13957 19146 13991
rect 19180 13988 19192 13991
rect 19180 13960 20484 13988
rect 19180 13957 19192 13960
rect 19134 13951 19192 13957
rect 19242 13880 19248 13932
rect 19300 13920 19306 13932
rect 19337 13923 19395 13929
rect 19337 13920 19349 13923
rect 19300 13892 19349 13920
rect 19300 13880 19306 13892
rect 19337 13889 19349 13892
rect 19383 13920 19395 13923
rect 20254 13920 20260 13932
rect 19383 13892 20260 13920
rect 19383 13889 19395 13892
rect 19337 13883 19395 13889
rect 20254 13880 20260 13892
rect 20312 13880 20318 13932
rect 18966 13852 18972 13864
rect 17788 13824 18000 13852
rect 18927 13824 18972 13852
rect 13265 13787 13323 13793
rect 13265 13753 13277 13787
rect 13311 13784 13323 13787
rect 13541 13787 13599 13793
rect 13541 13784 13553 13787
rect 13311 13756 13553 13784
rect 13311 13753 13323 13756
rect 13265 13747 13323 13753
rect 13541 13753 13553 13756
rect 13587 13784 13599 13787
rect 14001 13787 14059 13793
rect 14001 13784 14013 13787
rect 13587 13756 14013 13784
rect 13587 13753 13599 13756
rect 13541 13747 13599 13753
rect 14001 13753 14013 13756
rect 14047 13753 14059 13787
rect 14001 13747 14059 13753
rect 14369 13787 14427 13793
rect 14369 13753 14381 13787
rect 14415 13784 14427 13787
rect 14918 13784 14924 13796
rect 14415 13756 14924 13784
rect 14415 13753 14427 13756
rect 14369 13747 14427 13753
rect 13722 13716 13728 13728
rect 13188 13688 13728 13716
rect 13722 13676 13728 13688
rect 13780 13716 13786 13728
rect 13817 13719 13875 13725
rect 13817 13716 13829 13719
rect 13780 13688 13829 13716
rect 13780 13676 13786 13688
rect 13817 13685 13829 13688
rect 13863 13685 13875 13719
rect 14016 13716 14044 13747
rect 14918 13744 14924 13756
rect 14976 13744 14982 13796
rect 15105 13787 15163 13793
rect 15105 13753 15117 13787
rect 15151 13784 15163 13787
rect 15470 13784 15476 13796
rect 15151 13756 15476 13784
rect 15151 13753 15163 13756
rect 15105 13747 15163 13753
rect 15470 13744 15476 13756
rect 15528 13744 15534 13796
rect 17310 13744 17316 13796
rect 17368 13784 17374 13796
rect 17696 13784 17724 13812
rect 17972 13784 18000 13824
rect 18966 13812 18972 13824
rect 19024 13812 19030 13864
rect 19705 13855 19763 13861
rect 19705 13852 19717 13855
rect 19352 13824 19717 13852
rect 18598 13784 18604 13796
rect 17368 13756 17908 13784
rect 17972 13756 18604 13784
rect 17368 13744 17374 13756
rect 14182 13716 14188 13728
rect 14016 13688 14188 13716
rect 13817 13679 13875 13685
rect 14182 13676 14188 13688
rect 14240 13716 14246 13728
rect 15838 13716 15844 13728
rect 14240 13688 15844 13716
rect 14240 13676 14246 13688
rect 15838 13676 15844 13688
rect 15896 13676 15902 13728
rect 17681 13719 17739 13725
rect 17681 13685 17693 13719
rect 17727 13716 17739 13719
rect 17770 13716 17776 13728
rect 17727 13688 17776 13716
rect 17727 13685 17739 13688
rect 17681 13679 17739 13685
rect 17770 13676 17776 13688
rect 17828 13676 17834 13728
rect 17880 13716 17908 13756
rect 18598 13744 18604 13756
rect 18656 13744 18662 13796
rect 19058 13744 19064 13796
rect 19116 13784 19122 13796
rect 19352 13784 19380 13824
rect 19705 13821 19717 13824
rect 19751 13821 19763 13855
rect 20456 13852 20484 13960
rect 21358 13948 21364 14000
rect 21416 13988 21422 14000
rect 22373 13991 22431 13997
rect 22373 13988 22385 13991
rect 21416 13960 22385 13988
rect 21416 13948 21422 13960
rect 22373 13957 22385 13960
rect 22419 13957 22431 13991
rect 25866 13988 25872 14000
rect 25779 13960 25872 13988
rect 22373 13951 22431 13957
rect 25866 13948 25872 13960
rect 25924 13988 25930 14000
rect 26237 13991 26295 13997
rect 26237 13988 26249 13991
rect 25924 13960 26249 13988
rect 25924 13948 25930 13960
rect 26237 13957 26249 13960
rect 26283 13988 26295 13991
rect 26510 13988 26516 14000
rect 26283 13960 26516 13988
rect 26283 13957 26295 13960
rect 26237 13951 26295 13957
rect 26510 13948 26516 13960
rect 26568 13948 26574 14000
rect 29914 13948 29920 14000
rect 29972 13988 29978 14000
rect 30285 13991 30343 13997
rect 30285 13988 30297 13991
rect 29972 13960 30297 13988
rect 29972 13948 29978 13960
rect 30285 13957 30297 13960
rect 30331 13957 30343 13991
rect 30285 13951 30343 13957
rect 31938 13948 31944 14000
rect 31996 13948 32002 14000
rect 24026 13880 24032 13932
rect 24084 13920 24090 13932
rect 24084 13892 24532 13920
rect 24084 13880 24090 13892
rect 20533 13855 20591 13861
rect 20533 13852 20545 13855
rect 20456 13824 20545 13852
rect 19705 13815 19763 13821
rect 20533 13821 20545 13824
rect 20579 13852 20591 13855
rect 20622 13852 20628 13864
rect 20579 13824 20628 13852
rect 20579 13821 20591 13824
rect 20533 13815 20591 13821
rect 20622 13812 20628 13824
rect 20680 13812 20686 13864
rect 21637 13855 21695 13861
rect 21637 13821 21649 13855
rect 21683 13821 21695 13855
rect 21637 13815 21695 13821
rect 19116 13756 19380 13784
rect 19116 13744 19122 13756
rect 20717 13719 20775 13725
rect 20717 13716 20729 13719
rect 17880 13688 20729 13716
rect 20717 13685 20729 13688
rect 20763 13685 20775 13719
rect 20717 13679 20775 13685
rect 21453 13719 21511 13725
rect 21453 13685 21465 13719
rect 21499 13716 21511 13719
rect 21652 13716 21680 13815
rect 21726 13812 21732 13864
rect 21784 13852 21790 13864
rect 21913 13855 21971 13861
rect 21913 13852 21925 13855
rect 21784 13824 21925 13852
rect 21784 13812 21790 13824
rect 21913 13821 21925 13824
rect 21959 13821 21971 13855
rect 21913 13815 21971 13821
rect 22465 13855 22523 13861
rect 22465 13821 22477 13855
rect 22511 13852 22523 13855
rect 22554 13852 22560 13864
rect 22511 13824 22560 13852
rect 22511 13821 22523 13824
rect 22465 13815 22523 13821
rect 22554 13812 22560 13824
rect 22612 13812 22618 13864
rect 24394 13852 24400 13864
rect 24355 13824 24400 13852
rect 24394 13812 24400 13824
rect 24452 13812 24458 13864
rect 24504 13861 24532 13892
rect 25406 13880 25412 13932
rect 25464 13920 25470 13932
rect 26326 13920 26332 13932
rect 25464 13892 26332 13920
rect 25464 13880 25470 13892
rect 26326 13880 26332 13892
rect 26384 13880 26390 13932
rect 24489 13855 24547 13861
rect 24489 13821 24501 13855
rect 24535 13852 24547 13855
rect 25958 13852 25964 13864
rect 24535 13824 24808 13852
rect 25919 13824 25964 13852
rect 24535 13821 24547 13824
rect 24489 13815 24547 13821
rect 24780 13784 24808 13824
rect 25958 13812 25964 13824
rect 26016 13852 26022 13864
rect 26694 13852 26700 13864
rect 26016 13824 26700 13852
rect 26016 13812 26022 13824
rect 26694 13812 26700 13824
rect 26752 13812 26758 13864
rect 27430 13852 27436 13864
rect 27391 13824 27436 13852
rect 27430 13812 27436 13824
rect 27488 13852 27494 13864
rect 27525 13855 27583 13861
rect 27525 13852 27537 13855
rect 27488 13824 27537 13852
rect 27488 13812 27494 13824
rect 27525 13821 27537 13824
rect 27571 13821 27583 13855
rect 27525 13815 27583 13821
rect 28169 13855 28227 13861
rect 28169 13821 28181 13855
rect 28215 13852 28227 13855
rect 28442 13852 28448 13864
rect 28215 13824 28448 13852
rect 28215 13821 28227 13824
rect 28169 13815 28227 13821
rect 28442 13812 28448 13824
rect 28500 13852 28506 13864
rect 29270 13852 29276 13864
rect 28500 13824 29276 13852
rect 28500 13812 28506 13824
rect 29270 13812 29276 13824
rect 29328 13812 29334 13864
rect 29454 13852 29460 13864
rect 29415 13824 29460 13852
rect 29454 13812 29460 13824
rect 29512 13812 29518 13864
rect 29549 13855 29607 13861
rect 29549 13821 29561 13855
rect 29595 13852 29607 13855
rect 29932 13852 29960 13948
rect 31481 13923 31539 13929
rect 31481 13889 31493 13923
rect 31527 13920 31539 13923
rect 31956 13920 31984 13948
rect 34149 13923 34207 13929
rect 34149 13920 34161 13923
rect 31527 13892 31984 13920
rect 33612 13892 34161 13920
rect 31527 13889 31539 13892
rect 31481 13883 31539 13889
rect 33612 13864 33640 13892
rect 34149 13889 34161 13892
rect 34195 13889 34207 13923
rect 34149 13883 34207 13889
rect 30926 13852 30932 13864
rect 29595 13824 29960 13852
rect 30887 13824 30932 13852
rect 29595 13821 29607 13824
rect 29549 13815 29607 13821
rect 30926 13812 30932 13824
rect 30984 13812 30990 13864
rect 31386 13812 31392 13864
rect 31444 13852 31450 13864
rect 31757 13855 31815 13861
rect 31757 13852 31769 13855
rect 31444 13824 31769 13852
rect 31444 13812 31450 13824
rect 31757 13821 31769 13824
rect 31803 13821 31815 13855
rect 31941 13855 31999 13861
rect 31941 13852 31953 13855
rect 31757 13815 31815 13821
rect 31864 13824 31953 13852
rect 25038 13784 25044 13796
rect 24780 13756 25044 13784
rect 25038 13744 25044 13756
rect 25096 13744 25102 13796
rect 27890 13744 27896 13796
rect 27948 13784 27954 13796
rect 28810 13784 28816 13796
rect 27948 13756 28816 13784
rect 27948 13744 27954 13756
rect 28810 13744 28816 13756
rect 28868 13784 28874 13796
rect 28997 13787 29055 13793
rect 28997 13784 29009 13787
rect 28868 13756 29009 13784
rect 28868 13744 28874 13756
rect 28997 13753 29009 13756
rect 29043 13753 29055 13787
rect 29641 13787 29699 13793
rect 29641 13784 29653 13787
rect 28997 13747 29055 13753
rect 29380 13756 29653 13784
rect 21818 13716 21824 13728
rect 21499 13688 21824 13716
rect 21499 13685 21511 13688
rect 21453 13679 21511 13685
rect 21818 13676 21824 13688
rect 21876 13676 21882 13728
rect 23477 13719 23535 13725
rect 23477 13685 23489 13719
rect 23523 13716 23535 13719
rect 23750 13716 23756 13728
rect 23523 13688 23756 13716
rect 23523 13685 23535 13688
rect 23477 13679 23535 13685
rect 23750 13676 23756 13688
rect 23808 13716 23814 13728
rect 24210 13716 24216 13728
rect 23808 13688 24216 13716
rect 23808 13676 23814 13688
rect 24210 13676 24216 13688
rect 24268 13676 24274 13728
rect 29012 13716 29040 13747
rect 29380 13716 29408 13756
rect 29641 13753 29653 13756
rect 29687 13753 29699 13787
rect 30006 13784 30012 13796
rect 29967 13756 30012 13784
rect 29641 13747 29699 13753
rect 30006 13744 30012 13756
rect 30064 13744 30070 13796
rect 31570 13744 31576 13796
rect 31628 13784 31634 13796
rect 31864 13784 31892 13824
rect 31941 13821 31953 13824
rect 31987 13852 31999 13855
rect 32582 13852 32588 13864
rect 31987 13824 32588 13852
rect 31987 13821 31999 13824
rect 31941 13815 31999 13821
rect 32582 13812 32588 13824
rect 32640 13812 32646 13864
rect 32677 13855 32735 13861
rect 32677 13821 32689 13855
rect 32723 13852 32735 13855
rect 32769 13855 32827 13861
rect 32769 13852 32781 13855
rect 32723 13824 32781 13852
rect 32723 13821 32735 13824
rect 32677 13815 32735 13821
rect 32769 13821 32781 13824
rect 32815 13852 32827 13855
rect 32858 13852 32864 13864
rect 32815 13824 32864 13852
rect 32815 13821 32827 13824
rect 32769 13815 32827 13821
rect 32858 13812 32864 13824
rect 32916 13812 32922 13864
rect 33134 13852 33140 13864
rect 33095 13824 33140 13852
rect 33134 13812 33140 13824
rect 33192 13812 33198 13864
rect 33594 13852 33600 13864
rect 33555 13824 33600 13852
rect 33594 13812 33600 13824
rect 33652 13812 33658 13864
rect 33873 13855 33931 13861
rect 33873 13821 33885 13855
rect 33919 13852 33931 13855
rect 34422 13852 34428 13864
rect 33919 13824 34428 13852
rect 33919 13821 33931 13824
rect 33873 13815 33931 13821
rect 34422 13812 34428 13824
rect 34480 13812 34486 13864
rect 31628 13756 31892 13784
rect 31628 13744 31634 13756
rect 29012 13688 29408 13716
rect 1104 13626 38548 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 38548 13626
rect 1104 13552 38548 13574
rect 5258 13512 5264 13524
rect 5219 13484 5264 13512
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 5626 13512 5632 13524
rect 5587 13484 5632 13512
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 6914 13472 6920 13524
rect 6972 13512 6978 13524
rect 7469 13515 7527 13521
rect 7469 13512 7481 13515
rect 6972 13484 7481 13512
rect 6972 13472 6978 13484
rect 7469 13481 7481 13484
rect 7515 13512 7527 13515
rect 8110 13512 8116 13524
rect 7515 13484 8116 13512
rect 7515 13481 7527 13484
rect 7469 13475 7527 13481
rect 8110 13472 8116 13484
rect 8168 13472 8174 13524
rect 8205 13515 8263 13521
rect 8205 13481 8217 13515
rect 8251 13512 8263 13515
rect 8662 13512 8668 13524
rect 8251 13484 8668 13512
rect 8251 13481 8263 13484
rect 8205 13475 8263 13481
rect 8662 13472 8668 13484
rect 8720 13472 8726 13524
rect 9493 13515 9551 13521
rect 9493 13481 9505 13515
rect 9539 13512 9551 13515
rect 9766 13512 9772 13524
rect 9539 13484 9772 13512
rect 9539 13481 9551 13484
rect 9493 13475 9551 13481
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 10505 13515 10563 13521
rect 10505 13512 10517 13515
rect 10008 13484 10517 13512
rect 10008 13472 10014 13484
rect 10505 13481 10517 13484
rect 10551 13481 10563 13515
rect 10505 13475 10563 13481
rect 11057 13515 11115 13521
rect 11057 13481 11069 13515
rect 11103 13512 11115 13515
rect 11698 13512 11704 13524
rect 11103 13484 11704 13512
rect 11103 13481 11115 13484
rect 11057 13475 11115 13481
rect 3050 13444 3056 13456
rect 3011 13416 3056 13444
rect 3050 13404 3056 13416
rect 3108 13404 3114 13456
rect 1394 13376 1400 13388
rect 1355 13348 1400 13376
rect 1394 13336 1400 13348
rect 1452 13336 1458 13388
rect 5629 13379 5687 13385
rect 5629 13345 5641 13379
rect 5675 13376 5687 13379
rect 5718 13376 5724 13388
rect 5675 13348 5724 13376
rect 5675 13345 5687 13348
rect 5629 13339 5687 13345
rect 5718 13336 5724 13348
rect 5776 13376 5782 13388
rect 5902 13376 5908 13388
rect 5776 13348 5908 13376
rect 5776 13336 5782 13348
rect 5902 13336 5908 13348
rect 5960 13336 5966 13388
rect 6178 13376 6184 13388
rect 6139 13348 6184 13376
rect 6178 13336 6184 13348
rect 6236 13336 6242 13388
rect 6365 13379 6423 13385
rect 6365 13345 6377 13379
rect 6411 13376 6423 13379
rect 6454 13376 6460 13388
rect 6411 13348 6460 13376
rect 6411 13345 6423 13348
rect 6365 13339 6423 13345
rect 6454 13336 6460 13348
rect 6512 13376 6518 13388
rect 6932 13376 6960 13472
rect 7006 13404 7012 13456
rect 7064 13444 7070 13456
rect 8386 13444 8392 13456
rect 7064 13416 7109 13444
rect 8347 13416 8392 13444
rect 7064 13404 7070 13416
rect 8386 13404 8392 13416
rect 8444 13404 8450 13456
rect 10520 13444 10548 13475
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 12710 13472 12716 13524
rect 12768 13512 12774 13524
rect 13446 13512 13452 13524
rect 12768 13484 13452 13512
rect 12768 13472 12774 13484
rect 13446 13472 13452 13484
rect 13504 13472 13510 13524
rect 13906 13512 13912 13524
rect 13867 13484 13912 13512
rect 13906 13472 13912 13484
rect 13964 13472 13970 13524
rect 14366 13512 14372 13524
rect 14327 13484 14372 13512
rect 14366 13472 14372 13484
rect 14424 13472 14430 13524
rect 14737 13515 14795 13521
rect 14737 13481 14749 13515
rect 14783 13512 14795 13515
rect 15102 13512 15108 13524
rect 14783 13484 15108 13512
rect 14783 13481 14795 13484
rect 14737 13475 14795 13481
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 16485 13515 16543 13521
rect 16485 13481 16497 13515
rect 16531 13512 16543 13515
rect 17126 13512 17132 13524
rect 16531 13484 17132 13512
rect 16531 13481 16543 13484
rect 16485 13475 16543 13481
rect 17126 13472 17132 13484
rect 17184 13512 17190 13524
rect 17184 13484 17448 13512
rect 17184 13472 17190 13484
rect 10686 13444 10692 13456
rect 10520 13416 10692 13444
rect 10686 13404 10692 13416
rect 10744 13444 10750 13456
rect 10873 13447 10931 13453
rect 10873 13444 10885 13447
rect 10744 13416 10885 13444
rect 10744 13404 10750 13416
rect 10873 13413 10885 13416
rect 10919 13413 10931 13447
rect 10873 13407 10931 13413
rect 11241 13447 11299 13453
rect 11241 13413 11253 13447
rect 11287 13444 11299 13447
rect 12342 13444 12348 13456
rect 11287 13416 12348 13444
rect 11287 13413 11299 13416
rect 11241 13407 11299 13413
rect 12342 13404 12348 13416
rect 12400 13404 12406 13456
rect 14090 13404 14096 13456
rect 14148 13444 14154 13456
rect 15930 13444 15936 13456
rect 14148 13416 15936 13444
rect 14148 13404 14154 13416
rect 15930 13404 15936 13416
rect 15988 13404 15994 13456
rect 16022 13404 16028 13456
rect 16080 13444 16086 13456
rect 16574 13444 16580 13456
rect 16080 13416 16580 13444
rect 16080 13404 16086 13416
rect 16574 13404 16580 13416
rect 16632 13404 16638 13456
rect 16669 13447 16727 13453
rect 16669 13413 16681 13447
rect 16715 13444 16727 13447
rect 16758 13444 16764 13456
rect 16715 13416 16764 13444
rect 16715 13413 16727 13416
rect 16669 13407 16727 13413
rect 16758 13404 16764 13416
rect 16816 13404 16822 13456
rect 7926 13376 7932 13388
rect 6512 13348 6960 13376
rect 7839 13348 7932 13376
rect 6512 13336 6518 13348
rect 7926 13336 7932 13348
rect 7984 13376 7990 13388
rect 8297 13379 8355 13385
rect 8297 13376 8309 13379
rect 7984 13348 8309 13376
rect 7984 13336 7990 13348
rect 8297 13345 8309 13348
rect 8343 13376 8355 13379
rect 9677 13379 9735 13385
rect 8343 13348 8984 13376
rect 8343 13345 8355 13348
rect 8297 13339 8355 13345
rect 1578 13268 1584 13320
rect 1636 13308 1642 13320
rect 1673 13311 1731 13317
rect 1673 13308 1685 13311
rect 1636 13280 1685 13308
rect 1636 13268 1642 13280
rect 1673 13277 1685 13280
rect 1719 13277 1731 13311
rect 8018 13308 8024 13320
rect 7979 13280 8024 13308
rect 1673 13271 1731 13277
rect 8018 13268 8024 13280
rect 8076 13268 8082 13320
rect 8754 13308 8760 13320
rect 8715 13280 8760 13308
rect 8754 13268 8760 13280
rect 8812 13268 8818 13320
rect 8956 13308 8984 13348
rect 9677 13345 9689 13379
rect 9723 13376 9735 13379
rect 9858 13376 9864 13388
rect 9723 13348 9864 13376
rect 9723 13345 9735 13348
rect 9677 13339 9735 13345
rect 9858 13336 9864 13348
rect 9916 13376 9922 13388
rect 10318 13376 10324 13388
rect 9916 13348 10324 13376
rect 9916 13336 9922 13348
rect 10318 13336 10324 13348
rect 10376 13336 10382 13388
rect 11146 13376 11152 13388
rect 11059 13348 11152 13376
rect 11146 13336 11152 13348
rect 11204 13376 11210 13388
rect 11974 13376 11980 13388
rect 11204 13348 11980 13376
rect 11204 13336 11210 13348
rect 11974 13336 11980 13348
rect 12032 13336 12038 13388
rect 12710 13376 12716 13388
rect 12671 13348 12716 13376
rect 12710 13336 12716 13348
rect 12768 13336 12774 13388
rect 12894 13376 12900 13388
rect 12855 13348 12900 13376
rect 12894 13336 12900 13348
rect 12952 13336 12958 13388
rect 13078 13336 13084 13388
rect 13136 13376 13142 13388
rect 13265 13379 13323 13385
rect 13265 13376 13277 13379
rect 13136 13348 13277 13376
rect 13136 13336 13142 13348
rect 13265 13345 13277 13348
rect 13311 13376 13323 13379
rect 13722 13376 13728 13388
rect 13311 13348 13728 13376
rect 13311 13345 13323 13348
rect 13265 13339 13323 13345
rect 13722 13336 13728 13348
rect 13780 13336 13786 13388
rect 14182 13336 14188 13388
rect 14240 13376 14246 13388
rect 14734 13376 14740 13388
rect 14240 13348 14740 13376
rect 14240 13336 14246 13348
rect 14734 13336 14740 13348
rect 14792 13336 14798 13388
rect 15289 13379 15347 13385
rect 15289 13345 15301 13379
rect 15335 13376 15347 13379
rect 15378 13376 15384 13388
rect 15335 13348 15384 13376
rect 15335 13345 15347 13348
rect 15289 13339 15347 13345
rect 15378 13336 15384 13348
rect 15436 13336 15442 13388
rect 16301 13379 16359 13385
rect 16301 13345 16313 13379
rect 16347 13376 16359 13379
rect 17310 13376 17316 13388
rect 16347 13348 17316 13376
rect 16347 13345 16359 13348
rect 16301 13339 16359 13345
rect 17310 13336 17316 13348
rect 17368 13336 17374 13388
rect 17420 13385 17448 13484
rect 17494 13472 17500 13524
rect 17552 13512 17558 13524
rect 18141 13515 18199 13521
rect 18141 13512 18153 13515
rect 17552 13484 18153 13512
rect 17552 13472 17558 13484
rect 18141 13481 18153 13484
rect 18187 13481 18199 13515
rect 18141 13475 18199 13481
rect 19061 13515 19119 13521
rect 19061 13481 19073 13515
rect 19107 13512 19119 13515
rect 19242 13512 19248 13524
rect 19107 13484 19248 13512
rect 19107 13481 19119 13484
rect 19061 13475 19119 13481
rect 19242 13472 19248 13484
rect 19300 13472 19306 13524
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 19889 13515 19947 13521
rect 19889 13512 19901 13515
rect 19392 13484 19901 13512
rect 19392 13472 19398 13484
rect 19889 13481 19901 13484
rect 19935 13481 19947 13515
rect 20714 13512 20720 13524
rect 20675 13484 20720 13512
rect 19889 13475 19947 13481
rect 20714 13472 20720 13484
rect 20772 13472 20778 13524
rect 20990 13472 20996 13524
rect 21048 13512 21054 13524
rect 21177 13515 21235 13521
rect 21177 13512 21189 13515
rect 21048 13484 21189 13512
rect 21048 13472 21054 13484
rect 21177 13481 21189 13484
rect 21223 13481 21235 13515
rect 21177 13475 21235 13481
rect 22094 13472 22100 13524
rect 22152 13512 22158 13524
rect 22833 13515 22891 13521
rect 22833 13512 22845 13515
rect 22152 13484 22845 13512
rect 22152 13472 22158 13484
rect 22833 13481 22845 13484
rect 22879 13481 22891 13515
rect 22833 13475 22891 13481
rect 23201 13515 23259 13521
rect 23201 13481 23213 13515
rect 23247 13512 23259 13515
rect 23385 13515 23443 13521
rect 23385 13512 23397 13515
rect 23247 13484 23397 13512
rect 23247 13481 23259 13484
rect 23201 13475 23259 13481
rect 23385 13481 23397 13484
rect 23431 13512 23443 13515
rect 23569 13515 23627 13521
rect 23569 13512 23581 13515
rect 23431 13484 23581 13512
rect 23431 13481 23443 13484
rect 23385 13475 23443 13481
rect 23569 13481 23581 13484
rect 23615 13512 23627 13515
rect 23842 13512 23848 13524
rect 23615 13484 23848 13512
rect 23615 13481 23627 13484
rect 23569 13475 23627 13481
rect 23842 13472 23848 13484
rect 23900 13512 23906 13524
rect 24673 13515 24731 13521
rect 24673 13512 24685 13515
rect 23900 13484 24685 13512
rect 23900 13472 23906 13484
rect 24673 13481 24685 13484
rect 24719 13481 24731 13515
rect 25038 13512 25044 13524
rect 24999 13484 25044 13512
rect 24673 13475 24731 13481
rect 25038 13472 25044 13484
rect 25096 13472 25102 13524
rect 25406 13512 25412 13524
rect 25367 13484 25412 13512
rect 25406 13472 25412 13484
rect 25464 13512 25470 13524
rect 25961 13515 26019 13521
rect 25961 13512 25973 13515
rect 25464 13484 25973 13512
rect 25464 13472 25470 13484
rect 25961 13481 25973 13484
rect 26007 13481 26019 13515
rect 26694 13512 26700 13524
rect 26655 13484 26700 13512
rect 25961 13475 26019 13481
rect 26694 13472 26700 13484
rect 26752 13472 26758 13524
rect 26786 13472 26792 13524
rect 26844 13512 26850 13524
rect 27617 13515 27675 13521
rect 27617 13512 27629 13515
rect 26844 13484 27629 13512
rect 26844 13472 26850 13484
rect 27617 13481 27629 13484
rect 27663 13512 27675 13515
rect 27706 13512 27712 13524
rect 27663 13484 27712 13512
rect 27663 13481 27675 13484
rect 27617 13475 27675 13481
rect 27706 13472 27712 13484
rect 27764 13472 27770 13524
rect 29270 13512 29276 13524
rect 29231 13484 29276 13512
rect 29270 13472 29276 13484
rect 29328 13472 29334 13524
rect 30837 13515 30895 13521
rect 30837 13481 30849 13515
rect 30883 13512 30895 13515
rect 31018 13512 31024 13524
rect 30883 13484 31024 13512
rect 30883 13481 30895 13484
rect 30837 13475 30895 13481
rect 31018 13472 31024 13484
rect 31076 13472 31082 13524
rect 31570 13512 31576 13524
rect 31531 13484 31576 13512
rect 31570 13472 31576 13484
rect 31628 13472 31634 13524
rect 31938 13472 31944 13524
rect 31996 13512 32002 13524
rect 32217 13515 32275 13521
rect 32217 13512 32229 13515
rect 31996 13484 32229 13512
rect 31996 13472 32002 13484
rect 32217 13481 32229 13484
rect 32263 13481 32275 13515
rect 33134 13512 33140 13524
rect 33095 13484 33140 13512
rect 32217 13475 32275 13481
rect 33134 13472 33140 13484
rect 33192 13472 33198 13524
rect 33594 13512 33600 13524
rect 33555 13484 33600 13512
rect 33594 13472 33600 13484
rect 33652 13472 33658 13524
rect 33870 13512 33876 13524
rect 33831 13484 33876 13512
rect 33870 13472 33876 13484
rect 33928 13472 33934 13524
rect 17954 13404 17960 13456
rect 18012 13444 18018 13456
rect 18233 13447 18291 13453
rect 18233 13444 18245 13447
rect 18012 13416 18245 13444
rect 18012 13404 18018 13416
rect 18233 13413 18245 13416
rect 18279 13413 18291 13447
rect 18598 13444 18604 13456
rect 18559 13416 18604 13444
rect 18233 13407 18291 13413
rect 17405 13379 17463 13385
rect 17405 13345 17417 13379
rect 17451 13376 17463 13379
rect 18046 13376 18052 13388
rect 17451 13348 18052 13376
rect 17451 13345 17463 13348
rect 17405 13339 17463 13345
rect 18046 13336 18052 13348
rect 18104 13336 18110 13388
rect 18248 13376 18276 13407
rect 18598 13404 18604 13416
rect 18656 13404 18662 13456
rect 28258 13404 28264 13456
rect 28316 13444 28322 13456
rect 28905 13447 28963 13453
rect 28316 13416 28488 13444
rect 28316 13404 28322 13416
rect 18782 13376 18788 13388
rect 18248 13348 18788 13376
rect 18782 13336 18788 13348
rect 18840 13336 18846 13388
rect 18966 13336 18972 13388
rect 19024 13376 19030 13388
rect 19429 13379 19487 13385
rect 19429 13376 19441 13379
rect 19024 13348 19441 13376
rect 19024 13336 19030 13348
rect 19429 13345 19441 13348
rect 19475 13345 19487 13379
rect 19429 13339 19487 13345
rect 19886 13336 19892 13388
rect 19944 13376 19950 13388
rect 20257 13379 20315 13385
rect 20257 13376 20269 13379
rect 19944 13348 20269 13376
rect 19944 13336 19950 13348
rect 20257 13345 20269 13348
rect 20303 13345 20315 13379
rect 21450 13376 21456 13388
rect 21411 13348 21456 13376
rect 20257 13339 20315 13345
rect 21450 13336 21456 13348
rect 21508 13336 21514 13388
rect 22373 13379 22431 13385
rect 22373 13345 22385 13379
rect 22419 13376 22431 13379
rect 22554 13376 22560 13388
rect 22419 13348 22560 13376
rect 22419 13345 22431 13348
rect 22373 13339 22431 13345
rect 22554 13336 22560 13348
rect 22612 13336 22618 13388
rect 22649 13379 22707 13385
rect 22649 13345 22661 13379
rect 22695 13345 22707 13379
rect 22649 13339 22707 13345
rect 23385 13379 23443 13385
rect 23385 13345 23397 13379
rect 23431 13376 23443 13379
rect 23661 13379 23719 13385
rect 23661 13376 23673 13379
rect 23431 13348 23673 13376
rect 23431 13345 23443 13348
rect 23385 13339 23443 13345
rect 23661 13345 23673 13348
rect 23707 13345 23719 13379
rect 23661 13339 23719 13345
rect 23808 13379 23866 13385
rect 23808 13345 23820 13379
rect 23854 13376 23866 13379
rect 24118 13376 24124 13388
rect 23854 13348 24124 13376
rect 23854 13345 23866 13348
rect 23808 13339 23866 13345
rect 11164 13308 11192 13336
rect 11606 13308 11612 13320
rect 8956 13280 11192 13308
rect 11567 13280 11612 13308
rect 11606 13268 11612 13280
rect 11664 13308 11670 13320
rect 11885 13311 11943 13317
rect 11885 13308 11897 13311
rect 11664 13280 11897 13308
rect 11664 13268 11670 13280
rect 11885 13277 11897 13280
rect 11931 13277 11943 13311
rect 11885 13271 11943 13277
rect 16666 13268 16672 13320
rect 16724 13308 16730 13320
rect 17037 13311 17095 13317
rect 17037 13308 17049 13311
rect 16724 13280 17049 13308
rect 16724 13268 16730 13280
rect 17037 13277 17049 13280
rect 17083 13277 17095 13311
rect 17037 13271 17095 13277
rect 17770 13268 17776 13320
rect 17828 13308 17834 13320
rect 17865 13311 17923 13317
rect 17865 13308 17877 13311
rect 17828 13280 17877 13308
rect 17828 13268 17834 13280
rect 17865 13277 17877 13280
rect 17911 13277 17923 13311
rect 17865 13271 17923 13277
rect 4062 13200 4068 13252
rect 4120 13240 4126 13252
rect 4341 13243 4399 13249
rect 4341 13240 4353 13243
rect 4120 13212 4353 13240
rect 4120 13200 4126 13212
rect 4341 13209 4353 13212
rect 4387 13240 4399 13243
rect 5074 13240 5080 13252
rect 4387 13212 5080 13240
rect 4387 13209 4399 13212
rect 4341 13203 4399 13209
rect 5074 13200 5080 13212
rect 5132 13200 5138 13252
rect 8662 13200 8668 13252
rect 8720 13240 8726 13252
rect 9125 13243 9183 13249
rect 9125 13240 9137 13243
rect 8720 13212 9137 13240
rect 8720 13200 8726 13212
rect 9125 13209 9137 13212
rect 9171 13240 9183 13243
rect 13262 13240 13268 13252
rect 9171 13212 10272 13240
rect 13223 13212 13268 13240
rect 9171 13209 9183 13212
rect 9125 13203 9183 13209
rect 10244 13184 10272 13212
rect 13262 13200 13268 13212
rect 13320 13200 13326 13252
rect 14734 13200 14740 13252
rect 14792 13240 14798 13252
rect 15470 13240 15476 13252
rect 14792 13212 15476 13240
rect 14792 13200 14798 13212
rect 15470 13200 15476 13212
rect 15528 13200 15534 13252
rect 19426 13200 19432 13252
rect 19484 13240 19490 13252
rect 19613 13243 19671 13249
rect 19613 13240 19625 13243
rect 19484 13212 19625 13240
rect 19484 13200 19490 13212
rect 19613 13209 19625 13212
rect 19659 13209 19671 13243
rect 22664 13240 22692 13339
rect 24118 13336 24124 13348
rect 24176 13336 24182 13388
rect 25222 13376 25228 13388
rect 25183 13348 25228 13376
rect 25222 13336 25228 13348
rect 25280 13336 25286 13388
rect 26050 13336 26056 13388
rect 26108 13376 26114 13388
rect 26513 13379 26571 13385
rect 26513 13376 26525 13379
rect 26108 13348 26525 13376
rect 26108 13336 26114 13348
rect 26513 13345 26525 13348
rect 26559 13376 26571 13379
rect 26973 13379 27031 13385
rect 26973 13376 26985 13379
rect 26559 13348 26985 13376
rect 26559 13345 26571 13348
rect 26513 13339 26571 13345
rect 26973 13345 26985 13348
rect 27019 13345 27031 13379
rect 26973 13339 27031 13345
rect 27798 13336 27804 13388
rect 27856 13376 27862 13388
rect 28350 13376 28356 13388
rect 27856 13348 28356 13376
rect 27856 13336 27862 13348
rect 28350 13336 28356 13348
rect 28408 13336 28414 13388
rect 28460 13385 28488 13416
rect 28905 13413 28917 13447
rect 28951 13444 28963 13447
rect 29546 13444 29552 13456
rect 28951 13416 29552 13444
rect 28951 13413 28963 13416
rect 28905 13407 28963 13413
rect 29546 13404 29552 13416
rect 29604 13444 29610 13456
rect 30098 13444 30104 13456
rect 29604 13416 30104 13444
rect 29604 13404 29610 13416
rect 30098 13404 30104 13416
rect 30156 13404 30162 13456
rect 28445 13379 28503 13385
rect 28445 13345 28457 13379
rect 28491 13345 28503 13379
rect 28445 13339 28503 13345
rect 29733 13379 29791 13385
rect 29733 13345 29745 13379
rect 29779 13376 29791 13379
rect 29822 13376 29828 13388
rect 29779 13348 29828 13376
rect 29779 13345 29791 13348
rect 29733 13339 29791 13345
rect 29822 13336 29828 13348
rect 29880 13336 29886 13388
rect 30009 13379 30067 13385
rect 30009 13345 30021 13379
rect 30055 13376 30067 13379
rect 30190 13376 30196 13388
rect 30055 13348 30196 13376
rect 30055 13345 30067 13348
rect 30009 13339 30067 13345
rect 30190 13336 30196 13348
rect 30248 13336 30254 13388
rect 31754 13336 31760 13388
rect 31812 13376 31818 13388
rect 32401 13379 32459 13385
rect 32401 13376 32413 13379
rect 31812 13348 32413 13376
rect 31812 13336 31818 13348
rect 32401 13345 32413 13348
rect 32447 13376 32459 13379
rect 32490 13376 32496 13388
rect 32447 13348 32496 13376
rect 32447 13345 32459 13348
rect 32401 13339 32459 13345
rect 32490 13336 32496 13348
rect 32548 13336 32554 13388
rect 32585 13379 32643 13385
rect 32585 13345 32597 13379
rect 32631 13345 32643 13379
rect 32585 13339 32643 13345
rect 24029 13311 24087 13317
rect 24029 13277 24041 13311
rect 24075 13308 24087 13311
rect 24210 13308 24216 13320
rect 24075 13280 24216 13308
rect 24075 13277 24087 13280
rect 24029 13271 24087 13277
rect 24210 13268 24216 13280
rect 24268 13268 24274 13320
rect 27246 13268 27252 13320
rect 27304 13308 27310 13320
rect 28169 13311 28227 13317
rect 28169 13308 28181 13311
rect 27304 13280 28181 13308
rect 27304 13268 27310 13280
rect 28169 13277 28181 13280
rect 28215 13277 28227 13311
rect 28169 13271 28227 13277
rect 30469 13311 30527 13317
rect 30469 13277 30481 13311
rect 30515 13308 30527 13311
rect 31110 13308 31116 13320
rect 30515 13280 31116 13308
rect 30515 13277 30527 13280
rect 30469 13271 30527 13277
rect 31110 13268 31116 13280
rect 31168 13268 31174 13320
rect 32600 13308 32628 13339
rect 32858 13308 32864 13320
rect 31864 13280 32864 13308
rect 22922 13240 22928 13252
rect 22664 13212 22928 13240
rect 19613 13203 19671 13209
rect 22922 13200 22928 13212
rect 22980 13240 22986 13252
rect 24121 13243 24179 13249
rect 24121 13240 24133 13243
rect 22980 13212 24133 13240
rect 22980 13200 22986 13212
rect 24121 13209 24133 13212
rect 24167 13209 24179 13243
rect 24121 13203 24179 13209
rect 27614 13200 27620 13252
rect 27672 13240 27678 13252
rect 27985 13243 28043 13249
rect 27985 13240 27997 13243
rect 27672 13212 27997 13240
rect 27672 13200 27678 13212
rect 27985 13209 27997 13212
rect 28031 13209 28043 13243
rect 27985 13203 28043 13209
rect 29825 13243 29883 13249
rect 29825 13209 29837 13243
rect 29871 13240 29883 13243
rect 30006 13240 30012 13252
rect 29871 13212 30012 13240
rect 29871 13209 29883 13212
rect 29825 13203 29883 13209
rect 30006 13200 30012 13212
rect 30064 13240 30070 13252
rect 30558 13240 30564 13252
rect 30064 13212 30564 13240
rect 30064 13200 30070 13212
rect 30558 13200 30564 13212
rect 30616 13200 30622 13252
rect 31864 13184 31892 13280
rect 32858 13268 32864 13280
rect 32916 13268 32922 13320
rect 4890 13172 4896 13184
rect 4851 13144 4896 13172
rect 4890 13132 4896 13144
rect 4948 13132 4954 13184
rect 9858 13172 9864 13184
rect 9819 13144 9864 13172
rect 9858 13132 9864 13144
rect 9916 13132 9922 13184
rect 10226 13172 10232 13184
rect 10139 13144 10232 13172
rect 10226 13132 10232 13144
rect 10284 13172 10290 13184
rect 11330 13172 11336 13184
rect 10284 13144 11336 13172
rect 10284 13132 10290 13144
rect 11330 13132 11336 13144
rect 11388 13132 11394 13184
rect 12250 13172 12256 13184
rect 12211 13144 12256 13172
rect 12250 13132 12256 13144
rect 12308 13132 12314 13184
rect 15102 13172 15108 13184
rect 15063 13144 15108 13172
rect 15102 13132 15108 13144
rect 15160 13132 15166 13184
rect 17494 13132 17500 13184
rect 17552 13172 17558 13184
rect 17681 13175 17739 13181
rect 17681 13172 17693 13175
rect 17552 13144 17693 13172
rect 17552 13132 17558 13144
rect 17681 13141 17693 13144
rect 17727 13141 17739 13175
rect 17681 13135 17739 13141
rect 21910 13132 21916 13184
rect 21968 13172 21974 13184
rect 22005 13175 22063 13181
rect 22005 13172 22017 13175
rect 21968 13144 22017 13172
rect 21968 13132 21974 13144
rect 22005 13141 22017 13144
rect 22051 13172 22063 13175
rect 23385 13175 23443 13181
rect 23385 13172 23397 13175
rect 22051 13144 23397 13172
rect 22051 13141 22063 13144
rect 22005 13135 22063 13141
rect 23385 13141 23397 13144
rect 23431 13141 23443 13175
rect 23385 13135 23443 13141
rect 23750 13132 23756 13184
rect 23808 13172 23814 13184
rect 23937 13175 23995 13181
rect 23937 13172 23949 13175
rect 23808 13144 23949 13172
rect 23808 13132 23814 13144
rect 23937 13141 23949 13144
rect 23983 13141 23995 13175
rect 23937 13135 23995 13141
rect 28810 13132 28816 13184
rect 28868 13172 28874 13184
rect 29270 13172 29276 13184
rect 28868 13144 29276 13172
rect 28868 13132 28874 13144
rect 29270 13132 29276 13144
rect 29328 13132 29334 13184
rect 31846 13172 31852 13184
rect 31807 13144 31852 13172
rect 31846 13132 31852 13144
rect 31904 13132 31910 13184
rect 1104 13082 38548 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 38548 13082
rect 1104 13008 38548 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 5077 12971 5135 12977
rect 5077 12937 5089 12971
rect 5123 12968 5135 12971
rect 6178 12968 6184 12980
rect 5123 12940 6184 12968
rect 5123 12937 5135 12940
rect 5077 12931 5135 12937
rect 6178 12928 6184 12940
rect 6236 12928 6242 12980
rect 8113 12971 8171 12977
rect 8113 12937 8125 12971
rect 8159 12968 8171 12971
rect 8662 12968 8668 12980
rect 8159 12940 8668 12968
rect 8159 12937 8171 12940
rect 8113 12931 8171 12937
rect 5445 12903 5503 12909
rect 5445 12869 5457 12903
rect 5491 12900 5503 12903
rect 5718 12900 5724 12912
rect 5491 12872 5724 12900
rect 5491 12869 5503 12872
rect 5445 12863 5503 12869
rect 5718 12860 5724 12872
rect 5776 12860 5782 12912
rect 5813 12903 5871 12909
rect 5813 12869 5825 12903
rect 5859 12900 5871 12903
rect 6454 12900 6460 12912
rect 5859 12872 6460 12900
rect 5859 12869 5871 12872
rect 5813 12863 5871 12869
rect 6454 12860 6460 12872
rect 6512 12860 6518 12912
rect 1394 12792 1400 12844
rect 1452 12832 1458 12844
rect 1949 12835 2007 12841
rect 1949 12832 1961 12835
rect 1452 12804 1961 12832
rect 1452 12792 1458 12804
rect 1949 12801 1961 12804
rect 1995 12801 2007 12835
rect 1949 12795 2007 12801
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12832 6699 12835
rect 6914 12832 6920 12844
rect 6687 12804 6920 12832
rect 6687 12801 6699 12804
rect 6641 12795 6699 12801
rect 1964 12628 1992 12795
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 8128 12832 8156 12931
rect 8662 12928 8668 12940
rect 8720 12928 8726 12980
rect 10686 12968 10692 12980
rect 10647 12940 10692 12968
rect 10686 12928 10692 12940
rect 10744 12928 10750 12980
rect 10946 12971 11004 12977
rect 10946 12937 10958 12971
rect 10992 12968 11004 12971
rect 11606 12968 11612 12980
rect 10992 12940 11612 12968
rect 10992 12937 11004 12940
rect 10946 12931 11004 12937
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 11790 12968 11796 12980
rect 11751 12940 11796 12968
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 12158 12928 12164 12980
rect 12216 12968 12222 12980
rect 12253 12971 12311 12977
rect 12253 12968 12265 12971
rect 12216 12940 12265 12968
rect 12216 12928 12222 12940
rect 12253 12937 12265 12940
rect 12299 12968 12311 12971
rect 12299 12940 12572 12968
rect 12299 12937 12311 12940
rect 12253 12931 12311 12937
rect 9582 12860 9588 12912
rect 9640 12900 9646 12912
rect 9861 12903 9919 12909
rect 9861 12900 9873 12903
rect 9640 12872 9873 12900
rect 9640 12860 9646 12872
rect 9861 12869 9873 12872
rect 9907 12869 9919 12903
rect 10318 12900 10324 12912
rect 10279 12872 10324 12900
rect 9861 12863 9919 12869
rect 10318 12860 10324 12872
rect 10376 12860 10382 12912
rect 11054 12900 11060 12912
rect 11015 12872 11060 12900
rect 11054 12860 11060 12872
rect 11112 12860 11118 12912
rect 11238 12900 11244 12912
rect 11199 12872 11244 12900
rect 11238 12860 11244 12872
rect 11296 12860 11302 12912
rect 7116 12804 8156 12832
rect 7116 12773 7144 12804
rect 8846 12792 8852 12844
rect 8904 12832 8910 12844
rect 11146 12832 11152 12844
rect 8904 12804 10364 12832
rect 11107 12804 11152 12832
rect 8904 12792 8910 12804
rect 10336 12776 10364 12804
rect 11146 12792 11152 12804
rect 11204 12792 11210 12844
rect 11808 12832 11836 12928
rect 12544 12832 12572 12940
rect 12710 12928 12716 12980
rect 12768 12968 12774 12980
rect 12897 12971 12955 12977
rect 12897 12968 12909 12971
rect 12768 12940 12909 12968
rect 12768 12928 12774 12940
rect 12897 12937 12909 12940
rect 12943 12968 12955 12971
rect 13630 12968 13636 12980
rect 12943 12940 13636 12968
rect 12943 12937 12955 12940
rect 12897 12931 12955 12937
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 15102 12928 15108 12980
rect 15160 12968 15166 12980
rect 16209 12971 16267 12977
rect 16209 12968 16221 12971
rect 15160 12940 16221 12968
rect 15160 12928 15166 12940
rect 16209 12937 16221 12940
rect 16255 12968 16267 12971
rect 16298 12968 16304 12980
rect 16255 12940 16304 12968
rect 16255 12937 16267 12940
rect 16209 12931 16267 12937
rect 16298 12928 16304 12940
rect 16356 12928 16362 12980
rect 16574 12928 16580 12980
rect 16632 12968 16638 12980
rect 17313 12971 17371 12977
rect 17313 12968 17325 12971
rect 16632 12940 17325 12968
rect 16632 12928 16638 12940
rect 17313 12937 17325 12940
rect 17359 12937 17371 12971
rect 18966 12968 18972 12980
rect 18927 12940 18972 12968
rect 17313 12931 17371 12937
rect 18966 12928 18972 12940
rect 19024 12968 19030 12980
rect 19705 12971 19763 12977
rect 19705 12968 19717 12971
rect 19024 12940 19717 12968
rect 19024 12928 19030 12940
rect 19705 12937 19717 12940
rect 19751 12968 19763 12971
rect 20073 12971 20131 12977
rect 20073 12968 20085 12971
rect 19751 12940 20085 12968
rect 19751 12937 19763 12940
rect 19705 12931 19763 12937
rect 20073 12937 20085 12940
rect 20119 12937 20131 12971
rect 20073 12931 20131 12937
rect 20990 12928 20996 12980
rect 21048 12968 21054 12980
rect 21085 12971 21143 12977
rect 21085 12968 21097 12971
rect 21048 12940 21097 12968
rect 21048 12928 21054 12940
rect 21085 12937 21097 12940
rect 21131 12937 21143 12971
rect 21085 12931 21143 12937
rect 23109 12971 23167 12977
rect 23109 12937 23121 12971
rect 23155 12968 23167 12971
rect 24118 12968 24124 12980
rect 23155 12940 24124 12968
rect 23155 12937 23167 12940
rect 23109 12931 23167 12937
rect 24118 12928 24124 12940
rect 24176 12928 24182 12980
rect 25222 12968 25228 12980
rect 25183 12940 25228 12968
rect 25222 12928 25228 12940
rect 25280 12928 25286 12980
rect 26218 12971 26276 12977
rect 26218 12937 26230 12971
rect 26264 12968 26276 12971
rect 26694 12968 26700 12980
rect 26264 12940 26700 12968
rect 26264 12937 26276 12940
rect 26218 12931 26276 12937
rect 26694 12928 26700 12940
rect 26752 12968 26758 12980
rect 26970 12968 26976 12980
rect 26752 12940 26976 12968
rect 26752 12928 26758 12940
rect 26970 12928 26976 12940
rect 27028 12928 27034 12980
rect 27525 12971 27583 12977
rect 27525 12937 27537 12971
rect 27571 12968 27583 12971
rect 27890 12968 27896 12980
rect 27571 12940 27896 12968
rect 27571 12937 27583 12940
rect 27525 12931 27583 12937
rect 27890 12928 27896 12940
rect 27948 12928 27954 12980
rect 28626 12928 28632 12980
rect 28684 12968 28690 12980
rect 28997 12971 29055 12977
rect 28997 12968 29009 12971
rect 28684 12940 29009 12968
rect 28684 12928 28690 12940
rect 28997 12937 29009 12940
rect 29043 12937 29055 12971
rect 30190 12968 30196 12980
rect 30151 12940 30196 12968
rect 28997 12931 29055 12937
rect 30190 12928 30196 12940
rect 30248 12928 30254 12980
rect 30558 12968 30564 12980
rect 30519 12940 30564 12968
rect 30558 12928 30564 12940
rect 30616 12928 30622 12980
rect 32490 12968 32496 12980
rect 32451 12940 32496 12968
rect 32490 12928 32496 12940
rect 32548 12928 32554 12980
rect 32858 12968 32864 12980
rect 32819 12940 32864 12968
rect 32858 12928 32864 12940
rect 32916 12928 32922 12980
rect 13541 12903 13599 12909
rect 13541 12869 13553 12903
rect 13587 12900 13599 12903
rect 13587 12872 14044 12900
rect 13587 12869 13599 12872
rect 13541 12863 13599 12869
rect 12894 12832 12900 12844
rect 11808 12804 12480 12832
rect 12544 12804 12900 12832
rect 6273 12767 6331 12773
rect 6273 12733 6285 12767
rect 6319 12764 6331 12767
rect 7101 12767 7159 12773
rect 7101 12764 7113 12767
rect 6319 12736 7113 12764
rect 6319 12733 6331 12736
rect 6273 12727 6331 12733
rect 7101 12733 7113 12736
rect 7147 12733 7159 12767
rect 7101 12727 7159 12733
rect 7653 12767 7711 12773
rect 7653 12733 7665 12767
rect 7699 12764 7711 12767
rect 8481 12767 8539 12773
rect 8481 12764 8493 12767
rect 7699 12736 8493 12764
rect 7699 12733 7711 12736
rect 7653 12727 7711 12733
rect 8481 12733 8493 12736
rect 8527 12764 8539 12767
rect 8662 12764 8668 12776
rect 8527 12736 8668 12764
rect 8527 12733 8539 12736
rect 8481 12727 8539 12733
rect 8662 12724 8668 12736
rect 8720 12724 8726 12776
rect 8754 12724 8760 12776
rect 8812 12764 8818 12776
rect 8941 12767 8999 12773
rect 8941 12764 8953 12767
rect 8812 12736 8953 12764
rect 8812 12724 8818 12736
rect 8941 12733 8953 12736
rect 8987 12733 8999 12767
rect 8941 12727 8999 12733
rect 9493 12767 9551 12773
rect 9493 12733 9505 12767
rect 9539 12764 9551 12767
rect 9582 12764 9588 12776
rect 9539 12736 9588 12764
rect 9539 12733 9551 12736
rect 9493 12727 9551 12733
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 9766 12764 9772 12776
rect 9727 12736 9772 12764
rect 9766 12724 9772 12736
rect 9824 12724 9830 12776
rect 10318 12724 10324 12776
rect 10376 12724 10382 12776
rect 10781 12767 10839 12773
rect 10781 12733 10793 12767
rect 10827 12764 10839 12767
rect 12250 12764 12256 12776
rect 10827 12736 12256 12764
rect 10827 12733 10839 12736
rect 10781 12727 10839 12733
rect 12250 12724 12256 12736
rect 12308 12724 12314 12776
rect 12452 12773 12480 12804
rect 12894 12792 12900 12804
rect 12952 12792 12958 12844
rect 13906 12832 13912 12844
rect 13867 12804 13912 12832
rect 13906 12792 13912 12804
rect 13964 12792 13970 12844
rect 14016 12832 14044 12872
rect 15930 12860 15936 12912
rect 15988 12900 15994 12912
rect 16071 12903 16129 12909
rect 16071 12900 16083 12903
rect 15988 12872 16083 12900
rect 15988 12860 15994 12872
rect 16071 12869 16083 12872
rect 16117 12869 16129 12903
rect 22462 12900 22468 12912
rect 22423 12872 22468 12900
rect 16071 12863 16129 12869
rect 22462 12860 22468 12872
rect 22520 12860 22526 12912
rect 24026 12909 24032 12912
rect 24010 12903 24032 12909
rect 24010 12869 24022 12903
rect 24084 12900 24090 12912
rect 24670 12900 24676 12912
rect 24084 12872 24676 12900
rect 24010 12863 24032 12869
rect 24026 12860 24032 12863
rect 24084 12860 24090 12872
rect 24670 12860 24676 12872
rect 24728 12900 24734 12912
rect 24857 12903 24915 12909
rect 24857 12900 24869 12903
rect 24728 12872 24869 12900
rect 24728 12860 24734 12872
rect 24857 12869 24869 12872
rect 24903 12869 24915 12903
rect 26326 12900 26332 12912
rect 26287 12872 26332 12900
rect 24857 12863 24915 12869
rect 26326 12860 26332 12872
rect 26384 12860 26390 12912
rect 15102 12832 15108 12844
rect 14016 12804 15108 12832
rect 12437 12767 12495 12773
rect 12437 12733 12449 12767
rect 12483 12733 12495 12767
rect 12437 12727 12495 12733
rect 13446 12724 13452 12776
rect 13504 12764 13510 12776
rect 14016 12773 14044 12804
rect 15102 12792 15108 12804
rect 15160 12792 15166 12844
rect 15378 12792 15384 12844
rect 15436 12832 15442 12844
rect 16301 12835 16359 12841
rect 16301 12832 16313 12835
rect 15436 12804 16313 12832
rect 15436 12792 15442 12804
rect 16301 12801 16313 12804
rect 16347 12832 16359 12835
rect 17770 12832 17776 12844
rect 16347 12804 17776 12832
rect 16347 12801 16359 12804
rect 16301 12795 16359 12801
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 19061 12835 19119 12841
rect 19061 12801 19073 12835
rect 19107 12832 19119 12835
rect 19150 12832 19156 12844
rect 19107 12804 19156 12832
rect 19107 12801 19119 12804
rect 19061 12795 19119 12801
rect 19150 12792 19156 12804
rect 19208 12792 19214 12844
rect 19334 12792 19340 12844
rect 19392 12832 19398 12844
rect 24210 12832 24216 12844
rect 19392 12804 19437 12832
rect 24123 12804 24216 12832
rect 19392 12792 19398 12804
rect 24210 12792 24216 12804
rect 24268 12792 24274 12844
rect 25498 12792 25504 12844
rect 25556 12832 25562 12844
rect 25866 12832 25872 12844
rect 25556 12804 25872 12832
rect 25556 12792 25562 12804
rect 25866 12792 25872 12804
rect 25924 12832 25930 12844
rect 25961 12835 26019 12841
rect 25961 12832 25973 12835
rect 25924 12804 25973 12832
rect 25924 12792 25930 12804
rect 25961 12801 25973 12804
rect 26007 12832 26019 12835
rect 26421 12835 26479 12841
rect 26421 12832 26433 12835
rect 26007 12804 26433 12832
rect 26007 12801 26019 12804
rect 25961 12795 26019 12801
rect 26421 12801 26433 12804
rect 26467 12832 26479 12835
rect 27614 12832 27620 12844
rect 26467 12804 27620 12832
rect 26467 12801 26479 12804
rect 26421 12795 26479 12801
rect 27614 12792 27620 12804
rect 27672 12792 27678 12844
rect 27908 12832 27936 12928
rect 31389 12903 31447 12909
rect 31389 12869 31401 12903
rect 31435 12900 31447 12903
rect 32766 12900 32772 12912
rect 31435 12872 32772 12900
rect 31435 12869 31447 12872
rect 31389 12863 31447 12869
rect 32766 12860 32772 12872
rect 32824 12860 32830 12912
rect 27908 12804 28028 12832
rect 13633 12767 13691 12773
rect 13633 12764 13645 12767
rect 13504 12736 13645 12764
rect 13504 12724 13510 12736
rect 13633 12733 13645 12736
rect 13679 12733 13691 12767
rect 13633 12727 13691 12733
rect 14001 12767 14059 12773
rect 14001 12733 14013 12767
rect 14047 12733 14059 12767
rect 14001 12727 14059 12733
rect 7285 12699 7343 12705
rect 7285 12665 7297 12699
rect 7331 12696 7343 12699
rect 7466 12696 7472 12708
rect 7331 12668 7472 12696
rect 7331 12665 7343 12668
rect 7285 12659 7343 12665
rect 7466 12656 7472 12668
rect 7524 12656 7530 12708
rect 9306 12656 9312 12708
rect 9364 12696 9370 12708
rect 9858 12696 9864 12708
rect 9364 12668 9864 12696
rect 9364 12656 9370 12668
rect 9858 12656 9864 12668
rect 9916 12656 9922 12708
rect 10962 12656 10968 12708
rect 11020 12696 11026 12708
rect 12526 12696 12532 12708
rect 11020 12668 12532 12696
rect 11020 12656 11026 12668
rect 12526 12656 12532 12668
rect 12584 12656 12590 12708
rect 12894 12656 12900 12708
rect 12952 12696 12958 12708
rect 13078 12696 13084 12708
rect 12952 12668 13084 12696
rect 12952 12656 12958 12668
rect 13078 12656 13084 12668
rect 13136 12656 13142 12708
rect 5534 12628 5540 12640
rect 1964 12600 5540 12628
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 7006 12588 7012 12640
rect 7064 12628 7070 12640
rect 7193 12631 7251 12637
rect 7193 12628 7205 12631
rect 7064 12600 7205 12628
rect 7064 12588 7070 12600
rect 7193 12597 7205 12600
rect 7239 12597 7251 12631
rect 7193 12591 7251 12597
rect 11606 12588 11612 12640
rect 11664 12628 11670 12640
rect 11974 12628 11980 12640
rect 11664 12600 11980 12628
rect 11664 12588 11670 12600
rect 11974 12588 11980 12600
rect 12032 12628 12038 12640
rect 12621 12631 12679 12637
rect 12621 12628 12633 12631
rect 12032 12600 12633 12628
rect 12032 12588 12038 12600
rect 12621 12597 12633 12600
rect 12667 12597 12679 12631
rect 13648 12628 13676 12727
rect 14090 12724 14096 12776
rect 14148 12764 14154 12776
rect 14550 12764 14556 12776
rect 14148 12736 14556 12764
rect 14148 12724 14154 12736
rect 14550 12724 14556 12736
rect 14608 12724 14614 12776
rect 14734 12724 14740 12776
rect 14792 12764 14798 12776
rect 14921 12767 14979 12773
rect 14921 12764 14933 12767
rect 14792 12736 14933 12764
rect 14792 12724 14798 12736
rect 14921 12733 14933 12736
rect 14967 12733 14979 12767
rect 15838 12764 15844 12776
rect 15751 12736 15844 12764
rect 14921 12727 14979 12733
rect 15838 12724 15844 12736
rect 15896 12764 15902 12776
rect 15933 12767 15991 12773
rect 15933 12764 15945 12767
rect 15896 12736 15945 12764
rect 15896 12724 15902 12736
rect 15933 12733 15945 12736
rect 15979 12733 15991 12767
rect 15933 12727 15991 12733
rect 17037 12767 17095 12773
rect 17037 12733 17049 12767
rect 17083 12764 17095 12767
rect 17310 12764 17316 12776
rect 17083 12736 17316 12764
rect 17083 12733 17095 12736
rect 17037 12727 17095 12733
rect 17310 12724 17316 12736
rect 17368 12724 17374 12776
rect 18598 12724 18604 12776
rect 18656 12764 18662 12776
rect 18693 12767 18751 12773
rect 18693 12764 18705 12767
rect 18656 12736 18705 12764
rect 18656 12724 18662 12736
rect 18693 12733 18705 12736
rect 18739 12733 18751 12767
rect 18693 12727 18751 12733
rect 18840 12767 18898 12773
rect 18840 12733 18852 12767
rect 18886 12764 18898 12767
rect 19426 12764 19432 12776
rect 18886 12736 19432 12764
rect 18886 12733 18898 12736
rect 18840 12727 18898 12733
rect 15010 12656 15016 12708
rect 15068 12696 15074 12708
rect 18708 12696 18736 12727
rect 19426 12724 19432 12736
rect 19484 12724 19490 12776
rect 20441 12767 20499 12773
rect 20441 12733 20453 12767
rect 20487 12764 20499 12767
rect 20990 12764 20996 12776
rect 20487 12736 20996 12764
rect 20487 12733 20499 12736
rect 20441 12727 20499 12733
rect 20990 12724 20996 12736
rect 21048 12724 21054 12776
rect 21545 12767 21603 12773
rect 21545 12733 21557 12767
rect 21591 12764 21603 12767
rect 21818 12764 21824 12776
rect 21591 12736 21824 12764
rect 21591 12733 21603 12736
rect 21545 12727 21603 12733
rect 21818 12724 21824 12736
rect 21876 12724 21882 12776
rect 22094 12724 22100 12776
rect 22152 12764 22158 12776
rect 22554 12764 22560 12776
rect 22152 12736 22197 12764
rect 22515 12736 22560 12764
rect 22152 12724 22158 12736
rect 22554 12724 22560 12736
rect 22612 12724 22618 12776
rect 23842 12764 23848 12776
rect 23803 12736 23848 12764
rect 23842 12724 23848 12736
rect 23900 12724 23906 12776
rect 19978 12696 19984 12708
rect 15068 12668 15516 12696
rect 18708 12668 19984 12696
rect 15068 12656 15074 12668
rect 15488 12640 15516 12668
rect 19978 12656 19984 12668
rect 20036 12696 20042 12708
rect 20162 12696 20168 12708
rect 20036 12668 20168 12696
rect 20036 12656 20042 12668
rect 20162 12656 20168 12668
rect 20220 12696 20226 12708
rect 20257 12699 20315 12705
rect 20257 12696 20269 12699
rect 20220 12668 20269 12696
rect 20220 12656 20226 12668
rect 20257 12665 20269 12668
rect 20303 12665 20315 12699
rect 20806 12696 20812 12708
rect 20767 12668 20812 12696
rect 20257 12659 20315 12665
rect 20806 12656 20812 12668
rect 20864 12656 20870 12708
rect 23566 12656 23572 12708
rect 23624 12696 23630 12708
rect 23934 12696 23940 12708
rect 23624 12668 23940 12696
rect 23624 12656 23630 12668
rect 23934 12656 23940 12668
rect 23992 12656 23998 12708
rect 24228 12696 24256 12792
rect 26050 12764 26056 12776
rect 26011 12736 26056 12764
rect 26050 12724 26056 12736
rect 26108 12764 26114 12776
rect 26326 12764 26332 12776
rect 26108 12736 26332 12764
rect 26108 12724 26114 12736
rect 26326 12724 26332 12736
rect 26384 12724 26390 12776
rect 27706 12724 27712 12776
rect 27764 12764 27770 12776
rect 27893 12767 27951 12773
rect 27893 12764 27905 12767
rect 27764 12736 27905 12764
rect 27764 12724 27770 12736
rect 27893 12733 27905 12736
rect 27939 12733 27951 12767
rect 27893 12727 27951 12733
rect 26602 12696 26608 12708
rect 24228 12668 26608 12696
rect 14366 12628 14372 12640
rect 13648 12600 14372 12628
rect 12621 12591 12679 12597
rect 14366 12588 14372 12600
rect 14424 12588 14430 12640
rect 15378 12628 15384 12640
rect 15339 12600 15384 12628
rect 15378 12588 15384 12600
rect 15436 12588 15442 12640
rect 15470 12588 15476 12640
rect 15528 12588 15534 12640
rect 16022 12588 16028 12640
rect 16080 12628 16086 12640
rect 16577 12631 16635 12637
rect 16577 12628 16589 12631
rect 16080 12600 16589 12628
rect 16080 12588 16086 12600
rect 16577 12597 16589 12600
rect 16623 12597 16635 12631
rect 16577 12591 16635 12597
rect 17954 12588 17960 12640
rect 18012 12628 18018 12640
rect 18601 12631 18659 12637
rect 18601 12628 18613 12631
rect 18012 12600 18613 12628
rect 18012 12588 18018 12600
rect 18601 12597 18613 12600
rect 18647 12628 18659 12631
rect 19150 12628 19156 12640
rect 18647 12600 19156 12628
rect 18647 12597 18659 12600
rect 18601 12591 18659 12597
rect 19150 12588 19156 12600
rect 19208 12588 19214 12640
rect 23290 12588 23296 12640
rect 23348 12628 23354 12640
rect 23385 12631 23443 12637
rect 23385 12628 23397 12631
rect 23348 12600 23397 12628
rect 23348 12588 23354 12600
rect 23385 12597 23397 12600
rect 23431 12628 23443 12631
rect 24228 12628 24256 12668
rect 26602 12656 26608 12668
rect 26660 12656 26666 12708
rect 26786 12696 26792 12708
rect 26747 12668 26792 12696
rect 26786 12656 26792 12668
rect 26844 12656 26850 12708
rect 27157 12699 27215 12705
rect 27157 12665 27169 12699
rect 27203 12696 27215 12699
rect 27338 12696 27344 12708
rect 27203 12668 27344 12696
rect 27203 12665 27215 12668
rect 27157 12659 27215 12665
rect 27338 12656 27344 12668
rect 27396 12696 27402 12708
rect 27798 12696 27804 12708
rect 27396 12668 27568 12696
rect 27759 12668 27804 12696
rect 27396 12656 27402 12668
rect 24486 12628 24492 12640
rect 23431 12600 24256 12628
rect 24447 12600 24492 12628
rect 23431 12597 23443 12600
rect 23385 12591 23443 12597
rect 24486 12588 24492 12600
rect 24544 12588 24550 12640
rect 26234 12588 26240 12640
rect 26292 12628 26298 12640
rect 26510 12628 26516 12640
rect 26292 12600 26516 12628
rect 26292 12588 26298 12600
rect 26510 12588 26516 12600
rect 26568 12588 26574 12640
rect 27540 12628 27568 12668
rect 27798 12656 27804 12668
rect 27856 12656 27862 12708
rect 28000 12705 28028 12804
rect 28258 12792 28264 12844
rect 28316 12832 28322 12844
rect 28629 12835 28687 12841
rect 28629 12832 28641 12835
rect 28316 12804 28641 12832
rect 28316 12792 28322 12804
rect 28629 12801 28641 12804
rect 28675 12801 28687 12835
rect 28629 12795 28687 12801
rect 29917 12835 29975 12841
rect 29917 12801 29929 12835
rect 29963 12832 29975 12835
rect 30374 12832 30380 12844
rect 29963 12804 30380 12832
rect 29963 12801 29975 12804
rect 29917 12795 29975 12801
rect 30374 12792 30380 12804
rect 30432 12792 30438 12844
rect 31021 12835 31079 12841
rect 31021 12801 31033 12835
rect 31067 12832 31079 12835
rect 35713 12835 35771 12841
rect 31067 12804 31708 12832
rect 31067 12801 31079 12804
rect 31021 12795 31079 12801
rect 31680 12776 31708 12804
rect 35713 12801 35725 12835
rect 35759 12832 35771 12835
rect 37274 12832 37280 12844
rect 35759 12804 36124 12832
rect 37235 12804 37280 12832
rect 35759 12801 35771 12804
rect 35713 12795 35771 12801
rect 29546 12764 29552 12776
rect 29507 12736 29552 12764
rect 29546 12724 29552 12736
rect 29604 12724 29610 12776
rect 30650 12724 30656 12776
rect 30708 12764 30714 12776
rect 31110 12764 31116 12776
rect 30708 12736 31116 12764
rect 30708 12724 30714 12736
rect 31110 12724 31116 12736
rect 31168 12724 31174 12776
rect 31662 12764 31668 12776
rect 31623 12736 31668 12764
rect 31662 12724 31668 12736
rect 31720 12724 31726 12776
rect 31938 12764 31944 12776
rect 31899 12736 31944 12764
rect 31938 12724 31944 12736
rect 31996 12724 32002 12776
rect 35802 12764 35808 12776
rect 35763 12736 35808 12764
rect 35802 12724 35808 12736
rect 35860 12724 35866 12776
rect 36096 12773 36124 12804
rect 37274 12792 37280 12804
rect 37332 12792 37338 12844
rect 36081 12767 36139 12773
rect 36081 12733 36093 12767
rect 36127 12764 36139 12767
rect 37182 12764 37188 12776
rect 36127 12736 37188 12764
rect 36127 12733 36139 12736
rect 36081 12727 36139 12733
rect 37182 12724 37188 12736
rect 37240 12724 37246 12776
rect 27985 12699 28043 12705
rect 27985 12665 27997 12699
rect 28031 12665 28043 12699
rect 27985 12659 28043 12665
rect 28353 12699 28411 12705
rect 28353 12665 28365 12699
rect 28399 12696 28411 12699
rect 29365 12699 29423 12705
rect 29365 12696 29377 12699
rect 28399 12668 29377 12696
rect 28399 12665 28411 12668
rect 28353 12659 28411 12665
rect 29365 12665 29377 12668
rect 29411 12696 29423 12699
rect 30558 12696 30564 12708
rect 29411 12668 30564 12696
rect 29411 12665 29423 12668
rect 29365 12659 29423 12665
rect 30558 12656 30564 12668
rect 30616 12656 30622 12708
rect 27816 12628 27844 12656
rect 27540 12600 27844 12628
rect 28258 12588 28264 12640
rect 28316 12628 28322 12640
rect 28442 12628 28448 12640
rect 28316 12600 28448 12628
rect 28316 12588 28322 12600
rect 28442 12588 28448 12600
rect 28500 12588 28506 12640
rect 1104 12538 38548 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 38548 12538
rect 1104 12464 38548 12486
rect 5258 12424 5264 12436
rect 5219 12396 5264 12424
rect 5258 12384 5264 12396
rect 5316 12384 5322 12436
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 5721 12427 5779 12433
rect 5721 12424 5733 12427
rect 5592 12396 5733 12424
rect 5592 12384 5598 12396
rect 5721 12393 5733 12396
rect 5767 12393 5779 12427
rect 5721 12387 5779 12393
rect 6822 12384 6828 12436
rect 6880 12424 6886 12436
rect 7745 12427 7803 12433
rect 6880 12396 7328 12424
rect 6880 12384 6886 12396
rect 5810 12316 5816 12368
rect 5868 12356 5874 12368
rect 6365 12359 6423 12365
rect 6365 12356 6377 12359
rect 5868 12328 6377 12356
rect 5868 12316 5874 12328
rect 6365 12325 6377 12328
rect 6411 12325 6423 12359
rect 6365 12319 6423 12325
rect 6546 12316 6552 12368
rect 6604 12356 6610 12368
rect 6604 12328 7236 12356
rect 6604 12316 6610 12328
rect 1578 12248 1584 12300
rect 1636 12288 1642 12300
rect 1765 12291 1823 12297
rect 1765 12288 1777 12291
rect 1636 12260 1777 12288
rect 1636 12248 1642 12260
rect 1765 12257 1777 12260
rect 1811 12257 1823 12291
rect 3142 12288 3148 12300
rect 3103 12260 3148 12288
rect 1765 12251 1823 12257
rect 3142 12248 3148 12260
rect 3200 12248 3206 12300
rect 4157 12291 4215 12297
rect 4157 12257 4169 12291
rect 4203 12288 4215 12291
rect 4614 12288 4620 12300
rect 4203 12260 4620 12288
rect 4203 12257 4215 12260
rect 4157 12251 4215 12257
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 5905 12291 5963 12297
rect 5905 12257 5917 12291
rect 5951 12257 5963 12291
rect 5905 12251 5963 12257
rect 6181 12291 6239 12297
rect 6181 12257 6193 12291
rect 6227 12288 6239 12291
rect 6822 12288 6828 12300
rect 6227 12260 6828 12288
rect 6227 12257 6239 12260
rect 6181 12251 6239 12257
rect 1489 12223 1547 12229
rect 1489 12189 1501 12223
rect 1535 12220 1547 12223
rect 1946 12220 1952 12232
rect 1535 12192 1952 12220
rect 1535 12189 1547 12192
rect 1489 12183 1547 12189
rect 1946 12180 1952 12192
rect 2004 12180 2010 12232
rect 4341 12155 4399 12161
rect 4341 12121 4353 12155
rect 4387 12152 4399 12155
rect 4706 12152 4712 12164
rect 4387 12124 4712 12152
rect 4387 12121 4399 12124
rect 4341 12115 4399 12121
rect 4706 12112 4712 12124
rect 4764 12112 4770 12164
rect 5920 12152 5948 12251
rect 6822 12248 6828 12260
rect 6880 12248 6886 12300
rect 7208 12297 7236 12328
rect 7193 12291 7251 12297
rect 7193 12257 7205 12291
rect 7239 12257 7251 12291
rect 7300 12288 7328 12396
rect 7745 12393 7757 12427
rect 7791 12424 7803 12427
rect 7926 12424 7932 12436
rect 7791 12396 7932 12424
rect 7791 12393 7803 12396
rect 7745 12387 7803 12393
rect 7926 12384 7932 12396
rect 7984 12384 7990 12436
rect 8018 12384 8024 12436
rect 8076 12424 8082 12436
rect 8662 12424 8668 12436
rect 8076 12396 8121 12424
rect 8623 12396 8668 12424
rect 8076 12384 8082 12396
rect 8662 12384 8668 12396
rect 8720 12384 8726 12436
rect 8754 12384 8760 12436
rect 8812 12424 8818 12436
rect 9033 12427 9091 12433
rect 9033 12424 9045 12427
rect 8812 12396 9045 12424
rect 8812 12384 8818 12396
rect 9033 12393 9045 12396
rect 9079 12393 9091 12427
rect 9033 12387 9091 12393
rect 9861 12427 9919 12433
rect 9861 12393 9873 12427
rect 9907 12424 9919 12427
rect 9950 12424 9956 12436
rect 9907 12396 9956 12424
rect 9907 12393 9919 12396
rect 9861 12387 9919 12393
rect 9950 12384 9956 12396
rect 10008 12384 10014 12436
rect 11606 12424 11612 12436
rect 11567 12396 11612 12424
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 11790 12384 11796 12436
rect 11848 12424 11854 12436
rect 11885 12427 11943 12433
rect 11885 12424 11897 12427
rect 11848 12396 11897 12424
rect 11848 12384 11854 12396
rect 11885 12393 11897 12396
rect 11931 12393 11943 12427
rect 12618 12424 12624 12436
rect 12579 12396 12624 12424
rect 11885 12387 11943 12393
rect 12618 12384 12624 12396
rect 12676 12384 12682 12436
rect 14182 12384 14188 12436
rect 14240 12424 14246 12436
rect 14369 12427 14427 12433
rect 14369 12424 14381 12427
rect 14240 12396 14381 12424
rect 14240 12384 14246 12396
rect 14369 12393 14381 12396
rect 14415 12393 14427 12427
rect 14369 12387 14427 12393
rect 14829 12427 14887 12433
rect 14829 12393 14841 12427
rect 14875 12424 14887 12427
rect 15470 12424 15476 12436
rect 14875 12396 15476 12424
rect 14875 12393 14887 12396
rect 14829 12387 14887 12393
rect 14936 12368 14964 12396
rect 15470 12384 15476 12396
rect 15528 12384 15534 12436
rect 16574 12384 16580 12436
rect 16632 12424 16638 12436
rect 16850 12424 16856 12436
rect 16632 12396 16856 12424
rect 16632 12384 16638 12396
rect 16850 12384 16856 12396
rect 16908 12384 16914 12436
rect 17402 12384 17408 12436
rect 17460 12424 17466 12436
rect 17460 12396 17724 12424
rect 17460 12384 17466 12396
rect 10597 12359 10655 12365
rect 10597 12325 10609 12359
rect 10643 12356 10655 12359
rect 11146 12356 11152 12368
rect 10643 12328 11152 12356
rect 10643 12325 10655 12328
rect 10597 12319 10655 12325
rect 11146 12316 11152 12328
rect 11204 12356 11210 12368
rect 11241 12359 11299 12365
rect 11241 12356 11253 12359
rect 11204 12328 11253 12356
rect 11204 12316 11210 12328
rect 11241 12325 11253 12328
rect 11287 12325 11299 12359
rect 11241 12319 11299 12325
rect 12434 12316 12440 12368
rect 12492 12356 12498 12368
rect 13078 12356 13084 12368
rect 12492 12328 13084 12356
rect 12492 12316 12498 12328
rect 13078 12316 13084 12328
rect 13136 12356 13142 12368
rect 13265 12359 13323 12365
rect 13265 12356 13277 12359
rect 13136 12328 13277 12356
rect 13136 12316 13142 12328
rect 13265 12325 13277 12328
rect 13311 12325 13323 12359
rect 14090 12356 14096 12368
rect 14051 12328 14096 12356
rect 13265 12319 13323 12325
rect 14090 12316 14096 12328
rect 14148 12316 14154 12368
rect 14918 12316 14924 12368
rect 14976 12316 14982 12368
rect 8202 12288 8208 12300
rect 7300 12260 8208 12288
rect 7193 12251 7251 12257
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 9674 12248 9680 12300
rect 9732 12288 9738 12300
rect 10778 12288 10784 12300
rect 9732 12260 9777 12288
rect 10739 12260 10784 12288
rect 9732 12248 9738 12260
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 11882 12248 11888 12300
rect 11940 12288 11946 12300
rect 12069 12291 12127 12297
rect 12069 12288 12081 12291
rect 11940 12260 12081 12288
rect 11940 12248 11946 12260
rect 12069 12257 12081 12260
rect 12115 12288 12127 12291
rect 12158 12288 12164 12300
rect 12115 12260 12164 12288
rect 12115 12257 12127 12260
rect 12069 12251 12127 12257
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 14185 12291 14243 12297
rect 14185 12257 14197 12291
rect 14231 12288 14243 12291
rect 14550 12288 14556 12300
rect 14231 12260 14556 12288
rect 14231 12257 14243 12260
rect 14185 12251 14243 12257
rect 14550 12248 14556 12260
rect 14608 12248 14614 12300
rect 15289 12291 15347 12297
rect 15289 12257 15301 12291
rect 15335 12288 15347 12291
rect 15378 12288 15384 12300
rect 15335 12260 15384 12288
rect 15335 12257 15347 12260
rect 15289 12251 15347 12257
rect 15378 12248 15384 12260
rect 15436 12288 15442 12300
rect 16574 12288 16580 12300
rect 15436 12260 16068 12288
rect 16535 12260 16580 12288
rect 15436 12248 15442 12260
rect 6270 12180 6276 12232
rect 6328 12220 6334 12232
rect 7282 12220 7288 12232
rect 6328 12192 7288 12220
rect 6328 12180 6334 12192
rect 7282 12180 7288 12192
rect 7340 12180 7346 12232
rect 9950 12180 9956 12232
rect 10008 12220 10014 12232
rect 10689 12223 10747 12229
rect 10689 12220 10701 12223
rect 10008 12192 10701 12220
rect 10008 12180 10014 12192
rect 10689 12189 10701 12192
rect 10735 12220 10747 12223
rect 11974 12220 11980 12232
rect 10735 12192 11980 12220
rect 10735 12189 10747 12192
rect 10689 12183 10747 12189
rect 11974 12180 11980 12192
rect 12032 12180 12038 12232
rect 12894 12180 12900 12232
rect 12952 12220 12958 12232
rect 13354 12220 13360 12232
rect 12952 12192 13360 12220
rect 12952 12180 12958 12192
rect 13354 12180 13360 12192
rect 13412 12180 13418 12232
rect 14734 12220 14740 12232
rect 13648 12192 14740 12220
rect 6454 12152 6460 12164
rect 5920 12124 6460 12152
rect 6454 12112 6460 12124
rect 6512 12112 6518 12164
rect 8389 12155 8447 12161
rect 8389 12121 8401 12155
rect 8435 12152 8447 12155
rect 9490 12152 9496 12164
rect 8435 12124 9496 12152
rect 8435 12121 8447 12124
rect 8389 12115 8447 12121
rect 9490 12112 9496 12124
rect 9548 12112 9554 12164
rect 9766 12112 9772 12164
rect 9824 12152 9830 12164
rect 10229 12155 10287 12161
rect 10229 12152 10241 12155
rect 9824 12124 10241 12152
rect 9824 12112 9830 12124
rect 10229 12121 10241 12124
rect 10275 12152 10287 12155
rect 10962 12152 10968 12164
rect 10275 12124 10968 12152
rect 10275 12121 10287 12124
rect 10229 12115 10287 12121
rect 10962 12112 10968 12124
rect 11020 12112 11026 12164
rect 11330 12112 11336 12164
rect 11388 12152 11394 12164
rect 13648 12161 13676 12192
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 12253 12155 12311 12161
rect 12253 12152 12265 12155
rect 11388 12124 12265 12152
rect 11388 12112 11394 12124
rect 12253 12121 12265 12124
rect 12299 12121 12311 12155
rect 13633 12155 13691 12161
rect 13633 12152 13645 12155
rect 12253 12115 12311 12121
rect 12636 12124 13645 12152
rect 4614 12084 4620 12096
rect 4575 12056 4620 12084
rect 4614 12044 4620 12056
rect 4672 12044 4678 12096
rect 5074 12044 5080 12096
rect 5132 12084 5138 12096
rect 5629 12087 5687 12093
rect 5629 12084 5641 12087
rect 5132 12056 5641 12084
rect 5132 12044 5138 12056
rect 5629 12053 5641 12056
rect 5675 12084 5687 12087
rect 7466 12084 7472 12096
rect 5675 12056 7472 12084
rect 5675 12053 5687 12056
rect 5629 12047 5687 12053
rect 7466 12044 7472 12056
rect 7524 12044 7530 12096
rect 9401 12087 9459 12093
rect 9401 12053 9413 12087
rect 9447 12084 9459 12087
rect 9582 12084 9588 12096
rect 9447 12056 9588 12084
rect 9447 12053 9459 12056
rect 9401 12047 9459 12053
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 12636 12084 12664 12124
rect 13633 12121 13645 12124
rect 13679 12121 13691 12155
rect 13633 12115 13691 12121
rect 9732 12056 12664 12084
rect 12989 12087 13047 12093
rect 9732 12044 9738 12056
rect 12989 12053 13001 12087
rect 13035 12084 13047 12087
rect 13354 12084 13360 12096
rect 13035 12056 13360 12084
rect 13035 12053 13047 12056
rect 12989 12047 13047 12053
rect 13354 12044 13360 12056
rect 13412 12044 13418 12096
rect 14734 12044 14740 12096
rect 14792 12084 14798 12096
rect 16040 12093 16068 12260
rect 16574 12248 16580 12260
rect 16632 12288 16638 12300
rect 16942 12288 16948 12300
rect 16632 12260 16948 12288
rect 16632 12248 16638 12260
rect 16942 12248 16948 12260
rect 17000 12248 17006 12300
rect 17696 12297 17724 12396
rect 18046 12384 18052 12436
rect 18104 12424 18110 12436
rect 18141 12427 18199 12433
rect 18141 12424 18153 12427
rect 18104 12396 18153 12424
rect 18104 12384 18110 12396
rect 18141 12393 18153 12396
rect 18187 12393 18199 12427
rect 18141 12387 18199 12393
rect 18417 12427 18475 12433
rect 18417 12393 18429 12427
rect 18463 12424 18475 12427
rect 18506 12424 18512 12436
rect 18463 12396 18512 12424
rect 18463 12393 18475 12396
rect 18417 12387 18475 12393
rect 18506 12384 18512 12396
rect 18564 12384 18570 12436
rect 18690 12384 18696 12436
rect 18748 12384 18754 12436
rect 18782 12384 18788 12436
rect 18840 12424 18846 12436
rect 19521 12427 19579 12433
rect 19521 12424 19533 12427
rect 18840 12396 19533 12424
rect 18840 12384 18846 12396
rect 19521 12393 19533 12396
rect 19567 12393 19579 12427
rect 19521 12387 19579 12393
rect 20162 12384 20168 12436
rect 20220 12424 20226 12436
rect 20257 12427 20315 12433
rect 20257 12424 20269 12427
rect 20220 12396 20269 12424
rect 20220 12384 20226 12396
rect 20257 12393 20269 12396
rect 20303 12393 20315 12427
rect 20257 12387 20315 12393
rect 21085 12427 21143 12433
rect 21085 12393 21097 12427
rect 21131 12393 21143 12427
rect 21085 12387 21143 12393
rect 17313 12291 17371 12297
rect 17313 12257 17325 12291
rect 17359 12257 17371 12291
rect 17313 12251 17371 12257
rect 17681 12291 17739 12297
rect 17681 12257 17693 12291
rect 17727 12257 17739 12291
rect 17681 12251 17739 12257
rect 16482 12180 16488 12232
rect 16540 12180 16546 12232
rect 16666 12220 16672 12232
rect 16627 12192 16672 12220
rect 16666 12180 16672 12192
rect 16724 12180 16730 12232
rect 17126 12220 17132 12232
rect 17087 12192 17132 12220
rect 17126 12180 17132 12192
rect 17184 12180 17190 12232
rect 16500 12152 16528 12180
rect 16942 12152 16948 12164
rect 16500 12124 16948 12152
rect 16942 12112 16948 12124
rect 17000 12112 17006 12164
rect 17218 12112 17224 12164
rect 17276 12152 17282 12164
rect 17328 12152 17356 12251
rect 18046 12248 18052 12300
rect 18104 12288 18110 12300
rect 18708 12288 18736 12384
rect 21100 12356 21128 12387
rect 22094 12384 22100 12436
rect 22152 12424 22158 12436
rect 22922 12424 22928 12436
rect 22152 12396 22197 12424
rect 22883 12396 22928 12424
rect 22152 12384 22158 12396
rect 22922 12384 22928 12396
rect 22980 12384 22986 12436
rect 23198 12424 23204 12436
rect 23111 12396 23204 12424
rect 23198 12384 23204 12396
rect 23256 12424 23262 12436
rect 23569 12427 23627 12433
rect 23569 12424 23581 12427
rect 23256 12396 23581 12424
rect 23256 12384 23262 12396
rect 23569 12393 23581 12396
rect 23615 12393 23627 12427
rect 24670 12424 24676 12436
rect 24631 12396 24676 12424
rect 23569 12387 23627 12393
rect 24670 12384 24676 12396
rect 24728 12384 24734 12436
rect 24765 12427 24823 12433
rect 24765 12393 24777 12427
rect 24811 12424 24823 12427
rect 26326 12424 26332 12436
rect 24811 12396 26332 12424
rect 24811 12393 24823 12396
rect 24765 12387 24823 12393
rect 26326 12384 26332 12396
rect 26384 12384 26390 12436
rect 26694 12424 26700 12436
rect 26655 12396 26700 12424
rect 26694 12384 26700 12396
rect 26752 12384 26758 12436
rect 27430 12384 27436 12436
rect 27488 12424 27494 12436
rect 27709 12427 27767 12433
rect 27709 12424 27721 12427
rect 27488 12396 27721 12424
rect 27488 12384 27494 12396
rect 27709 12393 27721 12396
rect 27755 12393 27767 12427
rect 27709 12387 27767 12393
rect 28261 12427 28319 12433
rect 28261 12393 28273 12427
rect 28307 12424 28319 12427
rect 28350 12424 28356 12436
rect 28307 12396 28356 12424
rect 28307 12393 28319 12396
rect 28261 12387 28319 12393
rect 28350 12384 28356 12396
rect 28408 12384 28414 12436
rect 28810 12424 28816 12436
rect 28771 12396 28816 12424
rect 28810 12384 28816 12396
rect 28868 12384 28874 12436
rect 29457 12427 29515 12433
rect 29457 12393 29469 12427
rect 29503 12424 29515 12427
rect 29546 12424 29552 12436
rect 29503 12396 29552 12424
rect 29503 12393 29515 12396
rect 29457 12387 29515 12393
rect 29546 12384 29552 12396
rect 29604 12384 29610 12436
rect 30466 12424 30472 12436
rect 30427 12396 30472 12424
rect 30466 12384 30472 12396
rect 30524 12384 30530 12436
rect 30558 12384 30564 12436
rect 30616 12424 30622 12436
rect 30837 12427 30895 12433
rect 30837 12424 30849 12427
rect 30616 12396 30849 12424
rect 30616 12384 30622 12396
rect 30837 12393 30849 12396
rect 30883 12393 30895 12427
rect 30837 12387 30895 12393
rect 31205 12427 31263 12433
rect 31205 12393 31217 12427
rect 31251 12424 31263 12427
rect 32490 12424 32496 12436
rect 31251 12396 32496 12424
rect 31251 12393 31263 12396
rect 31205 12387 31263 12393
rect 32490 12384 32496 12396
rect 32548 12384 32554 12436
rect 35894 12384 35900 12436
rect 35952 12424 35958 12436
rect 36170 12424 36176 12436
rect 35952 12396 36176 12424
rect 35952 12384 35958 12396
rect 36170 12384 36176 12396
rect 36228 12384 36234 12436
rect 19260 12328 21128 12356
rect 21729 12359 21787 12365
rect 19260 12297 19288 12328
rect 21729 12325 21741 12359
rect 21775 12356 21787 12359
rect 22554 12356 22560 12368
rect 21775 12328 22560 12356
rect 21775 12325 21787 12328
rect 21729 12319 21787 12325
rect 22112 12300 22140 12328
rect 22554 12316 22560 12328
rect 22612 12316 22618 12368
rect 19245 12291 19303 12297
rect 19245 12288 19257 12291
rect 18104 12260 18736 12288
rect 18892 12260 19257 12288
rect 18104 12248 18110 12260
rect 18892 12232 18920 12260
rect 19245 12257 19257 12260
rect 19291 12257 19303 12291
rect 19518 12288 19524 12300
rect 19479 12260 19524 12288
rect 19245 12251 19303 12257
rect 19518 12248 19524 12260
rect 19576 12248 19582 12300
rect 20898 12288 20904 12300
rect 20859 12260 20904 12288
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 22094 12248 22100 12300
rect 22152 12248 22158 12300
rect 22370 12288 22376 12300
rect 22331 12260 22376 12288
rect 22370 12248 22376 12260
rect 22428 12248 22434 12300
rect 17586 12220 17592 12232
rect 17547 12192 17592 12220
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 18417 12223 18475 12229
rect 18417 12189 18429 12223
rect 18463 12220 18475 12223
rect 18601 12223 18659 12229
rect 18601 12220 18613 12223
rect 18463 12192 18613 12220
rect 18463 12189 18475 12192
rect 18417 12183 18475 12189
rect 18601 12189 18613 12192
rect 18647 12220 18659 12223
rect 18693 12223 18751 12229
rect 18693 12220 18705 12223
rect 18647 12192 18705 12220
rect 18647 12189 18659 12192
rect 18601 12183 18659 12189
rect 18693 12189 18705 12192
rect 18739 12189 18751 12223
rect 18693 12183 18751 12189
rect 18874 12180 18880 12232
rect 18932 12180 18938 12232
rect 22002 12180 22008 12232
rect 22060 12220 22066 12232
rect 23216 12220 23244 12384
rect 23750 12316 23756 12368
rect 23808 12356 23814 12368
rect 24305 12359 24363 12365
rect 24305 12356 24317 12359
rect 23808 12328 24317 12356
rect 23808 12316 23814 12328
rect 24305 12325 24317 12328
rect 24351 12356 24363 12359
rect 24351 12328 25360 12356
rect 24351 12325 24363 12328
rect 24305 12319 24363 12325
rect 23385 12291 23443 12297
rect 23385 12257 23397 12291
rect 23431 12288 23443 12291
rect 23474 12288 23480 12300
rect 23431 12260 23480 12288
rect 23431 12257 23443 12260
rect 23385 12251 23443 12257
rect 23474 12248 23480 12260
rect 23532 12288 23538 12300
rect 24486 12288 24492 12300
rect 23532 12260 24492 12288
rect 23532 12248 23538 12260
rect 24486 12248 24492 12260
rect 24544 12248 24550 12300
rect 24765 12291 24823 12297
rect 24765 12257 24777 12291
rect 24811 12288 24823 12291
rect 24854 12288 24860 12300
rect 24811 12260 24860 12288
rect 24811 12257 24823 12260
rect 24765 12251 24823 12257
rect 24854 12248 24860 12260
rect 24912 12248 24918 12300
rect 22060 12192 23244 12220
rect 22060 12180 22066 12192
rect 24946 12180 24952 12232
rect 25004 12220 25010 12232
rect 25225 12223 25283 12229
rect 25225 12220 25237 12223
rect 25004 12192 25237 12220
rect 25004 12180 25010 12192
rect 25225 12189 25237 12192
rect 25271 12189 25283 12223
rect 25332 12220 25360 12328
rect 25590 12288 25596 12300
rect 25551 12260 25596 12288
rect 25590 12248 25596 12260
rect 25648 12248 25654 12300
rect 26326 12248 26332 12300
rect 26384 12288 26390 12300
rect 26970 12288 26976 12300
rect 26384 12260 26976 12288
rect 26384 12248 26390 12260
rect 26970 12248 26976 12260
rect 27028 12288 27034 12300
rect 27065 12291 27123 12297
rect 27065 12288 27077 12291
rect 27028 12260 27077 12288
rect 27028 12248 27034 12260
rect 27065 12257 27077 12260
rect 27111 12257 27123 12291
rect 28626 12288 28632 12300
rect 27065 12251 27123 12257
rect 27448 12260 28632 12288
rect 25332 12192 25636 12220
rect 25225 12183 25283 12189
rect 18892 12152 18920 12180
rect 21450 12152 21456 12164
rect 17276 12124 18920 12152
rect 20640 12124 21456 12152
rect 17276 12112 17282 12124
rect 15473 12087 15531 12093
rect 15473 12084 15485 12087
rect 14792 12056 15485 12084
rect 14792 12044 14798 12056
rect 15473 12053 15485 12056
rect 15519 12053 15531 12087
rect 15473 12047 15531 12053
rect 16025 12087 16083 12093
rect 16025 12053 16037 12087
rect 16071 12084 16083 12087
rect 16114 12084 16120 12096
rect 16071 12056 16120 12084
rect 16071 12053 16083 12056
rect 16025 12047 16083 12053
rect 16114 12044 16120 12056
rect 16172 12044 16178 12096
rect 16393 12087 16451 12093
rect 16393 12053 16405 12087
rect 16439 12084 16451 12087
rect 16482 12084 16488 12096
rect 16439 12056 16488 12084
rect 16439 12053 16451 12056
rect 16393 12047 16451 12053
rect 16482 12044 16488 12056
rect 16540 12044 16546 12096
rect 18322 12044 18328 12096
rect 18380 12084 18386 12096
rect 19705 12087 19763 12093
rect 19705 12084 19717 12087
rect 18380 12056 19717 12084
rect 18380 12044 18386 12056
rect 19705 12053 19717 12056
rect 19751 12053 19763 12087
rect 19705 12047 19763 12053
rect 20530 12044 20536 12096
rect 20588 12084 20594 12096
rect 20640 12093 20668 12124
rect 21450 12112 21456 12124
rect 21508 12112 21514 12164
rect 23750 12112 23756 12164
rect 23808 12152 23814 12164
rect 24118 12152 24124 12164
rect 23808 12124 24124 12152
rect 23808 12112 23814 12124
rect 24118 12112 24124 12124
rect 24176 12112 24182 12164
rect 25130 12152 25136 12164
rect 25091 12124 25136 12152
rect 25130 12112 25136 12124
rect 25188 12112 25194 12164
rect 25608 12096 25636 12192
rect 26602 12180 26608 12232
rect 26660 12220 26666 12232
rect 27246 12220 27252 12232
rect 26660 12192 27252 12220
rect 26660 12180 26666 12192
rect 27246 12180 27252 12192
rect 27304 12220 27310 12232
rect 27448 12229 27476 12260
rect 28626 12248 28632 12260
rect 28684 12248 28690 12300
rect 29638 12288 29644 12300
rect 29599 12260 29644 12288
rect 29638 12248 29644 12260
rect 29696 12248 29702 12300
rect 30926 12248 30932 12300
rect 30984 12288 30990 12300
rect 31021 12291 31079 12297
rect 31021 12288 31033 12291
rect 30984 12260 31033 12288
rect 30984 12248 30990 12260
rect 31021 12257 31033 12260
rect 31067 12257 31079 12291
rect 31021 12251 31079 12257
rect 32490 12248 32496 12300
rect 32548 12288 32554 12300
rect 32769 12291 32827 12297
rect 32769 12288 32781 12291
rect 32548 12260 32781 12288
rect 32548 12248 32554 12260
rect 32769 12257 32781 12260
rect 32815 12288 32827 12291
rect 32858 12288 32864 12300
rect 32815 12260 32864 12288
rect 32815 12257 32827 12260
rect 32769 12251 32827 12257
rect 32858 12248 32864 12260
rect 32916 12248 32922 12300
rect 27433 12223 27491 12229
rect 27433 12220 27445 12223
rect 27304 12192 27445 12220
rect 27304 12180 27310 12192
rect 27433 12189 27445 12192
rect 27479 12189 27491 12223
rect 27433 12183 27491 12189
rect 27706 12152 27712 12164
rect 27218 12124 27712 12152
rect 20625 12087 20683 12093
rect 20625 12084 20637 12087
rect 20588 12056 20637 12084
rect 20588 12044 20594 12056
rect 20625 12053 20637 12056
rect 20671 12053 20683 12087
rect 20625 12047 20683 12053
rect 22557 12087 22615 12093
rect 22557 12053 22569 12087
rect 22603 12084 22615 12087
rect 23290 12084 23296 12096
rect 22603 12056 23296 12084
rect 22603 12053 22615 12056
rect 22557 12047 22615 12053
rect 23290 12044 23296 12056
rect 23348 12084 23354 12096
rect 25038 12093 25044 12096
rect 23845 12087 23903 12093
rect 23845 12084 23857 12087
rect 23348 12056 23857 12084
rect 23348 12044 23354 12056
rect 23845 12053 23857 12056
rect 23891 12053 23903 12087
rect 23845 12047 23903 12053
rect 25022 12087 25044 12093
rect 25022 12053 25034 12087
rect 25022 12047 25044 12053
rect 25038 12044 25044 12047
rect 25096 12044 25102 12096
rect 25590 12044 25596 12096
rect 25648 12084 25654 12096
rect 26053 12087 26111 12093
rect 26053 12084 26065 12087
rect 25648 12056 26065 12084
rect 25648 12044 25654 12056
rect 26053 12053 26065 12056
rect 26099 12084 26111 12087
rect 26142 12084 26148 12096
rect 26099 12056 26148 12084
rect 26099 12053 26111 12056
rect 26053 12047 26111 12053
rect 26142 12044 26148 12056
rect 26200 12044 26206 12096
rect 27218 12093 27246 12124
rect 27706 12112 27712 12124
rect 27764 12112 27770 12164
rect 29825 12155 29883 12161
rect 29825 12121 29837 12155
rect 29871 12152 29883 12155
rect 30193 12155 30251 12161
rect 30193 12152 30205 12155
rect 29871 12124 30205 12152
rect 29871 12121 29883 12124
rect 29825 12115 29883 12121
rect 30193 12121 30205 12124
rect 30239 12152 30251 12155
rect 31018 12152 31024 12164
rect 30239 12124 31024 12152
rect 30239 12121 30251 12124
rect 30193 12115 30251 12121
rect 31018 12112 31024 12124
rect 31076 12112 31082 12164
rect 27203 12087 27261 12093
rect 27203 12053 27215 12087
rect 27249 12053 27261 12087
rect 27338 12084 27344 12096
rect 27299 12056 27344 12084
rect 27203 12047 27261 12053
rect 27338 12044 27344 12056
rect 27396 12044 27402 12096
rect 31478 12084 31484 12096
rect 31439 12056 31484 12084
rect 31478 12044 31484 12056
rect 31536 12084 31542 12096
rect 31938 12084 31944 12096
rect 31536 12056 31944 12084
rect 31536 12044 31542 12056
rect 31938 12044 31944 12056
rect 31996 12084 32002 12096
rect 32401 12087 32459 12093
rect 32401 12084 32413 12087
rect 31996 12056 32413 12084
rect 31996 12044 32002 12056
rect 32401 12053 32413 12056
rect 32447 12053 32459 12087
rect 35802 12084 35808 12096
rect 35763 12056 35808 12084
rect 32401 12047 32459 12053
rect 35802 12044 35808 12056
rect 35860 12044 35866 12096
rect 1104 11994 38548 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 38548 11994
rect 1104 11920 38548 11942
rect 5997 11883 6055 11889
rect 5997 11849 6009 11883
rect 6043 11880 6055 11883
rect 6270 11880 6276 11892
rect 6043 11852 6276 11880
rect 6043 11849 6055 11852
rect 5997 11843 6055 11849
rect 6270 11840 6276 11852
rect 6328 11840 6334 11892
rect 7282 11880 7288 11892
rect 7243 11852 7288 11880
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 8202 11880 8208 11892
rect 8163 11852 8208 11880
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 9585 11883 9643 11889
rect 9585 11849 9597 11883
rect 9631 11880 9643 11883
rect 9674 11880 9680 11892
rect 9631 11852 9680 11880
rect 9631 11849 9643 11852
rect 9585 11843 9643 11849
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 11882 11880 11888 11892
rect 11843 11852 11888 11880
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 14277 11883 14335 11889
rect 14277 11849 14289 11883
rect 14323 11880 14335 11883
rect 14550 11880 14556 11892
rect 14323 11852 14556 11880
rect 14323 11849 14335 11852
rect 14277 11843 14335 11849
rect 14550 11840 14556 11852
rect 14608 11840 14614 11892
rect 16761 11883 16819 11889
rect 16761 11849 16773 11883
rect 16807 11880 16819 11883
rect 17402 11880 17408 11892
rect 16807 11852 17408 11880
rect 16807 11849 16819 11852
rect 16761 11843 16819 11849
rect 17402 11840 17408 11852
rect 17460 11840 17466 11892
rect 17497 11883 17555 11889
rect 17497 11849 17509 11883
rect 17543 11880 17555 11883
rect 17862 11880 17868 11892
rect 17543 11852 17868 11880
rect 17543 11849 17555 11852
rect 17497 11843 17555 11849
rect 4706 11772 4712 11824
rect 4764 11812 4770 11824
rect 5629 11815 5687 11821
rect 5629 11812 5641 11815
rect 4764 11784 5641 11812
rect 4764 11772 4770 11784
rect 5629 11781 5641 11784
rect 5675 11812 5687 11815
rect 6546 11812 6552 11824
rect 5675 11784 6552 11812
rect 5675 11781 5687 11784
rect 5629 11775 5687 11781
rect 6546 11772 6552 11784
rect 6604 11772 6610 11824
rect 11517 11815 11575 11821
rect 11517 11781 11529 11815
rect 11563 11812 11575 11815
rect 11974 11812 11980 11824
rect 11563 11784 11980 11812
rect 11563 11781 11575 11784
rect 11517 11775 11575 11781
rect 11974 11772 11980 11784
rect 12032 11772 12038 11824
rect 14645 11815 14703 11821
rect 14645 11781 14657 11815
rect 14691 11812 14703 11815
rect 16114 11812 16120 11824
rect 14691 11784 16120 11812
rect 14691 11781 14703 11784
rect 14645 11775 14703 11781
rect 16114 11772 16120 11784
rect 16172 11812 16178 11824
rect 17129 11815 17187 11821
rect 17129 11812 17141 11815
rect 16172 11784 17141 11812
rect 16172 11772 16178 11784
rect 17129 11781 17141 11784
rect 17175 11781 17187 11815
rect 17129 11775 17187 11781
rect 3050 11704 3056 11756
rect 3108 11744 3114 11756
rect 3329 11747 3387 11753
rect 3329 11744 3341 11747
rect 3108 11716 3341 11744
rect 3108 11704 3114 11716
rect 3329 11713 3341 11716
rect 3375 11744 3387 11747
rect 3697 11747 3755 11753
rect 3697 11744 3709 11747
rect 3375 11716 3709 11744
rect 3375 11713 3387 11716
rect 3329 11707 3387 11713
rect 3697 11713 3709 11716
rect 3743 11744 3755 11747
rect 4614 11744 4620 11756
rect 3743 11716 4620 11744
rect 3743 11713 3755 11716
rect 3697 11707 3755 11713
rect 4614 11704 4620 11716
rect 4672 11704 4678 11756
rect 7926 11704 7932 11756
rect 7984 11744 7990 11756
rect 8665 11747 8723 11753
rect 8665 11744 8677 11747
rect 7984 11716 8677 11744
rect 7984 11704 7990 11716
rect 8665 11713 8677 11716
rect 8711 11713 8723 11747
rect 8665 11707 8723 11713
rect 9217 11747 9275 11753
rect 9217 11713 9229 11747
rect 9263 11744 9275 11747
rect 9766 11744 9772 11756
rect 9263 11716 9772 11744
rect 9263 11713 9275 11716
rect 9217 11707 9275 11713
rect 9766 11704 9772 11716
rect 9824 11704 9830 11756
rect 12158 11704 12164 11756
rect 12216 11744 12222 11756
rect 12253 11747 12311 11753
rect 12253 11744 12265 11747
rect 12216 11716 12265 11744
rect 12216 11704 12222 11716
rect 12253 11713 12265 11716
rect 12299 11744 12311 11747
rect 12299 11716 12572 11744
rect 12299 11713 12311 11716
rect 12253 11707 12311 11713
rect 1946 11636 1952 11688
rect 2004 11676 2010 11688
rect 3418 11676 3424 11688
rect 2004 11648 3424 11676
rect 2004 11636 2010 11648
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 6638 11676 6644 11688
rect 6599 11648 6644 11676
rect 6638 11636 6644 11648
rect 6696 11636 6702 11688
rect 7469 11679 7527 11685
rect 7469 11645 7481 11679
rect 7515 11676 7527 11679
rect 8294 11676 8300 11688
rect 7515 11648 8300 11676
rect 7515 11645 7527 11648
rect 7469 11639 7527 11645
rect 5074 11608 5080 11620
rect 5035 11580 5080 11608
rect 5074 11568 5080 11580
rect 5132 11568 5138 11620
rect 6365 11611 6423 11617
rect 6365 11577 6377 11611
rect 6411 11608 6423 11611
rect 7484 11608 7512 11639
rect 8294 11636 8300 11648
rect 8352 11636 8358 11688
rect 8757 11679 8815 11685
rect 8757 11645 8769 11679
rect 8803 11676 8815 11679
rect 8938 11676 8944 11688
rect 8803 11648 8944 11676
rect 8803 11645 8815 11648
rect 8757 11639 8815 11645
rect 6411 11580 7512 11608
rect 7929 11611 7987 11617
rect 6411 11577 6423 11580
rect 6365 11571 6423 11577
rect 7929 11577 7941 11611
rect 7975 11608 7987 11611
rect 8772 11608 8800 11639
rect 8938 11636 8944 11648
rect 8996 11676 9002 11688
rect 9953 11679 10011 11685
rect 8996 11648 9444 11676
rect 8996 11636 9002 11648
rect 9416 11620 9444 11648
rect 9953 11645 9965 11679
rect 9999 11676 10011 11679
rect 10689 11679 10747 11685
rect 10689 11676 10701 11679
rect 9999 11648 10701 11676
rect 9999 11645 10011 11648
rect 9953 11639 10011 11645
rect 10689 11645 10701 11648
rect 10735 11676 10747 11679
rect 11330 11676 11336 11688
rect 10735 11648 11336 11676
rect 10735 11645 10747 11648
rect 10689 11639 10747 11645
rect 11330 11636 11336 11648
rect 11388 11636 11394 11688
rect 12544 11685 12572 11716
rect 13814 11704 13820 11756
rect 13872 11744 13878 11756
rect 14734 11744 14740 11756
rect 13872 11716 14740 11744
rect 13872 11704 13878 11716
rect 14734 11704 14740 11716
rect 14792 11704 14798 11756
rect 16022 11704 16028 11756
rect 16080 11704 16086 11756
rect 12529 11679 12587 11685
rect 12529 11645 12541 11679
rect 12575 11645 12587 11679
rect 13078 11676 13084 11688
rect 13039 11648 13084 11676
rect 12529 11639 12587 11645
rect 13078 11636 13084 11648
rect 13136 11636 13142 11688
rect 13262 11676 13268 11688
rect 13223 11648 13268 11676
rect 13262 11636 13268 11648
rect 13320 11636 13326 11688
rect 13354 11636 13360 11688
rect 13412 11676 13418 11688
rect 13725 11679 13783 11685
rect 13725 11676 13737 11679
rect 13412 11648 13737 11676
rect 13412 11636 13418 11648
rect 13725 11645 13737 11648
rect 13771 11645 13783 11679
rect 14918 11676 14924 11688
rect 14879 11648 14924 11676
rect 13725 11639 13783 11645
rect 7975 11580 8800 11608
rect 7975 11577 7987 11580
rect 7929 11571 7987 11577
rect 9398 11568 9404 11620
rect 9456 11608 9462 11620
rect 10045 11611 10103 11617
rect 10045 11608 10057 11611
rect 9456 11580 10057 11608
rect 9456 11568 9462 11580
rect 10045 11577 10057 11580
rect 10091 11577 10103 11611
rect 13740 11608 13768 11639
rect 14918 11636 14924 11648
rect 14976 11636 14982 11688
rect 15378 11676 15384 11688
rect 15339 11648 15384 11676
rect 15378 11636 15384 11648
rect 15436 11636 15442 11688
rect 15473 11679 15531 11685
rect 15473 11645 15485 11679
rect 15519 11676 15531 11679
rect 16040 11676 16068 11704
rect 15519 11648 16068 11676
rect 15519 11645 15531 11648
rect 15473 11639 15531 11645
rect 16758 11636 16764 11688
rect 16816 11636 16822 11688
rect 16945 11679 17003 11685
rect 16945 11645 16957 11679
rect 16991 11676 17003 11679
rect 17512 11676 17540 11843
rect 17862 11840 17868 11852
rect 17920 11840 17926 11892
rect 18874 11840 18880 11892
rect 18932 11880 18938 11892
rect 19061 11883 19119 11889
rect 19061 11880 19073 11883
rect 18932 11852 19073 11880
rect 18932 11840 18938 11852
rect 19061 11849 19073 11852
rect 19107 11849 19119 11883
rect 19518 11880 19524 11892
rect 19479 11852 19524 11880
rect 19061 11843 19119 11849
rect 19518 11840 19524 11852
rect 19576 11840 19582 11892
rect 20898 11880 20904 11892
rect 20859 11852 20904 11880
rect 20898 11840 20904 11852
rect 20956 11840 20962 11892
rect 23474 11880 23480 11892
rect 23435 11852 23480 11880
rect 23474 11840 23480 11852
rect 23532 11840 23538 11892
rect 23842 11840 23848 11892
rect 23900 11880 23906 11892
rect 24029 11883 24087 11889
rect 24029 11880 24041 11883
rect 23900 11852 24041 11880
rect 23900 11840 23906 11852
rect 24029 11849 24041 11852
rect 24075 11849 24087 11883
rect 24029 11843 24087 11849
rect 24118 11840 24124 11892
rect 24176 11880 24182 11892
rect 24949 11883 25007 11889
rect 24949 11880 24961 11883
rect 24176 11852 24961 11880
rect 24176 11840 24182 11852
rect 24949 11849 24961 11852
rect 24995 11880 25007 11883
rect 25130 11880 25136 11892
rect 24995 11852 25136 11880
rect 24995 11849 25007 11852
rect 24949 11843 25007 11849
rect 25130 11840 25136 11852
rect 25188 11840 25194 11892
rect 27246 11880 27252 11892
rect 27207 11852 27252 11880
rect 27246 11840 27252 11852
rect 27304 11840 27310 11892
rect 27706 11880 27712 11892
rect 27667 11852 27712 11880
rect 27706 11840 27712 11852
rect 27764 11840 27770 11892
rect 27985 11883 28043 11889
rect 27985 11849 27997 11883
rect 28031 11880 28043 11883
rect 28258 11880 28264 11892
rect 28031 11852 28264 11880
rect 28031 11849 28043 11852
rect 27985 11843 28043 11849
rect 28258 11840 28264 11852
rect 28316 11840 28322 11892
rect 28626 11880 28632 11892
rect 28587 11852 28632 11880
rect 28626 11840 28632 11852
rect 28684 11840 28690 11892
rect 29638 11880 29644 11892
rect 29599 11852 29644 11880
rect 29638 11840 29644 11852
rect 29696 11840 29702 11892
rect 30742 11840 30748 11892
rect 30800 11880 30806 11892
rect 31941 11883 31999 11889
rect 31941 11880 31953 11883
rect 30800 11852 31953 11880
rect 30800 11840 30806 11852
rect 31941 11849 31953 11852
rect 31987 11849 31999 11883
rect 32858 11880 32864 11892
rect 32819 11852 32864 11880
rect 31941 11843 31999 11849
rect 32858 11840 32864 11852
rect 32916 11840 32922 11892
rect 37274 11840 37280 11892
rect 37332 11880 37338 11892
rect 37369 11883 37427 11889
rect 37369 11880 37381 11883
rect 37332 11852 37381 11880
rect 37332 11840 37338 11852
rect 37369 11849 37381 11852
rect 37415 11849 37427 11883
rect 37369 11843 37427 11849
rect 22370 11772 22376 11824
rect 22428 11812 22434 11824
rect 23109 11815 23167 11821
rect 23109 11812 23121 11815
rect 22428 11784 23121 11812
rect 22428 11772 22434 11784
rect 23109 11781 23121 11784
rect 23155 11812 23167 11815
rect 25222 11812 25228 11824
rect 23155 11784 25228 11812
rect 23155 11781 23167 11784
rect 23109 11775 23167 11781
rect 25222 11772 25228 11784
rect 25280 11772 25286 11824
rect 19150 11704 19156 11756
rect 19208 11744 19214 11756
rect 19889 11747 19947 11753
rect 19889 11744 19901 11747
rect 19208 11716 19901 11744
rect 19208 11704 19214 11716
rect 19889 11713 19901 11716
rect 19935 11713 19947 11747
rect 22554 11744 22560 11756
rect 22515 11716 22560 11744
rect 19889 11707 19947 11713
rect 22554 11704 22560 11716
rect 22612 11704 22618 11756
rect 26786 11704 26792 11756
rect 26844 11744 26850 11756
rect 26973 11747 27031 11753
rect 26973 11744 26985 11747
rect 26844 11716 26985 11744
rect 26844 11704 26850 11716
rect 26973 11713 26985 11716
rect 27019 11744 27031 11747
rect 27724 11744 27752 11840
rect 30926 11772 30932 11824
rect 30984 11812 30990 11824
rect 31113 11815 31171 11821
rect 31113 11812 31125 11815
rect 30984 11784 31125 11812
rect 30984 11772 30990 11784
rect 31113 11781 31125 11784
rect 31159 11781 31171 11815
rect 31113 11775 31171 11781
rect 31662 11744 31668 11756
rect 27019 11716 27752 11744
rect 31575 11716 31668 11744
rect 27019 11713 27031 11716
rect 26973 11707 27031 11713
rect 31662 11704 31668 11716
rect 31720 11744 31726 11756
rect 32493 11747 32551 11753
rect 32493 11744 32505 11747
rect 31720 11716 32505 11744
rect 31720 11704 31726 11716
rect 32493 11713 32505 11716
rect 32539 11713 32551 11747
rect 32493 11707 32551 11713
rect 35713 11747 35771 11753
rect 35713 11713 35725 11747
rect 35759 11744 35771 11747
rect 35759 11716 36124 11744
rect 35759 11713 35771 11716
rect 35713 11707 35771 11713
rect 36096 11688 36124 11716
rect 18141 11679 18199 11685
rect 18141 11676 18153 11679
rect 16991 11648 17540 11676
rect 17880 11648 18153 11676
rect 16991 11645 17003 11648
rect 16945 11639 17003 11645
rect 16025 11611 16083 11617
rect 16025 11608 16037 11611
rect 13740 11580 16037 11608
rect 10045 11571 10103 11577
rect 16025 11577 16037 11580
rect 16071 11577 16083 11611
rect 16776 11608 16804 11636
rect 17880 11608 17908 11648
rect 18141 11645 18153 11648
rect 18187 11676 18199 11679
rect 18322 11676 18328 11688
rect 18187 11648 18328 11676
rect 18187 11645 18199 11648
rect 18141 11639 18199 11645
rect 18322 11636 18328 11648
rect 18380 11636 18386 11688
rect 20533 11679 20591 11685
rect 20533 11645 20545 11679
rect 20579 11676 20591 11679
rect 20622 11676 20628 11688
rect 20579 11648 20628 11676
rect 20579 11645 20591 11648
rect 20533 11639 20591 11645
rect 20622 11636 20628 11648
rect 20680 11636 20686 11688
rect 21545 11679 21603 11685
rect 21545 11645 21557 11679
rect 21591 11676 21603 11679
rect 21818 11676 21824 11688
rect 21591 11648 21824 11676
rect 21591 11645 21603 11648
rect 21545 11639 21603 11645
rect 21818 11636 21824 11648
rect 21876 11636 21882 11688
rect 22002 11676 22008 11688
rect 21963 11648 22008 11676
rect 22002 11636 22008 11648
rect 22060 11636 22066 11688
rect 22094 11636 22100 11688
rect 22152 11676 22158 11688
rect 22465 11679 22523 11685
rect 22465 11676 22477 11679
rect 22152 11648 22477 11676
rect 22152 11636 22158 11648
rect 22465 11645 22477 11648
rect 22511 11645 22523 11679
rect 22465 11639 22523 11645
rect 24026 11636 24032 11688
rect 24084 11676 24090 11688
rect 24397 11679 24455 11685
rect 24397 11676 24409 11679
rect 24084 11648 24409 11676
rect 24084 11636 24090 11648
rect 24397 11645 24409 11648
rect 24443 11676 24455 11679
rect 24854 11676 24860 11688
rect 24443 11648 24860 11676
rect 24443 11645 24455 11648
rect 24397 11639 24455 11645
rect 24854 11636 24860 11648
rect 24912 11636 24918 11688
rect 25038 11636 25044 11688
rect 25096 11676 25102 11688
rect 25685 11679 25743 11685
rect 25685 11676 25697 11679
rect 25096 11648 25697 11676
rect 25096 11636 25102 11648
rect 25685 11645 25697 11648
rect 25731 11676 25743 11679
rect 26145 11679 26203 11685
rect 26145 11676 26157 11679
rect 25731 11648 26157 11676
rect 25731 11645 25743 11648
rect 25685 11639 25743 11645
rect 26145 11645 26157 11648
rect 26191 11676 26203 11679
rect 26694 11676 26700 11688
rect 26191 11648 26700 11676
rect 26191 11645 26203 11648
rect 26145 11639 26203 11645
rect 26694 11636 26700 11648
rect 26752 11636 26758 11688
rect 27798 11676 27804 11688
rect 27759 11648 27804 11676
rect 27798 11636 27804 11648
rect 27856 11676 27862 11688
rect 28261 11679 28319 11685
rect 28261 11676 28273 11679
rect 27856 11648 28273 11676
rect 27856 11636 27862 11648
rect 28261 11645 28273 11648
rect 28307 11645 28319 11679
rect 28261 11639 28319 11645
rect 30745 11679 30803 11685
rect 30745 11645 30757 11679
rect 30791 11676 30803 11679
rect 31018 11676 31024 11688
rect 30791 11648 31024 11676
rect 30791 11645 30803 11648
rect 30745 11639 30803 11645
rect 31018 11636 31024 11648
rect 31076 11636 31082 11688
rect 31757 11679 31815 11685
rect 31757 11676 31769 11679
rect 31496 11648 31769 11676
rect 18046 11608 18052 11620
rect 16776 11580 17908 11608
rect 18007 11580 18052 11608
rect 16025 11571 16083 11577
rect 18046 11568 18052 11580
rect 18104 11568 18110 11620
rect 31496 11617 31524 11648
rect 31757 11645 31769 11648
rect 31803 11645 31815 11679
rect 35802 11676 35808 11688
rect 35763 11648 35808 11676
rect 31757 11639 31815 11645
rect 35802 11636 35808 11648
rect 35860 11636 35866 11688
rect 36078 11676 36084 11688
rect 36039 11648 36084 11676
rect 36078 11636 36084 11648
rect 36136 11636 36142 11688
rect 31481 11611 31539 11617
rect 31481 11608 31493 11611
rect 30392 11580 31493 11608
rect 30392 11552 30420 11580
rect 31481 11577 31493 11580
rect 31527 11577 31539 11611
rect 31481 11571 31539 11577
rect 1486 11500 1492 11552
rect 1544 11540 1550 11552
rect 1581 11543 1639 11549
rect 1581 11540 1593 11543
rect 1544 11512 1593 11540
rect 1544 11500 1550 11512
rect 1581 11509 1593 11512
rect 1627 11509 1639 11543
rect 1946 11540 1952 11552
rect 1907 11512 1952 11540
rect 1581 11503 1639 11509
rect 1946 11500 1952 11512
rect 2004 11500 2010 11552
rect 6454 11540 6460 11552
rect 6415 11512 6460 11540
rect 6454 11500 6460 11512
rect 6512 11500 6518 11552
rect 10778 11500 10784 11552
rect 10836 11540 10842 11552
rect 11054 11540 11060 11552
rect 10836 11512 11060 11540
rect 10836 11500 10842 11512
rect 11054 11500 11060 11512
rect 11112 11540 11118 11552
rect 11149 11543 11207 11549
rect 11149 11540 11161 11543
rect 11112 11512 11161 11540
rect 11112 11500 11118 11512
rect 11149 11509 11161 11512
rect 11195 11540 11207 11543
rect 11514 11540 11520 11552
rect 11195 11512 11520 11540
rect 11195 11509 11207 11512
rect 11149 11503 11207 11509
rect 11514 11500 11520 11512
rect 11572 11500 11578 11552
rect 12526 11540 12532 11552
rect 12487 11512 12532 11540
rect 12526 11500 12532 11512
rect 12584 11500 12590 11552
rect 16758 11500 16764 11552
rect 16816 11540 16822 11552
rect 17126 11540 17132 11552
rect 16816 11512 17132 11540
rect 16816 11500 16822 11512
rect 17126 11500 17132 11512
rect 17184 11540 17190 11552
rect 17773 11543 17831 11549
rect 17773 11540 17785 11543
rect 17184 11512 17785 11540
rect 17184 11500 17190 11512
rect 17773 11509 17785 11512
rect 17819 11509 17831 11543
rect 17773 11503 17831 11509
rect 24946 11500 24952 11552
rect 25004 11540 25010 11552
rect 25225 11543 25283 11549
rect 25225 11540 25237 11543
rect 25004 11512 25237 11540
rect 25004 11500 25010 11512
rect 25225 11509 25237 11512
rect 25271 11509 25283 11543
rect 30374 11540 30380 11552
rect 30335 11512 30380 11540
rect 25225 11503 25283 11509
rect 30374 11500 30380 11512
rect 30432 11500 30438 11552
rect 1104 11450 38548 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 38548 11450
rect 1104 11376 38548 11398
rect 5997 11339 6055 11345
rect 5997 11305 6009 11339
rect 6043 11336 6055 11339
rect 6638 11336 6644 11348
rect 6043 11308 6644 11336
rect 6043 11305 6055 11308
rect 5997 11299 6055 11305
rect 6638 11296 6644 11308
rect 6696 11296 6702 11348
rect 7653 11339 7711 11345
rect 7653 11305 7665 11339
rect 7699 11336 7711 11339
rect 8202 11336 8208 11348
rect 7699 11308 8208 11336
rect 7699 11305 7711 11308
rect 7653 11299 7711 11305
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 9398 11336 9404 11348
rect 9359 11308 9404 11336
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 9953 11339 10011 11345
rect 9953 11305 9965 11339
rect 9999 11336 10011 11339
rect 10042 11336 10048 11348
rect 9999 11308 10048 11336
rect 9999 11305 10011 11308
rect 9953 11299 10011 11305
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 10226 11296 10232 11348
rect 10284 11336 10290 11348
rect 10594 11336 10600 11348
rect 10284 11308 10600 11336
rect 10284 11296 10290 11308
rect 10594 11296 10600 11308
rect 10652 11296 10658 11348
rect 12989 11339 13047 11345
rect 12989 11305 13001 11339
rect 13035 11336 13047 11339
rect 13262 11336 13268 11348
rect 13035 11308 13268 11336
rect 13035 11305 13047 11308
rect 12989 11299 13047 11305
rect 13262 11296 13268 11308
rect 13320 11296 13326 11348
rect 14734 11336 14740 11348
rect 14695 11308 14740 11336
rect 14734 11296 14740 11308
rect 14792 11296 14798 11348
rect 15194 11296 15200 11348
rect 15252 11336 15258 11348
rect 16485 11339 16543 11345
rect 16485 11336 16497 11339
rect 15252 11308 16497 11336
rect 15252 11296 15258 11308
rect 16485 11305 16497 11308
rect 16531 11305 16543 11339
rect 16485 11299 16543 11305
rect 17037 11339 17095 11345
rect 17037 11305 17049 11339
rect 17083 11336 17095 11339
rect 17218 11336 17224 11348
rect 17083 11308 17224 11336
rect 17083 11305 17095 11308
rect 17037 11299 17095 11305
rect 17218 11296 17224 11308
rect 17276 11296 17282 11348
rect 18322 11296 18328 11348
rect 18380 11336 18386 11348
rect 18509 11339 18567 11345
rect 18509 11336 18521 11339
rect 18380 11308 18521 11336
rect 18380 11296 18386 11308
rect 18509 11305 18521 11308
rect 18555 11305 18567 11339
rect 18509 11299 18567 11305
rect 18598 11296 18604 11348
rect 18656 11336 18662 11348
rect 18877 11339 18935 11345
rect 18877 11336 18889 11339
rect 18656 11308 18889 11336
rect 18656 11296 18662 11308
rect 18877 11305 18889 11308
rect 18923 11305 18935 11339
rect 18877 11299 18935 11305
rect 19150 11296 19156 11348
rect 19208 11336 19214 11348
rect 19245 11339 19303 11345
rect 19245 11336 19257 11339
rect 19208 11308 19257 11336
rect 19208 11296 19214 11308
rect 19245 11305 19257 11308
rect 19291 11305 19303 11339
rect 19245 11299 19303 11305
rect 19981 11339 20039 11345
rect 19981 11305 19993 11339
rect 20027 11336 20039 11339
rect 20349 11339 20407 11345
rect 20349 11336 20361 11339
rect 20027 11308 20361 11336
rect 20027 11305 20039 11308
rect 19981 11299 20039 11305
rect 20349 11305 20361 11308
rect 20395 11336 20407 11339
rect 20622 11336 20628 11348
rect 20395 11308 20628 11336
rect 20395 11305 20407 11308
rect 20349 11299 20407 11305
rect 20622 11296 20628 11308
rect 20680 11296 20686 11348
rect 21729 11339 21787 11345
rect 21729 11305 21741 11339
rect 21775 11336 21787 11339
rect 22002 11336 22008 11348
rect 21775 11308 22008 11336
rect 21775 11305 21787 11308
rect 21729 11299 21787 11305
rect 22002 11296 22008 11308
rect 22060 11296 22066 11348
rect 22094 11296 22100 11348
rect 22152 11336 22158 11348
rect 23661 11339 23719 11345
rect 22152 11308 22197 11336
rect 22152 11296 22158 11308
rect 23661 11305 23673 11339
rect 23707 11336 23719 11339
rect 23750 11336 23756 11348
rect 23707 11308 23756 11336
rect 23707 11305 23719 11308
rect 23661 11299 23719 11305
rect 23750 11296 23756 11308
rect 23808 11296 23814 11348
rect 24026 11336 24032 11348
rect 23987 11308 24032 11336
rect 24026 11296 24032 11308
rect 24084 11296 24090 11348
rect 26234 11296 26240 11348
rect 26292 11336 26298 11348
rect 26789 11339 26847 11345
rect 26789 11336 26801 11339
rect 26292 11308 26801 11336
rect 26292 11296 26298 11308
rect 26789 11305 26801 11308
rect 26835 11305 26847 11339
rect 26789 11299 26847 11305
rect 3050 11268 3056 11280
rect 3011 11240 3056 11268
rect 3050 11228 3056 11240
rect 3108 11228 3114 11280
rect 3602 11228 3608 11280
rect 3660 11268 3666 11280
rect 6089 11271 6147 11277
rect 6089 11268 6101 11271
rect 3660 11240 6101 11268
rect 3660 11228 3666 11240
rect 6089 11237 6101 11240
rect 6135 11237 6147 11271
rect 8662 11268 8668 11280
rect 8623 11240 8668 11268
rect 6089 11231 6147 11237
rect 8662 11228 8668 11240
rect 8720 11228 8726 11280
rect 11330 11228 11336 11280
rect 11388 11228 11394 11280
rect 12158 11268 12164 11280
rect 12119 11240 12164 11268
rect 12158 11228 12164 11240
rect 12216 11228 12222 11280
rect 17405 11271 17463 11277
rect 17405 11268 17417 11271
rect 16224 11240 17417 11268
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 1946 11200 1952 11212
rect 1443 11172 1952 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 1946 11160 1952 11172
rect 2004 11160 2010 11212
rect 4709 11203 4767 11209
rect 4709 11169 4721 11203
rect 4755 11200 4767 11203
rect 4798 11200 4804 11212
rect 4755 11172 4804 11200
rect 4755 11169 4767 11172
rect 4709 11163 4767 11169
rect 4798 11160 4804 11172
rect 4856 11160 4862 11212
rect 5074 11200 5080 11212
rect 5035 11172 5080 11200
rect 5074 11160 5080 11172
rect 5132 11160 5138 11212
rect 5261 11203 5319 11209
rect 5261 11169 5273 11203
rect 5307 11200 5319 11203
rect 5442 11200 5448 11212
rect 5307 11172 5448 11200
rect 5307 11169 5319 11172
rect 5261 11163 5319 11169
rect 1578 11092 1584 11144
rect 1636 11132 1642 11144
rect 1673 11135 1731 11141
rect 1673 11132 1685 11135
rect 1636 11104 1685 11132
rect 1636 11092 1642 11104
rect 1673 11101 1685 11104
rect 1719 11101 1731 11135
rect 4154 11132 4160 11144
rect 4115 11104 4160 11132
rect 1673 11095 1731 11101
rect 4154 11092 4160 11104
rect 4212 11092 4218 11144
rect 4614 11132 4620 11144
rect 4575 11104 4620 11132
rect 4614 11092 4620 11104
rect 4672 11092 4678 11144
rect 3418 11024 3424 11076
rect 3476 11064 3482 11076
rect 3513 11067 3571 11073
rect 3513 11064 3525 11067
rect 3476 11036 3525 11064
rect 3476 11024 3482 11036
rect 3513 11033 3525 11036
rect 3559 11064 3571 11067
rect 3970 11064 3976 11076
rect 3559 11036 3976 11064
rect 3559 11033 3571 11036
rect 3513 11027 3571 11033
rect 3970 11024 3976 11036
rect 4028 11024 4034 11076
rect 5276 11064 5304 11163
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 6730 11200 6736 11212
rect 6691 11172 6736 11200
rect 6730 11160 6736 11172
rect 6788 11160 6794 11212
rect 6914 11160 6920 11212
rect 6972 11200 6978 11212
rect 7101 11203 7159 11209
rect 7101 11200 7113 11203
rect 6972 11172 7113 11200
rect 6972 11160 6978 11172
rect 7101 11169 7113 11172
rect 7147 11169 7159 11203
rect 8202 11200 8208 11212
rect 8163 11172 8208 11200
rect 7101 11163 7159 11169
rect 8202 11160 8208 11172
rect 8260 11160 8266 11212
rect 10318 11160 10324 11212
rect 10376 11200 10382 11212
rect 10873 11203 10931 11209
rect 10873 11200 10885 11203
rect 10376 11172 10885 11200
rect 10376 11160 10382 11172
rect 10873 11169 10885 11172
rect 10919 11169 10931 11203
rect 11054 11200 11060 11212
rect 11015 11172 11060 11200
rect 10873 11163 10931 11169
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 11348 11200 11376 11228
rect 11609 11203 11667 11209
rect 11609 11200 11621 11203
rect 11348 11172 11621 11200
rect 11609 11169 11621 11172
rect 11655 11169 11667 11203
rect 11790 11200 11796 11212
rect 11751 11172 11796 11200
rect 11609 11163 11667 11169
rect 11790 11160 11796 11172
rect 11848 11160 11854 11212
rect 13630 11200 13636 11212
rect 13591 11172 13636 11200
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 13814 11160 13820 11212
rect 13872 11200 13878 11212
rect 13909 11203 13967 11209
rect 13909 11200 13921 11203
rect 13872 11172 13921 11200
rect 13872 11160 13878 11172
rect 13909 11169 13921 11172
rect 13955 11169 13967 11203
rect 13909 11163 13967 11169
rect 15102 11160 15108 11212
rect 15160 11200 15166 11212
rect 15473 11203 15531 11209
rect 15473 11200 15485 11203
rect 15160 11172 15485 11200
rect 15160 11160 15166 11172
rect 15473 11169 15485 11172
rect 15519 11169 15531 11203
rect 15473 11163 15531 11169
rect 15565 11203 15623 11209
rect 15565 11169 15577 11203
rect 15611 11200 15623 11203
rect 15838 11200 15844 11212
rect 15611 11172 15844 11200
rect 15611 11169 15623 11172
rect 15565 11163 15623 11169
rect 15838 11160 15844 11172
rect 15896 11160 15902 11212
rect 16022 11200 16028 11212
rect 15983 11172 16028 11200
rect 16022 11160 16028 11172
rect 16080 11160 16086 11212
rect 16114 11160 16120 11212
rect 16172 11200 16178 11212
rect 16224 11209 16252 11240
rect 17405 11237 17417 11240
rect 17451 11268 17463 11271
rect 17494 11268 17500 11280
rect 17451 11240 17500 11268
rect 17451 11237 17463 11240
rect 17405 11231 17463 11237
rect 17494 11228 17500 11240
rect 17552 11228 17558 11280
rect 19426 11228 19432 11280
rect 19484 11268 19490 11280
rect 19613 11271 19671 11277
rect 19613 11268 19625 11271
rect 19484 11240 19625 11268
rect 19484 11228 19490 11240
rect 19613 11237 19625 11240
rect 19659 11268 19671 11271
rect 20530 11268 20536 11280
rect 19659 11240 20536 11268
rect 19659 11237 19671 11240
rect 19613 11231 19671 11237
rect 20530 11228 20536 11240
rect 20588 11228 20594 11280
rect 25222 11268 25228 11280
rect 25183 11240 25228 11268
rect 25222 11228 25228 11240
rect 25280 11228 25286 11280
rect 29917 11271 29975 11277
rect 29917 11237 29929 11271
rect 29963 11268 29975 11271
rect 31478 11268 31484 11280
rect 29963 11240 31484 11268
rect 29963 11237 29975 11240
rect 29917 11231 29975 11237
rect 16209 11203 16267 11209
rect 16209 11200 16221 11203
rect 16172 11172 16221 11200
rect 16172 11160 16178 11172
rect 16209 11169 16221 11172
rect 16255 11169 16267 11203
rect 16209 11163 16267 11169
rect 17589 11203 17647 11209
rect 17589 11169 17601 11203
rect 17635 11169 17647 11203
rect 17589 11163 17647 11169
rect 19061 11203 19119 11209
rect 19061 11169 19073 11203
rect 19107 11200 19119 11203
rect 19242 11200 19248 11212
rect 19107 11172 19248 11200
rect 19107 11169 19119 11172
rect 19061 11163 19119 11169
rect 6270 11092 6276 11144
rect 6328 11132 6334 11144
rect 6549 11135 6607 11141
rect 6549 11132 6561 11135
rect 6328 11104 6561 11132
rect 6328 11092 6334 11104
rect 6549 11101 6561 11104
rect 6595 11101 6607 11135
rect 6549 11095 6607 11101
rect 7009 11135 7067 11141
rect 7009 11101 7021 11135
rect 7055 11101 7067 11135
rect 7926 11132 7932 11144
rect 7887 11104 7932 11132
rect 7009 11095 7067 11101
rect 5537 11067 5595 11073
rect 5537 11064 5549 11067
rect 4080 11036 5304 11064
rect 5460 11036 5549 11064
rect 3694 10956 3700 11008
rect 3752 10996 3758 11008
rect 4080 10996 4108 11036
rect 3752 10968 4108 10996
rect 3752 10956 3758 10968
rect 4706 10956 4712 11008
rect 4764 10996 4770 11008
rect 5460 10996 5488 11036
rect 5537 11033 5549 11036
rect 5583 11064 5595 11067
rect 6454 11064 6460 11076
rect 5583 11036 6460 11064
rect 5583 11033 5595 11036
rect 5537 11027 5595 11033
rect 6454 11024 6460 11036
rect 6512 11024 6518 11076
rect 4764 10968 5488 10996
rect 4764 10956 4770 10968
rect 5626 10956 5632 11008
rect 5684 10996 5690 11008
rect 6546 10996 6552 11008
rect 5684 10968 6552 10996
rect 5684 10956 5690 10968
rect 6546 10956 6552 10968
rect 6604 10996 6610 11008
rect 7024 10996 7052 11095
rect 7926 11092 7932 11104
rect 7984 11092 7990 11144
rect 8110 11132 8116 11144
rect 8071 11104 8116 11132
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 10778 11132 10784 11144
rect 10739 11104 10784 11132
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 13170 11132 13176 11144
rect 13131 11104 13176 11132
rect 13170 11092 13176 11104
rect 13228 11092 13234 11144
rect 17402 11092 17408 11144
rect 17460 11132 17466 11144
rect 17604 11132 17632 11163
rect 19242 11160 19248 11172
rect 19300 11160 19306 11212
rect 23477 11203 23535 11209
rect 23477 11169 23489 11203
rect 23523 11200 23535 11203
rect 24118 11200 24124 11212
rect 23523 11172 24124 11200
rect 23523 11169 23535 11172
rect 23477 11163 23535 11169
rect 24118 11160 24124 11172
rect 24176 11160 24182 11212
rect 24854 11200 24860 11212
rect 24815 11172 24860 11200
rect 24854 11160 24860 11172
rect 24912 11160 24918 11212
rect 26234 11160 26240 11212
rect 26292 11200 26298 11212
rect 26605 11203 26663 11209
rect 26605 11200 26617 11203
rect 26292 11172 26617 11200
rect 26292 11160 26298 11172
rect 26605 11169 26617 11172
rect 26651 11200 26663 11203
rect 27798 11200 27804 11212
rect 26651 11172 27804 11200
rect 26651 11169 26663 11172
rect 26605 11163 26663 11169
rect 27798 11160 27804 11172
rect 27856 11160 27862 11212
rect 28534 11200 28540 11212
rect 28495 11172 28540 11200
rect 28534 11160 28540 11172
rect 28592 11160 28598 11212
rect 30650 11200 30656 11212
rect 30611 11172 30656 11200
rect 30650 11160 30656 11172
rect 30708 11160 30714 11212
rect 30742 11160 30748 11212
rect 30800 11200 30806 11212
rect 31018 11200 31024 11212
rect 30800 11172 30845 11200
rect 30979 11172 31024 11200
rect 30800 11160 30806 11172
rect 31018 11160 31024 11172
rect 31076 11160 31082 11212
rect 31128 11209 31156 11240
rect 31478 11228 31484 11240
rect 31536 11228 31542 11280
rect 31113 11203 31171 11209
rect 31113 11169 31125 11203
rect 31159 11169 31171 11203
rect 31113 11163 31171 11169
rect 17460 11104 17632 11132
rect 17460 11092 17466 11104
rect 23750 11092 23756 11144
rect 23808 11132 23814 11144
rect 27065 11135 27123 11141
rect 27065 11132 27077 11135
rect 23808 11104 27077 11132
rect 23808 11092 23814 11104
rect 27065 11101 27077 11104
rect 27111 11132 27123 11135
rect 27338 11132 27344 11144
rect 27111 11104 27344 11132
rect 27111 11101 27123 11104
rect 27065 11095 27123 11101
rect 27338 11092 27344 11104
rect 27396 11132 27402 11144
rect 27614 11132 27620 11144
rect 27396 11104 27620 11132
rect 27396 11092 27402 11104
rect 27614 11092 27620 11104
rect 27672 11092 27678 11144
rect 29914 11092 29920 11144
rect 29972 11132 29978 11144
rect 30009 11135 30067 11141
rect 30009 11132 30021 11135
rect 29972 11104 30021 11132
rect 29972 11092 29978 11104
rect 30009 11101 30021 11104
rect 30055 11101 30067 11135
rect 30009 11095 30067 11101
rect 12621 11067 12679 11073
rect 12621 11033 12633 11067
rect 12667 11064 12679 11067
rect 13078 11064 13084 11076
rect 12667 11036 13084 11064
rect 12667 11033 12679 11036
rect 12621 11027 12679 11033
rect 13078 11024 13084 11036
rect 13136 11064 13142 11076
rect 13909 11067 13967 11073
rect 13909 11064 13921 11067
rect 13136 11036 13921 11064
rect 13136 11024 13142 11036
rect 13909 11033 13921 11036
rect 13955 11033 13967 11067
rect 13909 11027 13967 11033
rect 25593 11067 25651 11073
rect 25593 11033 25605 11067
rect 25639 11064 25651 11067
rect 26145 11067 26203 11073
rect 26145 11064 26157 11067
rect 25639 11036 26157 11064
rect 25639 11033 25651 11036
rect 25593 11027 25651 11033
rect 26145 11033 26157 11036
rect 26191 11064 26203 11067
rect 26970 11064 26976 11076
rect 26191 11036 26976 11064
rect 26191 11033 26203 11036
rect 26145 11027 26203 11033
rect 26970 11024 26976 11036
rect 27028 11064 27034 11076
rect 27525 11067 27583 11073
rect 27525 11064 27537 11067
rect 27028 11036 27537 11064
rect 27028 11024 27034 11036
rect 27525 11033 27537 11036
rect 27571 11064 27583 11067
rect 28905 11067 28963 11073
rect 27571 11036 27660 11064
rect 27571 11033 27583 11036
rect 27525 11027 27583 11033
rect 6604 10968 7052 10996
rect 6604 10956 6610 10968
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 9033 10999 9091 11005
rect 9033 10996 9045 10999
rect 8352 10968 9045 10996
rect 8352 10956 8358 10968
rect 9033 10965 9045 10968
rect 9079 10996 9091 10999
rect 9490 10996 9496 11008
rect 9079 10968 9496 10996
rect 9079 10965 9091 10968
rect 9033 10959 9091 10965
rect 9490 10956 9496 10968
rect 9548 10956 9554 11008
rect 10134 10956 10140 11008
rect 10192 10996 10198 11008
rect 10229 10999 10287 11005
rect 10229 10996 10241 10999
rect 10192 10968 10241 10996
rect 10192 10956 10198 10968
rect 10229 10965 10241 10968
rect 10275 10965 10287 10999
rect 27632 10996 27660 11036
rect 28905 11033 28917 11067
rect 28951 11064 28963 11067
rect 28994 11064 29000 11076
rect 28951 11036 29000 11064
rect 28951 11033 28963 11036
rect 28905 11027 28963 11033
rect 28994 11024 29000 11036
rect 29052 11024 29058 11076
rect 27706 10996 27712 11008
rect 27632 10968 27712 10996
rect 10229 10959 10287 10965
rect 27706 10956 27712 10968
rect 27764 10956 27770 11008
rect 35342 10956 35348 11008
rect 35400 10996 35406 11008
rect 35802 10996 35808 11008
rect 35400 10968 35808 10996
rect 35400 10956 35406 10968
rect 35802 10956 35808 10968
rect 35860 10956 35866 11008
rect 1104 10906 38548 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 38548 10906
rect 1104 10832 38548 10854
rect 3694 10792 3700 10804
rect 3655 10764 3700 10792
rect 3694 10752 3700 10764
rect 3752 10752 3758 10804
rect 4525 10795 4583 10801
rect 4525 10761 4537 10795
rect 4571 10792 4583 10795
rect 4798 10792 4804 10804
rect 4571 10764 4804 10792
rect 4571 10761 4583 10764
rect 4525 10755 4583 10761
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 8202 10792 8208 10804
rect 8163 10764 8208 10792
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 8478 10792 8484 10804
rect 8439 10764 8484 10792
rect 8478 10752 8484 10764
rect 8536 10752 8542 10804
rect 10318 10752 10324 10804
rect 10376 10792 10382 10804
rect 10505 10795 10563 10801
rect 10505 10792 10517 10795
rect 10376 10764 10517 10792
rect 10376 10752 10382 10764
rect 10505 10761 10517 10764
rect 10551 10761 10563 10795
rect 13170 10792 13176 10804
rect 13131 10764 13176 10792
rect 10505 10755 10563 10761
rect 4157 10727 4215 10733
rect 4157 10693 4169 10727
rect 4203 10724 4215 10727
rect 4614 10724 4620 10736
rect 4203 10696 4620 10724
rect 4203 10693 4215 10696
rect 4157 10687 4215 10693
rect 4614 10684 4620 10696
rect 4672 10684 4678 10736
rect 9674 10684 9680 10736
rect 9732 10724 9738 10736
rect 9861 10727 9919 10733
rect 9861 10724 9873 10727
rect 9732 10696 9873 10724
rect 9732 10684 9738 10696
rect 9861 10693 9873 10696
rect 9907 10693 9919 10727
rect 10520 10724 10548 10755
rect 13170 10752 13176 10764
rect 13228 10792 13234 10804
rect 13906 10792 13912 10804
rect 13228 10764 13912 10792
rect 13228 10752 13234 10764
rect 13906 10752 13912 10764
rect 13964 10752 13970 10804
rect 14642 10792 14648 10804
rect 14603 10764 14648 10792
rect 14642 10752 14648 10764
rect 14700 10752 14706 10804
rect 15102 10752 15108 10804
rect 15160 10792 15166 10804
rect 15289 10795 15347 10801
rect 15289 10792 15301 10795
rect 15160 10764 15301 10792
rect 15160 10752 15166 10764
rect 15289 10761 15301 10764
rect 15335 10761 15347 10795
rect 15289 10755 15347 10761
rect 15749 10795 15807 10801
rect 15749 10761 15761 10795
rect 15795 10792 15807 10795
rect 16022 10792 16028 10804
rect 15795 10764 16028 10792
rect 15795 10761 15807 10764
rect 15749 10755 15807 10761
rect 16022 10752 16028 10764
rect 16080 10752 16086 10804
rect 16114 10752 16120 10804
rect 16172 10792 16178 10804
rect 16172 10764 16217 10792
rect 16172 10752 16178 10764
rect 19334 10752 19340 10804
rect 19392 10792 19398 10804
rect 20073 10795 20131 10801
rect 19392 10764 19437 10792
rect 19392 10752 19398 10764
rect 20073 10761 20085 10795
rect 20119 10792 20131 10795
rect 20254 10792 20260 10804
rect 20119 10764 20260 10792
rect 20119 10761 20131 10764
rect 20073 10755 20131 10761
rect 20254 10752 20260 10764
rect 20312 10752 20318 10804
rect 23937 10795 23995 10801
rect 23937 10761 23949 10795
rect 23983 10792 23995 10795
rect 24118 10792 24124 10804
rect 23983 10764 24124 10792
rect 23983 10761 23995 10764
rect 23937 10755 23995 10761
rect 24118 10752 24124 10764
rect 24176 10752 24182 10804
rect 25314 10792 25320 10804
rect 25275 10764 25320 10792
rect 25314 10752 25320 10764
rect 25372 10752 25378 10804
rect 25685 10795 25743 10801
rect 25685 10761 25697 10795
rect 25731 10792 25743 10795
rect 25866 10792 25872 10804
rect 25731 10764 25872 10792
rect 25731 10761 25743 10764
rect 25685 10755 25743 10761
rect 12526 10724 12532 10736
rect 10520 10696 12532 10724
rect 9861 10687 9919 10693
rect 12526 10684 12532 10696
rect 12584 10684 12590 10736
rect 12710 10684 12716 10736
rect 12768 10724 12774 10736
rect 12805 10727 12863 10733
rect 12805 10724 12817 10727
rect 12768 10696 12817 10724
rect 12768 10684 12774 10696
rect 12805 10693 12817 10696
rect 12851 10724 12863 10727
rect 13630 10724 13636 10736
rect 12851 10696 13636 10724
rect 12851 10693 12863 10696
rect 12805 10687 12863 10693
rect 13630 10684 13636 10696
rect 13688 10684 13694 10736
rect 13814 10684 13820 10736
rect 13872 10724 13878 10736
rect 14660 10724 14688 10752
rect 16666 10724 16672 10736
rect 13872 10696 14688 10724
rect 16627 10696 16672 10724
rect 13872 10684 13878 10696
rect 16666 10684 16672 10696
rect 16724 10684 16730 10736
rect 24305 10727 24363 10733
rect 24305 10693 24317 10727
rect 24351 10724 24363 10727
rect 24351 10696 25176 10724
rect 24351 10693 24363 10696
rect 24305 10687 24363 10693
rect 14369 10659 14427 10665
rect 14369 10625 14381 10659
rect 14415 10656 14427 10659
rect 15378 10656 15384 10668
rect 14415 10628 15384 10656
rect 14415 10625 14427 10628
rect 14369 10619 14427 10625
rect 15378 10616 15384 10628
rect 15436 10616 15442 10668
rect 4706 10548 4712 10600
rect 4764 10588 4770 10600
rect 4801 10591 4859 10597
rect 4801 10588 4813 10591
rect 4764 10560 4813 10588
rect 4764 10548 4770 10560
rect 4801 10557 4813 10560
rect 4847 10557 4859 10591
rect 4801 10551 4859 10557
rect 5813 10591 5871 10597
rect 5813 10557 5825 10591
rect 5859 10588 5871 10591
rect 6730 10588 6736 10600
rect 5859 10560 6736 10588
rect 5859 10557 5871 10560
rect 5813 10551 5871 10557
rect 6730 10548 6736 10560
rect 6788 10548 6794 10600
rect 8662 10588 8668 10600
rect 8623 10560 8668 10588
rect 8662 10548 8668 10560
rect 8720 10548 8726 10600
rect 8754 10548 8760 10600
rect 8812 10588 8818 10600
rect 8938 10588 8944 10600
rect 8812 10560 8857 10588
rect 8899 10560 8944 10588
rect 8812 10548 8818 10560
rect 8938 10548 8944 10560
rect 8996 10548 9002 10600
rect 9398 10588 9404 10600
rect 9359 10560 9404 10588
rect 9398 10548 9404 10560
rect 9456 10548 9462 10600
rect 9490 10548 9496 10600
rect 9548 10588 9554 10600
rect 12253 10591 12311 10597
rect 9548 10560 9593 10588
rect 9548 10548 9554 10560
rect 12253 10557 12265 10591
rect 12299 10588 12311 10591
rect 12802 10588 12808 10600
rect 12299 10560 12808 10588
rect 12299 10557 12311 10560
rect 12253 10551 12311 10557
rect 12802 10548 12808 10560
rect 12860 10588 12866 10600
rect 12989 10591 13047 10597
rect 12989 10588 13001 10591
rect 12860 10560 13001 10588
rect 12860 10548 12866 10560
rect 12989 10557 13001 10560
rect 13035 10557 13047 10591
rect 14458 10588 14464 10600
rect 14419 10560 14464 10588
rect 12989 10551 13047 10557
rect 14458 10548 14464 10560
rect 14516 10588 14522 10600
rect 14921 10591 14979 10597
rect 14921 10588 14933 10591
rect 14516 10560 14933 10588
rect 14516 10548 14522 10560
rect 14921 10557 14933 10560
rect 14967 10557 14979 10591
rect 14921 10551 14979 10557
rect 15930 10548 15936 10600
rect 15988 10588 15994 10600
rect 16301 10591 16359 10597
rect 16301 10588 16313 10591
rect 15988 10560 16313 10588
rect 15988 10548 15994 10560
rect 16301 10557 16313 10560
rect 16347 10557 16359 10591
rect 16301 10551 16359 10557
rect 17865 10591 17923 10597
rect 17865 10557 17877 10591
rect 17911 10588 17923 10591
rect 18414 10588 18420 10600
rect 17911 10560 18420 10588
rect 17911 10557 17923 10560
rect 17865 10551 17923 10557
rect 18414 10548 18420 10560
rect 18472 10588 18478 10600
rect 19889 10591 19947 10597
rect 19889 10588 19901 10591
rect 18472 10560 19901 10588
rect 18472 10548 18478 10560
rect 19889 10557 19901 10560
rect 19935 10588 19947 10591
rect 20349 10591 20407 10597
rect 20349 10588 20361 10591
rect 19935 10560 20361 10588
rect 19935 10557 19947 10560
rect 19889 10551 19947 10557
rect 20349 10557 20361 10560
rect 20395 10557 20407 10591
rect 24118 10588 24124 10600
rect 24079 10560 24124 10588
rect 20349 10551 20407 10557
rect 24118 10548 24124 10560
rect 24176 10588 24182 10600
rect 24581 10591 24639 10597
rect 24581 10588 24593 10591
rect 24176 10560 24593 10588
rect 24176 10548 24182 10560
rect 24581 10557 24593 10560
rect 24627 10588 24639 10591
rect 24854 10588 24860 10600
rect 24627 10560 24860 10588
rect 24627 10557 24639 10560
rect 24581 10551 24639 10557
rect 24854 10548 24860 10560
rect 24912 10588 24918 10600
rect 25148 10597 25176 10696
rect 24949 10591 25007 10597
rect 24949 10588 24961 10591
rect 24912 10560 24961 10588
rect 24912 10548 24918 10560
rect 24949 10557 24961 10560
rect 24995 10557 25007 10591
rect 24949 10551 25007 10557
rect 25133 10591 25191 10597
rect 25133 10557 25145 10591
rect 25179 10588 25191 10591
rect 25700 10588 25728 10755
rect 25866 10752 25872 10764
rect 25924 10752 25930 10804
rect 27706 10752 27712 10804
rect 27764 10792 27770 10804
rect 28077 10795 28135 10801
rect 28077 10792 28089 10795
rect 27764 10764 28089 10792
rect 27764 10752 27770 10764
rect 28077 10761 28089 10764
rect 28123 10761 28135 10795
rect 28077 10755 28135 10761
rect 28534 10752 28540 10804
rect 28592 10792 28598 10804
rect 28629 10795 28687 10801
rect 28629 10792 28641 10795
rect 28592 10764 28641 10792
rect 28592 10752 28598 10764
rect 28629 10761 28641 10764
rect 28675 10761 28687 10795
rect 28629 10755 28687 10761
rect 28994 10752 29000 10804
rect 29052 10792 29058 10804
rect 29641 10795 29699 10801
rect 29641 10792 29653 10795
rect 29052 10764 29653 10792
rect 29052 10752 29058 10764
rect 29641 10761 29653 10764
rect 29687 10792 29699 10795
rect 30190 10792 30196 10804
rect 29687 10764 30196 10792
rect 29687 10761 29699 10764
rect 29641 10755 29699 10761
rect 30190 10752 30196 10764
rect 30248 10792 30254 10804
rect 31018 10792 31024 10804
rect 30248 10764 31024 10792
rect 30248 10752 30254 10764
rect 31018 10752 31024 10764
rect 31076 10752 31082 10804
rect 30101 10727 30159 10733
rect 30101 10693 30113 10727
rect 30147 10724 30159 10727
rect 30374 10724 30380 10736
rect 30147 10696 30380 10724
rect 30147 10693 30159 10696
rect 30101 10687 30159 10693
rect 30374 10684 30380 10696
rect 30432 10724 30438 10736
rect 30432 10696 30972 10724
rect 30432 10684 30438 10696
rect 26605 10659 26663 10665
rect 26605 10625 26617 10659
rect 26651 10656 26663 10659
rect 30742 10656 30748 10668
rect 26651 10628 27016 10656
rect 30703 10628 30748 10656
rect 26651 10625 26663 10628
rect 26605 10619 26663 10625
rect 26988 10600 27016 10628
rect 30742 10616 30748 10628
rect 30800 10616 30806 10668
rect 25179 10560 25728 10588
rect 26697 10591 26755 10597
rect 25179 10557 25191 10560
rect 25133 10551 25191 10557
rect 26697 10557 26709 10591
rect 26743 10557 26755 10591
rect 26970 10588 26976 10600
rect 26931 10560 26976 10588
rect 26697 10551 26755 10557
rect 5445 10523 5503 10529
rect 5445 10489 5457 10523
rect 5491 10520 5503 10523
rect 6822 10520 6828 10532
rect 5491 10492 6828 10520
rect 5491 10489 5503 10492
rect 5445 10483 5503 10489
rect 6822 10480 6828 10492
rect 6880 10480 6886 10532
rect 10965 10523 11023 10529
rect 10965 10489 10977 10523
rect 11011 10520 11023 10523
rect 11790 10520 11796 10532
rect 11011 10492 11796 10520
rect 11011 10489 11023 10492
rect 10965 10483 11023 10489
rect 11790 10480 11796 10492
rect 11848 10480 11854 10532
rect 18322 10520 18328 10532
rect 18283 10492 18328 10520
rect 18322 10480 18328 10492
rect 18380 10480 18386 10532
rect 1578 10452 1584 10464
rect 1539 10424 1584 10452
rect 1578 10412 1584 10424
rect 1636 10412 1642 10464
rect 1946 10452 1952 10464
rect 1907 10424 1952 10452
rect 1946 10412 1952 10424
rect 2004 10412 2010 10464
rect 3970 10412 3976 10464
rect 4028 10452 4034 10464
rect 4614 10452 4620 10464
rect 4028 10424 4620 10452
rect 4028 10412 4034 10424
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 6181 10455 6239 10461
rect 6181 10421 6193 10455
rect 6227 10452 6239 10455
rect 6270 10452 6276 10464
rect 6227 10424 6276 10452
rect 6227 10421 6239 10424
rect 6181 10415 6239 10421
rect 6270 10412 6276 10424
rect 6328 10412 6334 10464
rect 6546 10452 6552 10464
rect 6507 10424 6552 10452
rect 6546 10412 6552 10424
rect 6604 10412 6610 10464
rect 7837 10455 7895 10461
rect 7837 10421 7849 10455
rect 7883 10452 7895 10455
rect 8110 10452 8116 10464
rect 7883 10424 8116 10452
rect 7883 10421 7895 10424
rect 7837 10415 7895 10421
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 11330 10452 11336 10464
rect 11291 10424 11336 10452
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 11514 10412 11520 10464
rect 11572 10452 11578 10464
rect 11701 10455 11759 10461
rect 11701 10452 11713 10455
rect 11572 10424 11713 10452
rect 11572 10412 11578 10424
rect 11701 10421 11713 10424
rect 11747 10452 11759 10455
rect 15102 10452 15108 10464
rect 11747 10424 15108 10452
rect 11747 10421 11759 10424
rect 11701 10415 11759 10421
rect 15102 10412 15108 10424
rect 15160 10412 15166 10464
rect 17402 10452 17408 10464
rect 17363 10424 17408 10452
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 26142 10452 26148 10464
rect 26103 10424 26148 10452
rect 26142 10412 26148 10424
rect 26200 10412 26206 10464
rect 26712 10452 26740 10551
rect 26970 10548 26976 10560
rect 27028 10548 27034 10600
rect 30650 10548 30656 10600
rect 30708 10588 30714 10600
rect 30837 10591 30895 10597
rect 30837 10588 30849 10591
rect 30708 10560 30849 10588
rect 30708 10548 30714 10560
rect 30837 10557 30849 10560
rect 30883 10557 30895 10591
rect 30944 10588 30972 10696
rect 31036 10656 31064 10752
rect 31297 10659 31355 10665
rect 31297 10656 31309 10659
rect 31036 10628 31309 10656
rect 31297 10625 31309 10628
rect 31343 10625 31355 10659
rect 31297 10619 31355 10625
rect 31205 10591 31263 10597
rect 31205 10588 31217 10591
rect 30944 10560 31217 10588
rect 30837 10551 30895 10557
rect 31205 10557 31217 10560
rect 31251 10557 31263 10591
rect 31205 10551 31263 10557
rect 30193 10523 30251 10529
rect 30193 10489 30205 10523
rect 30239 10520 30251 10523
rect 31386 10520 31392 10532
rect 30239 10492 31392 10520
rect 30239 10489 30251 10492
rect 30193 10483 30251 10489
rect 31386 10480 31392 10492
rect 31444 10480 31450 10532
rect 27338 10452 27344 10464
rect 26712 10424 27344 10452
rect 27338 10412 27344 10424
rect 27396 10412 27402 10464
rect 30650 10412 30656 10464
rect 30708 10452 30714 10464
rect 31665 10455 31723 10461
rect 31665 10452 31677 10455
rect 30708 10424 31677 10452
rect 30708 10412 30714 10424
rect 31665 10421 31677 10424
rect 31711 10421 31723 10455
rect 31665 10415 31723 10421
rect 1104 10362 38548 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 38548 10362
rect 1104 10288 38548 10310
rect 4341 10251 4399 10257
rect 4341 10217 4353 10251
rect 4387 10248 4399 10251
rect 5074 10248 5080 10260
rect 4387 10220 5080 10248
rect 4387 10217 4399 10220
rect 4341 10211 4399 10217
rect 5074 10208 5080 10220
rect 5132 10208 5138 10260
rect 6822 10248 6828 10260
rect 6783 10220 6828 10248
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 8481 10251 8539 10257
rect 8481 10217 8493 10251
rect 8527 10248 8539 10251
rect 8662 10248 8668 10260
rect 8527 10220 8668 10248
rect 8527 10217 8539 10220
rect 8481 10211 8539 10217
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 9125 10251 9183 10257
rect 9125 10217 9137 10251
rect 9171 10248 9183 10251
rect 9398 10248 9404 10260
rect 9171 10220 9404 10248
rect 9171 10217 9183 10220
rect 9125 10211 9183 10217
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 11698 10208 11704 10260
rect 11756 10248 11762 10260
rect 11977 10251 12035 10257
rect 11977 10248 11989 10251
rect 11756 10220 11989 10248
rect 11756 10208 11762 10220
rect 11977 10217 11989 10220
rect 12023 10217 12035 10251
rect 11977 10211 12035 10217
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 13173 10251 13231 10257
rect 12492 10220 12537 10248
rect 12492 10208 12498 10220
rect 13173 10217 13185 10251
rect 13219 10248 13231 10251
rect 13722 10248 13728 10260
rect 13219 10220 13728 10248
rect 13219 10217 13231 10220
rect 13173 10211 13231 10217
rect 13722 10208 13728 10220
rect 13780 10208 13786 10260
rect 14829 10251 14887 10257
rect 14829 10217 14841 10251
rect 14875 10248 14887 10251
rect 16022 10248 16028 10260
rect 14875 10220 16028 10248
rect 14875 10217 14887 10220
rect 14829 10211 14887 10217
rect 16022 10208 16028 10220
rect 16080 10208 16086 10260
rect 16574 10248 16580 10260
rect 16535 10220 16580 10248
rect 16574 10208 16580 10220
rect 16632 10208 16638 10260
rect 17681 10251 17739 10257
rect 17681 10217 17693 10251
rect 17727 10248 17739 10251
rect 17862 10248 17868 10260
rect 17727 10220 17868 10248
rect 17727 10217 17739 10220
rect 17681 10211 17739 10217
rect 17862 10208 17868 10220
rect 17920 10208 17926 10260
rect 19150 10248 19156 10260
rect 19111 10220 19156 10248
rect 19150 10208 19156 10220
rect 19208 10208 19214 10260
rect 19521 10251 19579 10257
rect 19521 10217 19533 10251
rect 19567 10248 19579 10251
rect 20254 10248 20260 10260
rect 19567 10220 20260 10248
rect 19567 10217 19579 10220
rect 19521 10211 19579 10217
rect 19904 10192 19932 10220
rect 20254 10208 20260 10220
rect 20312 10208 20318 10260
rect 20346 10208 20352 10260
rect 20404 10248 20410 10260
rect 21729 10251 21787 10257
rect 21729 10248 21741 10251
rect 20404 10220 21741 10248
rect 20404 10208 20410 10220
rect 21729 10217 21741 10220
rect 21775 10248 21787 10251
rect 25590 10248 25596 10260
rect 21775 10220 22324 10248
rect 25551 10220 25596 10248
rect 21775 10217 21787 10220
rect 21729 10211 21787 10217
rect 4706 10180 4712 10192
rect 4667 10152 4712 10180
rect 4706 10140 4712 10152
rect 4764 10140 4770 10192
rect 12805 10183 12863 10189
rect 12805 10149 12817 10183
rect 12851 10180 12863 10183
rect 13262 10180 13268 10192
rect 12851 10152 13268 10180
rect 12851 10149 12863 10152
rect 12805 10143 12863 10149
rect 13262 10140 13268 10152
rect 13320 10180 13326 10192
rect 14366 10180 14372 10192
rect 13320 10152 14372 10180
rect 13320 10140 13326 10152
rect 14366 10140 14372 10152
rect 14424 10140 14430 10192
rect 15838 10180 15844 10192
rect 15799 10152 15844 10180
rect 15838 10140 15844 10152
rect 15896 10140 15902 10192
rect 15930 10140 15936 10192
rect 15988 10180 15994 10192
rect 16209 10183 16267 10189
rect 16209 10180 16221 10183
rect 15988 10152 16221 10180
rect 15988 10140 15994 10152
rect 16209 10149 16221 10152
rect 16255 10180 16267 10183
rect 16298 10180 16304 10192
rect 16255 10152 16304 10180
rect 16255 10149 16267 10152
rect 16209 10143 16267 10149
rect 16298 10140 16304 10152
rect 16356 10140 16362 10192
rect 19886 10140 19892 10192
rect 19944 10140 19950 10192
rect 5534 10112 5540 10124
rect 5495 10084 5540 10112
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 7098 10072 7104 10124
rect 7156 10112 7162 10124
rect 8573 10115 8631 10121
rect 7156 10084 8340 10112
rect 7156 10072 7162 10084
rect 4614 10004 4620 10056
rect 4672 10044 4678 10056
rect 5261 10047 5319 10053
rect 5261 10044 5273 10047
rect 4672 10016 5273 10044
rect 4672 10004 4678 10016
rect 5261 10013 5273 10016
rect 5307 10044 5319 10047
rect 5442 10044 5448 10056
rect 5307 10016 5448 10044
rect 5307 10013 5319 10016
rect 5261 10007 5319 10013
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 6546 10004 6552 10056
rect 6604 10044 6610 10056
rect 7377 10047 7435 10053
rect 7377 10044 7389 10047
rect 6604 10016 7389 10044
rect 6604 10004 6610 10016
rect 7377 10013 7389 10016
rect 7423 10044 7435 10047
rect 8202 10044 8208 10056
rect 7423 10016 8208 10044
rect 7423 10013 7435 10016
rect 7377 10007 7435 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 8312 10044 8340 10084
rect 8573 10081 8585 10115
rect 8619 10112 8631 10115
rect 8754 10112 8760 10124
rect 8619 10084 8760 10112
rect 8619 10081 8631 10084
rect 8573 10075 8631 10081
rect 8754 10072 8760 10084
rect 8812 10112 8818 10124
rect 9490 10112 9496 10124
rect 8812 10084 9496 10112
rect 8812 10072 8818 10084
rect 9490 10072 9496 10084
rect 9548 10072 9554 10124
rect 11422 10112 11428 10124
rect 11383 10084 11428 10112
rect 11422 10072 11428 10084
rect 11480 10072 11486 10124
rect 13446 10112 13452 10124
rect 13359 10084 13452 10112
rect 13446 10072 13452 10084
rect 13504 10112 13510 10124
rect 14458 10112 14464 10124
rect 13504 10084 14464 10112
rect 13504 10072 13510 10084
rect 14458 10072 14464 10084
rect 14516 10072 14522 10124
rect 15286 10112 15292 10124
rect 15247 10084 15292 10112
rect 15286 10072 15292 10084
rect 15344 10072 15350 10124
rect 16945 10115 17003 10121
rect 16945 10081 16957 10115
rect 16991 10112 17003 10115
rect 17957 10115 18015 10121
rect 17957 10112 17969 10115
rect 16991 10084 17969 10112
rect 16991 10081 17003 10084
rect 16945 10075 17003 10081
rect 17957 10081 17969 10084
rect 18003 10112 18015 10115
rect 18322 10112 18328 10124
rect 18003 10084 18328 10112
rect 18003 10081 18015 10084
rect 17957 10075 18015 10081
rect 18322 10072 18328 10084
rect 18380 10072 18386 10124
rect 18969 10115 19027 10121
rect 18969 10081 18981 10115
rect 19015 10112 19027 10115
rect 19058 10112 19064 10124
rect 19015 10084 19064 10112
rect 19015 10081 19027 10084
rect 18969 10075 19027 10081
rect 19058 10072 19064 10084
rect 19116 10072 19122 10124
rect 21910 10112 21916 10124
rect 21871 10084 21916 10112
rect 21910 10072 21916 10084
rect 21968 10072 21974 10124
rect 9582 10044 9588 10056
rect 8312 10016 9588 10044
rect 9582 10004 9588 10016
rect 9640 10004 9646 10056
rect 9674 10004 9680 10056
rect 9732 10004 9738 10056
rect 11701 10047 11759 10053
rect 11701 10013 11713 10047
rect 11747 10044 11759 10047
rect 11790 10044 11796 10056
rect 11747 10016 11796 10044
rect 11747 10013 11759 10016
rect 11701 10007 11759 10013
rect 11790 10004 11796 10016
rect 11848 10004 11854 10056
rect 12526 10004 12532 10056
rect 12584 10044 12590 10056
rect 13357 10047 13415 10053
rect 13357 10044 13369 10047
rect 12584 10016 13369 10044
rect 12584 10004 12590 10016
rect 13357 10013 13369 10016
rect 13403 10013 13415 10047
rect 13357 10007 13415 10013
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 22296 10053 22324 10220
rect 25590 10208 25596 10220
rect 25648 10208 25654 10260
rect 26973 10251 27031 10257
rect 26973 10217 26985 10251
rect 27019 10248 27031 10251
rect 27062 10248 27068 10260
rect 27019 10220 27068 10248
rect 27019 10217 27031 10220
rect 26973 10211 27031 10217
rect 27062 10208 27068 10220
rect 27120 10208 27126 10260
rect 27985 10251 28043 10257
rect 27985 10217 27997 10251
rect 28031 10248 28043 10251
rect 28074 10248 28080 10260
rect 28031 10220 28080 10248
rect 28031 10217 28043 10220
rect 27985 10211 28043 10217
rect 28074 10208 28080 10220
rect 28132 10208 28138 10260
rect 30190 10248 30196 10260
rect 30151 10220 30196 10248
rect 30190 10208 30196 10220
rect 30248 10208 30254 10260
rect 30653 10251 30711 10257
rect 30653 10217 30665 10251
rect 30699 10248 30711 10251
rect 30742 10248 30748 10260
rect 30699 10220 30748 10248
rect 30699 10217 30711 10220
rect 30653 10211 30711 10217
rect 30742 10208 30748 10220
rect 30800 10248 30806 10260
rect 30929 10251 30987 10257
rect 30929 10248 30941 10251
rect 30800 10220 30941 10248
rect 30800 10208 30806 10220
rect 30929 10217 30941 10220
rect 30975 10217 30987 10251
rect 30929 10211 30987 10217
rect 36078 10208 36084 10260
rect 36136 10248 36142 10260
rect 36541 10251 36599 10257
rect 36541 10248 36553 10251
rect 36136 10220 36553 10248
rect 36136 10208 36142 10220
rect 36541 10217 36553 10220
rect 36587 10217 36599 10251
rect 36541 10211 36599 10217
rect 23937 10183 23995 10189
rect 23937 10149 23949 10183
rect 23983 10180 23995 10183
rect 24118 10180 24124 10192
rect 23983 10152 24124 10180
rect 23983 10149 23995 10152
rect 23937 10143 23995 10149
rect 24118 10140 24124 10152
rect 24176 10140 24182 10192
rect 22370 10072 22376 10124
rect 22428 10112 22434 10124
rect 22557 10115 22615 10121
rect 22557 10112 22569 10115
rect 22428 10084 22569 10112
rect 22428 10072 22434 10084
rect 22557 10081 22569 10084
rect 22603 10081 22615 10115
rect 22557 10075 22615 10081
rect 24394 10072 24400 10124
rect 24452 10112 24458 10124
rect 25409 10115 25467 10121
rect 25409 10112 25421 10115
rect 24452 10084 25421 10112
rect 24452 10072 24458 10084
rect 25409 10081 25421 10084
rect 25455 10112 25467 10115
rect 25498 10112 25504 10124
rect 25455 10084 25504 10112
rect 25455 10081 25467 10084
rect 25409 10075 25467 10081
rect 25498 10072 25504 10084
rect 25556 10112 25562 10124
rect 26142 10112 26148 10124
rect 25556 10084 26148 10112
rect 25556 10072 25562 10084
rect 26142 10072 26148 10084
rect 26200 10072 26206 10124
rect 26786 10112 26792 10124
rect 26747 10084 26792 10112
rect 26786 10072 26792 10084
rect 26844 10072 26850 10124
rect 27614 10072 27620 10124
rect 27672 10112 27678 10124
rect 27801 10115 27859 10121
rect 27801 10112 27813 10115
rect 27672 10084 27813 10112
rect 27672 10072 27678 10084
rect 27801 10081 27813 10084
rect 27847 10081 27859 10115
rect 27801 10075 27859 10081
rect 29917 10115 29975 10121
rect 29917 10081 29929 10115
rect 29963 10112 29975 10115
rect 30650 10112 30656 10124
rect 29963 10084 30656 10112
rect 29963 10081 29975 10084
rect 29917 10075 29975 10081
rect 30650 10072 30656 10084
rect 30708 10072 30714 10124
rect 35250 10072 35256 10124
rect 35308 10112 35314 10124
rect 35437 10115 35495 10121
rect 35437 10112 35449 10115
rect 35308 10084 35449 10112
rect 35308 10072 35314 10084
rect 35437 10081 35449 10084
rect 35483 10081 35495 10115
rect 35437 10075 35495 10081
rect 13909 10047 13967 10053
rect 13909 10044 13921 10047
rect 13872 10016 13921 10044
rect 13872 10004 13878 10016
rect 13909 10013 13921 10016
rect 13955 10013 13967 10047
rect 13909 10007 13967 10013
rect 22281 10047 22339 10053
rect 22281 10013 22293 10047
rect 22327 10044 22339 10047
rect 22646 10044 22652 10056
rect 22327 10016 22652 10044
rect 22327 10013 22339 10016
rect 22281 10007 22339 10013
rect 22646 10004 22652 10016
rect 22704 10004 22710 10056
rect 35161 10047 35219 10053
rect 35161 10013 35173 10047
rect 35207 10044 35219 10047
rect 35342 10044 35348 10056
rect 35207 10016 35348 10044
rect 35207 10013 35219 10016
rect 35161 10007 35219 10013
rect 35342 10004 35348 10016
rect 35400 10004 35406 10056
rect 8110 9936 8116 9988
rect 8168 9976 8174 9988
rect 8754 9976 8760 9988
rect 8168 9948 8760 9976
rect 8168 9936 8174 9948
rect 8754 9936 8760 9948
rect 8812 9936 8818 9988
rect 9692 9976 9720 10004
rect 17126 9976 17132 9988
rect 9692 9948 17132 9976
rect 17126 9936 17132 9948
rect 17184 9936 17190 9988
rect 7745 9911 7803 9917
rect 7745 9877 7757 9911
rect 7791 9908 7803 9911
rect 8294 9908 8300 9920
rect 7791 9880 8300 9908
rect 7791 9877 7803 9880
rect 7745 9871 7803 9877
rect 8294 9868 8300 9880
rect 8352 9868 8358 9920
rect 9490 9908 9496 9920
rect 9451 9880 9496 9908
rect 9490 9868 9496 9880
rect 9548 9868 9554 9920
rect 14274 9908 14280 9920
rect 14235 9880 14280 9908
rect 14274 9868 14280 9880
rect 14332 9908 14338 9920
rect 15473 9911 15531 9917
rect 15473 9908 15485 9911
rect 14332 9880 15485 9908
rect 14332 9868 14338 9880
rect 15473 9877 15485 9880
rect 15519 9908 15531 9911
rect 15654 9908 15660 9920
rect 15519 9880 15660 9908
rect 15519 9877 15531 9880
rect 15473 9871 15531 9877
rect 15654 9868 15660 9880
rect 15712 9868 15718 9920
rect 18138 9908 18144 9920
rect 18099 9880 18144 9908
rect 18138 9868 18144 9880
rect 18196 9868 18202 9920
rect 18598 9868 18604 9920
rect 18656 9908 18662 9920
rect 18785 9911 18843 9917
rect 18785 9908 18797 9911
rect 18656 9880 18797 9908
rect 18656 9868 18662 9880
rect 18785 9877 18797 9880
rect 18831 9877 18843 9911
rect 18785 9871 18843 9877
rect 19518 9868 19524 9920
rect 19576 9908 19582 9920
rect 19797 9911 19855 9917
rect 19797 9908 19809 9911
rect 19576 9880 19809 9908
rect 19576 9868 19582 9880
rect 19797 9877 19809 9880
rect 19843 9877 19855 9911
rect 27338 9908 27344 9920
rect 27299 9880 27344 9908
rect 19797 9871 19855 9877
rect 27338 9868 27344 9880
rect 27396 9868 27402 9920
rect 1104 9818 38548 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 38548 9818
rect 1104 9744 38548 9766
rect 2590 9664 2596 9716
rect 2648 9704 2654 9716
rect 3878 9704 3884 9716
rect 2648 9676 3884 9704
rect 2648 9664 2654 9676
rect 3878 9664 3884 9676
rect 3936 9664 3942 9716
rect 11057 9707 11115 9713
rect 11057 9673 11069 9707
rect 11103 9704 11115 9707
rect 11422 9704 11428 9716
rect 11103 9676 11428 9704
rect 11103 9673 11115 9676
rect 11057 9667 11115 9673
rect 11422 9664 11428 9676
rect 11480 9664 11486 9716
rect 12526 9664 12532 9716
rect 12584 9704 12590 9716
rect 12621 9707 12679 9713
rect 12621 9704 12633 9707
rect 12584 9676 12633 9704
rect 12584 9664 12590 9676
rect 12621 9673 12633 9676
rect 12667 9673 12679 9707
rect 13446 9704 13452 9716
rect 13407 9676 13452 9704
rect 12621 9667 12679 9673
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 15286 9664 15292 9716
rect 15344 9704 15350 9716
rect 15381 9707 15439 9713
rect 15381 9704 15393 9707
rect 15344 9676 15393 9704
rect 15344 9664 15350 9676
rect 15381 9673 15393 9676
rect 15427 9673 15439 9707
rect 15381 9667 15439 9673
rect 17497 9707 17555 9713
rect 17497 9673 17509 9707
rect 17543 9704 17555 9707
rect 18322 9704 18328 9716
rect 17543 9676 18328 9704
rect 17543 9673 17555 9676
rect 17497 9667 17555 9673
rect 5353 9639 5411 9645
rect 5353 9605 5365 9639
rect 5399 9636 5411 9639
rect 5534 9636 5540 9648
rect 5399 9608 5540 9636
rect 5399 9605 5411 9608
rect 5353 9599 5411 9605
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 7193 9639 7251 9645
rect 7193 9605 7205 9639
rect 7239 9636 7251 9639
rect 11977 9639 12035 9645
rect 7239 9608 8064 9636
rect 7239 9605 7251 9608
rect 7193 9599 7251 9605
rect 1857 9571 1915 9577
rect 1857 9537 1869 9571
rect 1903 9568 1915 9571
rect 1903 9540 2268 9568
rect 1903 9537 1915 9540
rect 1857 9531 1915 9537
rect 1946 9500 1952 9512
rect 1907 9472 1952 9500
rect 1946 9460 1952 9472
rect 2004 9460 2010 9512
rect 2240 9509 2268 9540
rect 2866 9528 2872 9580
rect 2924 9568 2930 9580
rect 3329 9571 3387 9577
rect 3329 9568 3341 9571
rect 2924 9540 3341 9568
rect 2924 9528 2930 9540
rect 3329 9537 3341 9540
rect 3375 9537 3387 9571
rect 3329 9531 3387 9537
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 6730 9568 6736 9580
rect 6687 9540 6736 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 6730 9528 6736 9540
rect 6788 9568 6794 9580
rect 8036 9577 8064 9608
rect 11977 9605 11989 9639
rect 12023 9636 12035 9639
rect 12066 9636 12072 9648
rect 12023 9608 12072 9636
rect 12023 9605 12035 9608
rect 11977 9599 12035 9605
rect 12066 9596 12072 9608
rect 12124 9596 12130 9648
rect 14366 9636 14372 9648
rect 13832 9608 14372 9636
rect 8021 9571 8079 9577
rect 6788 9540 7972 9568
rect 6788 9528 6794 9540
rect 7944 9512 7972 9540
rect 8021 9537 8033 9571
rect 8067 9568 8079 9571
rect 8110 9568 8116 9580
rect 8067 9540 8116 9568
rect 8067 9537 8079 9540
rect 8021 9531 8079 9537
rect 8110 9528 8116 9540
rect 8168 9528 8174 9580
rect 8202 9528 8208 9580
rect 8260 9568 8266 9580
rect 13832 9577 13860 9608
rect 14366 9596 14372 9608
rect 14424 9596 14430 9648
rect 16485 9639 16543 9645
rect 16485 9605 16497 9639
rect 16531 9636 16543 9639
rect 17512 9636 17540 9667
rect 18322 9664 18328 9676
rect 18380 9664 18386 9716
rect 18877 9707 18935 9713
rect 18877 9673 18889 9707
rect 18923 9704 18935 9707
rect 19058 9704 19064 9716
rect 18923 9676 19064 9704
rect 18923 9673 18935 9676
rect 18877 9667 18935 9673
rect 19058 9664 19064 9676
rect 19116 9664 19122 9716
rect 20898 9664 20904 9716
rect 20956 9704 20962 9716
rect 21634 9704 21640 9716
rect 20956 9676 21640 9704
rect 20956 9664 20962 9676
rect 21634 9664 21640 9676
rect 21692 9664 21698 9716
rect 21821 9707 21879 9713
rect 21821 9673 21833 9707
rect 21867 9704 21879 9707
rect 21910 9704 21916 9716
rect 21867 9676 21916 9704
rect 21867 9673 21879 9676
rect 21821 9667 21879 9673
rect 21910 9664 21916 9676
rect 21968 9664 21974 9716
rect 26786 9704 26792 9716
rect 26747 9676 26792 9704
rect 26786 9664 26792 9676
rect 26844 9664 26850 9716
rect 27614 9664 27620 9716
rect 27672 9704 27678 9716
rect 27801 9707 27859 9713
rect 27801 9704 27813 9707
rect 27672 9676 27813 9704
rect 27672 9664 27678 9676
rect 27801 9673 27813 9676
rect 27847 9673 27859 9707
rect 27801 9667 27859 9673
rect 16531 9608 17540 9636
rect 16531 9605 16543 9608
rect 16485 9599 16543 9605
rect 13817 9571 13875 9577
rect 8260 9540 8305 9568
rect 8260 9528 8266 9540
rect 13817 9537 13829 9571
rect 13863 9537 13875 9571
rect 13817 9531 13875 9537
rect 2225 9503 2283 9509
rect 2225 9469 2237 9503
rect 2271 9500 2283 9503
rect 2314 9500 2320 9512
rect 2271 9472 2320 9500
rect 2271 9469 2283 9472
rect 2225 9463 2283 9469
rect 2314 9460 2320 9472
rect 2372 9460 2378 9512
rect 5442 9460 5448 9512
rect 5500 9500 5506 9512
rect 5721 9503 5779 9509
rect 5721 9500 5733 9503
rect 5500 9472 5733 9500
rect 5500 9460 5506 9472
rect 5721 9469 5733 9472
rect 5767 9500 5779 9503
rect 7098 9500 7104 9512
rect 5767 9472 7104 9500
rect 5767 9469 5779 9472
rect 5721 9463 5779 9469
rect 7098 9460 7104 9472
rect 7156 9460 7162 9512
rect 7926 9500 7932 9512
rect 7887 9472 7932 9500
rect 7926 9460 7932 9472
rect 7984 9460 7990 9512
rect 8294 9500 8300 9512
rect 8255 9472 8300 9500
rect 8294 9460 8300 9472
rect 8352 9460 8358 9512
rect 8846 9500 8852 9512
rect 8759 9472 8852 9500
rect 8846 9460 8852 9472
rect 8904 9500 8910 9512
rect 9490 9500 9496 9512
rect 8904 9472 9496 9500
rect 8904 9460 8910 9472
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 13909 9503 13967 9509
rect 13909 9469 13921 9503
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 7282 9432 7288 9444
rect 7243 9404 7288 9432
rect 7282 9392 7288 9404
rect 7340 9392 7346 9444
rect 13924 9432 13952 9463
rect 14090 9460 14096 9512
rect 14148 9500 14154 9512
rect 14369 9503 14427 9509
rect 14369 9500 14381 9503
rect 14148 9472 14381 9500
rect 14148 9460 14154 9472
rect 14369 9469 14381 9472
rect 14415 9469 14427 9503
rect 14369 9463 14427 9469
rect 14461 9503 14519 9509
rect 14461 9469 14473 9503
rect 14507 9469 14519 9503
rect 14461 9463 14519 9469
rect 15933 9503 15991 9509
rect 15933 9469 15945 9503
rect 15979 9500 15991 9503
rect 16500 9500 16528 9599
rect 19886 9596 19892 9648
rect 19944 9596 19950 9648
rect 25774 9636 25780 9648
rect 25735 9608 25780 9636
rect 25774 9596 25780 9608
rect 25832 9596 25838 9648
rect 35250 9636 35256 9648
rect 35211 9608 35256 9636
rect 35250 9596 35256 9608
rect 35308 9596 35314 9648
rect 18598 9528 18604 9580
rect 18656 9568 18662 9580
rect 19904 9568 19932 9596
rect 24305 9571 24363 9577
rect 18656 9540 19748 9568
rect 19904 9540 20208 9568
rect 18656 9528 18662 9540
rect 15979 9472 16528 9500
rect 16945 9503 17003 9509
rect 15979 9469 15991 9472
rect 15933 9463 15991 9469
rect 16945 9469 16957 9503
rect 16991 9500 17003 9503
rect 17221 9503 17279 9509
rect 17221 9500 17233 9503
rect 16991 9472 17233 9500
rect 16991 9469 17003 9472
rect 16945 9463 17003 9469
rect 17221 9469 17233 9472
rect 17267 9469 17279 9503
rect 17221 9463 17279 9469
rect 19429 9503 19487 9509
rect 19429 9469 19441 9503
rect 19475 9500 19487 9503
rect 19518 9500 19524 9512
rect 19475 9472 19524 9500
rect 19475 9469 19487 9472
rect 19429 9463 19487 9469
rect 14274 9432 14280 9444
rect 13924 9404 14280 9432
rect 12986 9364 12992 9376
rect 12947 9336 12992 9364
rect 12986 9324 12992 9336
rect 13044 9364 13050 9376
rect 13924 9364 13952 9404
rect 14274 9392 14280 9404
rect 14332 9432 14338 9444
rect 14476 9432 14504 9463
rect 15010 9432 15016 9444
rect 14332 9404 14504 9432
rect 14971 9404 15016 9432
rect 14332 9392 14338 9404
rect 15010 9392 15016 9404
rect 15068 9392 15074 9444
rect 19058 9432 19064 9444
rect 17144 9404 19064 9432
rect 16114 9364 16120 9376
rect 13044 9336 13952 9364
rect 16075 9336 16120 9364
rect 13044 9324 13050 9336
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 17144 9373 17172 9404
rect 19058 9392 19064 9404
rect 19116 9432 19122 9444
rect 19444 9432 19472 9463
rect 19518 9460 19524 9472
rect 19576 9460 19582 9512
rect 19613 9503 19671 9509
rect 19613 9469 19625 9503
rect 19659 9469 19671 9503
rect 19720 9500 19748 9540
rect 20180 9509 20208 9540
rect 24305 9537 24317 9571
rect 24351 9568 24363 9571
rect 24351 9540 24716 9568
rect 24351 9537 24363 9540
rect 24305 9531 24363 9537
rect 24688 9512 24716 9540
rect 35066 9528 35072 9580
rect 35124 9568 35130 9580
rect 35342 9568 35348 9580
rect 35124 9540 35348 9568
rect 35124 9528 35130 9540
rect 35342 9528 35348 9540
rect 35400 9568 35406 9580
rect 35529 9571 35587 9577
rect 35529 9568 35541 9571
rect 35400 9540 35541 9568
rect 35400 9528 35406 9540
rect 35529 9537 35541 9540
rect 35575 9537 35587 9571
rect 35529 9531 35587 9537
rect 19935 9503 19993 9509
rect 19935 9500 19947 9503
rect 19720 9472 19947 9500
rect 19613 9463 19671 9469
rect 19935 9469 19947 9472
rect 19981 9469 19993 9503
rect 19935 9463 19993 9469
rect 20165 9503 20223 9509
rect 20165 9469 20177 9503
rect 20211 9469 20223 9503
rect 20165 9463 20223 9469
rect 23477 9503 23535 9509
rect 23477 9469 23489 9503
rect 23523 9469 23535 9503
rect 24394 9500 24400 9512
rect 24355 9472 24400 9500
rect 23477 9463 23535 9469
rect 19116 9404 19472 9432
rect 19628 9432 19656 9463
rect 20441 9435 20499 9441
rect 20441 9432 20453 9435
rect 19628 9404 20453 9432
rect 19116 9392 19122 9404
rect 19996 9376 20024 9404
rect 20441 9401 20453 9404
rect 20487 9401 20499 9435
rect 20441 9395 20499 9401
rect 21910 9392 21916 9444
rect 21968 9432 21974 9444
rect 21968 9404 23336 9432
rect 21968 9392 21974 9404
rect 23308 9376 23336 9404
rect 23492 9376 23520 9463
rect 24394 9460 24400 9472
rect 24452 9460 24458 9512
rect 24670 9500 24676 9512
rect 24631 9472 24676 9500
rect 24670 9460 24676 9472
rect 24728 9460 24734 9512
rect 17129 9367 17187 9373
rect 17129 9333 17141 9367
rect 17175 9333 17187 9367
rect 17129 9327 17187 9333
rect 17221 9367 17279 9373
rect 17221 9333 17233 9367
rect 17267 9364 17279 9367
rect 17865 9367 17923 9373
rect 17865 9364 17877 9367
rect 17267 9336 17877 9364
rect 17267 9333 17279 9336
rect 17221 9327 17279 9333
rect 17865 9333 17877 9336
rect 17911 9364 17923 9367
rect 18230 9364 18236 9376
rect 17911 9336 18236 9364
rect 17911 9333 17923 9336
rect 17865 9327 17923 9333
rect 18230 9324 18236 9336
rect 18288 9324 18294 9376
rect 19242 9364 19248 9376
rect 19203 9336 19248 9364
rect 19242 9324 19248 9336
rect 19300 9324 19306 9376
rect 19978 9324 19984 9376
rect 20036 9324 20042 9376
rect 22278 9364 22284 9376
rect 22239 9336 22284 9364
rect 22278 9324 22284 9336
rect 22336 9324 22342 9376
rect 22646 9364 22652 9376
rect 22607 9336 22652 9364
rect 22646 9324 22652 9336
rect 22704 9324 22710 9376
rect 23290 9364 23296 9376
rect 23203 9336 23296 9364
rect 23290 9324 23296 9336
rect 23348 9324 23354 9376
rect 23474 9324 23480 9376
rect 23532 9364 23538 9376
rect 23845 9367 23903 9373
rect 23845 9364 23857 9367
rect 23532 9336 23857 9364
rect 23532 9324 23538 9336
rect 23845 9333 23857 9336
rect 23891 9333 23903 9367
rect 23845 9327 23903 9333
rect 1104 9274 38548 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 38548 9274
rect 1104 9200 38548 9222
rect 1946 9160 1952 9172
rect 1907 9132 1952 9160
rect 1946 9120 1952 9132
rect 2004 9120 2010 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 8481 9163 8539 9169
rect 8481 9160 8493 9163
rect 8352 9132 8493 9160
rect 8352 9120 8358 9132
rect 8481 9129 8493 9132
rect 8527 9129 8539 9163
rect 8481 9123 8539 9129
rect 9674 9120 9680 9172
rect 9732 9160 9738 9172
rect 9950 9160 9956 9172
rect 9732 9132 9956 9160
rect 9732 9120 9738 9132
rect 9950 9120 9956 9132
rect 10008 9160 10014 9172
rect 10045 9163 10103 9169
rect 10045 9160 10057 9163
rect 10008 9132 10057 9160
rect 10008 9120 10014 9132
rect 10045 9129 10057 9132
rect 10091 9160 10103 9163
rect 11146 9160 11152 9172
rect 10091 9132 11152 9160
rect 10091 9129 10103 9132
rect 10045 9123 10103 9129
rect 11146 9120 11152 9132
rect 11204 9120 11210 9172
rect 12618 9160 12624 9172
rect 12579 9132 12624 9160
rect 12618 9120 12624 9132
rect 12676 9160 12682 9172
rect 13906 9160 13912 9172
rect 12676 9132 13400 9160
rect 13867 9132 13912 9160
rect 12676 9120 12682 9132
rect 12986 9092 12992 9104
rect 11624 9064 12992 9092
rect 11624 9036 11652 9064
rect 12986 9052 12992 9064
rect 13044 9052 13050 9104
rect 13372 9092 13400 9132
rect 13906 9120 13912 9132
rect 13964 9120 13970 9172
rect 24394 9120 24400 9172
rect 24452 9160 24458 9172
rect 24489 9163 24547 9169
rect 24489 9160 24501 9163
rect 24452 9132 24501 9160
rect 24452 9120 24458 9132
rect 24489 9129 24501 9132
rect 24535 9160 24547 9163
rect 25958 9160 25964 9172
rect 24535 9132 25964 9160
rect 24535 9129 24547 9132
rect 24489 9123 24547 9129
rect 25958 9120 25964 9132
rect 26016 9120 26022 9172
rect 14645 9095 14703 9101
rect 14645 9092 14657 9095
rect 13372 9064 14657 9092
rect 14645 9061 14657 9064
rect 14691 9061 14703 9095
rect 14645 9055 14703 9061
rect 15378 9052 15384 9104
rect 15436 9092 15442 9104
rect 19978 9092 19984 9104
rect 15436 9064 16252 9092
rect 19939 9064 19984 9092
rect 15436 9052 15442 9064
rect 5534 8984 5540 9036
rect 5592 9024 5598 9036
rect 6086 9024 6092 9036
rect 5592 8996 6092 9024
rect 5592 8984 5598 8996
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 7190 8984 7196 9036
rect 7248 9024 7254 9036
rect 7377 9027 7435 9033
rect 7377 9024 7389 9027
rect 7248 8996 7389 9024
rect 7248 8984 7254 8996
rect 7377 8993 7389 8996
rect 7423 9024 7435 9027
rect 8846 9024 8852 9036
rect 7423 8996 8852 9024
rect 7423 8993 7435 8996
rect 7377 8987 7435 8993
rect 8846 8984 8852 8996
rect 8904 8984 8910 9036
rect 9858 9024 9864 9036
rect 9819 8996 9864 9024
rect 9858 8984 9864 8996
rect 9916 9024 9922 9036
rect 10321 9027 10379 9033
rect 10321 9024 10333 9027
rect 9916 8996 10333 9024
rect 9916 8984 9922 8996
rect 10321 8993 10333 8996
rect 10367 8993 10379 9027
rect 10870 9024 10876 9036
rect 10831 8996 10876 9024
rect 10321 8987 10379 8993
rect 10870 8984 10876 8996
rect 10928 8984 10934 9036
rect 11057 9027 11115 9033
rect 11057 8993 11069 9027
rect 11103 9024 11115 9027
rect 11606 9024 11612 9036
rect 11103 8996 11612 9024
rect 11103 8993 11115 8996
rect 11057 8987 11115 8993
rect 11606 8984 11612 8996
rect 11664 8984 11670 9036
rect 11790 9024 11796 9036
rect 11751 8996 11796 9024
rect 11790 8984 11796 8996
rect 11848 8984 11854 9036
rect 13170 9024 13176 9036
rect 13083 8996 13176 9024
rect 13170 8984 13176 8996
rect 13228 9024 13234 9036
rect 13722 9024 13728 9036
rect 13228 8996 13728 9024
rect 13228 8984 13234 8996
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 14826 8984 14832 9036
rect 14884 9024 14890 9036
rect 15470 9024 15476 9036
rect 14884 8996 15476 9024
rect 14884 8984 14890 8996
rect 15470 8984 15476 8996
rect 15528 8984 15534 9036
rect 15654 8984 15660 9036
rect 15712 9024 15718 9036
rect 16224 9033 16252 9064
rect 19978 9052 19984 9064
rect 20036 9052 20042 9104
rect 25498 9092 25504 9104
rect 25459 9064 25504 9092
rect 25498 9052 25504 9064
rect 25556 9052 25562 9104
rect 16025 9027 16083 9033
rect 16025 9024 16037 9027
rect 15712 8996 16037 9024
rect 15712 8984 15718 8996
rect 16025 8993 16037 8996
rect 16071 8993 16083 9027
rect 16025 8987 16083 8993
rect 16209 9027 16267 9033
rect 16209 8993 16221 9027
rect 16255 8993 16267 9027
rect 16209 8987 16267 8993
rect 18325 9027 18383 9033
rect 18325 8993 18337 9027
rect 18371 9024 18383 9027
rect 18414 9024 18420 9036
rect 18371 8996 18420 9024
rect 18371 8993 18383 8996
rect 18325 8987 18383 8993
rect 18414 8984 18420 8996
rect 18472 8984 18478 9036
rect 18598 9024 18604 9036
rect 18559 8996 18604 9024
rect 18598 8984 18604 8996
rect 18656 8984 18662 9036
rect 26142 9024 26148 9036
rect 26103 8996 26148 9024
rect 26142 8984 26148 8996
rect 26200 8984 26206 9036
rect 7098 8956 7104 8968
rect 7059 8928 7104 8956
rect 7098 8916 7104 8928
rect 7156 8916 7162 8968
rect 13078 8956 13084 8968
rect 13039 8928 13084 8956
rect 13078 8916 13084 8928
rect 13136 8956 13142 8968
rect 13354 8956 13360 8968
rect 13136 8928 13360 8956
rect 13136 8916 13142 8928
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 15194 8916 15200 8968
rect 15252 8956 15258 8968
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 15252 8928 15301 8956
rect 15252 8916 15258 8928
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 6270 8888 6276 8900
rect 6231 8860 6276 8888
rect 6270 8848 6276 8860
rect 6328 8848 6334 8900
rect 9125 8823 9183 8829
rect 9125 8789 9137 8823
rect 9171 8820 9183 8823
rect 9950 8820 9956 8832
rect 9171 8792 9956 8820
rect 9171 8789 9183 8792
rect 9125 8783 9183 8789
rect 9950 8780 9956 8792
rect 10008 8780 10014 8832
rect 12069 8823 12127 8829
rect 12069 8789 12081 8823
rect 12115 8820 12127 8823
rect 12342 8820 12348 8832
rect 12115 8792 12348 8820
rect 12115 8789 12127 8792
rect 12069 8783 12127 8789
rect 12342 8780 12348 8792
rect 12400 8780 12406 8832
rect 13354 8820 13360 8832
rect 13315 8792 13360 8820
rect 13354 8780 13360 8792
rect 13412 8780 13418 8832
rect 14366 8820 14372 8832
rect 14279 8792 14372 8820
rect 14366 8780 14372 8792
rect 14424 8820 14430 8832
rect 15194 8820 15200 8832
rect 14424 8792 15200 8820
rect 14424 8780 14430 8792
rect 15194 8780 15200 8792
rect 15252 8780 15258 8832
rect 16482 8820 16488 8832
rect 16443 8792 16488 8820
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 1104 8730 38548 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 38548 8730
rect 1104 8656 38548 8678
rect 6086 8616 6092 8628
rect 6047 8588 6092 8616
rect 6086 8576 6092 8588
rect 6144 8576 6150 8628
rect 7098 8576 7104 8628
rect 7156 8616 7162 8628
rect 7469 8619 7527 8625
rect 7469 8616 7481 8619
rect 7156 8588 7481 8616
rect 7156 8576 7162 8588
rect 7469 8585 7481 8588
rect 7515 8585 7527 8619
rect 7469 8579 7527 8585
rect 10597 8619 10655 8625
rect 10597 8585 10609 8619
rect 10643 8616 10655 8619
rect 11606 8616 11612 8628
rect 10643 8588 11612 8616
rect 10643 8585 10655 8588
rect 10597 8579 10655 8585
rect 11606 8576 11612 8588
rect 11664 8576 11670 8628
rect 12805 8619 12863 8625
rect 12805 8585 12817 8619
rect 12851 8616 12863 8619
rect 12894 8616 12900 8628
rect 12851 8588 12900 8616
rect 12851 8585 12863 8588
rect 12805 8579 12863 8585
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 13170 8616 13176 8628
rect 13131 8588 13176 8616
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 14274 8576 14280 8628
rect 14332 8616 14338 8628
rect 14921 8619 14979 8625
rect 14921 8616 14933 8619
rect 14332 8588 14933 8616
rect 14332 8576 14338 8588
rect 14921 8585 14933 8588
rect 14967 8585 14979 8619
rect 15378 8616 15384 8628
rect 15339 8588 15384 8616
rect 14921 8579 14979 8585
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15470 8576 15476 8628
rect 15528 8616 15534 8628
rect 15657 8619 15715 8625
rect 15657 8616 15669 8619
rect 15528 8588 15669 8616
rect 15528 8576 15534 8588
rect 15657 8585 15669 8588
rect 15703 8585 15715 8619
rect 18230 8616 18236 8628
rect 18191 8588 18236 8616
rect 15657 8579 15715 8585
rect 18230 8576 18236 8588
rect 18288 8576 18294 8628
rect 18322 8576 18328 8628
rect 18380 8616 18386 8628
rect 18509 8619 18567 8625
rect 18509 8616 18521 8619
rect 18380 8588 18521 8616
rect 18380 8576 18386 8588
rect 18509 8585 18521 8588
rect 18555 8585 18567 8619
rect 18509 8579 18567 8585
rect 18598 8576 18604 8628
rect 18656 8616 18662 8628
rect 18877 8619 18935 8625
rect 18877 8616 18889 8619
rect 18656 8588 18889 8616
rect 18656 8576 18662 8588
rect 18877 8585 18889 8588
rect 18923 8585 18935 8619
rect 18877 8579 18935 8585
rect 26053 8619 26111 8625
rect 26053 8585 26065 8619
rect 26099 8616 26111 8619
rect 26142 8616 26148 8628
rect 26099 8588 26148 8616
rect 26099 8585 26111 8588
rect 26053 8579 26111 8585
rect 26142 8576 26148 8588
rect 26200 8576 26206 8628
rect 7190 8548 7196 8560
rect 7151 8520 7196 8548
rect 7190 8508 7196 8520
rect 7248 8508 7254 8560
rect 8849 8551 8907 8557
rect 8849 8517 8861 8551
rect 8895 8548 8907 8551
rect 10965 8551 11023 8557
rect 8895 8520 9720 8548
rect 8895 8517 8907 8520
rect 8849 8511 8907 8517
rect 9692 8492 9720 8520
rect 10965 8517 10977 8551
rect 11011 8548 11023 8551
rect 11790 8548 11796 8560
rect 11011 8520 11796 8548
rect 11011 8517 11023 8520
rect 10965 8511 11023 8517
rect 11790 8508 11796 8520
rect 11848 8508 11854 8560
rect 16942 8548 16948 8560
rect 16592 8520 16948 8548
rect 7926 8440 7932 8492
rect 7984 8480 7990 8492
rect 8481 8483 8539 8489
rect 8481 8480 8493 8483
rect 7984 8452 8493 8480
rect 7984 8440 7990 8452
rect 8481 8449 8493 8452
rect 8527 8480 8539 8483
rect 8527 8452 9628 8480
rect 8527 8449 8539 8452
rect 8481 8443 8539 8449
rect 9600 8424 9628 8452
rect 9674 8440 9680 8492
rect 9732 8480 9738 8492
rect 9732 8452 9777 8480
rect 9732 8440 9738 8452
rect 10870 8440 10876 8492
rect 10928 8480 10934 8492
rect 11241 8483 11299 8489
rect 11241 8480 11253 8483
rect 10928 8452 11253 8480
rect 10928 8440 10934 8452
rect 11241 8449 11253 8452
rect 11287 8449 11299 8483
rect 11241 8443 11299 8449
rect 12894 8440 12900 8492
rect 12952 8480 12958 8492
rect 14185 8483 14243 8489
rect 12952 8452 14136 8480
rect 12952 8440 12958 8452
rect 9582 8412 9588 8424
rect 9543 8384 9588 8412
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 9950 8412 9956 8424
rect 9911 8384 9956 8412
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 10134 8412 10140 8424
rect 10095 8384 10140 8412
rect 10134 8372 10140 8384
rect 10192 8372 10198 8424
rect 13722 8412 13728 8424
rect 13683 8384 13728 8412
rect 13722 8372 13728 8384
rect 13780 8372 13786 8424
rect 14108 8421 14136 8452
rect 14185 8449 14197 8483
rect 14231 8480 14243 8483
rect 14826 8480 14832 8492
rect 14231 8452 14832 8480
rect 14231 8449 14243 8452
rect 14185 8443 14243 8449
rect 14093 8415 14151 8421
rect 14093 8381 14105 8415
rect 14139 8381 14151 8415
rect 14093 8375 14151 8381
rect 1486 8304 1492 8356
rect 1544 8344 1550 8356
rect 8941 8347 8999 8353
rect 8941 8344 8953 8347
rect 1544 8316 8953 8344
rect 1544 8304 1550 8316
rect 8941 8313 8953 8316
rect 8987 8313 8999 8347
rect 9968 8344 9996 8372
rect 11054 8344 11060 8356
rect 9968 8316 11060 8344
rect 8941 8307 8999 8313
rect 11054 8304 11060 8316
rect 11112 8304 11118 8356
rect 13262 8344 13268 8356
rect 13223 8316 13268 8344
rect 13262 8304 13268 8316
rect 13320 8304 13326 8356
rect 13630 8304 13636 8356
rect 13688 8344 13694 8356
rect 14200 8344 14228 8443
rect 14826 8440 14832 8452
rect 14884 8440 14890 8492
rect 15746 8440 15752 8492
rect 15804 8480 15810 8492
rect 15933 8483 15991 8489
rect 15933 8480 15945 8483
rect 15804 8452 15945 8480
rect 15804 8440 15810 8452
rect 15933 8449 15945 8452
rect 15979 8449 15991 8483
rect 15933 8443 15991 8449
rect 16298 8440 16304 8492
rect 16356 8480 16362 8492
rect 16393 8483 16451 8489
rect 16393 8480 16405 8483
rect 16356 8452 16405 8480
rect 16356 8440 16362 8452
rect 16393 8449 16405 8452
rect 16439 8449 16451 8483
rect 16393 8443 16451 8449
rect 16592 8421 16620 8520
rect 16942 8508 16948 8520
rect 17000 8508 17006 8560
rect 17865 8551 17923 8557
rect 17865 8517 17877 8551
rect 17911 8548 17923 8551
rect 18414 8548 18420 8560
rect 17911 8520 18420 8548
rect 17911 8517 17923 8520
rect 17865 8511 17923 8517
rect 18414 8508 18420 8520
rect 18472 8508 18478 8560
rect 16850 8480 16856 8492
rect 16811 8452 16856 8480
rect 16850 8440 16856 8452
rect 16908 8480 16914 8492
rect 17405 8483 17463 8489
rect 17405 8480 17417 8483
rect 16908 8452 17417 8480
rect 16908 8440 16914 8452
rect 17405 8449 17417 8452
rect 17451 8449 17463 8483
rect 17405 8443 17463 8449
rect 16577 8415 16635 8421
rect 16577 8381 16589 8415
rect 16623 8381 16635 8415
rect 16577 8375 16635 8381
rect 14642 8344 14648 8356
rect 13688 8316 14228 8344
rect 14603 8316 14648 8344
rect 13688 8304 13694 8316
rect 14642 8304 14648 8316
rect 14700 8304 14706 8356
rect 16592 8344 16620 8375
rect 16666 8372 16672 8424
rect 16724 8412 16730 8424
rect 16945 8415 17003 8421
rect 16945 8412 16957 8415
rect 16724 8384 16957 8412
rect 16724 8372 16730 8384
rect 16945 8381 16957 8384
rect 16991 8381 17003 8415
rect 16945 8375 17003 8381
rect 18049 8415 18107 8421
rect 18049 8381 18061 8415
rect 18095 8412 18107 8415
rect 18322 8412 18328 8424
rect 18095 8384 18328 8412
rect 18095 8381 18107 8384
rect 18049 8375 18107 8381
rect 18322 8372 18328 8384
rect 18380 8372 18386 8424
rect 16500 8316 16620 8344
rect 9950 8236 9956 8288
rect 10008 8276 10014 8288
rect 12161 8279 12219 8285
rect 12161 8276 12173 8279
rect 10008 8248 12173 8276
rect 10008 8236 10014 8248
rect 12161 8245 12173 8248
rect 12207 8276 12219 8279
rect 13078 8276 13084 8288
rect 12207 8248 13084 8276
rect 12207 8245 12219 8248
rect 12161 8239 12219 8245
rect 13078 8236 13084 8248
rect 13136 8236 13142 8288
rect 16022 8236 16028 8288
rect 16080 8276 16086 8288
rect 16500 8276 16528 8316
rect 16080 8248 16528 8276
rect 16080 8236 16086 8248
rect 1104 8186 38548 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 38548 8186
rect 1104 8112 38548 8134
rect 9030 8072 9036 8084
rect 8991 8044 9036 8072
rect 9030 8032 9036 8044
rect 9088 8032 9094 8084
rect 11054 8072 11060 8084
rect 11015 8044 11060 8072
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 13541 8075 13599 8081
rect 13541 8041 13553 8075
rect 13587 8072 13599 8075
rect 13630 8072 13636 8084
rect 13587 8044 13636 8072
rect 13587 8041 13599 8044
rect 13541 8035 13599 8041
rect 13354 8004 13360 8016
rect 12636 7976 13360 8004
rect 12636 7948 12664 7976
rect 13354 7964 13360 7976
rect 13412 7964 13418 8016
rect 12618 7936 12624 7948
rect 12531 7908 12624 7936
rect 12618 7896 12624 7908
rect 12676 7896 12682 7948
rect 12710 7896 12716 7948
rect 12768 7936 12774 7948
rect 12989 7939 13047 7945
rect 12989 7936 13001 7939
rect 12768 7908 13001 7936
rect 12768 7896 12774 7908
rect 12989 7905 13001 7908
rect 13035 7905 13047 7939
rect 12989 7899 13047 7905
rect 13081 7939 13139 7945
rect 13081 7905 13093 7939
rect 13127 7936 13139 7939
rect 13556 7936 13584 8035
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 13814 8072 13820 8084
rect 13775 8044 13820 8072
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 15102 8072 15108 8084
rect 15063 8044 15108 8072
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 16666 8072 16672 8084
rect 16627 8044 16672 8072
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 20257 8075 20315 8081
rect 20257 8041 20269 8075
rect 20303 8072 20315 8075
rect 20346 8072 20352 8084
rect 20303 8044 20352 8072
rect 20303 8041 20315 8044
rect 20257 8035 20315 8041
rect 20346 8032 20352 8044
rect 20404 8032 20410 8084
rect 19702 7964 19708 8016
rect 19760 8004 19766 8016
rect 21082 8004 21088 8016
rect 19760 7976 21088 8004
rect 19760 7964 19766 7976
rect 21082 7964 21088 7976
rect 21140 7964 21146 8016
rect 13127 7908 13584 7936
rect 13127 7905 13139 7908
rect 13081 7899 13139 7905
rect 9674 7828 9680 7880
rect 9732 7868 9738 7880
rect 9732 7840 9777 7868
rect 9732 7828 9738 7840
rect 9858 7828 9864 7880
rect 9916 7868 9922 7880
rect 9953 7871 10011 7877
rect 9953 7868 9965 7871
rect 9916 7840 9965 7868
rect 9916 7828 9922 7840
rect 9953 7837 9965 7840
rect 9999 7837 10011 7871
rect 9953 7831 10011 7837
rect 11330 7828 11336 7880
rect 11388 7868 11394 7880
rect 12161 7871 12219 7877
rect 12161 7868 12173 7871
rect 11388 7840 12173 7868
rect 11388 7828 11394 7840
rect 12161 7837 12173 7840
rect 12207 7837 12219 7871
rect 12161 7831 12219 7837
rect 12802 7828 12808 7880
rect 12860 7868 12866 7880
rect 13096 7868 13124 7899
rect 15194 7896 15200 7948
rect 15252 7936 15258 7948
rect 15565 7939 15623 7945
rect 15565 7936 15577 7939
rect 15252 7908 15577 7936
rect 15252 7896 15258 7908
rect 15565 7905 15577 7908
rect 15611 7936 15623 7939
rect 16298 7936 16304 7948
rect 15611 7908 16304 7936
rect 15611 7905 15623 7908
rect 15565 7899 15623 7905
rect 16298 7896 16304 7908
rect 16356 7896 16362 7948
rect 16574 7896 16580 7948
rect 16632 7936 16638 7948
rect 17862 7936 17868 7948
rect 16632 7908 17868 7936
rect 16632 7896 16638 7908
rect 17862 7896 17868 7908
rect 17920 7936 17926 7948
rect 18049 7939 18107 7945
rect 18049 7936 18061 7939
rect 17920 7908 18061 7936
rect 17920 7896 17926 7908
rect 18049 7905 18061 7908
rect 18095 7905 18107 7939
rect 18049 7899 18107 7905
rect 21174 7896 21180 7948
rect 21232 7936 21238 7948
rect 21232 7908 21496 7936
rect 21232 7896 21238 7908
rect 12860 7840 13124 7868
rect 12860 7828 12866 7840
rect 15010 7828 15016 7880
rect 15068 7868 15074 7880
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 15068 7840 15301 7868
rect 15068 7828 15074 7840
rect 15289 7837 15301 7840
rect 15335 7868 15347 7871
rect 17773 7871 17831 7877
rect 17773 7868 17785 7871
rect 15335 7840 17785 7868
rect 15335 7837 15347 7840
rect 15289 7831 15347 7837
rect 17773 7837 17785 7840
rect 17819 7868 17831 7871
rect 18414 7868 18420 7880
rect 17819 7840 18420 7868
rect 17819 7837 17831 7840
rect 17773 7831 17831 7837
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 20346 7828 20352 7880
rect 20404 7868 20410 7880
rect 21361 7871 21419 7877
rect 21361 7868 21373 7871
rect 20404 7840 21373 7868
rect 20404 7828 20410 7840
rect 21361 7837 21373 7840
rect 21407 7837 21419 7871
rect 21468 7868 21496 7908
rect 21542 7896 21548 7948
rect 21600 7936 21606 7948
rect 21910 7936 21916 7948
rect 21600 7908 21645 7936
rect 21871 7908 21916 7936
rect 21600 7896 21606 7908
rect 21910 7896 21916 7908
rect 21968 7896 21974 7948
rect 23106 7936 23112 7948
rect 23067 7908 23112 7936
rect 23106 7896 23112 7908
rect 23164 7896 23170 7948
rect 21821 7871 21879 7877
rect 21821 7868 21833 7871
rect 21468 7840 21833 7868
rect 21361 7831 21419 7837
rect 21821 7837 21833 7840
rect 21867 7837 21879 7871
rect 21821 7831 21879 7837
rect 19334 7732 19340 7744
rect 19295 7704 19340 7732
rect 19334 7692 19340 7704
rect 19392 7692 19398 7744
rect 21174 7732 21180 7744
rect 21135 7704 21180 7732
rect 21174 7692 21180 7704
rect 21232 7692 21238 7744
rect 22925 7735 22983 7741
rect 22925 7701 22937 7735
rect 22971 7732 22983 7735
rect 23474 7732 23480 7744
rect 22971 7704 23480 7732
rect 22971 7701 22983 7704
rect 22925 7695 22983 7701
rect 23474 7692 23480 7704
rect 23532 7692 23538 7744
rect 1104 7642 38548 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 38548 7642
rect 1104 7568 38548 7590
rect 8478 7528 8484 7540
rect 8439 7500 8484 7528
rect 8478 7488 8484 7500
rect 8536 7488 8542 7540
rect 9493 7531 9551 7537
rect 9493 7497 9505 7531
rect 9539 7528 9551 7531
rect 9858 7528 9864 7540
rect 9539 7500 9864 7528
rect 9539 7497 9551 7500
rect 9493 7491 9551 7497
rect 9858 7488 9864 7500
rect 9916 7488 9922 7540
rect 10042 7488 10048 7540
rect 10100 7528 10106 7540
rect 10137 7531 10195 7537
rect 10137 7528 10149 7531
rect 10100 7500 10149 7528
rect 10100 7488 10106 7500
rect 10137 7497 10149 7500
rect 10183 7528 10195 7531
rect 11885 7531 11943 7537
rect 10183 7500 11100 7528
rect 10183 7497 10195 7500
rect 10137 7491 10195 7497
rect 10870 7392 10876 7404
rect 10831 7364 10876 7392
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 11072 7392 11100 7500
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 12618 7528 12624 7540
rect 11931 7500 12624 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 15010 7528 15016 7540
rect 14971 7500 15016 7528
rect 15010 7488 15016 7500
rect 15068 7488 15074 7540
rect 15381 7531 15439 7537
rect 15381 7497 15393 7531
rect 15427 7528 15439 7531
rect 16298 7528 16304 7540
rect 15427 7500 16304 7528
rect 15427 7497 15439 7500
rect 15381 7491 15439 7497
rect 16298 7488 16304 7500
rect 16356 7488 16362 7540
rect 17862 7528 17868 7540
rect 17823 7500 17868 7528
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 19426 7488 19432 7540
rect 19484 7528 19490 7540
rect 20073 7531 20131 7537
rect 20073 7528 20085 7531
rect 19484 7500 20085 7528
rect 19484 7488 19490 7500
rect 20073 7497 20085 7500
rect 20119 7528 20131 7531
rect 21542 7528 21548 7540
rect 20119 7500 21548 7528
rect 20119 7497 20131 7500
rect 20073 7491 20131 7497
rect 21542 7488 21548 7500
rect 21600 7488 21606 7540
rect 21729 7531 21787 7537
rect 21729 7497 21741 7531
rect 21775 7528 21787 7531
rect 21910 7528 21916 7540
rect 21775 7500 21916 7528
rect 21775 7497 21787 7500
rect 21729 7491 21787 7497
rect 21910 7488 21916 7500
rect 21968 7488 21974 7540
rect 23017 7531 23075 7537
rect 23017 7497 23029 7531
rect 23063 7528 23075 7531
rect 23106 7528 23112 7540
rect 23063 7500 23112 7528
rect 23063 7497 23075 7500
rect 23017 7491 23075 7497
rect 23106 7488 23112 7500
rect 23164 7488 23170 7540
rect 11146 7420 11152 7472
rect 11204 7460 11210 7472
rect 12161 7463 12219 7469
rect 12161 7460 12173 7463
rect 11204 7432 12173 7460
rect 11204 7420 11210 7432
rect 12161 7429 12173 7432
rect 12207 7460 12219 7463
rect 12710 7460 12716 7472
rect 12207 7432 12716 7460
rect 12207 7429 12219 7432
rect 12161 7423 12219 7429
rect 12710 7420 12716 7432
rect 12768 7420 12774 7472
rect 16022 7460 16028 7472
rect 15983 7432 16028 7460
rect 16022 7420 16028 7432
rect 16080 7420 16086 7472
rect 11238 7392 11244 7404
rect 11072 7364 11244 7392
rect 11238 7352 11244 7364
rect 11296 7352 11302 7404
rect 13173 7395 13231 7401
rect 13173 7361 13185 7395
rect 13219 7392 13231 7395
rect 13262 7392 13268 7404
rect 13219 7364 13268 7392
rect 13219 7361 13231 7364
rect 13173 7355 13231 7361
rect 13262 7352 13268 7364
rect 13320 7352 13326 7404
rect 20346 7352 20352 7404
rect 20404 7392 20410 7404
rect 20441 7395 20499 7401
rect 20441 7392 20453 7395
rect 20404 7364 20453 7392
rect 20404 7352 20410 7364
rect 20441 7361 20453 7364
rect 20487 7392 20499 7395
rect 22097 7395 22155 7401
rect 22097 7392 22109 7395
rect 20487 7364 22109 7392
rect 20487 7361 20499 7364
rect 20441 7355 20499 7361
rect 22097 7361 22109 7364
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 8478 7284 8484 7336
rect 8536 7324 8542 7336
rect 8849 7327 8907 7333
rect 8849 7324 8861 7327
rect 8536 7296 8861 7324
rect 8536 7284 8542 7296
rect 8849 7293 8861 7296
rect 8895 7293 8907 7327
rect 10962 7324 10968 7336
rect 10923 7296 10968 7324
rect 8849 7287 8907 7293
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 11330 7324 11336 7336
rect 11291 7296 11336 7324
rect 11330 7284 11336 7296
rect 11388 7284 11394 7336
rect 12526 7284 12532 7336
rect 12584 7324 12590 7336
rect 12897 7327 12955 7333
rect 12897 7324 12909 7327
rect 12584 7296 12909 7324
rect 12584 7284 12590 7296
rect 12897 7293 12909 7296
rect 12943 7293 12955 7327
rect 12897 7287 12955 7293
rect 18325 7327 18383 7333
rect 18325 7293 18337 7327
rect 18371 7324 18383 7327
rect 18414 7324 18420 7336
rect 18371 7296 18420 7324
rect 18371 7293 18383 7296
rect 18325 7287 18383 7293
rect 18414 7284 18420 7296
rect 18472 7324 18478 7336
rect 20165 7327 20223 7333
rect 20165 7324 20177 7327
rect 18472 7296 20177 7324
rect 18472 7284 18478 7296
rect 20165 7293 20177 7296
rect 20211 7324 20223 7327
rect 20254 7324 20260 7336
rect 20211 7296 20260 7324
rect 20211 7293 20223 7296
rect 20165 7287 20223 7293
rect 20254 7284 20260 7296
rect 20312 7284 20318 7336
rect 9861 7259 9919 7265
rect 9861 7225 9873 7259
rect 9907 7256 9919 7259
rect 10980 7256 11008 7284
rect 9907 7228 11008 7256
rect 9907 7225 9919 7228
rect 9861 7219 9919 7225
rect 8662 7188 8668 7200
rect 8623 7160 8668 7188
rect 8662 7148 8668 7160
rect 8720 7148 8726 7200
rect 10226 7148 10232 7200
rect 10284 7188 10290 7200
rect 10413 7191 10471 7197
rect 10413 7188 10425 7191
rect 10284 7160 10425 7188
rect 10284 7148 10290 7160
rect 10413 7157 10425 7160
rect 10459 7157 10471 7191
rect 10413 7151 10471 7157
rect 10962 7148 10968 7200
rect 11020 7188 11026 7200
rect 11348 7188 11376 7284
rect 12713 7259 12771 7265
rect 12713 7225 12725 7259
rect 12759 7256 12771 7259
rect 12802 7256 12808 7268
rect 12759 7228 12808 7256
rect 12759 7225 12771 7228
rect 12713 7219 12771 7225
rect 12802 7216 12808 7228
rect 12860 7216 12866 7268
rect 11020 7160 11376 7188
rect 11020 7148 11026 7160
rect 13630 7148 13636 7200
rect 13688 7188 13694 7200
rect 14277 7191 14335 7197
rect 14277 7188 14289 7191
rect 13688 7160 14289 7188
rect 13688 7148 13694 7160
rect 14277 7157 14289 7160
rect 14323 7157 14335 7191
rect 14277 7151 14335 7157
rect 1104 7098 38548 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 38548 7098
rect 1104 7024 38548 7046
rect 10413 6987 10471 6993
rect 10413 6953 10425 6987
rect 10459 6984 10471 6987
rect 10870 6984 10876 6996
rect 10459 6956 10876 6984
rect 10459 6953 10471 6956
rect 10413 6947 10471 6953
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 12710 6944 12716 6996
rect 12768 6984 12774 6996
rect 12989 6987 13047 6993
rect 12989 6984 13001 6987
rect 12768 6956 13001 6984
rect 12768 6944 12774 6956
rect 12989 6953 13001 6956
rect 13035 6984 13047 6987
rect 13262 6984 13268 6996
rect 13035 6956 13268 6984
rect 13035 6953 13047 6956
rect 12989 6947 13047 6953
rect 13262 6944 13268 6956
rect 13320 6944 13326 6996
rect 20257 6987 20315 6993
rect 20257 6953 20269 6987
rect 20303 6984 20315 6987
rect 20346 6984 20352 6996
rect 20303 6956 20352 6984
rect 20303 6953 20315 6956
rect 20257 6947 20315 6953
rect 20346 6944 20352 6956
rect 20404 6944 20410 6996
rect 21082 6984 21088 6996
rect 21043 6956 21088 6984
rect 21082 6944 21088 6956
rect 21140 6944 21146 6996
rect 21545 6987 21603 6993
rect 21545 6953 21557 6987
rect 21591 6984 21603 6987
rect 21910 6984 21916 6996
rect 21591 6956 21916 6984
rect 21591 6953 21603 6956
rect 21545 6947 21603 6953
rect 21910 6944 21916 6956
rect 21968 6944 21974 6996
rect 13280 6916 13308 6944
rect 13280 6888 13860 6916
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6848 9551 6851
rect 9674 6848 9680 6860
rect 9539 6820 9680 6848
rect 9539 6817 9551 6820
rect 9493 6811 9551 6817
rect 9674 6808 9680 6820
rect 9732 6808 9738 6860
rect 10045 6851 10103 6857
rect 10045 6817 10057 6851
rect 10091 6848 10103 6851
rect 10091 6820 10824 6848
rect 10091 6817 10103 6820
rect 10045 6811 10103 6817
rect 9692 6780 9720 6808
rect 10796 6789 10824 6820
rect 11054 6808 11060 6860
rect 11112 6848 11118 6860
rect 11112 6820 11928 6848
rect 11112 6808 11118 6820
rect 10505 6783 10563 6789
rect 10505 6780 10517 6783
rect 9692 6752 10517 6780
rect 10505 6749 10517 6752
rect 10551 6749 10563 6783
rect 10505 6743 10563 6749
rect 10781 6783 10839 6789
rect 10781 6749 10793 6783
rect 10827 6780 10839 6783
rect 10962 6780 10968 6792
rect 10827 6752 10968 6780
rect 10827 6749 10839 6752
rect 10781 6743 10839 6749
rect 10962 6740 10968 6752
rect 11020 6740 11026 6792
rect 11900 6789 11928 6820
rect 13630 6808 13636 6860
rect 13688 6848 13694 6860
rect 13725 6851 13783 6857
rect 13725 6848 13737 6851
rect 13688 6820 13737 6848
rect 13688 6808 13694 6820
rect 13725 6817 13737 6820
rect 13771 6817 13783 6851
rect 13832 6848 13860 6888
rect 17862 6876 17868 6928
rect 17920 6916 17926 6928
rect 18874 6916 18880 6928
rect 17920 6888 18880 6916
rect 17920 6876 17926 6888
rect 18874 6876 18880 6888
rect 18932 6916 18938 6928
rect 18932 6888 19380 6916
rect 18932 6876 18938 6888
rect 14093 6851 14151 6857
rect 14093 6848 14105 6851
rect 13832 6820 14105 6848
rect 13725 6811 13783 6817
rect 14093 6817 14105 6820
rect 14139 6817 14151 6851
rect 14093 6811 14151 6817
rect 16761 6851 16819 6857
rect 16761 6817 16773 6851
rect 16807 6848 16819 6851
rect 16850 6848 16856 6860
rect 16807 6820 16856 6848
rect 16807 6817 16819 6820
rect 16761 6811 16819 6817
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 16942 6808 16948 6860
rect 17000 6848 17006 6860
rect 17129 6851 17187 6857
rect 17129 6848 17141 6851
rect 17000 6820 17141 6848
rect 17000 6808 17006 6820
rect 17129 6817 17141 6820
rect 17175 6817 17187 6851
rect 17129 6811 17187 6817
rect 17218 6808 17224 6860
rect 17276 6848 17282 6860
rect 19153 6851 19211 6857
rect 17276 6820 17321 6848
rect 17276 6808 17282 6820
rect 19153 6817 19165 6851
rect 19199 6848 19211 6851
rect 19242 6848 19248 6860
rect 19199 6820 19248 6848
rect 19199 6817 19211 6820
rect 19153 6811 19211 6817
rect 19242 6808 19248 6820
rect 19300 6808 19306 6860
rect 19352 6848 19380 6888
rect 19521 6851 19579 6857
rect 19521 6848 19533 6851
rect 19352 6820 19533 6848
rect 19521 6817 19533 6820
rect 19567 6817 19579 6851
rect 19521 6811 19579 6817
rect 27154 6808 27160 6860
rect 27212 6848 27218 6860
rect 27341 6851 27399 6857
rect 27341 6848 27353 6851
rect 27212 6820 27353 6848
rect 27212 6808 27218 6820
rect 27341 6817 27353 6820
rect 27387 6817 27399 6851
rect 28718 6848 28724 6860
rect 28679 6820 28724 6848
rect 27341 6811 27399 6817
rect 28718 6808 28724 6820
rect 28776 6808 28782 6860
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6749 11943 6783
rect 11885 6743 11943 6749
rect 12434 6740 12440 6792
rect 12492 6780 12498 6792
rect 13081 6783 13139 6789
rect 13081 6780 13093 6783
rect 12492 6752 13093 6780
rect 12492 6740 12498 6752
rect 13081 6749 13093 6752
rect 13127 6749 13139 6783
rect 13814 6780 13820 6792
rect 13775 6752 13820 6780
rect 13081 6743 13139 6749
rect 13814 6740 13820 6752
rect 13872 6740 13878 6792
rect 13998 6780 14004 6792
rect 13959 6752 14004 6780
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 16114 6780 16120 6792
rect 16075 6752 16120 6780
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 16666 6780 16672 6792
rect 16627 6752 16672 6780
rect 16666 6740 16672 6752
rect 16724 6740 16730 6792
rect 19058 6780 19064 6792
rect 19019 6752 19064 6780
rect 19058 6740 19064 6752
rect 19116 6740 19122 6792
rect 19429 6783 19487 6789
rect 19429 6749 19441 6783
rect 19475 6780 19487 6783
rect 19886 6780 19892 6792
rect 19475 6752 19892 6780
rect 19475 6749 19487 6752
rect 19429 6743 19487 6749
rect 12342 6672 12348 6724
rect 12400 6712 12406 6724
rect 14921 6715 14979 6721
rect 14921 6712 14933 6715
rect 12400 6684 14933 6712
rect 12400 6672 12406 6684
rect 14921 6681 14933 6684
rect 14967 6712 14979 6715
rect 15102 6712 15108 6724
rect 14967 6684 15108 6712
rect 14967 6681 14979 6684
rect 14921 6675 14979 6681
rect 15102 6672 15108 6684
rect 15160 6672 15166 6724
rect 18506 6672 18512 6724
rect 18564 6712 18570 6724
rect 19444 6712 19472 6743
rect 19886 6740 19892 6752
rect 19944 6740 19950 6792
rect 22186 6780 22192 6792
rect 22147 6752 22192 6780
rect 22186 6740 22192 6752
rect 22244 6740 22250 6792
rect 22462 6780 22468 6792
rect 22423 6752 22468 6780
rect 22462 6740 22468 6752
rect 22520 6740 22526 6792
rect 23566 6780 23572 6792
rect 23527 6752 23572 6780
rect 23566 6740 23572 6752
rect 23624 6740 23630 6792
rect 27065 6783 27123 6789
rect 27065 6749 27077 6783
rect 27111 6780 27123 6783
rect 27246 6780 27252 6792
rect 27111 6752 27252 6780
rect 27111 6749 27123 6752
rect 27065 6743 27123 6749
rect 27246 6740 27252 6752
rect 27304 6740 27310 6792
rect 18564 6684 19472 6712
rect 18564 6672 18570 6684
rect 12526 6644 12532 6656
rect 12487 6616 12532 6644
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 14550 6644 14556 6656
rect 14511 6616 14556 6644
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 18782 6644 18788 6656
rect 18743 6616 18788 6644
rect 18782 6604 18788 6616
rect 18840 6604 18846 6656
rect 1104 6554 38548 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 38548 6554
rect 1104 6480 38548 6502
rect 9674 6400 9680 6452
rect 9732 6440 9738 6452
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 9732 6412 10057 6440
rect 9732 6400 9738 6412
rect 10045 6409 10057 6412
rect 10091 6409 10103 6443
rect 10045 6403 10103 6409
rect 10597 6443 10655 6449
rect 10597 6409 10609 6443
rect 10643 6440 10655 6443
rect 10962 6440 10968 6452
rect 10643 6412 10968 6440
rect 10643 6409 10655 6412
rect 10597 6403 10655 6409
rect 7653 6375 7711 6381
rect 7653 6341 7665 6375
rect 7699 6372 7711 6375
rect 8202 6372 8208 6384
rect 7699 6344 8208 6372
rect 7699 6341 7711 6344
rect 7653 6335 7711 6341
rect 8202 6332 8208 6344
rect 8260 6332 8266 6384
rect 10060 6372 10088 6403
rect 10962 6400 10968 6412
rect 11020 6400 11026 6452
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6440 12311 6443
rect 12710 6440 12716 6452
rect 12299 6412 12716 6440
rect 12299 6409 12311 6412
rect 12253 6403 12311 6409
rect 12710 6400 12716 6412
rect 12768 6400 12774 6452
rect 12805 6443 12863 6449
rect 12805 6409 12817 6443
rect 12851 6440 12863 6443
rect 13630 6440 13636 6452
rect 12851 6412 13636 6440
rect 12851 6409 12863 6412
rect 12805 6403 12863 6409
rect 13630 6400 13636 6412
rect 13688 6400 13694 6452
rect 13906 6440 13912 6452
rect 13867 6412 13912 6440
rect 13906 6400 13912 6412
rect 13964 6400 13970 6452
rect 16577 6443 16635 6449
rect 16577 6409 16589 6443
rect 16623 6440 16635 6443
rect 17218 6440 17224 6452
rect 16623 6412 17224 6440
rect 16623 6409 16635 6412
rect 16577 6403 16635 6409
rect 17218 6400 17224 6412
rect 17276 6400 17282 6452
rect 17865 6443 17923 6449
rect 17865 6409 17877 6443
rect 17911 6440 17923 6443
rect 19242 6440 19248 6452
rect 17911 6412 19248 6440
rect 17911 6409 17923 6412
rect 17865 6403 17923 6409
rect 19242 6400 19248 6412
rect 19300 6400 19306 6452
rect 20346 6400 20352 6452
rect 20404 6440 20410 6452
rect 20441 6443 20499 6449
rect 20441 6440 20453 6443
rect 20404 6412 20453 6440
rect 20404 6400 20410 6412
rect 20441 6409 20453 6412
rect 20487 6409 20499 6443
rect 20441 6403 20499 6409
rect 22186 6400 22192 6452
rect 22244 6440 22250 6452
rect 22557 6443 22615 6449
rect 22557 6440 22569 6443
rect 22244 6412 22569 6440
rect 22244 6400 22250 6412
rect 22557 6409 22569 6412
rect 22603 6440 22615 6443
rect 22646 6440 22652 6452
rect 22603 6412 22652 6440
rect 22603 6409 22615 6412
rect 22557 6403 22615 6409
rect 22646 6400 22652 6412
rect 22704 6400 22710 6452
rect 27246 6400 27252 6452
rect 27304 6440 27310 6452
rect 27433 6443 27491 6449
rect 27433 6440 27445 6443
rect 27304 6412 27445 6440
rect 27304 6400 27310 6412
rect 27433 6409 27445 6412
rect 27479 6409 27491 6443
rect 27433 6403 27491 6409
rect 11241 6375 11299 6381
rect 11241 6372 11253 6375
rect 10060 6344 11253 6372
rect 11241 6341 11253 6344
rect 11287 6372 11299 6375
rect 12526 6372 12532 6384
rect 11287 6344 12532 6372
rect 11287 6341 11299 6344
rect 11241 6335 11299 6341
rect 12526 6332 12532 6344
rect 12584 6332 12590 6384
rect 13924 6304 13952 6400
rect 15841 6375 15899 6381
rect 15841 6341 15853 6375
rect 15887 6372 15899 6375
rect 15930 6372 15936 6384
rect 15887 6344 15936 6372
rect 15887 6341 15899 6344
rect 15841 6335 15899 6341
rect 15930 6332 15936 6344
rect 15988 6372 15994 6384
rect 16666 6372 16672 6384
rect 15988 6344 16672 6372
rect 15988 6332 15994 6344
rect 16666 6332 16672 6344
rect 16724 6332 16730 6384
rect 18506 6372 18512 6384
rect 18467 6344 18512 6372
rect 18506 6332 18512 6344
rect 18564 6332 18570 6384
rect 15013 6307 15071 6313
rect 15013 6304 15025 6307
rect 13924 6276 15025 6304
rect 15013 6273 15025 6276
rect 15059 6273 15071 6307
rect 15013 6267 15071 6273
rect 16209 6307 16267 6313
rect 16209 6273 16221 6307
rect 16255 6304 16267 6307
rect 16850 6304 16856 6316
rect 16255 6276 16856 6304
rect 16255 6273 16267 6276
rect 16209 6267 16267 6273
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 18969 6307 19027 6313
rect 18969 6273 18981 6307
rect 19015 6304 19027 6307
rect 19015 6276 19380 6304
rect 19015 6273 19027 6276
rect 18969 6267 19027 6273
rect 19352 6248 19380 6276
rect 7837 6239 7895 6245
rect 7837 6205 7849 6239
rect 7883 6236 7895 6239
rect 8205 6239 8263 6245
rect 8205 6236 8217 6239
rect 7883 6208 8217 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 8205 6205 8217 6208
rect 8251 6236 8263 6239
rect 8662 6236 8668 6248
rect 8251 6208 8668 6236
rect 8251 6205 8263 6208
rect 8205 6199 8263 6205
rect 8662 6196 8668 6208
rect 8720 6236 8726 6248
rect 10229 6239 10287 6245
rect 10229 6236 10241 6239
rect 8720 6208 10241 6236
rect 8720 6196 8726 6208
rect 10229 6205 10241 6208
rect 10275 6236 10287 6239
rect 10873 6239 10931 6245
rect 10873 6236 10885 6239
rect 10275 6208 10885 6236
rect 10275 6205 10287 6208
rect 10229 6199 10287 6205
rect 10873 6205 10885 6208
rect 10919 6205 10931 6239
rect 10873 6199 10931 6205
rect 13541 6239 13599 6245
rect 13541 6205 13553 6239
rect 13587 6236 13599 6239
rect 13814 6236 13820 6248
rect 13587 6208 13820 6236
rect 13587 6205 13599 6208
rect 13541 6199 13599 6205
rect 13814 6196 13820 6208
rect 13872 6236 13878 6248
rect 14550 6236 14556 6248
rect 13872 6208 14556 6236
rect 13872 6196 13878 6208
rect 14550 6196 14556 6208
rect 14608 6196 14614 6248
rect 14734 6236 14740 6248
rect 14695 6208 14740 6236
rect 14734 6196 14740 6208
rect 14792 6196 14798 6248
rect 15102 6236 15108 6248
rect 15063 6208 15108 6236
rect 15102 6196 15108 6208
rect 15160 6196 15166 6248
rect 19061 6239 19119 6245
rect 19061 6205 19073 6239
rect 19107 6236 19119 6239
rect 19150 6236 19156 6248
rect 19107 6208 19156 6236
rect 19107 6205 19119 6208
rect 19061 6199 19119 6205
rect 19150 6196 19156 6208
rect 19208 6196 19214 6248
rect 19334 6236 19340 6248
rect 19295 6208 19340 6236
rect 19334 6196 19340 6208
rect 19392 6196 19398 6248
rect 13173 6171 13231 6177
rect 13173 6137 13185 6171
rect 13219 6168 13231 6171
rect 13998 6168 14004 6180
rect 13219 6140 14004 6168
rect 13219 6137 13231 6140
rect 13173 6131 13231 6137
rect 13998 6128 14004 6140
rect 14056 6128 14062 6180
rect 22281 6171 22339 6177
rect 22281 6137 22293 6171
rect 22327 6168 22339 6171
rect 22462 6168 22468 6180
rect 22327 6140 22468 6168
rect 22327 6137 22339 6140
rect 22281 6131 22339 6137
rect 22462 6128 22468 6140
rect 22520 6168 22526 6180
rect 23014 6168 23020 6180
rect 22520 6140 23020 6168
rect 22520 6128 22526 6140
rect 23014 6128 23020 6140
rect 23072 6128 23078 6180
rect 14366 6100 14372 6112
rect 14327 6072 14372 6100
rect 14366 6060 14372 6072
rect 14424 6060 14430 6112
rect 16942 6100 16948 6112
rect 16903 6072 16948 6100
rect 16942 6060 16948 6072
rect 17000 6060 17006 6112
rect 27062 6100 27068 6112
rect 27023 6072 27068 6100
rect 27062 6060 27068 6072
rect 27120 6060 27126 6112
rect 1104 6010 38548 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 38548 6010
rect 1104 5936 38548 5958
rect 14277 5899 14335 5905
rect 14277 5865 14289 5899
rect 14323 5896 14335 5899
rect 14734 5896 14740 5908
rect 14323 5868 14740 5896
rect 14323 5865 14335 5868
rect 14277 5859 14335 5865
rect 14734 5856 14740 5868
rect 14792 5856 14798 5908
rect 16942 5856 16948 5908
rect 17000 5896 17006 5908
rect 17037 5899 17095 5905
rect 17037 5896 17049 5899
rect 17000 5868 17049 5896
rect 17000 5856 17006 5868
rect 17037 5865 17049 5868
rect 17083 5865 17095 5899
rect 18874 5896 18880 5908
rect 18835 5868 18880 5896
rect 17037 5859 17095 5865
rect 18874 5856 18880 5868
rect 18932 5856 18938 5908
rect 18601 5831 18659 5837
rect 18601 5797 18613 5831
rect 18647 5828 18659 5831
rect 19058 5828 19064 5840
rect 18647 5800 19064 5828
rect 18647 5797 18659 5800
rect 18601 5791 18659 5797
rect 19058 5788 19064 5800
rect 19116 5788 19122 5840
rect 12342 5720 12348 5772
rect 12400 5760 12406 5772
rect 12802 5760 12808 5772
rect 12400 5732 12808 5760
rect 12400 5720 12406 5732
rect 12802 5720 12808 5732
rect 12860 5760 12866 5772
rect 12989 5763 13047 5769
rect 12989 5760 13001 5763
rect 12860 5732 13001 5760
rect 12860 5720 12866 5732
rect 12989 5729 13001 5732
rect 13035 5729 13047 5763
rect 15930 5760 15936 5772
rect 15891 5732 15936 5760
rect 12989 5723 13047 5729
rect 15930 5720 15936 5732
rect 15988 5720 15994 5772
rect 23474 5720 23480 5772
rect 23532 5760 23538 5772
rect 23661 5763 23719 5769
rect 23661 5760 23673 5763
rect 23532 5732 23673 5760
rect 23532 5720 23538 5732
rect 23661 5729 23673 5732
rect 23707 5760 23719 5763
rect 23842 5760 23848 5772
rect 23707 5732 23848 5760
rect 23707 5729 23719 5732
rect 23661 5723 23719 5729
rect 23842 5720 23848 5732
rect 23900 5720 23906 5772
rect 12526 5652 12532 5704
rect 12584 5692 12590 5704
rect 12713 5695 12771 5701
rect 12713 5692 12725 5695
rect 12584 5664 12725 5692
rect 12584 5652 12590 5664
rect 12713 5661 12725 5664
rect 12759 5661 12771 5695
rect 12713 5655 12771 5661
rect 15657 5695 15715 5701
rect 15657 5661 15669 5695
rect 15703 5692 15715 5695
rect 16022 5692 16028 5704
rect 15703 5664 16028 5692
rect 15703 5661 15715 5664
rect 15657 5655 15715 5661
rect 16022 5652 16028 5664
rect 16080 5652 16086 5704
rect 18138 5516 18144 5568
rect 18196 5556 18202 5568
rect 19150 5556 19156 5568
rect 18196 5528 19156 5556
rect 18196 5516 18202 5528
rect 19150 5516 19156 5528
rect 19208 5556 19214 5568
rect 19245 5559 19303 5565
rect 19245 5556 19257 5559
rect 19208 5528 19257 5556
rect 19208 5516 19214 5528
rect 19245 5525 19257 5528
rect 19291 5525 19303 5559
rect 23474 5556 23480 5568
rect 23435 5528 23480 5556
rect 19245 5519 19303 5525
rect 23474 5516 23480 5528
rect 23532 5516 23538 5568
rect 1104 5466 38548 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 38548 5466
rect 1104 5392 38548 5414
rect 10413 5355 10471 5361
rect 10413 5321 10425 5355
rect 10459 5352 10471 5355
rect 10502 5352 10508 5364
rect 10459 5324 10508 5352
rect 10459 5321 10471 5324
rect 10413 5315 10471 5321
rect 10502 5312 10508 5324
rect 10560 5312 10566 5364
rect 12802 5352 12808 5364
rect 12763 5324 12808 5352
rect 12802 5312 12808 5324
rect 12860 5312 12866 5364
rect 16022 5352 16028 5364
rect 15983 5324 16028 5352
rect 16022 5312 16028 5324
rect 16080 5312 16086 5364
rect 23842 5352 23848 5364
rect 23803 5324 23848 5352
rect 23842 5312 23848 5324
rect 23900 5312 23906 5364
rect 12526 5244 12532 5296
rect 12584 5284 12590 5296
rect 13081 5287 13139 5293
rect 13081 5284 13093 5287
rect 12584 5256 13093 5284
rect 12584 5244 12590 5256
rect 13081 5253 13093 5256
rect 13127 5253 13139 5287
rect 13081 5247 13139 5253
rect 15749 5287 15807 5293
rect 15749 5253 15761 5287
rect 15795 5284 15807 5287
rect 15930 5284 15936 5296
rect 15795 5256 15936 5284
rect 15795 5253 15807 5256
rect 15749 5247 15807 5253
rect 15930 5244 15936 5256
rect 15988 5244 15994 5296
rect 8757 5219 8815 5225
rect 8757 5185 8769 5219
rect 8803 5216 8815 5219
rect 8803 5188 9168 5216
rect 8803 5185 8815 5188
rect 8757 5179 8815 5185
rect 8294 5108 8300 5160
rect 8352 5148 8358 5160
rect 8846 5148 8852 5160
rect 8352 5120 8852 5148
rect 8352 5108 8358 5120
rect 8846 5108 8852 5120
rect 8904 5108 8910 5160
rect 9140 5157 9168 5188
rect 9125 5151 9183 5157
rect 9125 5117 9137 5151
rect 9171 5148 9183 5151
rect 9214 5148 9220 5160
rect 9171 5120 9220 5148
rect 9171 5117 9183 5120
rect 9125 5111 9183 5117
rect 9214 5108 9220 5120
rect 9272 5108 9278 5160
rect 21821 5151 21879 5157
rect 21821 5117 21833 5151
rect 21867 5148 21879 5151
rect 22189 5151 22247 5157
rect 22189 5148 22201 5151
rect 21867 5120 22201 5148
rect 21867 5117 21879 5120
rect 21821 5111 21879 5117
rect 22189 5117 22201 5120
rect 22235 5148 22247 5151
rect 23474 5148 23480 5160
rect 22235 5120 23480 5148
rect 22235 5117 22247 5120
rect 22189 5111 22247 5117
rect 23474 5108 23480 5120
rect 23532 5148 23538 5160
rect 25593 5151 25651 5157
rect 25593 5148 25605 5151
rect 23532 5120 25605 5148
rect 23532 5108 23538 5120
rect 25593 5117 25605 5120
rect 25639 5148 25651 5151
rect 25869 5151 25927 5157
rect 25869 5148 25881 5151
rect 25639 5120 25881 5148
rect 25639 5117 25651 5120
rect 25593 5111 25651 5117
rect 25869 5117 25881 5120
rect 25915 5117 25927 5151
rect 25869 5111 25927 5117
rect 21634 5012 21640 5024
rect 21595 4984 21640 5012
rect 21634 4972 21640 4984
rect 21692 4972 21698 5024
rect 25406 5012 25412 5024
rect 25367 4984 25412 5012
rect 25406 4972 25412 4984
rect 25464 4972 25470 5024
rect 1104 4922 38548 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 38548 4922
rect 1104 4848 38548 4870
rect 8846 4808 8852 4820
rect 8807 4780 8852 4808
rect 8846 4768 8852 4780
rect 8904 4768 8910 4820
rect 12158 4808 12164 4820
rect 12119 4780 12164 4808
rect 12158 4768 12164 4780
rect 12216 4768 12222 4820
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 17310 4808 17316 4820
rect 13872 4780 17316 4808
rect 13872 4768 13878 4780
rect 17310 4768 17316 4780
rect 17368 4768 17374 4820
rect 33502 4808 33508 4820
rect 33463 4780 33508 4808
rect 33502 4768 33508 4780
rect 33560 4768 33566 4820
rect 19426 4740 19432 4752
rect 19387 4712 19432 4740
rect 19426 4700 19432 4712
rect 19484 4700 19490 4752
rect 28169 4743 28227 4749
rect 28169 4709 28181 4743
rect 28215 4740 28227 4743
rect 28902 4740 28908 4752
rect 28215 4712 28908 4740
rect 28215 4709 28227 4712
rect 28169 4703 28227 4709
rect 28902 4700 28908 4712
rect 28960 4700 28966 4752
rect 10781 4675 10839 4681
rect 10781 4641 10793 4675
rect 10827 4672 10839 4675
rect 11330 4672 11336 4684
rect 10827 4644 11336 4672
rect 10827 4641 10839 4644
rect 10781 4635 10839 4641
rect 11330 4632 11336 4644
rect 11388 4672 11394 4684
rect 12526 4672 12532 4684
rect 11388 4644 12532 4672
rect 11388 4632 11394 4644
rect 12526 4632 12532 4644
rect 12584 4632 12590 4684
rect 16022 4632 16028 4684
rect 16080 4672 16086 4684
rect 17773 4675 17831 4681
rect 17773 4672 17785 4675
rect 16080 4644 17785 4672
rect 16080 4632 16086 4644
rect 17773 4641 17785 4644
rect 17819 4672 17831 4675
rect 18138 4672 18144 4684
rect 17819 4644 18144 4672
rect 17819 4641 17831 4644
rect 17773 4635 17831 4641
rect 18138 4632 18144 4644
rect 18196 4632 18202 4684
rect 32401 4675 32459 4681
rect 32401 4641 32413 4675
rect 32447 4672 32459 4675
rect 32674 4672 32680 4684
rect 32447 4644 32680 4672
rect 32447 4641 32459 4644
rect 32401 4635 32459 4641
rect 32674 4632 32680 4644
rect 32732 4632 32738 4684
rect 11054 4604 11060 4616
rect 11015 4576 11060 4604
rect 11054 4564 11060 4576
rect 11112 4564 11118 4616
rect 17954 4564 17960 4616
rect 18012 4604 18018 4616
rect 18049 4607 18107 4613
rect 18049 4604 18061 4607
rect 18012 4576 18061 4604
rect 18012 4564 18018 4576
rect 18049 4573 18061 4576
rect 18095 4573 18107 4607
rect 26510 4604 26516 4616
rect 26471 4576 26516 4604
rect 18049 4567 18107 4573
rect 26510 4564 26516 4576
rect 26568 4564 26574 4616
rect 26786 4604 26792 4616
rect 26747 4576 26792 4604
rect 26786 4564 26792 4576
rect 26844 4564 26850 4616
rect 32122 4604 32128 4616
rect 32083 4576 32128 4604
rect 32122 4564 32128 4576
rect 32180 4564 32186 4616
rect 1104 4378 38548 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 38548 4378
rect 1104 4304 38548 4326
rect 9950 4264 9956 4276
rect 9911 4236 9956 4264
rect 9950 4224 9956 4236
rect 10008 4224 10014 4276
rect 11241 4267 11299 4273
rect 11241 4233 11253 4267
rect 11287 4264 11299 4267
rect 11330 4264 11336 4276
rect 11287 4236 11336 4264
rect 11287 4233 11299 4236
rect 11241 4227 11299 4233
rect 11330 4224 11336 4236
rect 11388 4224 11394 4276
rect 18138 4224 18144 4276
rect 18196 4264 18202 4276
rect 18233 4267 18291 4273
rect 18233 4264 18245 4267
rect 18196 4236 18245 4264
rect 18196 4224 18202 4236
rect 18233 4233 18245 4236
rect 18279 4233 18291 4267
rect 18233 4227 18291 4233
rect 8294 4088 8300 4140
rect 8352 4128 8358 4140
rect 8389 4131 8447 4137
rect 8389 4128 8401 4131
rect 8352 4100 8401 4128
rect 8352 4088 8358 4100
rect 8389 4097 8401 4100
rect 8435 4097 8447 4131
rect 8389 4091 8447 4097
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 8496 4032 8677 4060
rect 8496 3992 8524 4032
rect 8665 4029 8677 4032
rect 8711 4029 8723 4063
rect 17862 4060 17868 4072
rect 17823 4032 17868 4060
rect 8665 4023 8723 4029
rect 17862 4020 17868 4032
rect 17920 4020 17926 4072
rect 18248 4060 18276 4227
rect 26786 4224 26792 4276
rect 26844 4264 26850 4276
rect 27341 4267 27399 4273
rect 27341 4264 27353 4267
rect 26844 4236 27353 4264
rect 26844 4224 26850 4236
rect 27341 4233 27353 4236
rect 27387 4233 27399 4267
rect 27341 4227 27399 4233
rect 19061 4131 19119 4137
rect 19061 4097 19073 4131
rect 19107 4128 19119 4131
rect 19429 4131 19487 4137
rect 19429 4128 19441 4131
rect 19107 4100 19441 4128
rect 19107 4097 19119 4100
rect 19061 4091 19119 4097
rect 19429 4097 19441 4100
rect 19475 4128 19487 4131
rect 20530 4128 20536 4140
rect 19475 4100 20536 4128
rect 19475 4097 19487 4100
rect 19429 4091 19487 4097
rect 20530 4088 20536 4100
rect 20588 4088 20594 4140
rect 20809 4131 20867 4137
rect 20809 4097 20821 4131
rect 20855 4128 20867 4131
rect 21266 4128 21272 4140
rect 20855 4100 21272 4128
rect 20855 4097 20867 4100
rect 20809 4091 20867 4097
rect 21266 4088 21272 4100
rect 21324 4088 21330 4140
rect 25317 4131 25375 4137
rect 25317 4097 25329 4131
rect 25363 4128 25375 4131
rect 26878 4128 26884 4140
rect 25363 4100 25728 4128
rect 26839 4100 26884 4128
rect 25363 4097 25375 4100
rect 25317 4091 25375 4097
rect 19150 4060 19156 4072
rect 18248 4032 19156 4060
rect 19150 4020 19156 4032
rect 19208 4020 19214 4072
rect 25406 4060 25412 4072
rect 25367 4032 25412 4060
rect 25406 4020 25412 4032
rect 25464 4020 25470 4072
rect 25700 4069 25728 4100
rect 26878 4088 26884 4100
rect 26936 4088 26942 4140
rect 25685 4063 25743 4069
rect 25685 4029 25697 4063
rect 25731 4060 25743 4063
rect 25774 4060 25780 4072
rect 25731 4032 25780 4060
rect 25731 4029 25743 4032
rect 25685 4023 25743 4029
rect 25774 4020 25780 4032
rect 25832 4020 25838 4072
rect 8312 3964 8524 3992
rect 7834 3884 7840 3936
rect 7892 3924 7898 3936
rect 8312 3933 8340 3964
rect 9674 3952 9680 4004
rect 9732 3992 9738 4004
rect 10781 3995 10839 4001
rect 10781 3992 10793 3995
rect 9732 3964 10793 3992
rect 9732 3952 9738 3964
rect 10781 3961 10793 3964
rect 10827 3992 10839 3995
rect 10962 3992 10968 4004
rect 10827 3964 10968 3992
rect 10827 3961 10839 3964
rect 10781 3955 10839 3961
rect 10962 3952 10968 3964
rect 11020 3952 11026 4004
rect 32217 3995 32275 4001
rect 32217 3961 32229 3995
rect 32263 3992 32275 3995
rect 32674 3992 32680 4004
rect 32263 3964 32680 3992
rect 32263 3961 32275 3964
rect 32217 3955 32275 3961
rect 32674 3952 32680 3964
rect 32732 3952 32738 4004
rect 8297 3927 8355 3933
rect 8297 3924 8309 3927
rect 7892 3896 8309 3924
rect 7892 3884 7898 3896
rect 8297 3893 8309 3896
rect 8343 3893 8355 3927
rect 8297 3887 8355 3893
rect 32122 3884 32128 3936
rect 32180 3924 32186 3936
rect 32493 3927 32551 3933
rect 32493 3924 32505 3927
rect 32180 3896 32505 3924
rect 32180 3884 32186 3896
rect 32493 3893 32505 3896
rect 32539 3893 32551 3927
rect 32493 3887 32551 3893
rect 1104 3834 38548 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 38548 3834
rect 1104 3760 38548 3782
rect 8294 3680 8300 3732
rect 8352 3720 8358 3732
rect 8389 3723 8447 3729
rect 8389 3720 8401 3723
rect 8352 3692 8401 3720
rect 8352 3680 8358 3692
rect 8389 3689 8401 3692
rect 8435 3689 8447 3723
rect 11514 3720 11520 3732
rect 11475 3692 11520 3720
rect 8389 3683 8447 3689
rect 11514 3680 11520 3692
rect 11572 3680 11578 3732
rect 19150 3720 19156 3732
rect 19111 3692 19156 3720
rect 19150 3680 19156 3692
rect 19208 3720 19214 3732
rect 19978 3720 19984 3732
rect 19208 3692 19984 3720
rect 19208 3680 19214 3692
rect 19978 3680 19984 3692
rect 20036 3680 20042 3732
rect 24670 3720 24676 3732
rect 24631 3692 24676 3720
rect 24670 3680 24676 3692
rect 24728 3680 24734 3732
rect 33134 3680 33140 3732
rect 33192 3720 33198 3732
rect 33505 3723 33563 3729
rect 33505 3720 33517 3723
rect 33192 3692 33517 3720
rect 33192 3680 33198 3692
rect 33505 3689 33517 3692
rect 33551 3689 33563 3723
rect 33505 3683 33563 3689
rect 16945 3655 17003 3661
rect 16945 3621 16957 3655
rect 16991 3652 17003 3655
rect 17034 3652 17040 3664
rect 16991 3624 17040 3652
rect 16991 3621 17003 3624
rect 16945 3615 17003 3621
rect 17034 3612 17040 3624
rect 17092 3612 17098 3664
rect 1762 3584 1768 3596
rect 1723 3556 1768 3584
rect 1762 3544 1768 3556
rect 1820 3544 1826 3596
rect 4341 3587 4399 3593
rect 4341 3553 4353 3587
rect 4387 3584 4399 3587
rect 4614 3584 4620 3596
rect 4387 3556 4620 3584
rect 4387 3553 4399 3556
rect 4341 3547 4399 3553
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 10137 3587 10195 3593
rect 10137 3553 10149 3587
rect 10183 3584 10195 3587
rect 10778 3584 10784 3596
rect 10183 3556 10784 3584
rect 10183 3553 10195 3556
rect 10137 3547 10195 3553
rect 10778 3544 10784 3556
rect 10836 3584 10842 3596
rect 11330 3584 11336 3596
rect 10836 3556 11336 3584
rect 10836 3544 10842 3556
rect 11330 3544 11336 3556
rect 11388 3544 11394 3596
rect 15289 3587 15347 3593
rect 15289 3553 15301 3587
rect 15335 3584 15347 3587
rect 15378 3584 15384 3596
rect 15335 3556 15384 3584
rect 15335 3553 15347 3556
rect 15289 3547 15347 3553
rect 15378 3544 15384 3556
rect 15436 3544 15442 3596
rect 23198 3544 23204 3596
rect 23256 3584 23262 3596
rect 23385 3587 23443 3593
rect 23385 3584 23397 3587
rect 23256 3556 23397 3584
rect 23256 3544 23262 3556
rect 23385 3553 23397 3556
rect 23431 3553 23443 3587
rect 23385 3547 23443 3553
rect 1486 3516 1492 3528
rect 1447 3488 1492 3516
rect 1486 3476 1492 3488
rect 1544 3476 1550 3528
rect 3142 3516 3148 3528
rect 3103 3488 3148 3516
rect 3142 3476 3148 3488
rect 3200 3476 3206 3528
rect 3418 3476 3424 3528
rect 3476 3516 3482 3528
rect 4065 3519 4123 3525
rect 4065 3516 4077 3519
rect 3476 3488 4077 3516
rect 3476 3476 3482 3488
rect 4065 3485 4077 3488
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 10413 3519 10471 3525
rect 10413 3485 10425 3519
rect 10459 3516 10471 3519
rect 10502 3516 10508 3528
rect 10459 3488 10508 3516
rect 10459 3485 10471 3488
rect 10413 3479 10471 3485
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 15562 3516 15568 3528
rect 15523 3488 15568 3516
rect 15562 3476 15568 3488
rect 15620 3476 15626 3528
rect 23106 3516 23112 3528
rect 23067 3488 23112 3516
rect 23106 3476 23112 3488
rect 23164 3476 23170 3528
rect 32122 3516 32128 3528
rect 32083 3488 32128 3516
rect 32122 3476 32128 3488
rect 32180 3476 32186 3528
rect 32398 3516 32404 3528
rect 32359 3488 32404 3516
rect 32398 3476 32404 3488
rect 32456 3476 32462 3528
rect 4706 3340 4712 3392
rect 4764 3380 4770 3392
rect 5445 3383 5503 3389
rect 5445 3380 5457 3383
rect 4764 3352 5457 3380
rect 4764 3340 4770 3352
rect 5445 3349 5457 3352
rect 5491 3349 5503 3383
rect 19978 3380 19984 3392
rect 19939 3352 19984 3380
rect 5445 3343 5503 3349
rect 19978 3340 19984 3352
rect 20036 3340 20042 3392
rect 25406 3340 25412 3392
rect 25464 3380 25470 3392
rect 25501 3383 25559 3389
rect 25501 3380 25513 3383
rect 25464 3352 25513 3380
rect 25464 3340 25470 3352
rect 25501 3349 25513 3352
rect 25547 3380 25559 3383
rect 26510 3380 26516 3392
rect 25547 3352 26516 3380
rect 25547 3349 25559 3352
rect 25501 3343 25559 3349
rect 26510 3340 26516 3352
rect 26568 3380 26574 3392
rect 26789 3383 26847 3389
rect 26789 3380 26801 3383
rect 26568 3352 26801 3380
rect 26568 3340 26574 3352
rect 26789 3349 26801 3352
rect 26835 3380 26847 3383
rect 27338 3380 27344 3392
rect 26835 3352 27344 3380
rect 26835 3349 26847 3352
rect 26789 3343 26847 3349
rect 27338 3340 27344 3352
rect 27396 3340 27402 3392
rect 35802 3380 35808 3392
rect 35763 3352 35808 3380
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 1104 3290 38548 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 38548 3290
rect 1104 3216 38548 3238
rect 1486 3136 1492 3188
rect 1544 3176 1550 3188
rect 1949 3179 2007 3185
rect 1949 3176 1961 3179
rect 1544 3148 1961 3176
rect 1544 3136 1550 3148
rect 1949 3145 1961 3148
rect 1995 3176 2007 3179
rect 3418 3176 3424 3188
rect 1995 3148 3424 3176
rect 1995 3145 2007 3148
rect 1949 3139 2007 3145
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 4157 3179 4215 3185
rect 4157 3145 4169 3179
rect 4203 3176 4215 3179
rect 4614 3176 4620 3188
rect 4203 3148 4620 3176
rect 4203 3145 4215 3148
rect 4157 3139 4215 3145
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 10045 3179 10103 3185
rect 10045 3145 10057 3179
rect 10091 3176 10103 3179
rect 10686 3176 10692 3188
rect 10091 3148 10692 3176
rect 10091 3145 10103 3148
rect 10045 3139 10103 3145
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 10778 3136 10784 3188
rect 10836 3176 10842 3188
rect 10836 3148 10881 3176
rect 10836 3136 10842 3148
rect 14734 3136 14740 3188
rect 14792 3176 14798 3188
rect 15289 3179 15347 3185
rect 15289 3176 15301 3179
rect 14792 3148 15301 3176
rect 14792 3136 14798 3148
rect 15289 3145 15301 3148
rect 15335 3176 15347 3179
rect 15562 3176 15568 3188
rect 15335 3148 15568 3176
rect 15335 3145 15347 3148
rect 15289 3139 15347 3145
rect 15562 3136 15568 3148
rect 15620 3136 15626 3188
rect 16945 3179 17003 3185
rect 16945 3145 16957 3179
rect 16991 3176 17003 3179
rect 17678 3176 17684 3188
rect 16991 3148 17684 3176
rect 16991 3145 17003 3148
rect 16945 3139 17003 3145
rect 17678 3136 17684 3148
rect 17736 3136 17742 3188
rect 21266 3176 21272 3188
rect 21227 3148 21272 3176
rect 21266 3136 21272 3148
rect 21324 3136 21330 3188
rect 23106 3136 23112 3188
rect 23164 3176 23170 3188
rect 23845 3179 23903 3185
rect 23845 3176 23857 3179
rect 23164 3148 23857 3176
rect 23164 3136 23170 3148
rect 23845 3145 23857 3148
rect 23891 3145 23903 3179
rect 24578 3176 24584 3188
rect 24539 3148 24584 3176
rect 23845 3139 23903 3145
rect 24578 3136 24584 3148
rect 24636 3136 24642 3188
rect 26329 3179 26387 3185
rect 26329 3145 26341 3179
rect 26375 3176 26387 3179
rect 26418 3176 26424 3188
rect 26375 3148 26424 3176
rect 26375 3145 26387 3148
rect 26329 3139 26387 3145
rect 26418 3136 26424 3148
rect 26476 3136 26482 3188
rect 29089 3179 29147 3185
rect 29089 3145 29101 3179
rect 29135 3176 29147 3179
rect 29546 3176 29552 3188
rect 29135 3148 29552 3176
rect 29135 3145 29147 3148
rect 29089 3139 29147 3145
rect 29546 3136 29552 3148
rect 29604 3136 29610 3188
rect 32766 3136 32772 3188
rect 32824 3176 32830 3188
rect 33137 3179 33195 3185
rect 33137 3176 33149 3179
rect 32824 3148 33149 3176
rect 32824 3136 32830 3148
rect 33137 3145 33149 3148
rect 33183 3145 33195 3179
rect 37366 3176 37372 3188
rect 37327 3148 37372 3176
rect 33137 3139 33195 3145
rect 37366 3136 37372 3148
rect 37424 3136 37430 3188
rect 1673 3111 1731 3117
rect 1673 3077 1685 3111
rect 1719 3108 1731 3111
rect 1762 3108 1768 3120
rect 1719 3080 1768 3108
rect 1719 3077 1731 3080
rect 1673 3071 1731 3077
rect 1762 3068 1768 3080
rect 1820 3068 1826 3120
rect 23198 3108 23204 3120
rect 23159 3080 23204 3108
rect 23198 3068 23204 3080
rect 23256 3068 23262 3120
rect 4614 3000 4620 3052
rect 4672 3040 4678 3052
rect 4798 3040 4804 3052
rect 4672 3012 4804 3040
rect 4672 3000 4678 3012
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 8389 3043 8447 3049
rect 8389 3009 8401 3043
rect 8435 3040 8447 3043
rect 8754 3040 8760 3052
rect 8435 3012 8760 3040
rect 8435 3009 8447 3012
rect 8389 3003 8447 3009
rect 8754 3000 8760 3012
rect 8812 3000 8818 3052
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3040 14611 3043
rect 15378 3040 15384 3052
rect 14599 3012 15384 3040
rect 14599 3009 14611 3012
rect 14553 3003 14611 3009
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 15654 3040 15660 3052
rect 15615 3012 15660 3040
rect 15654 3000 15660 3012
rect 15712 3000 15718 3052
rect 19797 3043 19855 3049
rect 19797 3009 19809 3043
rect 19843 3040 19855 3043
rect 24596 3040 24624 3136
rect 25041 3043 25099 3049
rect 25041 3040 25053 3043
rect 19843 3012 20208 3040
rect 24596 3012 25053 3040
rect 19843 3009 19855 3012
rect 19797 3003 19855 3009
rect 8294 2932 8300 2984
rect 8352 2972 8358 2984
rect 8478 2972 8484 2984
rect 8352 2944 8484 2972
rect 8352 2932 8358 2944
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 10502 2972 10508 2984
rect 10463 2944 10508 2972
rect 10502 2932 10508 2944
rect 10560 2932 10566 2984
rect 14921 2975 14979 2981
rect 14921 2941 14933 2975
rect 14967 2972 14979 2975
rect 15672 2972 15700 3000
rect 20180 2984 20208 3012
rect 25041 3009 25053 3012
rect 25087 3009 25099 3043
rect 25041 3003 25099 3009
rect 29273 3043 29331 3049
rect 29273 3009 29285 3043
rect 29319 3040 29331 3043
rect 31665 3043 31723 3049
rect 29319 3012 31248 3040
rect 29319 3009 29331 3012
rect 29273 3003 29331 3009
rect 29380 2984 29408 3012
rect 14967 2944 15700 2972
rect 19889 2975 19947 2981
rect 14967 2941 14979 2944
rect 14921 2935 14979 2941
rect 19889 2941 19901 2975
rect 19935 2972 19947 2975
rect 19978 2972 19984 2984
rect 19935 2944 19984 2972
rect 19935 2941 19947 2944
rect 19889 2935 19947 2941
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 20162 2972 20168 2984
rect 20123 2944 20168 2972
rect 20162 2932 20168 2944
rect 20220 2932 20226 2984
rect 24765 2975 24823 2981
rect 24765 2941 24777 2975
rect 24811 2972 24823 2975
rect 24854 2972 24860 2984
rect 24811 2944 24860 2972
rect 24811 2941 24823 2944
rect 24765 2935 24823 2941
rect 24854 2932 24860 2944
rect 24912 2932 24918 2984
rect 29362 2932 29368 2984
rect 29420 2932 29426 2984
rect 29546 2972 29552 2984
rect 29507 2944 29552 2972
rect 29546 2932 29552 2944
rect 29604 2932 29610 2984
rect 31220 2981 31248 3012
rect 31665 3009 31677 3043
rect 31711 3040 31723 3043
rect 32033 3043 32091 3049
rect 32033 3040 32045 3043
rect 31711 3012 32045 3040
rect 31711 3009 31723 3012
rect 31665 3003 31723 3009
rect 32033 3009 32045 3012
rect 32079 3040 32091 3043
rect 32214 3040 32220 3052
rect 32079 3012 32220 3040
rect 32079 3009 32091 3012
rect 32033 3003 32091 3009
rect 32214 3000 32220 3012
rect 32272 3000 32278 3052
rect 31205 2975 31263 2981
rect 31205 2941 31217 2975
rect 31251 2972 31263 2975
rect 31757 2975 31815 2981
rect 31757 2972 31769 2975
rect 31251 2944 31769 2972
rect 31251 2941 31263 2944
rect 31205 2935 31263 2941
rect 31757 2941 31769 2944
rect 31803 2972 31815 2975
rect 32122 2972 32128 2984
rect 31803 2944 32128 2972
rect 31803 2941 31815 2944
rect 31757 2935 31815 2941
rect 32122 2932 32128 2944
rect 32180 2972 32186 2984
rect 35802 2972 35808 2984
rect 32180 2944 35808 2972
rect 32180 2932 32186 2944
rect 35802 2932 35808 2944
rect 35860 2932 35866 2984
rect 36081 2975 36139 2981
rect 36081 2972 36093 2975
rect 35912 2944 36093 2972
rect 30929 2907 30987 2913
rect 30929 2873 30941 2907
rect 30975 2904 30987 2907
rect 31294 2904 31300 2916
rect 30975 2876 31300 2904
rect 30975 2873 30987 2876
rect 30929 2867 30987 2873
rect 31294 2864 31300 2876
rect 31352 2864 31358 2916
rect 3418 2796 3424 2848
rect 3476 2836 3482 2848
rect 4338 2836 4344 2848
rect 3476 2808 4344 2836
rect 3476 2796 3482 2808
rect 4338 2796 4344 2808
rect 4396 2836 4402 2848
rect 4433 2839 4491 2845
rect 4433 2836 4445 2839
rect 4396 2808 4445 2836
rect 4396 2796 4402 2808
rect 4433 2805 4445 2808
rect 4479 2805 4491 2839
rect 4433 2799 4491 2805
rect 19426 2796 19432 2848
rect 19484 2836 19490 2848
rect 27522 2836 27528 2848
rect 19484 2808 27528 2836
rect 19484 2796 19490 2808
rect 27522 2796 27528 2808
rect 27580 2796 27586 2848
rect 35618 2836 35624 2848
rect 35579 2808 35624 2836
rect 35618 2796 35624 2808
rect 35676 2836 35682 2848
rect 35912 2836 35940 2944
rect 36081 2941 36093 2944
rect 36127 2941 36139 2975
rect 36081 2935 36139 2941
rect 35676 2808 35940 2836
rect 35676 2796 35682 2808
rect 1104 2746 38548 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 38548 2746
rect 1104 2672 38548 2694
rect 3418 2632 3424 2644
rect 3379 2604 3424 2632
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 8478 2632 8484 2644
rect 8439 2604 8484 2632
rect 8478 2592 8484 2604
rect 8536 2592 8542 2644
rect 11422 2632 11428 2644
rect 11383 2604 11428 2632
rect 11422 2592 11428 2604
rect 11480 2592 11486 2644
rect 12437 2635 12495 2641
rect 12437 2601 12449 2635
rect 12483 2632 12495 2635
rect 12526 2632 12532 2644
rect 12483 2604 12532 2632
rect 12483 2601 12495 2604
rect 12437 2595 12495 2601
rect 12526 2592 12532 2604
rect 12584 2592 12590 2644
rect 15378 2592 15384 2644
rect 15436 2632 15442 2644
rect 15749 2635 15807 2641
rect 15749 2632 15761 2635
rect 15436 2604 15761 2632
rect 15436 2592 15442 2604
rect 15749 2601 15761 2604
rect 15795 2632 15807 2635
rect 17773 2635 17831 2641
rect 17773 2632 17785 2635
rect 15795 2604 17785 2632
rect 15795 2601 15807 2604
rect 15749 2595 15807 2601
rect 17773 2601 17785 2604
rect 17819 2632 17831 2635
rect 18322 2632 18328 2644
rect 17819 2604 18328 2632
rect 17819 2601 17831 2604
rect 17773 2595 17831 2601
rect 18322 2592 18328 2604
rect 18380 2632 18386 2644
rect 19978 2632 19984 2644
rect 18380 2604 19984 2632
rect 18380 2592 18386 2604
rect 19978 2592 19984 2604
rect 20036 2592 20042 2644
rect 22830 2632 22836 2644
rect 22791 2604 22836 2632
rect 22830 2592 22836 2604
rect 22888 2592 22894 2644
rect 29362 2632 29368 2644
rect 29323 2604 29368 2632
rect 29362 2592 29368 2604
rect 29420 2592 29426 2644
rect 31849 2635 31907 2641
rect 31849 2601 31861 2635
rect 31895 2632 31907 2635
rect 32122 2632 32128 2644
rect 31895 2604 32128 2632
rect 31895 2601 31907 2604
rect 31849 2595 31907 2601
rect 32122 2592 32128 2604
rect 32180 2592 32186 2644
rect 35158 2632 35164 2644
rect 35119 2604 35164 2632
rect 35158 2592 35164 2604
rect 35216 2592 35222 2644
rect 5997 2567 6055 2573
rect 5997 2533 6009 2567
rect 6043 2564 6055 2567
rect 6178 2564 6184 2576
rect 6043 2536 6184 2564
rect 6043 2533 6055 2536
rect 5997 2527 6055 2533
rect 6178 2524 6184 2536
rect 6236 2524 6242 2576
rect 11330 2524 11336 2576
rect 11388 2564 11394 2576
rect 11977 2567 12035 2573
rect 11977 2564 11989 2567
rect 11388 2536 11989 2564
rect 11388 2524 11394 2536
rect 11977 2533 11989 2536
rect 12023 2533 12035 2567
rect 11977 2527 12035 2533
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 3804 2468 4629 2496
rect 3694 2252 3700 2304
rect 3752 2292 3758 2304
rect 3804 2301 3832 2468
rect 4617 2465 4629 2468
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 9585 2499 9643 2505
rect 9585 2465 9597 2499
rect 9631 2496 9643 2499
rect 10318 2496 10324 2508
rect 9631 2468 10324 2496
rect 9631 2465 9643 2468
rect 9585 2459 9643 2465
rect 10318 2456 10324 2468
rect 10376 2456 10382 2508
rect 4338 2428 4344 2440
rect 4299 2400 4344 2428
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2428 9275 2431
rect 10045 2431 10103 2437
rect 10045 2428 10057 2431
rect 9263 2400 10057 2428
rect 9263 2397 9275 2400
rect 9217 2391 9275 2397
rect 10045 2397 10057 2400
rect 10091 2428 10103 2431
rect 11348 2428 11376 2524
rect 10091 2400 11376 2428
rect 11992 2428 12020 2527
rect 12544 2496 12572 2592
rect 28813 2567 28871 2573
rect 28813 2533 28825 2567
rect 28859 2564 28871 2567
rect 29178 2564 29184 2576
rect 28859 2536 29184 2564
rect 28859 2533 28871 2536
rect 28813 2527 28871 2533
rect 29178 2524 29184 2536
rect 29236 2524 29242 2576
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12544 2468 13185 2496
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 18601 2499 18659 2505
rect 18601 2496 18613 2499
rect 13173 2459 13231 2465
rect 18064 2468 18613 2496
rect 12897 2431 12955 2437
rect 12897 2428 12909 2431
rect 11992 2400 12909 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 12897 2397 12909 2400
rect 12943 2397 12955 2431
rect 12897 2391 12955 2397
rect 14553 2431 14611 2437
rect 14553 2397 14565 2431
rect 14599 2428 14611 2431
rect 16114 2428 16120 2440
rect 14599 2400 16120 2428
rect 14599 2397 14611 2400
rect 14553 2391 14611 2397
rect 16114 2388 16120 2400
rect 16172 2388 16178 2440
rect 18064 2372 18092 2468
rect 18601 2465 18613 2468
rect 18647 2465 18659 2499
rect 18601 2459 18659 2465
rect 20993 2499 21051 2505
rect 20993 2465 21005 2499
rect 21039 2496 21051 2499
rect 21729 2499 21787 2505
rect 21729 2496 21741 2499
rect 21039 2468 21741 2496
rect 21039 2465 21051 2468
rect 20993 2459 21051 2465
rect 21729 2465 21741 2468
rect 21775 2496 21787 2499
rect 21818 2496 21824 2508
rect 21775 2468 21824 2496
rect 21775 2465 21787 2468
rect 21729 2459 21787 2465
rect 21818 2456 21824 2468
rect 21876 2456 21882 2508
rect 26697 2499 26755 2505
rect 26697 2465 26709 2499
rect 26743 2496 26755 2499
rect 34885 2499 34943 2505
rect 26743 2468 27476 2496
rect 26743 2465 26755 2468
rect 26697 2459 26755 2465
rect 18322 2428 18328 2440
rect 18283 2400 18328 2428
rect 18322 2388 18328 2400
rect 18380 2388 18386 2440
rect 19978 2388 19984 2440
rect 20036 2428 20042 2440
rect 20625 2431 20683 2437
rect 20625 2428 20637 2431
rect 20036 2400 20637 2428
rect 20036 2388 20042 2400
rect 20625 2397 20637 2400
rect 20671 2428 20683 2431
rect 21453 2431 21511 2437
rect 21453 2428 21465 2431
rect 20671 2400 21465 2428
rect 20671 2397 20683 2400
rect 20625 2391 20683 2397
rect 21453 2397 21465 2400
rect 21499 2428 21511 2431
rect 21634 2428 21640 2440
rect 21499 2400 21640 2428
rect 21499 2397 21511 2400
rect 21453 2391 21511 2397
rect 21634 2388 21640 2400
rect 21692 2428 21698 2440
rect 23106 2428 23112 2440
rect 21692 2400 23112 2428
rect 21692 2388 21698 2400
rect 23106 2388 23112 2400
rect 23164 2388 23170 2440
rect 24854 2428 24860 2440
rect 24767 2400 24860 2428
rect 24854 2388 24860 2400
rect 24912 2428 24918 2440
rect 26329 2431 26387 2437
rect 26329 2428 26341 2431
rect 24912 2400 26341 2428
rect 24912 2388 24918 2400
rect 26329 2397 26341 2400
rect 26375 2428 26387 2431
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 26375 2400 27169 2428
rect 26375 2397 26387 2400
rect 26329 2391 26387 2397
rect 27157 2397 27169 2400
rect 27203 2428 27215 2431
rect 27338 2428 27344 2440
rect 27203 2400 27344 2428
rect 27203 2397 27215 2400
rect 27157 2391 27215 2397
rect 27338 2388 27344 2400
rect 27396 2388 27402 2440
rect 27448 2437 27476 2468
rect 34885 2465 34897 2499
rect 34931 2496 34943 2499
rect 35437 2499 35495 2505
rect 35437 2496 35449 2499
rect 34931 2468 35449 2496
rect 34931 2465 34943 2468
rect 34885 2459 34943 2465
rect 35437 2465 35449 2468
rect 35483 2496 35495 2499
rect 35802 2496 35808 2508
rect 35483 2468 35808 2496
rect 35483 2465 35495 2468
rect 35437 2459 35495 2465
rect 35802 2456 35808 2468
rect 35860 2456 35866 2508
rect 27433 2431 27491 2437
rect 27433 2397 27445 2431
rect 27479 2428 27491 2431
rect 27522 2428 27528 2440
rect 27479 2400 27528 2428
rect 27479 2397 27491 2400
rect 27433 2391 27491 2397
rect 27522 2388 27528 2400
rect 27580 2388 27586 2440
rect 35158 2388 35164 2440
rect 35216 2428 35222 2440
rect 35713 2431 35771 2437
rect 35713 2428 35725 2431
rect 35216 2400 35725 2428
rect 35216 2388 35222 2400
rect 35713 2397 35725 2400
rect 35759 2397 35771 2431
rect 35713 2391 35771 2397
rect 18046 2360 18052 2372
rect 18007 2332 18052 2360
rect 18046 2320 18052 2332
rect 18104 2320 18110 2372
rect 3789 2295 3847 2301
rect 3789 2292 3801 2295
rect 3752 2264 3801 2292
rect 3752 2252 3758 2264
rect 3789 2261 3801 2264
rect 3835 2261 3847 2295
rect 3789 2255 3847 2261
rect 19794 2252 19800 2304
rect 19852 2292 19858 2304
rect 19889 2295 19947 2301
rect 19889 2292 19901 2295
rect 19852 2264 19901 2292
rect 19852 2252 19858 2264
rect 19889 2261 19901 2264
rect 19935 2261 19947 2295
rect 19889 2255 19947 2261
rect 32217 2295 32275 2301
rect 32217 2261 32229 2295
rect 32263 2292 32275 2295
rect 32398 2292 32404 2304
rect 32263 2264 32404 2292
rect 32263 2261 32275 2264
rect 32217 2255 32275 2261
rect 32398 2252 32404 2264
rect 32456 2252 32462 2304
rect 36354 2252 36360 2304
rect 36412 2292 36418 2304
rect 36817 2295 36875 2301
rect 36817 2292 36829 2295
rect 36412 2264 36829 2292
rect 36412 2252 36418 2264
rect 36817 2261 36829 2264
rect 36863 2261 36875 2295
rect 36817 2255 36875 2261
rect 1104 2202 38548 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 38548 2202
rect 1104 2128 38548 2150
rect 29086 2048 29092 2100
rect 29144 2088 29150 2100
rect 37274 2088 37280 2100
rect 29144 2060 37280 2088
rect 29144 2048 29150 2060
rect 37274 2048 37280 2060
rect 37332 2048 37338 2100
rect 15654 1776 15660 1828
rect 15712 1816 15718 1828
rect 16390 1816 16396 1828
rect 15712 1788 16396 1816
rect 15712 1776 15718 1788
rect 16390 1776 16396 1788
rect 16448 1776 16454 1828
rect 32398 1708 32404 1760
rect 32456 1748 32462 1760
rect 33042 1748 33048 1760
rect 32456 1720 33048 1748
rect 32456 1708 32462 1720
rect 33042 1708 33048 1720
rect 33100 1708 33106 1760
rect 8294 1572 8300 1624
rect 8352 1612 8358 1624
rect 17862 1612 17868 1624
rect 8352 1584 17868 1612
rect 8352 1572 8358 1584
rect 17862 1572 17868 1584
rect 17920 1572 17926 1624
rect 17034 1164 17040 1216
rect 17092 1204 17098 1216
rect 17770 1204 17776 1216
rect 17092 1176 17776 1204
rect 17092 1164 17098 1176
rect 17770 1164 17776 1176
rect 17828 1164 17834 1216
<< via1 >>
rect 3424 40196 3476 40248
rect 7012 40196 7064 40248
rect 2964 40128 3016 40180
rect 19156 40128 19208 40180
rect 3240 40060 3292 40112
rect 20076 40060 20128 40112
rect 26884 40060 26936 40112
rect 35256 40060 35308 40112
rect 15752 39380 15804 39432
rect 33600 39380 33652 39432
rect 4160 39312 4212 39364
rect 5172 39312 5224 39364
rect 8852 39312 8904 39364
rect 22928 39312 22980 39364
rect 11428 39244 11480 39296
rect 34520 39244 34572 39296
rect 4246 39142 4298 39194
rect 4310 39142 4362 39194
rect 4374 39142 4426 39194
rect 4438 39142 4490 39194
rect 34966 39142 35018 39194
rect 35030 39142 35082 39194
rect 35094 39142 35146 39194
rect 35158 39142 35210 39194
rect 2780 39040 2832 39092
rect 8852 39040 8904 39092
rect 9680 39040 9732 39092
rect 11428 39083 11480 39092
rect 11428 39049 11437 39083
rect 11437 39049 11471 39083
rect 11471 39049 11480 39083
rect 11428 39040 11480 39049
rect 26240 39040 26292 39092
rect 27344 39040 27396 39092
rect 6460 38972 6512 39024
rect 12900 38904 12952 38956
rect 19984 38972 20036 39024
rect 15752 38947 15804 38956
rect 15752 38913 15761 38947
rect 15761 38913 15795 38947
rect 15795 38913 15804 38947
rect 15752 38904 15804 38913
rect 35256 38904 35308 38956
rect 2780 38700 2832 38752
rect 5448 38836 5500 38888
rect 9680 38836 9732 38888
rect 13360 38836 13412 38888
rect 13636 38836 13688 38888
rect 14372 38879 14424 38888
rect 14372 38845 14381 38879
rect 14381 38845 14415 38879
rect 14415 38845 14424 38879
rect 14372 38836 14424 38845
rect 15292 38768 15344 38820
rect 26148 38768 26200 38820
rect 17868 38700 17920 38752
rect 26056 38700 26108 38752
rect 27344 38879 27396 38888
rect 27344 38845 27353 38879
rect 27353 38845 27387 38879
rect 27387 38845 27396 38879
rect 27344 38836 27396 38845
rect 28724 38811 28776 38820
rect 28724 38777 28733 38811
rect 28733 38777 28767 38811
rect 28767 38777 28776 38811
rect 28724 38768 28776 38777
rect 19606 38598 19658 38650
rect 19670 38598 19722 38650
rect 19734 38598 19786 38650
rect 19798 38598 19850 38650
rect 5540 38496 5592 38548
rect 6736 38496 6788 38548
rect 13360 38496 13412 38548
rect 13636 38539 13688 38548
rect 13636 38505 13645 38539
rect 13645 38505 13679 38539
rect 13679 38505 13688 38539
rect 13636 38496 13688 38505
rect 19432 38496 19484 38548
rect 24584 38496 24636 38548
rect 31484 38496 31536 38548
rect 37740 38496 37792 38548
rect 20 38428 72 38480
rect 480 38428 532 38480
rect 3700 38428 3752 38480
rect 4620 38360 4672 38412
rect 5540 38360 5592 38412
rect 13360 38403 13412 38412
rect 13360 38369 13369 38403
rect 13369 38369 13403 38403
rect 13403 38369 13412 38403
rect 13360 38360 13412 38369
rect 17316 38360 17368 38412
rect 23204 38403 23256 38412
rect 23204 38369 23213 38403
rect 23213 38369 23247 38403
rect 23247 38369 23256 38403
rect 23204 38360 23256 38369
rect 26792 38403 26844 38412
rect 26792 38369 26801 38403
rect 26801 38369 26835 38403
rect 26835 38369 26844 38403
rect 26792 38360 26844 38369
rect 29460 38360 29512 38412
rect 31760 38360 31812 38412
rect 1492 38335 1544 38344
rect 1492 38301 1501 38335
rect 1501 38301 1535 38335
rect 1535 38301 1544 38335
rect 1492 38292 1544 38301
rect 1676 38292 1728 38344
rect 5448 38335 5500 38344
rect 5448 38301 5457 38335
rect 5457 38301 5491 38335
rect 5491 38301 5500 38335
rect 5448 38292 5500 38301
rect 7656 38292 7708 38344
rect 11704 38335 11756 38344
rect 7380 38199 7432 38208
rect 7380 38165 7389 38199
rect 7389 38165 7423 38199
rect 7423 38165 7432 38199
rect 7380 38156 7432 38165
rect 9680 38156 9732 38208
rect 11704 38301 11713 38335
rect 11713 38301 11747 38335
rect 11747 38301 11756 38335
rect 11704 38292 11756 38301
rect 11888 38292 11940 38344
rect 17224 38335 17276 38344
rect 17224 38301 17233 38335
rect 17233 38301 17267 38335
rect 17267 38301 17276 38335
rect 17224 38292 17276 38301
rect 23388 38292 23440 38344
rect 26056 38292 26108 38344
rect 30012 38292 30064 38344
rect 32128 38335 32180 38344
rect 32128 38301 32137 38335
rect 32137 38301 32171 38335
rect 32171 38301 32180 38335
rect 32128 38292 32180 38301
rect 15292 38156 15344 38208
rect 18236 38156 18288 38208
rect 19432 38199 19484 38208
rect 19432 38165 19441 38199
rect 19441 38165 19475 38199
rect 19475 38165 19484 38199
rect 19432 38156 19484 38165
rect 24308 38199 24360 38208
rect 24308 38165 24317 38199
rect 24317 38165 24351 38199
rect 24351 38165 24360 38199
rect 24308 38156 24360 38165
rect 27896 38199 27948 38208
rect 27896 38165 27905 38199
rect 27905 38165 27939 38199
rect 27939 38165 27948 38199
rect 27896 38156 27948 38165
rect 31024 38156 31076 38208
rect 33232 38156 33284 38208
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 34966 38054 35018 38106
rect 35030 38054 35082 38106
rect 35094 38054 35146 38106
rect 35158 38054 35210 38106
rect 1492 37952 1544 38004
rect 2688 37952 2740 38004
rect 5540 37995 5592 38004
rect 5540 37961 5549 37995
rect 5549 37961 5583 37995
rect 5583 37961 5592 37995
rect 5540 37952 5592 37961
rect 7012 37952 7064 38004
rect 11888 37995 11940 38004
rect 5448 37816 5500 37868
rect 11888 37961 11897 37995
rect 11897 37961 11931 37995
rect 11931 37961 11940 37995
rect 11888 37952 11940 37961
rect 23204 37952 23256 38004
rect 25228 37952 25280 38004
rect 29460 37952 29512 38004
rect 30012 37995 30064 38004
rect 30012 37961 30021 37995
rect 30021 37961 30055 37995
rect 30055 37961 30064 37995
rect 30012 37952 30064 37961
rect 31392 37995 31444 38004
rect 31392 37961 31401 37995
rect 31401 37961 31435 37995
rect 31435 37961 31444 37995
rect 31392 37952 31444 37961
rect 31760 37952 31812 38004
rect 33232 37884 33284 37936
rect 19984 37816 20036 37868
rect 26700 37816 26752 37868
rect 32404 37859 32456 37868
rect 32404 37825 32413 37859
rect 32413 37825 32447 37859
rect 32447 37825 32456 37859
rect 32404 37816 32456 37825
rect 7380 37791 7432 37800
rect 7380 37757 7389 37791
rect 7389 37757 7423 37791
rect 7423 37757 7432 37791
rect 7380 37748 7432 37757
rect 17316 37791 17368 37800
rect 9036 37723 9088 37732
rect 9036 37689 9045 37723
rect 9045 37689 9079 37723
rect 9079 37689 9088 37723
rect 9036 37680 9088 37689
rect 17316 37757 17325 37791
rect 17325 37757 17359 37791
rect 17359 37757 17368 37791
rect 17316 37748 17368 37757
rect 19432 37748 19484 37800
rect 36084 37859 36136 37868
rect 36084 37825 36093 37859
rect 36093 37825 36127 37859
rect 36127 37825 36136 37859
rect 36084 37816 36136 37825
rect 33232 37791 33284 37800
rect 33232 37757 33241 37791
rect 33241 37757 33275 37791
rect 33275 37757 33284 37791
rect 33232 37748 33284 37757
rect 35716 37680 35768 37732
rect 1676 37655 1728 37664
rect 1676 37621 1685 37655
rect 1685 37621 1719 37655
rect 1719 37621 1728 37655
rect 1676 37612 1728 37621
rect 10416 37655 10468 37664
rect 10416 37621 10425 37655
rect 10425 37621 10459 37655
rect 10459 37621 10468 37655
rect 10416 37612 10468 37621
rect 10968 37612 11020 37664
rect 11704 37612 11756 37664
rect 12164 37655 12216 37664
rect 12164 37621 12173 37655
rect 12173 37621 12207 37655
rect 12207 37621 12216 37655
rect 12164 37612 12216 37621
rect 17224 37612 17276 37664
rect 18144 37612 18196 37664
rect 20720 37655 20772 37664
rect 20720 37621 20729 37655
rect 20729 37621 20763 37655
rect 20763 37621 20772 37655
rect 20720 37612 20772 37621
rect 23388 37655 23440 37664
rect 23388 37621 23397 37655
rect 23397 37621 23431 37655
rect 23431 37621 23440 37655
rect 23388 37612 23440 37621
rect 26056 37612 26108 37664
rect 31852 37612 31904 37664
rect 36544 37612 36596 37664
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 1584 37408 1636 37460
rect 2320 37408 2372 37460
rect 26792 37451 26844 37460
rect 26792 37417 26801 37451
rect 26801 37417 26835 37451
rect 26835 37417 26844 37451
rect 26792 37408 26844 37417
rect 34796 37408 34848 37460
rect 32128 37340 32180 37392
rect 5448 37272 5500 37324
rect 6000 37272 6052 37324
rect 9680 37315 9732 37324
rect 9680 37281 9689 37315
rect 9689 37281 9723 37315
rect 9723 37281 9732 37315
rect 9680 37272 9732 37281
rect 9956 37315 10008 37324
rect 9956 37281 9965 37315
rect 9965 37281 9999 37315
rect 9999 37281 10008 37315
rect 9956 37272 10008 37281
rect 12440 37315 12492 37324
rect 12440 37281 12449 37315
rect 12449 37281 12483 37315
rect 12483 37281 12492 37315
rect 12440 37272 12492 37281
rect 13820 37272 13872 37324
rect 15016 37272 15068 37324
rect 15568 37315 15620 37324
rect 15568 37281 15577 37315
rect 15577 37281 15611 37315
rect 15611 37281 15620 37315
rect 15568 37272 15620 37281
rect 17592 37272 17644 37324
rect 18604 37315 18656 37324
rect 18604 37281 18613 37315
rect 18613 37281 18647 37315
rect 18647 37281 18656 37315
rect 18604 37272 18656 37281
rect 26056 37272 26108 37324
rect 33232 37272 33284 37324
rect 33600 37272 33652 37324
rect 10048 37204 10100 37256
rect 12164 37247 12216 37256
rect 12164 37213 12173 37247
rect 12173 37213 12207 37247
rect 12207 37213 12216 37247
rect 12164 37204 12216 37213
rect 12624 37204 12676 37256
rect 15292 37247 15344 37256
rect 15292 37213 15301 37247
rect 15301 37213 15335 37247
rect 15335 37213 15344 37247
rect 15292 37204 15344 37213
rect 18144 37204 18196 37256
rect 33876 37272 33928 37324
rect 34428 37272 34480 37324
rect 34520 37272 34572 37324
rect 35716 37272 35768 37324
rect 7012 37111 7064 37120
rect 7012 37077 7021 37111
rect 7021 37077 7055 37111
rect 7055 37077 7064 37111
rect 7012 37068 7064 37077
rect 11244 37111 11296 37120
rect 11244 37077 11253 37111
rect 11253 37077 11287 37111
rect 11287 37077 11296 37111
rect 11244 37068 11296 37077
rect 13544 37111 13596 37120
rect 13544 37077 13553 37111
rect 13553 37077 13587 37111
rect 13587 37077 13596 37111
rect 13544 37068 13596 37077
rect 19432 37068 19484 37120
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 1676 36907 1728 36916
rect 1676 36873 1685 36907
rect 1685 36873 1719 36907
rect 1719 36873 1728 36907
rect 1676 36864 1728 36873
rect 2320 36907 2372 36916
rect 2320 36873 2329 36907
rect 2329 36873 2363 36907
rect 2363 36873 2372 36907
rect 2320 36864 2372 36873
rect 6000 36864 6052 36916
rect 9956 36864 10008 36916
rect 10048 36907 10100 36916
rect 10048 36873 10057 36907
rect 10057 36873 10091 36907
rect 10091 36873 10100 36907
rect 10048 36864 10100 36873
rect 11060 36864 11112 36916
rect 12348 36864 12400 36916
rect 12624 36907 12676 36916
rect 12624 36873 12633 36907
rect 12633 36873 12667 36907
rect 12667 36873 12676 36907
rect 12624 36864 12676 36873
rect 15568 36864 15620 36916
rect 18604 36864 18656 36916
rect 27528 36864 27580 36916
rect 33876 36907 33928 36916
rect 33876 36873 33885 36907
rect 33885 36873 33919 36907
rect 33919 36873 33928 36907
rect 33876 36864 33928 36873
rect 34428 36864 34480 36916
rect 36544 36864 36596 36916
rect 5448 36728 5500 36780
rect 19432 36771 19484 36780
rect 19432 36737 19441 36771
rect 19441 36737 19475 36771
rect 19475 36737 19484 36771
rect 19432 36728 19484 36737
rect 25136 36771 25188 36780
rect 25136 36737 25145 36771
rect 25145 36737 25179 36771
rect 25179 36737 25188 36771
rect 25136 36728 25188 36737
rect 35808 36771 35860 36780
rect 35808 36737 35817 36771
rect 35817 36737 35851 36771
rect 35851 36737 35860 36771
rect 35808 36728 35860 36737
rect 1768 36660 1820 36712
rect 18144 36660 18196 36712
rect 20812 36635 20864 36644
rect 20812 36601 20821 36635
rect 20821 36601 20855 36635
rect 20855 36601 20864 36635
rect 20812 36592 20864 36601
rect 25136 36592 25188 36644
rect 26056 36660 26108 36712
rect 35532 36592 35584 36644
rect 36544 36703 36596 36712
rect 36544 36669 36553 36703
rect 36553 36669 36587 36703
rect 36587 36669 36596 36703
rect 36544 36660 36596 36669
rect 15292 36524 15344 36576
rect 16488 36524 16540 36576
rect 35440 36567 35492 36576
rect 35440 36533 35449 36567
rect 35449 36533 35483 36567
rect 35483 36533 35492 36567
rect 35440 36524 35492 36533
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 10048 36320 10100 36372
rect 22836 36320 22888 36372
rect 23020 36320 23072 36372
rect 37464 36320 37516 36372
rect 38660 36320 38712 36372
rect 5172 36227 5224 36236
rect 5172 36193 5181 36227
rect 5181 36193 5215 36227
rect 5215 36193 5224 36227
rect 5172 36184 5224 36193
rect 5448 36184 5500 36236
rect 10600 36227 10652 36236
rect 10600 36193 10609 36227
rect 10609 36193 10643 36227
rect 10643 36193 10652 36227
rect 10600 36184 10652 36193
rect 16488 36184 16540 36236
rect 16672 36159 16724 36168
rect 16672 36125 16681 36159
rect 16681 36125 16715 36159
rect 16715 36125 16724 36159
rect 16672 36116 16724 36125
rect 18052 36159 18104 36168
rect 18052 36125 18061 36159
rect 18061 36125 18095 36159
rect 18095 36125 18104 36159
rect 18052 36116 18104 36125
rect 1768 35980 1820 36032
rect 6920 35980 6972 36032
rect 18144 35980 18196 36032
rect 25136 35980 25188 36032
rect 35532 35980 35584 36032
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 5172 35776 5224 35828
rect 5448 35776 5500 35828
rect 10600 35776 10652 35828
rect 24952 35819 25004 35828
rect 24952 35785 24961 35819
rect 24961 35785 24995 35819
rect 24995 35785 25004 35819
rect 24952 35776 25004 35785
rect 36084 35683 36136 35692
rect 36084 35649 36093 35683
rect 36093 35649 36127 35683
rect 36127 35649 36136 35683
rect 36084 35640 36136 35649
rect 18052 35615 18104 35624
rect 18052 35581 18061 35615
rect 18061 35581 18095 35615
rect 18095 35581 18104 35615
rect 18052 35572 18104 35581
rect 16488 35504 16540 35556
rect 17776 35547 17828 35556
rect 15936 35436 15988 35488
rect 16672 35436 16724 35488
rect 17776 35513 17785 35547
rect 17785 35513 17819 35547
rect 17819 35513 17828 35547
rect 25136 35615 25188 35624
rect 25136 35581 25145 35615
rect 25145 35581 25179 35615
rect 25179 35581 25188 35615
rect 25136 35572 25188 35581
rect 35900 35572 35952 35624
rect 17776 35504 17828 35513
rect 19892 35504 19944 35556
rect 26792 35547 26844 35556
rect 26792 35513 26801 35547
rect 26801 35513 26835 35547
rect 26835 35513 26844 35547
rect 26792 35504 26844 35513
rect 18144 35436 18196 35488
rect 36084 35436 36136 35488
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 10600 35232 10652 35284
rect 29276 35232 29328 35284
rect 30012 35232 30064 35284
rect 14004 35164 14056 35216
rect 6920 35096 6972 35148
rect 11888 35139 11940 35148
rect 11888 35105 11897 35139
rect 11897 35105 11931 35139
rect 11931 35105 11940 35139
rect 11888 35096 11940 35105
rect 7380 35028 7432 35080
rect 9772 34892 9824 34944
rect 14740 34935 14792 34944
rect 14740 34901 14749 34935
rect 14749 34901 14783 34935
rect 14783 34901 14792 34935
rect 14740 34892 14792 34901
rect 18144 34935 18196 34944
rect 18144 34901 18153 34935
rect 18153 34901 18187 34935
rect 18187 34901 18196 34935
rect 18144 34892 18196 34901
rect 24584 34892 24636 34944
rect 25136 34935 25188 34944
rect 25136 34901 25145 34935
rect 25145 34901 25179 34935
rect 25179 34901 25188 34935
rect 25136 34892 25188 34901
rect 35900 34935 35952 34944
rect 35900 34901 35909 34935
rect 35909 34901 35943 34935
rect 35943 34901 35952 34935
rect 35900 34892 35952 34901
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 6920 34688 6972 34740
rect 7380 34731 7432 34740
rect 7380 34697 7389 34731
rect 7389 34697 7423 34731
rect 7423 34697 7432 34731
rect 7380 34688 7432 34697
rect 11060 34688 11112 34740
rect 11888 34688 11940 34740
rect 14004 34731 14056 34740
rect 14004 34697 14013 34731
rect 14013 34697 14047 34731
rect 14047 34697 14056 34731
rect 14004 34688 14056 34697
rect 25136 34688 25188 34740
rect 37372 34731 37424 34740
rect 14740 34595 14792 34604
rect 14740 34561 14749 34595
rect 14749 34561 14783 34595
rect 14783 34561 14792 34595
rect 14740 34552 14792 34561
rect 20076 34595 20128 34604
rect 20076 34561 20085 34595
rect 20085 34561 20119 34595
rect 20119 34561 20128 34595
rect 20076 34552 20128 34561
rect 20904 34552 20956 34604
rect 15292 34484 15344 34536
rect 19432 34484 19484 34536
rect 24584 34527 24636 34536
rect 24584 34493 24593 34527
rect 24593 34493 24627 34527
rect 24627 34493 24636 34527
rect 24584 34484 24636 34493
rect 37372 34697 37381 34731
rect 37381 34697 37415 34731
rect 37415 34697 37424 34731
rect 37372 34688 37424 34697
rect 30656 34663 30708 34672
rect 30656 34629 30665 34663
rect 30665 34629 30699 34663
rect 30699 34629 30708 34663
rect 30656 34620 30708 34629
rect 26884 34552 26936 34604
rect 29920 34552 29972 34604
rect 36084 34595 36136 34604
rect 36084 34561 36093 34595
rect 36093 34561 36127 34595
rect 36127 34561 36136 34595
rect 36084 34552 36136 34561
rect 27160 34484 27212 34536
rect 29276 34527 29328 34536
rect 29276 34493 29285 34527
rect 29285 34493 29319 34527
rect 29319 34493 29328 34527
rect 29276 34484 29328 34493
rect 35900 34484 35952 34536
rect 14556 34459 14608 34468
rect 14556 34425 14565 34459
rect 14565 34425 14599 34459
rect 14599 34425 14608 34459
rect 14556 34416 14608 34425
rect 15108 34348 15160 34400
rect 16488 34348 16540 34400
rect 24400 34391 24452 34400
rect 24400 34357 24409 34391
rect 24409 34357 24443 34391
rect 24443 34357 24452 34391
rect 24400 34348 24452 34357
rect 26424 34348 26476 34400
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 15108 34187 15160 34196
rect 15108 34153 15117 34187
rect 15117 34153 15151 34187
rect 15151 34153 15160 34187
rect 15108 34144 15160 34153
rect 15752 34187 15804 34196
rect 15752 34153 15761 34187
rect 15761 34153 15795 34187
rect 15795 34153 15804 34187
rect 15752 34144 15804 34153
rect 27160 34144 27212 34196
rect 27896 34144 27948 34196
rect 9772 34008 9824 34060
rect 15660 34008 15712 34060
rect 16488 34051 16540 34060
rect 16488 34017 16497 34051
rect 16497 34017 16531 34051
rect 16531 34017 16540 34051
rect 16488 34008 16540 34017
rect 17132 34008 17184 34060
rect 17960 34051 18012 34060
rect 17960 34017 17969 34051
rect 17969 34017 18003 34051
rect 18003 34017 18012 34051
rect 17960 34008 18012 34017
rect 21824 34008 21876 34060
rect 22468 34051 22520 34060
rect 22468 34017 22477 34051
rect 22477 34017 22511 34051
rect 22511 34017 22520 34051
rect 22468 34008 22520 34017
rect 23664 34008 23716 34060
rect 24400 34008 24452 34060
rect 27988 34008 28040 34060
rect 30288 34051 30340 34060
rect 10048 33940 10100 33992
rect 14556 33940 14608 33992
rect 15108 33940 15160 33992
rect 18144 33940 18196 33992
rect 19432 33940 19484 33992
rect 21732 33983 21784 33992
rect 21732 33949 21741 33983
rect 21741 33949 21775 33983
rect 21775 33949 21784 33983
rect 21732 33940 21784 33949
rect 23756 33940 23808 33992
rect 29644 33983 29696 33992
rect 29644 33949 29653 33983
rect 29653 33949 29687 33983
rect 29687 33949 29696 33983
rect 29644 33940 29696 33949
rect 30288 34017 30297 34051
rect 30297 34017 30331 34051
rect 30331 34017 30340 34051
rect 30288 34008 30340 34017
rect 30196 33940 30248 33992
rect 30380 33983 30432 33992
rect 30380 33949 30389 33983
rect 30389 33949 30423 33983
rect 30423 33949 30432 33983
rect 30380 33940 30432 33949
rect 22376 33915 22428 33924
rect 22376 33881 22385 33915
rect 22385 33881 22419 33915
rect 22419 33881 22428 33915
rect 22376 33872 22428 33881
rect 11980 33804 12032 33856
rect 16672 33804 16724 33856
rect 19064 33847 19116 33856
rect 19064 33813 19073 33847
rect 19073 33813 19107 33847
rect 19107 33813 19116 33847
rect 19064 33804 19116 33813
rect 20352 33847 20404 33856
rect 20352 33813 20361 33847
rect 20361 33813 20395 33847
rect 20395 33813 20404 33847
rect 20352 33804 20404 33813
rect 25412 33847 25464 33856
rect 25412 33813 25421 33847
rect 25421 33813 25455 33847
rect 25455 33813 25464 33847
rect 25412 33804 25464 33813
rect 27988 33804 28040 33856
rect 29000 33804 29052 33856
rect 30104 33804 30156 33856
rect 35900 33847 35952 33856
rect 35900 33813 35909 33847
rect 35909 33813 35943 33847
rect 35943 33813 35952 33847
rect 35900 33804 35952 33813
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 9772 33643 9824 33652
rect 9772 33609 9781 33643
rect 9781 33609 9815 33643
rect 9815 33609 9824 33643
rect 9772 33600 9824 33609
rect 10048 33643 10100 33652
rect 10048 33609 10057 33643
rect 10057 33609 10091 33643
rect 10091 33609 10100 33643
rect 10048 33600 10100 33609
rect 14556 33600 14608 33652
rect 16212 33643 16264 33652
rect 16212 33609 16221 33643
rect 16221 33609 16255 33643
rect 16255 33609 16264 33643
rect 16212 33600 16264 33609
rect 17960 33600 18012 33652
rect 21732 33600 21784 33652
rect 24400 33600 24452 33652
rect 26240 33600 26292 33652
rect 22468 33575 22520 33584
rect 22468 33541 22477 33575
rect 22477 33541 22511 33575
rect 22511 33541 22520 33575
rect 22468 33532 22520 33541
rect 16672 33507 16724 33516
rect 16672 33473 16681 33507
rect 16681 33473 16715 33507
rect 16715 33473 16724 33507
rect 16672 33464 16724 33473
rect 20444 33507 20496 33516
rect 20444 33473 20453 33507
rect 20453 33473 20487 33507
rect 20487 33473 20496 33507
rect 20444 33464 20496 33473
rect 20536 33507 20588 33516
rect 20536 33473 20545 33507
rect 20545 33473 20579 33507
rect 20579 33473 20588 33507
rect 25504 33507 25556 33516
rect 20536 33464 20588 33473
rect 25504 33473 25513 33507
rect 25513 33473 25547 33507
rect 25547 33473 25556 33507
rect 25504 33464 25556 33473
rect 16948 33439 17000 33448
rect 16948 33405 16957 33439
rect 16957 33405 16991 33439
rect 16991 33405 17000 33439
rect 16948 33396 17000 33405
rect 17132 33439 17184 33448
rect 17132 33405 17141 33439
rect 17141 33405 17175 33439
rect 17175 33405 17184 33439
rect 17132 33396 17184 33405
rect 20352 33396 20404 33448
rect 21364 33439 21416 33448
rect 21364 33405 21373 33439
rect 21373 33405 21407 33439
rect 21407 33405 21416 33439
rect 21364 33396 21416 33405
rect 22376 33396 22428 33448
rect 25412 33439 25464 33448
rect 25412 33405 25421 33439
rect 25421 33405 25455 33439
rect 25455 33405 25464 33439
rect 25412 33396 25464 33405
rect 26424 33464 26476 33516
rect 27068 33464 27120 33516
rect 17960 33328 18012 33380
rect 23664 33328 23716 33380
rect 27252 33396 27304 33448
rect 27528 33396 27580 33448
rect 27896 33396 27948 33448
rect 30104 33396 30156 33448
rect 30196 33396 30248 33448
rect 17132 33260 17184 33312
rect 18144 33260 18196 33312
rect 19064 33303 19116 33312
rect 19064 33269 19073 33303
rect 19073 33269 19107 33303
rect 19107 33269 19116 33303
rect 19064 33260 19116 33269
rect 21824 33303 21876 33312
rect 21824 33269 21833 33303
rect 21833 33269 21867 33303
rect 21867 33269 21876 33303
rect 21824 33260 21876 33269
rect 23756 33260 23808 33312
rect 29644 33328 29696 33380
rect 30012 33371 30064 33380
rect 30012 33337 30021 33371
rect 30021 33337 30055 33371
rect 30055 33337 30064 33371
rect 30012 33328 30064 33337
rect 27160 33303 27212 33312
rect 27160 33269 27169 33303
rect 27169 33269 27203 33303
rect 27203 33269 27212 33303
rect 27160 33260 27212 33269
rect 28264 33260 28316 33312
rect 32036 33260 32088 33312
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 10968 33056 11020 33108
rect 16948 33056 17000 33108
rect 21364 33056 21416 33108
rect 24584 33056 24636 33108
rect 25412 33056 25464 33108
rect 28172 33056 28224 33108
rect 28908 33056 28960 33108
rect 29276 33056 29328 33108
rect 15476 32988 15528 33040
rect 15660 32988 15712 33040
rect 20352 32988 20404 33040
rect 30288 32988 30340 33040
rect 6092 32920 6144 32972
rect 11060 32963 11112 32972
rect 11060 32929 11069 32963
rect 11069 32929 11103 32963
rect 11103 32929 11112 32963
rect 11060 32920 11112 32929
rect 15844 32920 15896 32972
rect 16672 32920 16724 32972
rect 24952 32963 25004 32972
rect 6368 32852 6420 32904
rect 12624 32895 12676 32904
rect 12624 32861 12633 32895
rect 12633 32861 12667 32895
rect 12667 32861 12676 32895
rect 12624 32852 12676 32861
rect 12808 32852 12860 32904
rect 15660 32852 15712 32904
rect 16488 32852 16540 32904
rect 18144 32852 18196 32904
rect 18604 32895 18656 32904
rect 18604 32861 18613 32895
rect 18613 32861 18647 32895
rect 18647 32861 18656 32895
rect 18604 32852 18656 32861
rect 21364 32852 21416 32904
rect 21916 32895 21968 32904
rect 21916 32861 21925 32895
rect 21925 32861 21959 32895
rect 21959 32861 21968 32895
rect 21916 32852 21968 32861
rect 24952 32929 24961 32963
rect 24961 32929 24995 32963
rect 24995 32929 25004 32963
rect 24952 32920 25004 32929
rect 25320 32920 25372 32972
rect 26976 32963 27028 32972
rect 26976 32929 26985 32963
rect 26985 32929 27019 32963
rect 27019 32929 27028 32963
rect 26976 32920 27028 32929
rect 27344 32963 27396 32972
rect 27344 32929 27353 32963
rect 27353 32929 27387 32963
rect 27387 32929 27396 32963
rect 27344 32920 27396 32929
rect 28356 32963 28408 32972
rect 28356 32929 28365 32963
rect 28365 32929 28399 32963
rect 28399 32929 28408 32963
rect 28356 32920 28408 32929
rect 29000 32920 29052 32972
rect 30104 32963 30156 32972
rect 30104 32929 30113 32963
rect 30113 32929 30147 32963
rect 30147 32929 30156 32963
rect 30104 32920 30156 32929
rect 23296 32852 23348 32904
rect 27436 32895 27488 32904
rect 27436 32861 27445 32895
rect 27445 32861 27479 32895
rect 27479 32861 27488 32895
rect 27436 32852 27488 32861
rect 27252 32784 27304 32836
rect 29828 32852 29880 32904
rect 30564 32852 30616 32904
rect 30748 32895 30800 32904
rect 30748 32861 30757 32895
rect 30757 32861 30791 32895
rect 30791 32861 30800 32895
rect 30748 32852 30800 32861
rect 31208 32895 31260 32904
rect 31208 32861 31217 32895
rect 31217 32861 31251 32895
rect 31251 32861 31260 32895
rect 31208 32852 31260 32861
rect 7932 32716 7984 32768
rect 14004 32759 14056 32768
rect 14004 32725 14013 32759
rect 14013 32725 14047 32759
rect 14047 32725 14056 32759
rect 14004 32716 14056 32725
rect 23296 32716 23348 32768
rect 27804 32759 27856 32768
rect 27804 32725 27813 32759
rect 27813 32725 27847 32759
rect 27847 32725 27856 32759
rect 27804 32716 27856 32725
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 6000 32555 6052 32564
rect 6000 32521 6009 32555
rect 6009 32521 6043 32555
rect 6043 32521 6052 32555
rect 6000 32512 6052 32521
rect 6368 32555 6420 32564
rect 6368 32521 6377 32555
rect 6377 32521 6411 32555
rect 6411 32521 6420 32555
rect 6368 32512 6420 32521
rect 12624 32512 12676 32564
rect 16488 32512 16540 32564
rect 16304 32444 16356 32496
rect 17684 32512 17736 32564
rect 17960 32512 18012 32564
rect 18972 32555 19024 32564
rect 18972 32521 18981 32555
rect 18981 32521 19015 32555
rect 19015 32521 19024 32555
rect 18972 32512 19024 32521
rect 21916 32512 21968 32564
rect 25320 32555 25372 32564
rect 25320 32521 25329 32555
rect 25329 32521 25363 32555
rect 25363 32521 25372 32555
rect 25320 32512 25372 32521
rect 27344 32512 27396 32564
rect 28356 32512 28408 32564
rect 29552 32512 29604 32564
rect 29828 32512 29880 32564
rect 30104 32512 30156 32564
rect 18144 32444 18196 32496
rect 13728 32376 13780 32428
rect 19340 32419 19392 32428
rect 19340 32385 19349 32419
rect 19349 32385 19383 32419
rect 19383 32385 19392 32419
rect 25228 32444 25280 32496
rect 29000 32487 29052 32496
rect 29000 32453 29009 32487
rect 29009 32453 29043 32487
rect 29043 32453 29052 32487
rect 29000 32444 29052 32453
rect 23756 32419 23808 32428
rect 19340 32376 19392 32385
rect 23756 32385 23765 32419
rect 23765 32385 23799 32419
rect 23799 32385 23808 32419
rect 23756 32376 23808 32385
rect 13636 32308 13688 32360
rect 15292 32308 15344 32360
rect 16028 32351 16080 32360
rect 16028 32317 16037 32351
rect 16037 32317 16071 32351
rect 16071 32317 16080 32351
rect 16028 32308 16080 32317
rect 11060 32172 11112 32224
rect 12808 32172 12860 32224
rect 13360 32215 13412 32224
rect 13360 32181 13369 32215
rect 13369 32181 13403 32215
rect 13403 32181 13412 32215
rect 18420 32308 18472 32360
rect 18972 32308 19024 32360
rect 19064 32351 19116 32360
rect 19064 32317 19073 32351
rect 19073 32317 19107 32351
rect 19107 32317 19116 32351
rect 19064 32308 19116 32317
rect 17960 32240 18012 32292
rect 18604 32240 18656 32292
rect 13360 32172 13412 32181
rect 18144 32172 18196 32224
rect 26976 32308 27028 32360
rect 27804 32351 27856 32360
rect 27804 32317 27813 32351
rect 27813 32317 27847 32351
rect 27847 32317 27856 32351
rect 27804 32308 27856 32317
rect 28172 32351 28224 32360
rect 28172 32317 28181 32351
rect 28181 32317 28215 32351
rect 28215 32317 28224 32351
rect 28172 32308 28224 32317
rect 27436 32240 27488 32292
rect 28724 32308 28776 32360
rect 29552 32308 29604 32360
rect 30748 32240 30800 32292
rect 20076 32172 20128 32224
rect 21364 32172 21416 32224
rect 24952 32215 25004 32224
rect 24952 32181 24961 32215
rect 24961 32181 24995 32215
rect 24995 32181 25004 32215
rect 24952 32172 25004 32181
rect 31392 32172 31444 32224
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 13636 32011 13688 32020
rect 13636 31977 13645 32011
rect 13645 31977 13679 32011
rect 13679 31977 13688 32011
rect 13636 31968 13688 31977
rect 15384 31968 15436 32020
rect 16028 31968 16080 32020
rect 18512 31968 18564 32020
rect 19340 31968 19392 32020
rect 19432 31968 19484 32020
rect 26424 31968 26476 32020
rect 15752 31943 15804 31952
rect 15752 31909 15761 31943
rect 15761 31909 15795 31943
rect 15795 31909 15804 31943
rect 15752 31900 15804 31909
rect 16580 31943 16632 31952
rect 16580 31909 16589 31943
rect 16589 31909 16623 31943
rect 16623 31909 16632 31943
rect 16580 31900 16632 31909
rect 17500 31900 17552 31952
rect 18144 31900 18196 31952
rect 24400 31943 24452 31952
rect 24400 31909 24409 31943
rect 24409 31909 24443 31943
rect 24443 31909 24452 31943
rect 27988 31968 28040 32020
rect 24400 31900 24452 31909
rect 26976 31900 27028 31952
rect 28724 31900 28776 31952
rect 30012 31968 30064 32020
rect 31208 31968 31260 32020
rect 14004 31832 14056 31884
rect 17040 31875 17092 31884
rect 17040 31841 17049 31875
rect 17049 31841 17083 31875
rect 17083 31841 17092 31875
rect 17040 31832 17092 31841
rect 17224 31875 17276 31884
rect 17224 31841 17233 31875
rect 17233 31841 17267 31875
rect 17267 31841 17276 31875
rect 17224 31832 17276 31841
rect 18420 31875 18472 31884
rect 13820 31807 13872 31816
rect 13820 31773 13829 31807
rect 13829 31773 13863 31807
rect 13863 31773 13872 31807
rect 13820 31764 13872 31773
rect 16396 31764 16448 31816
rect 18420 31841 18429 31875
rect 18429 31841 18463 31875
rect 18463 31841 18472 31875
rect 18420 31832 18472 31841
rect 19340 31832 19392 31884
rect 24676 31875 24728 31884
rect 24676 31841 24685 31875
rect 24685 31841 24719 31875
rect 24719 31841 24728 31875
rect 24676 31832 24728 31841
rect 25412 31875 25464 31884
rect 25412 31841 25421 31875
rect 25421 31841 25455 31875
rect 25455 31841 25464 31875
rect 25412 31832 25464 31841
rect 25504 31875 25556 31884
rect 25504 31841 25513 31875
rect 25513 31841 25547 31875
rect 25547 31841 25556 31875
rect 26700 31875 26752 31884
rect 25504 31832 25556 31841
rect 26700 31841 26709 31875
rect 26709 31841 26743 31875
rect 26743 31841 26752 31875
rect 26700 31832 26752 31841
rect 27436 31832 27488 31884
rect 28264 31875 28316 31884
rect 28264 31841 28273 31875
rect 28273 31841 28307 31875
rect 28307 31841 28316 31875
rect 28264 31832 28316 31841
rect 28816 31875 28868 31884
rect 28816 31841 28825 31875
rect 28825 31841 28859 31875
rect 28859 31841 28868 31875
rect 28816 31832 28868 31841
rect 30104 31900 30156 31952
rect 29184 31875 29236 31884
rect 29184 31841 29193 31875
rect 29193 31841 29227 31875
rect 29227 31841 29236 31875
rect 29184 31832 29236 31841
rect 12532 31696 12584 31748
rect 16120 31696 16172 31748
rect 19248 31696 19300 31748
rect 20444 31764 20496 31816
rect 24584 31807 24636 31816
rect 24584 31773 24593 31807
rect 24593 31773 24627 31807
rect 24627 31773 24636 31807
rect 24584 31764 24636 31773
rect 26516 31807 26568 31816
rect 26516 31773 26525 31807
rect 26525 31773 26559 31807
rect 26559 31773 26568 31807
rect 26516 31764 26568 31773
rect 29736 31696 29788 31748
rect 3792 31628 3844 31680
rect 12900 31671 12952 31680
rect 12900 31637 12909 31671
rect 12909 31637 12943 31671
rect 12943 31637 12952 31671
rect 12900 31628 12952 31637
rect 23664 31671 23716 31680
rect 23664 31637 23673 31671
rect 23673 31637 23707 31671
rect 23707 31637 23716 31671
rect 23664 31628 23716 31637
rect 25964 31628 26016 31680
rect 27252 31628 27304 31680
rect 30932 31671 30984 31680
rect 30932 31637 30941 31671
rect 30941 31637 30975 31671
rect 30975 31637 30984 31671
rect 30932 31628 30984 31637
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 3056 31399 3108 31408
rect 3056 31365 3065 31399
rect 3065 31365 3099 31399
rect 3099 31365 3108 31399
rect 3056 31356 3108 31365
rect 2780 31288 2832 31340
rect 7748 31356 7800 31408
rect 4068 31331 4120 31340
rect 4068 31297 4077 31331
rect 4077 31297 4111 31331
rect 4111 31297 4120 31331
rect 4068 31288 4120 31297
rect 3792 31263 3844 31272
rect 3792 31229 3801 31263
rect 3801 31229 3835 31263
rect 3835 31229 3844 31263
rect 3792 31220 3844 31229
rect 10968 31424 11020 31476
rect 17040 31424 17092 31476
rect 25412 31424 25464 31476
rect 28724 31424 28776 31476
rect 30932 31424 30984 31476
rect 35624 31467 35676 31476
rect 16396 31399 16448 31408
rect 16396 31365 16405 31399
rect 16405 31365 16439 31399
rect 16439 31365 16448 31399
rect 16396 31356 16448 31365
rect 17592 31356 17644 31408
rect 18880 31356 18932 31408
rect 19156 31356 19208 31408
rect 23664 31356 23716 31408
rect 12900 31331 12952 31340
rect 12900 31297 12909 31331
rect 12909 31297 12943 31331
rect 12943 31297 12952 31331
rect 12900 31288 12952 31297
rect 20076 31288 20128 31340
rect 23848 31331 23900 31340
rect 23848 31297 23857 31331
rect 23857 31297 23891 31331
rect 23891 31297 23900 31331
rect 23848 31288 23900 31297
rect 4620 31152 4672 31204
rect 16396 31220 16448 31272
rect 14556 31195 14608 31204
rect 14556 31161 14565 31195
rect 14565 31161 14599 31195
rect 14599 31161 14608 31195
rect 14556 31152 14608 31161
rect 16672 31263 16724 31272
rect 16672 31229 16681 31263
rect 16681 31229 16715 31263
rect 16715 31229 16724 31263
rect 16672 31220 16724 31229
rect 16948 31220 17000 31272
rect 17868 31220 17920 31272
rect 18144 31220 18196 31272
rect 18880 31263 18932 31272
rect 18880 31229 18889 31263
rect 18889 31229 18923 31263
rect 18923 31229 18932 31263
rect 18880 31220 18932 31229
rect 19248 31263 19300 31272
rect 19248 31229 19257 31263
rect 19257 31229 19291 31263
rect 19291 31229 19300 31263
rect 19248 31220 19300 31229
rect 20260 31220 20312 31272
rect 23756 31263 23808 31272
rect 23756 31229 23765 31263
rect 23765 31229 23799 31263
rect 23799 31229 23808 31263
rect 23756 31220 23808 31229
rect 26516 31288 26568 31340
rect 27804 31288 27856 31340
rect 30012 31331 30064 31340
rect 30012 31297 30021 31331
rect 30021 31297 30055 31331
rect 30055 31297 30064 31331
rect 30012 31288 30064 31297
rect 30564 31288 30616 31340
rect 30932 31331 30984 31340
rect 30932 31297 30941 31331
rect 30941 31297 30975 31331
rect 30975 31297 30984 31331
rect 35624 31433 35633 31467
rect 35633 31433 35667 31467
rect 35667 31433 35676 31467
rect 35624 31424 35676 31433
rect 32128 31331 32180 31340
rect 30932 31288 30984 31297
rect 2688 31127 2740 31136
rect 2688 31093 2697 31127
rect 2697 31093 2731 31127
rect 2731 31093 2740 31127
rect 2688 31084 2740 31093
rect 10324 31127 10376 31136
rect 10324 31093 10333 31127
rect 10333 31093 10367 31127
rect 10367 31093 10376 31127
rect 10324 31084 10376 31093
rect 12992 31084 13044 31136
rect 18512 31152 18564 31204
rect 28816 31220 28868 31272
rect 29736 31263 29788 31272
rect 25964 31195 26016 31204
rect 25964 31161 25973 31195
rect 25973 31161 26007 31195
rect 26007 31161 26016 31195
rect 25964 31152 26016 31161
rect 27528 31195 27580 31204
rect 18052 31084 18104 31136
rect 18420 31084 18472 31136
rect 18696 31084 18748 31136
rect 19064 31127 19116 31136
rect 19064 31093 19073 31127
rect 19073 31093 19107 31127
rect 19107 31093 19116 31127
rect 19064 31084 19116 31093
rect 20996 31127 21048 31136
rect 20996 31093 21005 31127
rect 21005 31093 21039 31127
rect 21039 31093 21048 31127
rect 20996 31084 21048 31093
rect 23664 31084 23716 31136
rect 25044 31127 25096 31136
rect 25044 31093 25053 31127
rect 25053 31093 25087 31127
rect 25087 31093 25096 31127
rect 25044 31084 25096 31093
rect 26056 31084 26108 31136
rect 26516 31084 26568 31136
rect 26976 31127 27028 31136
rect 26976 31093 26985 31127
rect 26985 31093 27019 31127
rect 27019 31093 27028 31127
rect 27528 31161 27537 31195
rect 27537 31161 27571 31195
rect 27571 31161 27580 31195
rect 27528 31152 27580 31161
rect 29736 31229 29745 31263
rect 29745 31229 29779 31263
rect 29779 31229 29788 31263
rect 29736 31220 29788 31229
rect 31484 31220 31536 31272
rect 32128 31297 32137 31331
rect 32137 31297 32171 31331
rect 32171 31297 32180 31331
rect 32128 31288 32180 31297
rect 35900 31220 35952 31272
rect 30748 31152 30800 31204
rect 26976 31084 27028 31093
rect 27252 31084 27304 31136
rect 27436 31127 27488 31136
rect 27436 31093 27445 31127
rect 27445 31093 27479 31127
rect 27479 31093 27488 31127
rect 28172 31127 28224 31136
rect 27436 31084 27488 31093
rect 28172 31093 28181 31127
rect 28181 31093 28215 31127
rect 28215 31093 28224 31127
rect 28172 31084 28224 31093
rect 31668 31084 31720 31136
rect 37280 31084 37332 31136
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 4068 30880 4120 30932
rect 13820 30880 13872 30932
rect 13728 30812 13780 30864
rect 14004 30880 14056 30932
rect 16672 30923 16724 30932
rect 16672 30889 16681 30923
rect 16681 30889 16715 30923
rect 16715 30889 16724 30923
rect 16672 30880 16724 30889
rect 17224 30923 17276 30932
rect 17224 30889 17233 30923
rect 17233 30889 17267 30923
rect 17267 30889 17276 30923
rect 17224 30880 17276 30889
rect 18880 30880 18932 30932
rect 19340 30880 19392 30932
rect 20076 30880 20128 30932
rect 23756 30923 23808 30932
rect 23756 30889 23765 30923
rect 23765 30889 23799 30923
rect 23799 30889 23808 30923
rect 23756 30880 23808 30889
rect 24584 30923 24636 30932
rect 24584 30889 24593 30923
rect 24593 30889 24627 30923
rect 24627 30889 24636 30923
rect 24584 30880 24636 30889
rect 27528 30880 27580 30932
rect 28540 30880 28592 30932
rect 29736 30923 29788 30932
rect 29736 30889 29745 30923
rect 29745 30889 29779 30923
rect 29779 30889 29788 30923
rect 29736 30880 29788 30889
rect 35900 30923 35952 30932
rect 35900 30889 35909 30923
rect 35909 30889 35943 30923
rect 35943 30889 35952 30923
rect 35900 30880 35952 30889
rect 14740 30812 14792 30864
rect 17592 30812 17644 30864
rect 13176 30787 13228 30796
rect 13176 30753 13185 30787
rect 13185 30753 13219 30787
rect 13219 30753 13228 30787
rect 13176 30744 13228 30753
rect 18420 30744 18472 30796
rect 18604 30744 18656 30796
rect 20260 30787 20312 30796
rect 20260 30753 20269 30787
rect 20269 30753 20303 30787
rect 20303 30753 20312 30787
rect 21364 30787 21416 30796
rect 20260 30744 20312 30753
rect 21364 30753 21373 30787
rect 21373 30753 21407 30787
rect 21407 30753 21416 30787
rect 21364 30744 21416 30753
rect 23020 30787 23072 30796
rect 23020 30753 23029 30787
rect 23029 30753 23063 30787
rect 23063 30753 23072 30787
rect 23020 30744 23072 30753
rect 12072 30719 12124 30728
rect 12072 30685 12081 30719
rect 12081 30685 12115 30719
rect 12115 30685 12124 30719
rect 12072 30676 12124 30685
rect 15476 30676 15528 30728
rect 15568 30719 15620 30728
rect 15568 30685 15577 30719
rect 15577 30685 15611 30719
rect 15611 30685 15620 30719
rect 15568 30676 15620 30685
rect 21272 30676 21324 30728
rect 4068 30608 4120 30660
rect 9588 30608 9640 30660
rect 18328 30651 18380 30660
rect 18328 30617 18337 30651
rect 18337 30617 18371 30651
rect 18371 30617 18380 30651
rect 18328 30608 18380 30617
rect 6920 30583 6972 30592
rect 6920 30549 6929 30583
rect 6929 30549 6963 30583
rect 6963 30549 6972 30583
rect 6920 30540 6972 30549
rect 10416 30583 10468 30592
rect 10416 30549 10425 30583
rect 10425 30549 10459 30583
rect 10459 30549 10468 30583
rect 10416 30540 10468 30549
rect 12716 30540 12768 30592
rect 13360 30583 13412 30592
rect 13360 30549 13369 30583
rect 13369 30549 13403 30583
rect 13403 30549 13412 30583
rect 13360 30540 13412 30549
rect 23204 30540 23256 30592
rect 27344 30855 27396 30864
rect 27344 30821 27353 30855
rect 27353 30821 27387 30855
rect 27387 30821 27396 30855
rect 27344 30812 27396 30821
rect 25044 30787 25096 30796
rect 25044 30753 25053 30787
rect 25053 30753 25087 30787
rect 25087 30753 25096 30787
rect 25044 30744 25096 30753
rect 27252 30787 27304 30796
rect 24860 30719 24912 30728
rect 24860 30685 24869 30719
rect 24869 30685 24903 30719
rect 24903 30685 24912 30719
rect 24860 30676 24912 30685
rect 27252 30753 27261 30787
rect 27261 30753 27295 30787
rect 27295 30753 27304 30787
rect 27252 30744 27304 30753
rect 28816 30812 28868 30864
rect 25596 30719 25648 30728
rect 25596 30685 25605 30719
rect 25605 30685 25639 30719
rect 25639 30685 25648 30719
rect 25596 30676 25648 30685
rect 26976 30676 27028 30728
rect 26792 30608 26844 30660
rect 27528 30744 27580 30796
rect 30012 30787 30064 30796
rect 30012 30753 30021 30787
rect 30021 30753 30055 30787
rect 30055 30753 30064 30787
rect 30012 30744 30064 30753
rect 30748 30787 30800 30796
rect 30748 30753 30757 30787
rect 30757 30753 30791 30787
rect 30791 30753 30800 30787
rect 30748 30744 30800 30753
rect 31484 30787 31536 30796
rect 31484 30753 31493 30787
rect 31493 30753 31527 30787
rect 31527 30753 31536 30787
rect 31484 30744 31536 30753
rect 27804 30719 27856 30728
rect 27804 30685 27813 30719
rect 27813 30685 27847 30719
rect 27847 30685 27856 30719
rect 27804 30676 27856 30685
rect 26056 30540 26108 30592
rect 26700 30583 26752 30592
rect 26700 30549 26709 30583
rect 26709 30549 26743 30583
rect 26743 30549 26752 30583
rect 26700 30540 26752 30549
rect 29276 30583 29328 30592
rect 29276 30549 29285 30583
rect 29285 30549 29319 30583
rect 29319 30549 29328 30583
rect 29276 30540 29328 30549
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 3792 30336 3844 30388
rect 10324 30336 10376 30388
rect 12900 30336 12952 30388
rect 13452 30336 13504 30388
rect 14556 30379 14608 30388
rect 14556 30345 14565 30379
rect 14565 30345 14599 30379
rect 14599 30345 14608 30379
rect 14556 30336 14608 30345
rect 15568 30336 15620 30388
rect 17224 30336 17276 30388
rect 17592 30336 17644 30388
rect 18328 30379 18380 30388
rect 2780 30200 2832 30252
rect 3240 30132 3292 30184
rect 6920 30200 6972 30252
rect 4620 30132 4672 30184
rect 7380 30175 7432 30184
rect 7380 30141 7389 30175
rect 7389 30141 7423 30175
rect 7423 30141 7432 30175
rect 7380 30132 7432 30141
rect 7104 30064 7156 30116
rect 8024 30132 8076 30184
rect 9680 30268 9732 30320
rect 10508 30268 10560 30320
rect 12532 30311 12584 30320
rect 12532 30277 12541 30311
rect 12541 30277 12575 30311
rect 12575 30277 12584 30311
rect 13912 30311 13964 30320
rect 12532 30268 12584 30277
rect 13912 30277 13921 30311
rect 13921 30277 13955 30311
rect 13955 30277 13964 30311
rect 13912 30268 13964 30277
rect 10416 30175 10468 30184
rect 10416 30141 10425 30175
rect 10425 30141 10459 30175
rect 10459 30141 10468 30175
rect 10416 30132 10468 30141
rect 12072 30200 12124 30252
rect 13176 30200 13228 30252
rect 18328 30345 18337 30379
rect 18337 30345 18371 30379
rect 18371 30345 18380 30379
rect 18328 30336 18380 30345
rect 21272 30336 21324 30388
rect 28172 30336 28224 30388
rect 32128 30336 32180 30388
rect 18420 30268 18472 30320
rect 27160 30268 27212 30320
rect 27896 30268 27948 30320
rect 28356 30268 28408 30320
rect 28816 30311 28868 30320
rect 28816 30277 28825 30311
rect 28825 30277 28859 30311
rect 28859 30277 28868 30311
rect 28816 30268 28868 30277
rect 15292 30243 15344 30252
rect 11704 30132 11756 30184
rect 12716 30175 12768 30184
rect 12716 30141 12725 30175
rect 12725 30141 12759 30175
rect 12759 30141 12768 30175
rect 12716 30132 12768 30141
rect 14188 30175 14240 30184
rect 14188 30141 14197 30175
rect 14197 30141 14231 30175
rect 14231 30141 14240 30175
rect 14188 30132 14240 30141
rect 14740 30175 14792 30184
rect 14740 30141 14749 30175
rect 14749 30141 14783 30175
rect 14783 30141 14792 30175
rect 14740 30132 14792 30141
rect 15292 30209 15301 30243
rect 15301 30209 15335 30243
rect 15335 30209 15344 30243
rect 15292 30200 15344 30209
rect 18052 30243 18104 30252
rect 18052 30209 18061 30243
rect 18061 30209 18095 30243
rect 18095 30209 18104 30243
rect 18052 30200 18104 30209
rect 18604 30200 18656 30252
rect 19156 30200 19208 30252
rect 20168 30200 20220 30252
rect 21088 30243 21140 30252
rect 21088 30209 21097 30243
rect 21097 30209 21131 30243
rect 21131 30209 21140 30243
rect 21088 30200 21140 30209
rect 24860 30200 24912 30252
rect 26608 30200 26660 30252
rect 28264 30200 28316 30252
rect 29276 30200 29328 30252
rect 29736 30200 29788 30252
rect 35808 30268 35860 30320
rect 13268 30064 13320 30116
rect 16396 30064 16448 30116
rect 22284 30175 22336 30184
rect 22284 30141 22293 30175
rect 22293 30141 22327 30175
rect 22327 30141 22336 30175
rect 22284 30132 22336 30141
rect 22192 30064 22244 30116
rect 24216 30132 24268 30184
rect 25596 30132 25648 30184
rect 26148 30132 26200 30184
rect 27712 30132 27764 30184
rect 27896 30132 27948 30184
rect 29000 30175 29052 30184
rect 29000 30141 29009 30175
rect 29009 30141 29043 30175
rect 29043 30141 29052 30175
rect 29000 30132 29052 30141
rect 27528 30064 27580 30116
rect 29368 30064 29420 30116
rect 30012 30132 30064 30184
rect 32036 30132 32088 30184
rect 32864 30132 32916 30184
rect 32956 30132 33008 30184
rect 35900 30132 35952 30184
rect 33416 30064 33468 30116
rect 8576 29996 8628 30048
rect 11428 29996 11480 30048
rect 12164 30039 12216 30048
rect 12164 30005 12173 30039
rect 12173 30005 12207 30039
rect 12207 30005 12216 30039
rect 12164 29996 12216 30005
rect 17592 29996 17644 30048
rect 19340 30039 19392 30048
rect 19340 30005 19349 30039
rect 19349 30005 19383 30039
rect 19383 30005 19392 30039
rect 19340 29996 19392 30005
rect 22284 30039 22336 30048
rect 22284 30005 22293 30039
rect 22293 30005 22327 30039
rect 22327 30005 22336 30039
rect 22284 29996 22336 30005
rect 23480 30039 23532 30048
rect 23480 30005 23489 30039
rect 23489 30005 23523 30039
rect 23523 30005 23532 30039
rect 23480 29996 23532 30005
rect 24124 30039 24176 30048
rect 24124 30005 24133 30039
rect 24133 30005 24167 30039
rect 24167 30005 24176 30039
rect 24124 29996 24176 30005
rect 26424 30039 26476 30048
rect 26424 30005 26433 30039
rect 26433 30005 26467 30039
rect 26467 30005 26476 30039
rect 26424 29996 26476 30005
rect 27252 29996 27304 30048
rect 30748 30039 30800 30048
rect 30748 30005 30757 30039
rect 30757 30005 30791 30039
rect 30791 30005 30800 30039
rect 30748 29996 30800 30005
rect 37372 30039 37424 30048
rect 37372 30005 37381 30039
rect 37381 30005 37415 30039
rect 37415 30005 37424 30039
rect 37372 29996 37424 30005
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 3424 29835 3476 29844
rect 3424 29801 3433 29835
rect 3433 29801 3467 29835
rect 3467 29801 3476 29835
rect 3424 29792 3476 29801
rect 7380 29792 7432 29844
rect 12532 29835 12584 29844
rect 12532 29801 12541 29835
rect 12541 29801 12575 29835
rect 12575 29801 12584 29835
rect 12532 29792 12584 29801
rect 12716 29792 12768 29844
rect 14188 29792 14240 29844
rect 15476 29835 15528 29844
rect 15476 29801 15485 29835
rect 15485 29801 15519 29835
rect 15519 29801 15528 29835
rect 15476 29792 15528 29801
rect 17592 29835 17644 29844
rect 17592 29801 17601 29835
rect 17601 29801 17635 29835
rect 17635 29801 17644 29835
rect 17592 29792 17644 29801
rect 18328 29792 18380 29844
rect 18512 29835 18564 29844
rect 18512 29801 18521 29835
rect 18521 29801 18555 29835
rect 18555 29801 18564 29835
rect 18512 29792 18564 29801
rect 19156 29835 19208 29844
rect 19156 29801 19165 29835
rect 19165 29801 19199 29835
rect 19199 29801 19208 29835
rect 19156 29792 19208 29801
rect 21364 29835 21416 29844
rect 21364 29801 21373 29835
rect 21373 29801 21407 29835
rect 21407 29801 21416 29835
rect 21364 29792 21416 29801
rect 22192 29792 22244 29844
rect 23296 29792 23348 29844
rect 24216 29835 24268 29844
rect 12164 29724 12216 29776
rect 13176 29724 13228 29776
rect 1676 29699 1728 29708
rect 1676 29665 1685 29699
rect 1685 29665 1719 29699
rect 1719 29665 1728 29699
rect 1676 29656 1728 29665
rect 7564 29699 7616 29708
rect 7564 29665 7573 29699
rect 7573 29665 7607 29699
rect 7607 29665 7616 29699
rect 7564 29656 7616 29665
rect 8024 29656 8076 29708
rect 10324 29656 10376 29708
rect 10416 29656 10468 29708
rect 11428 29699 11480 29708
rect 11428 29665 11437 29699
rect 11437 29665 11471 29699
rect 11471 29665 11480 29699
rect 11428 29656 11480 29665
rect 11704 29699 11756 29708
rect 11704 29665 11713 29699
rect 11713 29665 11747 29699
rect 11747 29665 11756 29699
rect 13636 29699 13688 29708
rect 11704 29656 11756 29665
rect 13636 29665 13645 29699
rect 13645 29665 13679 29699
rect 13679 29665 13688 29699
rect 13636 29656 13688 29665
rect 16304 29656 16356 29708
rect 19892 29699 19944 29708
rect 19892 29665 19901 29699
rect 19901 29665 19935 29699
rect 19935 29665 19944 29699
rect 19892 29656 19944 29665
rect 22560 29699 22612 29708
rect 22560 29665 22569 29699
rect 22569 29665 22603 29699
rect 22603 29665 22612 29699
rect 22560 29656 22612 29665
rect 22744 29656 22796 29708
rect 23204 29656 23256 29708
rect 2044 29588 2096 29640
rect 7196 29631 7248 29640
rect 7196 29597 7205 29631
rect 7205 29597 7239 29631
rect 7239 29597 7248 29631
rect 7196 29588 7248 29597
rect 10600 29631 10652 29640
rect 7840 29563 7892 29572
rect 7840 29529 7849 29563
rect 7849 29529 7883 29563
rect 7883 29529 7892 29563
rect 7840 29520 7892 29529
rect 10600 29597 10609 29631
rect 10609 29597 10643 29631
rect 10643 29597 10652 29631
rect 10600 29588 10652 29597
rect 11244 29588 11296 29640
rect 15476 29588 15528 29640
rect 20352 29588 20404 29640
rect 22284 29588 22336 29640
rect 10140 29520 10192 29572
rect 12072 29520 12124 29572
rect 22836 29588 22888 29640
rect 23664 29656 23716 29708
rect 24216 29801 24225 29835
rect 24225 29801 24259 29835
rect 24259 29801 24268 29835
rect 24216 29792 24268 29801
rect 27804 29835 27856 29844
rect 27804 29801 27813 29835
rect 27813 29801 27847 29835
rect 27847 29801 27856 29835
rect 27804 29792 27856 29801
rect 28264 29835 28316 29844
rect 28264 29801 28273 29835
rect 28273 29801 28307 29835
rect 28307 29801 28316 29835
rect 28264 29792 28316 29801
rect 29736 29835 29788 29844
rect 29736 29801 29745 29835
rect 29745 29801 29779 29835
rect 29779 29801 29788 29835
rect 29736 29792 29788 29801
rect 31760 29792 31812 29844
rect 32956 29792 33008 29844
rect 26516 29699 26568 29708
rect 26516 29665 26525 29699
rect 26525 29665 26559 29699
rect 26559 29665 26568 29699
rect 26516 29656 26568 29665
rect 28264 29699 28316 29708
rect 28264 29665 28273 29699
rect 28273 29665 28307 29699
rect 28307 29665 28316 29699
rect 28264 29656 28316 29665
rect 23480 29588 23532 29640
rect 24584 29588 24636 29640
rect 24768 29588 24820 29640
rect 27988 29588 28040 29640
rect 29736 29656 29788 29708
rect 30472 29699 30524 29708
rect 29276 29588 29328 29640
rect 29920 29631 29972 29640
rect 29920 29597 29929 29631
rect 29929 29597 29963 29631
rect 29963 29597 29972 29631
rect 29920 29588 29972 29597
rect 30472 29665 30481 29699
rect 30481 29665 30515 29699
rect 30515 29665 30524 29699
rect 30472 29656 30524 29665
rect 33692 29656 33744 29708
rect 36544 29656 36596 29708
rect 32956 29588 33008 29640
rect 33968 29588 34020 29640
rect 34152 29631 34204 29640
rect 34152 29597 34161 29631
rect 34161 29597 34195 29631
rect 34195 29597 34204 29631
rect 34152 29588 34204 29597
rect 34336 29588 34388 29640
rect 25136 29520 25188 29572
rect 26056 29520 26108 29572
rect 27436 29563 27488 29572
rect 27436 29529 27445 29563
rect 27445 29529 27479 29563
rect 27479 29529 27488 29563
rect 27436 29520 27488 29529
rect 2780 29495 2832 29504
rect 2780 29461 2789 29495
rect 2789 29461 2823 29495
rect 2823 29461 2832 29495
rect 8576 29495 8628 29504
rect 2780 29452 2832 29461
rect 8576 29461 8585 29495
rect 8585 29461 8619 29495
rect 8619 29461 8628 29495
rect 8576 29452 8628 29461
rect 11704 29452 11756 29504
rect 12716 29452 12768 29504
rect 21272 29452 21324 29504
rect 22928 29452 22980 29504
rect 23296 29452 23348 29504
rect 26148 29495 26200 29504
rect 26148 29461 26157 29495
rect 26157 29461 26191 29495
rect 26191 29461 26200 29495
rect 26148 29452 26200 29461
rect 26332 29452 26384 29504
rect 26976 29452 27028 29504
rect 29460 29495 29512 29504
rect 29460 29461 29469 29495
rect 29469 29461 29503 29495
rect 29503 29461 29512 29495
rect 29460 29452 29512 29461
rect 31208 29495 31260 29504
rect 31208 29461 31217 29495
rect 31217 29461 31251 29495
rect 31251 29461 31260 29495
rect 31208 29452 31260 29461
rect 35900 29495 35952 29504
rect 35900 29461 35909 29495
rect 35909 29461 35943 29495
rect 35943 29461 35952 29495
rect 35900 29452 35952 29461
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 1676 29291 1728 29300
rect 1676 29257 1685 29291
rect 1685 29257 1719 29291
rect 1719 29257 1728 29291
rect 1676 29248 1728 29257
rect 4896 29291 4948 29300
rect 4896 29257 4905 29291
rect 4905 29257 4939 29291
rect 4939 29257 4948 29291
rect 4896 29248 4948 29257
rect 8024 29248 8076 29300
rect 10140 29291 10192 29300
rect 10140 29257 10149 29291
rect 10149 29257 10183 29291
rect 10183 29257 10192 29291
rect 10140 29248 10192 29257
rect 11244 29291 11296 29300
rect 11244 29257 11253 29291
rect 11253 29257 11287 29291
rect 11287 29257 11296 29291
rect 11244 29248 11296 29257
rect 12164 29291 12216 29300
rect 12164 29257 12173 29291
rect 12173 29257 12207 29291
rect 12207 29257 12216 29291
rect 12164 29248 12216 29257
rect 13268 29291 13320 29300
rect 13268 29257 13277 29291
rect 13277 29257 13311 29291
rect 13311 29257 13320 29291
rect 13268 29248 13320 29257
rect 15200 29291 15252 29300
rect 15200 29257 15209 29291
rect 15209 29257 15243 29291
rect 15243 29257 15252 29291
rect 15200 29248 15252 29257
rect 16304 29291 16356 29300
rect 16304 29257 16313 29291
rect 16313 29257 16347 29291
rect 16347 29257 16356 29291
rect 16304 29248 16356 29257
rect 22744 29248 22796 29300
rect 23480 29291 23532 29300
rect 23480 29257 23489 29291
rect 23489 29257 23523 29291
rect 23523 29257 23532 29291
rect 23480 29248 23532 29257
rect 27988 29291 28040 29300
rect 27988 29257 27997 29291
rect 27997 29257 28031 29291
rect 28031 29257 28040 29291
rect 27988 29248 28040 29257
rect 28908 29291 28960 29300
rect 28908 29257 28917 29291
rect 28917 29257 28951 29291
rect 28951 29257 28960 29291
rect 28908 29248 28960 29257
rect 33692 29291 33744 29300
rect 33692 29257 33701 29291
rect 33701 29257 33735 29291
rect 33735 29257 33744 29291
rect 33692 29248 33744 29257
rect 33968 29291 34020 29300
rect 33968 29257 33977 29291
rect 33977 29257 34011 29291
rect 34011 29257 34020 29291
rect 33968 29248 34020 29257
rect 34336 29291 34388 29300
rect 34336 29257 34345 29291
rect 34345 29257 34379 29291
rect 34379 29257 34388 29291
rect 34336 29248 34388 29257
rect 36544 29291 36596 29300
rect 36544 29257 36553 29291
rect 36553 29257 36587 29291
rect 36587 29257 36596 29291
rect 36544 29248 36596 29257
rect 2044 29155 2096 29164
rect 2044 29121 2053 29155
rect 2053 29121 2087 29155
rect 2087 29121 2096 29155
rect 3332 29155 3384 29164
rect 2044 29112 2096 29121
rect 3332 29121 3341 29155
rect 3341 29121 3375 29155
rect 3375 29121 3384 29155
rect 3332 29112 3384 29121
rect 3148 29019 3200 29028
rect 3148 28985 3157 29019
rect 3157 28985 3191 29019
rect 3191 28985 3200 29019
rect 8576 29087 8628 29096
rect 8576 29053 8585 29087
rect 8585 29053 8619 29087
rect 8619 29053 8628 29087
rect 8576 29044 8628 29053
rect 8944 29044 8996 29096
rect 11520 29223 11572 29232
rect 11520 29189 11529 29223
rect 11529 29189 11563 29223
rect 11563 29189 11572 29223
rect 11520 29180 11572 29189
rect 21180 29223 21232 29232
rect 21180 29189 21189 29223
rect 21189 29189 21223 29223
rect 21223 29189 21232 29223
rect 21180 29180 21232 29189
rect 24860 29180 24912 29232
rect 28172 29180 28224 29232
rect 18604 29112 18656 29164
rect 13452 29044 13504 29096
rect 13912 29044 13964 29096
rect 14096 29087 14148 29096
rect 14096 29053 14105 29087
rect 14105 29053 14139 29087
rect 14139 29053 14148 29087
rect 14096 29044 14148 29053
rect 14464 29044 14516 29096
rect 15752 29044 15804 29096
rect 3148 28976 3200 28985
rect 7196 28976 7248 29028
rect 7564 28976 7616 29028
rect 10416 28976 10468 29028
rect 12072 28976 12124 29028
rect 12348 28976 12400 29028
rect 13636 28976 13688 29028
rect 15108 28976 15160 29028
rect 15844 28976 15896 29028
rect 16028 28976 16080 29028
rect 16304 28976 16356 29028
rect 19248 29044 19300 29096
rect 20352 29087 20404 29096
rect 20352 29053 20361 29087
rect 20361 29053 20395 29087
rect 20395 29053 20404 29087
rect 20352 29044 20404 29053
rect 21456 29112 21508 29164
rect 21824 29112 21876 29164
rect 24124 29112 24176 29164
rect 25044 29112 25096 29164
rect 21272 29087 21324 29096
rect 21272 29053 21281 29087
rect 21281 29053 21315 29087
rect 21315 29053 21324 29087
rect 21272 29044 21324 29053
rect 24860 29087 24912 29096
rect 24860 29053 24869 29087
rect 24869 29053 24903 29087
rect 24903 29053 24912 29087
rect 24860 29044 24912 29053
rect 24952 29044 25004 29096
rect 26056 29044 26108 29096
rect 26516 29112 26568 29164
rect 27804 29112 27856 29164
rect 29276 29155 29328 29164
rect 29276 29121 29285 29155
rect 29285 29121 29319 29155
rect 29319 29121 29328 29155
rect 29276 29112 29328 29121
rect 27436 29087 27488 29096
rect 7748 28908 7800 28960
rect 9588 28908 9640 28960
rect 12900 28908 12952 28960
rect 17500 28908 17552 28960
rect 19248 28908 19300 28960
rect 23112 28976 23164 29028
rect 24032 28976 24084 29028
rect 24768 28976 24820 29028
rect 25044 29019 25096 29028
rect 25044 28985 25053 29019
rect 25053 28985 25087 29019
rect 25087 28985 25096 29019
rect 25044 28976 25096 28985
rect 25228 29019 25280 29028
rect 25228 28985 25237 29019
rect 25237 28985 25271 29019
rect 25271 28985 25280 29019
rect 25228 28976 25280 28985
rect 27436 29053 27445 29087
rect 27445 29053 27479 29087
rect 27479 29053 27488 29087
rect 27436 29044 27488 29053
rect 29184 29044 29236 29096
rect 29920 29180 29972 29232
rect 29460 29112 29512 29164
rect 30380 29112 30432 29164
rect 30104 29087 30156 29096
rect 30104 29053 30113 29087
rect 30113 29053 30147 29087
rect 30147 29053 30156 29087
rect 30104 29044 30156 29053
rect 26700 28976 26752 29028
rect 27160 28976 27212 29028
rect 31300 29155 31352 29164
rect 31300 29121 31309 29155
rect 31309 29121 31343 29155
rect 31343 29121 31352 29155
rect 31300 29112 31352 29121
rect 35440 29155 35492 29164
rect 35440 29121 35449 29155
rect 35449 29121 35483 29155
rect 35483 29121 35492 29155
rect 35440 29112 35492 29121
rect 31208 29087 31260 29096
rect 31208 29053 31217 29087
rect 31217 29053 31251 29087
rect 31251 29053 31260 29087
rect 31208 29044 31260 29053
rect 31760 29044 31812 29096
rect 32220 29044 32272 29096
rect 35900 29044 35952 29096
rect 22744 28908 22796 28960
rect 25136 28951 25188 28960
rect 25136 28917 25145 28951
rect 25145 28917 25179 28951
rect 25179 28917 25188 28951
rect 25136 28908 25188 28917
rect 26424 28908 26476 28960
rect 28908 28951 28960 28960
rect 28908 28917 28917 28951
rect 28917 28917 28951 28951
rect 28951 28917 28960 28951
rect 28908 28908 28960 28917
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 3976 28704 4028 28756
rect 4988 28704 5040 28756
rect 11704 28704 11756 28756
rect 14372 28704 14424 28756
rect 16672 28747 16724 28756
rect 16672 28713 16681 28747
rect 16681 28713 16715 28747
rect 16715 28713 16724 28747
rect 16672 28704 16724 28713
rect 19340 28747 19392 28756
rect 19340 28713 19349 28747
rect 19349 28713 19383 28747
rect 19383 28713 19392 28747
rect 19340 28704 19392 28713
rect 20352 28747 20404 28756
rect 20352 28713 20361 28747
rect 20361 28713 20395 28747
rect 20395 28713 20404 28747
rect 20352 28704 20404 28713
rect 26240 28747 26292 28756
rect 26240 28713 26249 28747
rect 26249 28713 26283 28747
rect 26283 28713 26292 28747
rect 26240 28704 26292 28713
rect 28264 28704 28316 28756
rect 30380 28704 30432 28756
rect 31208 28704 31260 28756
rect 35440 28704 35492 28756
rect 26608 28636 26660 28688
rect 26884 28679 26936 28688
rect 26884 28645 26893 28679
rect 26893 28645 26927 28679
rect 26927 28645 26936 28679
rect 26884 28636 26936 28645
rect 30564 28636 30616 28688
rect 31852 28636 31904 28688
rect 1400 28568 1452 28620
rect 2044 28568 2096 28620
rect 4712 28611 4764 28620
rect 4712 28577 4721 28611
rect 4721 28577 4755 28611
rect 4755 28577 4764 28611
rect 4712 28568 4764 28577
rect 5356 28568 5408 28620
rect 7012 28611 7064 28620
rect 7012 28577 7021 28611
rect 7021 28577 7055 28611
rect 7055 28577 7064 28611
rect 7012 28568 7064 28577
rect 7840 28568 7892 28620
rect 8668 28611 8720 28620
rect 8668 28577 8677 28611
rect 8677 28577 8711 28611
rect 8711 28577 8720 28611
rect 8668 28568 8720 28577
rect 10600 28611 10652 28620
rect 10600 28577 10609 28611
rect 10609 28577 10643 28611
rect 10643 28577 10652 28611
rect 10600 28568 10652 28577
rect 10876 28568 10928 28620
rect 12900 28611 12952 28620
rect 12900 28577 12909 28611
rect 12909 28577 12943 28611
rect 12943 28577 12952 28611
rect 12900 28568 12952 28577
rect 13820 28611 13872 28620
rect 13820 28577 13829 28611
rect 13829 28577 13863 28611
rect 13863 28577 13872 28611
rect 13820 28568 13872 28577
rect 15384 28568 15436 28620
rect 22192 28611 22244 28620
rect 22192 28577 22201 28611
rect 22201 28577 22235 28611
rect 22235 28577 22244 28611
rect 22192 28568 22244 28577
rect 22928 28611 22980 28620
rect 22928 28577 22937 28611
rect 22937 28577 22971 28611
rect 22971 28577 22980 28611
rect 22928 28568 22980 28577
rect 24952 28611 25004 28620
rect 24952 28577 24961 28611
rect 24961 28577 24995 28611
rect 24995 28577 25004 28611
rect 24952 28568 25004 28577
rect 25320 28611 25372 28620
rect 25320 28577 25329 28611
rect 25329 28577 25363 28611
rect 25363 28577 25372 28611
rect 25320 28568 25372 28577
rect 25412 28611 25464 28620
rect 25412 28577 25421 28611
rect 25421 28577 25455 28611
rect 25455 28577 25464 28611
rect 25412 28568 25464 28577
rect 26424 28568 26476 28620
rect 28172 28568 28224 28620
rect 28632 28611 28684 28620
rect 28632 28577 28641 28611
rect 28641 28577 28675 28611
rect 28675 28577 28684 28611
rect 28632 28568 28684 28577
rect 28724 28568 28776 28620
rect 30288 28611 30340 28620
rect 30288 28577 30297 28611
rect 30297 28577 30331 28611
rect 30331 28577 30340 28611
rect 30288 28568 30340 28577
rect 33784 28611 33836 28620
rect 7104 28543 7156 28552
rect 7104 28509 7113 28543
rect 7113 28509 7147 28543
rect 7147 28509 7156 28543
rect 7104 28500 7156 28509
rect 8024 28543 8076 28552
rect 8024 28509 8033 28543
rect 8033 28509 8067 28543
rect 8067 28509 8076 28543
rect 8024 28500 8076 28509
rect 11244 28500 11296 28552
rect 13268 28500 13320 28552
rect 13912 28500 13964 28552
rect 15476 28500 15528 28552
rect 17500 28500 17552 28552
rect 18052 28543 18104 28552
rect 18052 28509 18061 28543
rect 18061 28509 18095 28543
rect 18095 28509 18104 28543
rect 18052 28500 18104 28509
rect 22100 28543 22152 28552
rect 22100 28509 22109 28543
rect 22109 28509 22143 28543
rect 22143 28509 22152 28543
rect 22100 28500 22152 28509
rect 22744 28500 22796 28552
rect 23020 28543 23072 28552
rect 23020 28509 23029 28543
rect 23029 28509 23063 28543
rect 23063 28509 23072 28543
rect 23020 28500 23072 28509
rect 24216 28500 24268 28552
rect 26332 28500 26384 28552
rect 26884 28500 26936 28552
rect 10416 28475 10468 28484
rect 10416 28441 10425 28475
rect 10425 28441 10459 28475
rect 10459 28441 10468 28475
rect 10416 28432 10468 28441
rect 33784 28577 33793 28611
rect 33793 28577 33827 28611
rect 33827 28577 33836 28611
rect 33784 28568 33836 28577
rect 34796 28568 34848 28620
rect 33692 28543 33744 28552
rect 33692 28509 33701 28543
rect 33701 28509 33735 28543
rect 33735 28509 33744 28543
rect 33692 28500 33744 28509
rect 31668 28432 31720 28484
rect 33140 28432 33192 28484
rect 3056 28407 3108 28416
rect 3056 28373 3065 28407
rect 3065 28373 3099 28407
rect 3099 28373 3108 28407
rect 3056 28364 3108 28373
rect 6092 28407 6144 28416
rect 6092 28373 6101 28407
rect 6101 28373 6135 28407
rect 6135 28373 6144 28407
rect 6092 28364 6144 28373
rect 9036 28364 9088 28416
rect 9404 28364 9456 28416
rect 14004 28407 14056 28416
rect 14004 28373 14013 28407
rect 14013 28373 14047 28407
rect 14047 28373 14056 28407
rect 14004 28364 14056 28373
rect 19800 28407 19852 28416
rect 19800 28373 19809 28407
rect 19809 28373 19843 28407
rect 19843 28373 19852 28407
rect 19800 28364 19852 28373
rect 27344 28364 27396 28416
rect 30840 28364 30892 28416
rect 31208 28407 31260 28416
rect 31208 28373 31217 28407
rect 31217 28373 31251 28407
rect 31251 28373 31260 28407
rect 31208 28364 31260 28373
rect 32220 28364 32272 28416
rect 33232 28407 33284 28416
rect 33232 28373 33241 28407
rect 33241 28373 33275 28407
rect 33275 28373 33284 28407
rect 33232 28364 33284 28373
rect 35808 28407 35860 28416
rect 35808 28373 35817 28407
rect 35817 28373 35851 28407
rect 35851 28373 35860 28407
rect 35808 28364 35860 28373
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 1400 28160 1452 28212
rect 2044 28203 2096 28212
rect 2044 28169 2053 28203
rect 2053 28169 2087 28203
rect 2087 28169 2096 28203
rect 2044 28160 2096 28169
rect 3700 28160 3752 28212
rect 4712 28203 4764 28212
rect 4712 28169 4721 28203
rect 4721 28169 4755 28203
rect 4755 28169 4764 28203
rect 4712 28160 4764 28169
rect 7012 28160 7064 28212
rect 8668 28160 8720 28212
rect 10600 28203 10652 28212
rect 10600 28169 10609 28203
rect 10609 28169 10643 28203
rect 10643 28169 10652 28203
rect 10600 28160 10652 28169
rect 11244 28203 11296 28212
rect 11244 28169 11253 28203
rect 11253 28169 11287 28203
rect 11287 28169 11296 28203
rect 11244 28160 11296 28169
rect 11704 28160 11756 28212
rect 23204 28160 23256 28212
rect 25412 28160 25464 28212
rect 28172 28203 28224 28212
rect 28172 28169 28181 28203
rect 28181 28169 28215 28203
rect 28215 28169 28224 28203
rect 28172 28160 28224 28169
rect 28264 28160 28316 28212
rect 28724 28160 28776 28212
rect 31668 28203 31720 28212
rect 31668 28169 31677 28203
rect 31677 28169 31711 28203
rect 31711 28169 31720 28203
rect 31668 28160 31720 28169
rect 31760 28160 31812 28212
rect 7104 28092 7156 28144
rect 9772 28092 9824 28144
rect 10876 28092 10928 28144
rect 19064 28135 19116 28144
rect 8944 28067 8996 28076
rect 8944 28033 8953 28067
rect 8953 28033 8987 28067
rect 8987 28033 8996 28067
rect 8944 28024 8996 28033
rect 11244 28024 11296 28076
rect 7472 27999 7524 28008
rect 7472 27965 7481 27999
rect 7481 27965 7515 27999
rect 7515 27965 7524 27999
rect 7472 27956 7524 27965
rect 8024 27956 8076 28008
rect 8852 27999 8904 28008
rect 8852 27965 8861 27999
rect 8861 27965 8895 27999
rect 8895 27965 8904 27999
rect 8852 27956 8904 27965
rect 9772 27999 9824 28008
rect 9772 27965 9781 27999
rect 9781 27965 9815 27999
rect 9815 27965 9824 27999
rect 9772 27956 9824 27965
rect 10232 27956 10284 28008
rect 14372 28067 14424 28076
rect 14372 28033 14381 28067
rect 14381 28033 14415 28067
rect 14415 28033 14424 28067
rect 14372 28024 14424 28033
rect 19064 28101 19073 28135
rect 19073 28101 19107 28135
rect 19107 28101 19116 28135
rect 19064 28092 19116 28101
rect 19432 28092 19484 28144
rect 22008 28092 22060 28144
rect 27620 28092 27672 28144
rect 30288 28135 30340 28144
rect 30288 28101 30297 28135
rect 30297 28101 30331 28135
rect 30331 28101 30340 28135
rect 30288 28092 30340 28101
rect 30748 28092 30800 28144
rect 13452 27999 13504 28008
rect 13452 27965 13461 27999
rect 13461 27965 13495 27999
rect 13495 27965 13504 27999
rect 13452 27956 13504 27965
rect 13636 27956 13688 28008
rect 14188 27956 14240 28008
rect 19248 27999 19300 28008
rect 19248 27965 19257 27999
rect 19257 27965 19291 27999
rect 19291 27965 19300 27999
rect 19248 27956 19300 27965
rect 5356 27863 5408 27872
rect 5356 27829 5365 27863
rect 5365 27829 5399 27863
rect 5399 27829 5408 27863
rect 5356 27820 5408 27829
rect 7656 27863 7708 27872
rect 7656 27829 7665 27863
rect 7665 27829 7699 27863
rect 7699 27829 7708 27863
rect 7656 27820 7708 27829
rect 8392 27820 8444 27872
rect 12900 27888 12952 27940
rect 13360 27888 13412 27940
rect 16856 27888 16908 27940
rect 18052 27888 18104 27940
rect 19892 27956 19944 28008
rect 21088 27956 21140 28008
rect 23020 28024 23072 28076
rect 24860 28024 24912 28076
rect 24216 27999 24268 28008
rect 21272 27888 21324 27940
rect 21364 27888 21416 27940
rect 23480 27931 23532 27940
rect 23480 27897 23489 27931
rect 23489 27897 23523 27931
rect 23523 27897 23532 27931
rect 24216 27965 24225 27999
rect 24225 27965 24259 27999
rect 24259 27965 24268 27999
rect 24216 27956 24268 27965
rect 23480 27888 23532 27897
rect 25412 27956 25464 28008
rect 26424 27956 26476 28008
rect 27344 27999 27396 28008
rect 27344 27965 27353 27999
rect 27353 27965 27387 27999
rect 27387 27965 27396 27999
rect 27344 27956 27396 27965
rect 27712 27956 27764 28008
rect 28172 27956 28224 28008
rect 28816 27956 28868 28008
rect 29644 27956 29696 28008
rect 30472 27999 30524 28008
rect 30472 27965 30481 27999
rect 30481 27965 30515 27999
rect 30515 27965 30524 27999
rect 30472 27956 30524 27965
rect 30564 27956 30616 28008
rect 30840 27999 30892 28008
rect 30840 27965 30849 27999
rect 30849 27965 30883 27999
rect 30883 27965 30892 27999
rect 30840 27956 30892 27965
rect 31116 27956 31168 28008
rect 34796 28160 34848 28212
rect 33784 28024 33836 28076
rect 36084 28067 36136 28076
rect 36084 28033 36093 28067
rect 36093 28033 36127 28067
rect 36127 28033 36136 28067
rect 36084 28024 36136 28033
rect 32680 27999 32732 28008
rect 32680 27965 32689 27999
rect 32689 27965 32723 27999
rect 32723 27965 32732 27999
rect 32680 27956 32732 27965
rect 33140 27999 33192 28008
rect 33140 27965 33149 27999
rect 33149 27965 33183 27999
rect 33183 27965 33192 27999
rect 33140 27956 33192 27965
rect 35808 27999 35860 28008
rect 35808 27965 35817 27999
rect 35817 27965 35851 27999
rect 35851 27965 35860 27999
rect 35808 27956 35860 27965
rect 25504 27888 25556 27940
rect 10968 27863 11020 27872
rect 10968 27829 10977 27863
rect 10977 27829 11011 27863
rect 11011 27829 11020 27863
rect 10968 27820 11020 27829
rect 15384 27863 15436 27872
rect 15384 27829 15393 27863
rect 15393 27829 15427 27863
rect 15427 27829 15436 27863
rect 15384 27820 15436 27829
rect 15476 27820 15528 27872
rect 16304 27820 16356 27872
rect 17500 27863 17552 27872
rect 17500 27829 17509 27863
rect 17509 27829 17543 27863
rect 17543 27829 17552 27863
rect 17500 27820 17552 27829
rect 22100 27820 22152 27872
rect 23756 27863 23808 27872
rect 23756 27829 23765 27863
rect 23765 27829 23799 27863
rect 23799 27829 23808 27863
rect 23756 27820 23808 27829
rect 25320 27820 25372 27872
rect 26332 27820 26384 27872
rect 27252 27888 27304 27940
rect 28632 27888 28684 27940
rect 30104 27888 30156 27940
rect 33692 27863 33744 27872
rect 33692 27829 33701 27863
rect 33701 27829 33735 27863
rect 33735 27829 33744 27863
rect 33692 27820 33744 27829
rect 37372 27863 37424 27872
rect 37372 27829 37381 27863
rect 37381 27829 37415 27863
rect 37415 27829 37424 27863
rect 37372 27820 37424 27829
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 7472 27659 7524 27668
rect 7472 27625 7481 27659
rect 7481 27625 7515 27659
rect 7515 27625 7524 27659
rect 7472 27616 7524 27625
rect 8852 27659 8904 27668
rect 6092 27548 6144 27600
rect 8852 27625 8861 27659
rect 8861 27625 8895 27659
rect 8895 27625 8904 27659
rect 8852 27616 8904 27625
rect 14188 27659 14240 27668
rect 14188 27625 14197 27659
rect 14197 27625 14231 27659
rect 14231 27625 14240 27659
rect 14188 27616 14240 27625
rect 20352 27616 20404 27668
rect 21364 27616 21416 27668
rect 21732 27616 21784 27668
rect 22008 27616 22060 27668
rect 22928 27616 22980 27668
rect 1492 27480 1544 27532
rect 5724 27523 5776 27532
rect 5724 27489 5733 27523
rect 5733 27489 5767 27523
rect 5767 27489 5776 27523
rect 5724 27480 5776 27489
rect 5816 27480 5868 27532
rect 6644 27523 6696 27532
rect 6644 27489 6653 27523
rect 6653 27489 6687 27523
rect 6687 27489 6696 27523
rect 6644 27480 6696 27489
rect 12348 27548 12400 27600
rect 13820 27591 13872 27600
rect 13820 27557 13829 27591
rect 13829 27557 13863 27591
rect 13863 27557 13872 27591
rect 13820 27548 13872 27557
rect 8024 27523 8076 27532
rect 2044 27412 2096 27464
rect 3056 27455 3108 27464
rect 3056 27421 3065 27455
rect 3065 27421 3099 27455
rect 3099 27421 3108 27455
rect 3056 27412 3108 27421
rect 8024 27489 8033 27523
rect 8033 27489 8067 27523
rect 8067 27489 8076 27523
rect 8024 27480 8076 27489
rect 8116 27480 8168 27532
rect 11060 27523 11112 27532
rect 11060 27489 11069 27523
rect 11069 27489 11103 27523
rect 11103 27489 11112 27523
rect 11060 27480 11112 27489
rect 11520 27480 11572 27532
rect 13360 27523 13412 27532
rect 13360 27489 13369 27523
rect 13369 27489 13403 27523
rect 13403 27489 13412 27523
rect 13360 27480 13412 27489
rect 15292 27523 15344 27532
rect 15292 27489 15301 27523
rect 15301 27489 15335 27523
rect 15335 27489 15344 27523
rect 15292 27480 15344 27489
rect 16396 27480 16448 27532
rect 17040 27480 17092 27532
rect 17684 27480 17736 27532
rect 18696 27480 18748 27532
rect 22836 27523 22888 27532
rect 22836 27489 22845 27523
rect 22845 27489 22879 27523
rect 22879 27489 22888 27523
rect 23480 27616 23532 27668
rect 23940 27591 23992 27600
rect 23940 27557 23949 27591
rect 23949 27557 23983 27591
rect 23983 27557 23992 27591
rect 23940 27548 23992 27557
rect 27252 27616 27304 27668
rect 27712 27659 27764 27668
rect 27712 27625 27721 27659
rect 27721 27625 27755 27659
rect 27755 27625 27764 27659
rect 27712 27616 27764 27625
rect 28264 27616 28316 27668
rect 28632 27616 28684 27668
rect 29000 27616 29052 27668
rect 29368 27616 29420 27668
rect 29644 27659 29696 27668
rect 29644 27625 29653 27659
rect 29653 27625 29687 27659
rect 29687 27625 29696 27659
rect 29644 27616 29696 27625
rect 22836 27480 22888 27489
rect 23756 27480 23808 27532
rect 24676 27523 24728 27532
rect 24676 27489 24685 27523
rect 24685 27489 24719 27523
rect 24719 27489 24728 27523
rect 24676 27480 24728 27489
rect 26608 27480 26660 27532
rect 11704 27412 11756 27464
rect 16304 27455 16356 27464
rect 16304 27421 16313 27455
rect 16313 27421 16347 27455
rect 16347 27421 16356 27455
rect 16304 27412 16356 27421
rect 17500 27412 17552 27464
rect 22192 27455 22244 27464
rect 22192 27421 22201 27455
rect 22201 27421 22235 27455
rect 22235 27421 22244 27455
rect 22192 27412 22244 27421
rect 24768 27455 24820 27464
rect 24768 27421 24777 27455
rect 24777 27421 24811 27455
rect 24811 27421 24820 27455
rect 24768 27412 24820 27421
rect 3424 27319 3476 27328
rect 3424 27285 3433 27319
rect 3433 27285 3467 27319
rect 3467 27285 3476 27319
rect 3424 27276 3476 27285
rect 4896 27276 4948 27328
rect 10508 27344 10560 27396
rect 18604 27344 18656 27396
rect 18880 27344 18932 27396
rect 26792 27344 26844 27396
rect 8208 27276 8260 27328
rect 9312 27319 9364 27328
rect 9312 27285 9321 27319
rect 9321 27285 9355 27319
rect 9355 27285 9364 27319
rect 9312 27276 9364 27285
rect 10324 27319 10376 27328
rect 10324 27285 10333 27319
rect 10333 27285 10367 27319
rect 10367 27285 10376 27319
rect 10324 27276 10376 27285
rect 10784 27319 10836 27328
rect 10784 27285 10793 27319
rect 10793 27285 10827 27319
rect 10827 27285 10836 27319
rect 10784 27276 10836 27285
rect 11704 27276 11756 27328
rect 12072 27319 12124 27328
rect 12072 27285 12081 27319
rect 12081 27285 12115 27319
rect 12115 27285 12124 27319
rect 12072 27276 12124 27285
rect 13544 27319 13596 27328
rect 13544 27285 13553 27319
rect 13553 27285 13587 27319
rect 13587 27285 13596 27319
rect 13544 27276 13596 27285
rect 15476 27319 15528 27328
rect 15476 27285 15485 27319
rect 15485 27285 15519 27319
rect 15519 27285 15528 27319
rect 15476 27276 15528 27285
rect 17684 27319 17736 27328
rect 17684 27285 17693 27319
rect 17693 27285 17727 27319
rect 17727 27285 17736 27319
rect 17684 27276 17736 27285
rect 19340 27319 19392 27328
rect 19340 27285 19349 27319
rect 19349 27285 19383 27319
rect 19383 27285 19392 27319
rect 19340 27276 19392 27285
rect 25412 27319 25464 27328
rect 25412 27285 25421 27319
rect 25421 27285 25455 27319
rect 25455 27285 25464 27319
rect 25412 27276 25464 27285
rect 26424 27276 26476 27328
rect 26976 27344 27028 27396
rect 32680 27591 32732 27600
rect 32680 27557 32689 27591
rect 32689 27557 32723 27591
rect 32723 27557 32732 27591
rect 32680 27548 32732 27557
rect 33600 27548 33652 27600
rect 36084 27548 36136 27600
rect 27988 27523 28040 27532
rect 27988 27489 27997 27523
rect 27997 27489 28031 27523
rect 28031 27489 28040 27523
rect 27988 27480 28040 27489
rect 28816 27523 28868 27532
rect 28816 27489 28825 27523
rect 28825 27489 28859 27523
rect 28859 27489 28868 27523
rect 28816 27480 28868 27489
rect 29000 27480 29052 27532
rect 29368 27480 29420 27532
rect 31116 27523 31168 27532
rect 31116 27489 31125 27523
rect 31125 27489 31159 27523
rect 31159 27489 31168 27523
rect 31116 27480 31168 27489
rect 32220 27480 32272 27532
rect 34520 27523 34572 27532
rect 28080 27455 28132 27464
rect 28080 27421 28089 27455
rect 28089 27421 28123 27455
rect 28123 27421 28132 27455
rect 28080 27412 28132 27421
rect 27896 27344 27948 27396
rect 31852 27412 31904 27464
rect 34520 27489 34529 27523
rect 34529 27489 34563 27523
rect 34563 27489 34572 27523
rect 34520 27480 34572 27489
rect 35624 27480 35676 27532
rect 35992 27412 36044 27464
rect 37188 27480 37240 27532
rect 29736 27276 29788 27328
rect 29828 27276 29880 27328
rect 30472 27276 30524 27328
rect 30840 27276 30892 27328
rect 31208 27276 31260 27328
rect 33140 27319 33192 27328
rect 33140 27285 33149 27319
rect 33149 27285 33183 27319
rect 33183 27285 33192 27319
rect 33140 27276 33192 27285
rect 33600 27276 33652 27328
rect 34796 27276 34848 27328
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 2044 27115 2096 27124
rect 2044 27081 2053 27115
rect 2053 27081 2087 27115
rect 2087 27081 2096 27115
rect 2044 27072 2096 27081
rect 4620 27072 4672 27124
rect 5816 27072 5868 27124
rect 6092 27072 6144 27124
rect 7104 27115 7156 27124
rect 7104 27081 7113 27115
rect 7113 27081 7147 27115
rect 7147 27081 7156 27115
rect 7104 27072 7156 27081
rect 12072 27072 12124 27124
rect 13360 27115 13412 27124
rect 13360 27081 13369 27115
rect 13369 27081 13403 27115
rect 13403 27081 13412 27115
rect 13360 27072 13412 27081
rect 21088 27072 21140 27124
rect 22836 27115 22888 27124
rect 22836 27081 22845 27115
rect 22845 27081 22879 27115
rect 22879 27081 22888 27115
rect 22836 27072 22888 27081
rect 24768 27072 24820 27124
rect 26976 27072 27028 27124
rect 27896 27115 27948 27124
rect 27896 27081 27905 27115
rect 27905 27081 27939 27115
rect 27939 27081 27948 27115
rect 27896 27072 27948 27081
rect 29552 27072 29604 27124
rect 31852 27115 31904 27124
rect 31852 27081 31861 27115
rect 31861 27081 31895 27115
rect 31895 27081 31904 27115
rect 31852 27072 31904 27081
rect 32496 27072 32548 27124
rect 34336 27072 34388 27124
rect 36268 27115 36320 27124
rect 36268 27081 36277 27115
rect 36277 27081 36311 27115
rect 36311 27081 36320 27115
rect 36268 27072 36320 27081
rect 5724 27004 5776 27056
rect 6276 27047 6328 27056
rect 6276 27013 6285 27047
rect 6285 27013 6319 27047
rect 6319 27013 6328 27047
rect 6276 27004 6328 27013
rect 8116 27047 8168 27056
rect 8116 27013 8125 27047
rect 8125 27013 8159 27047
rect 8159 27013 8168 27047
rect 8116 27004 8168 27013
rect 10324 27004 10376 27056
rect 3424 26979 3476 26988
rect 3424 26945 3433 26979
rect 3433 26945 3467 26979
rect 3467 26945 3476 26979
rect 3424 26936 3476 26945
rect 3332 26868 3384 26920
rect 3884 26868 3936 26920
rect 6460 26868 6512 26920
rect 8852 26911 8904 26920
rect 4528 26800 4580 26852
rect 6644 26800 6696 26852
rect 1492 26732 1544 26784
rect 8852 26877 8861 26911
rect 8861 26877 8895 26911
rect 8895 26877 8904 26911
rect 8852 26868 8904 26877
rect 9128 26911 9180 26920
rect 9128 26877 9137 26911
rect 9137 26877 9171 26911
rect 9171 26877 9180 26911
rect 9128 26868 9180 26877
rect 9680 26843 9732 26852
rect 9680 26809 9689 26843
rect 9689 26809 9723 26843
rect 9723 26809 9732 26843
rect 9680 26800 9732 26809
rect 10784 26868 10836 26920
rect 15016 27004 15068 27056
rect 15752 27004 15804 27056
rect 18880 27004 18932 27056
rect 15476 26936 15528 26988
rect 14004 26911 14056 26920
rect 11428 26843 11480 26852
rect 11428 26809 11437 26843
rect 11437 26809 11471 26843
rect 11471 26809 11480 26843
rect 11428 26800 11480 26809
rect 14004 26877 14013 26911
rect 14013 26877 14047 26911
rect 14047 26877 14056 26911
rect 14464 26911 14516 26920
rect 14004 26868 14056 26877
rect 14464 26877 14473 26911
rect 14473 26877 14507 26911
rect 14507 26877 14516 26911
rect 14464 26868 14516 26877
rect 15844 26868 15896 26920
rect 19340 26936 19392 26988
rect 19432 26868 19484 26920
rect 19892 26911 19944 26920
rect 19892 26877 19901 26911
rect 19901 26877 19935 26911
rect 19935 26877 19944 26911
rect 19892 26868 19944 26877
rect 22008 27004 22060 27056
rect 28724 27047 28776 27056
rect 28724 27013 28733 27047
rect 28733 27013 28767 27047
rect 28767 27013 28776 27047
rect 28724 27004 28776 27013
rect 30472 27004 30524 27056
rect 21732 26936 21784 26988
rect 23756 26979 23808 26988
rect 22192 26868 22244 26920
rect 23756 26945 23765 26979
rect 23765 26945 23799 26979
rect 23799 26945 23808 26979
rect 23756 26936 23808 26945
rect 22468 26911 22520 26920
rect 22468 26877 22477 26911
rect 22477 26877 22511 26911
rect 22511 26877 22520 26911
rect 22468 26868 22520 26877
rect 24492 26868 24544 26920
rect 25228 26936 25280 26988
rect 25412 26936 25464 26988
rect 24860 26868 24912 26920
rect 25964 26868 26016 26920
rect 27620 26936 27672 26988
rect 15292 26843 15344 26852
rect 15292 26809 15301 26843
rect 15301 26809 15335 26843
rect 15335 26809 15344 26843
rect 15292 26800 15344 26809
rect 7380 26732 7432 26784
rect 10140 26775 10192 26784
rect 10140 26741 10149 26775
rect 10149 26741 10183 26775
rect 10183 26741 10192 26775
rect 10140 26732 10192 26741
rect 11704 26732 11756 26784
rect 12532 26732 12584 26784
rect 13544 26732 13596 26784
rect 15568 26732 15620 26784
rect 16580 26843 16632 26852
rect 16580 26809 16589 26843
rect 16589 26809 16623 26843
rect 16623 26809 16632 26843
rect 16580 26800 16632 26809
rect 17500 26800 17552 26852
rect 18328 26800 18380 26852
rect 19248 26800 19300 26852
rect 21088 26800 21140 26852
rect 26884 26868 26936 26920
rect 26976 26911 27028 26920
rect 26976 26877 26985 26911
rect 26985 26877 27019 26911
rect 27019 26877 27028 26911
rect 26976 26868 27028 26877
rect 30840 26979 30892 26988
rect 30840 26945 30849 26979
rect 30849 26945 30883 26979
rect 30883 26945 30892 26979
rect 30840 26936 30892 26945
rect 30748 26911 30800 26920
rect 18052 26732 18104 26784
rect 18696 26732 18748 26784
rect 23756 26732 23808 26784
rect 26148 26732 26200 26784
rect 26240 26732 26292 26784
rect 30748 26877 30757 26911
rect 30757 26877 30791 26911
rect 30791 26877 30800 26911
rect 30748 26868 30800 26877
rect 31116 26911 31168 26920
rect 31116 26877 31125 26911
rect 31125 26877 31159 26911
rect 31159 26877 31168 26911
rect 31116 26868 31168 26877
rect 32404 26911 32456 26920
rect 32404 26877 32413 26911
rect 32413 26877 32447 26911
rect 32447 26877 32456 26911
rect 32404 26868 32456 26877
rect 34888 26911 34940 26920
rect 30840 26800 30892 26852
rect 32956 26843 33008 26852
rect 32956 26809 32965 26843
rect 32965 26809 32999 26843
rect 32999 26809 33008 26843
rect 32956 26800 33008 26809
rect 34888 26877 34897 26911
rect 34897 26877 34931 26911
rect 34931 26877 34940 26911
rect 34888 26868 34940 26877
rect 36176 26868 36228 26920
rect 27436 26732 27488 26784
rect 32220 26775 32272 26784
rect 32220 26741 32229 26775
rect 32229 26741 32263 26775
rect 32263 26741 32272 26775
rect 32220 26732 32272 26741
rect 34520 26732 34572 26784
rect 37188 26732 37240 26784
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 1400 26528 1452 26580
rect 2044 26528 2096 26580
rect 3332 26571 3384 26580
rect 3332 26537 3341 26571
rect 3341 26537 3375 26571
rect 3375 26537 3384 26571
rect 3332 26528 3384 26537
rect 4528 26571 4580 26580
rect 4528 26537 4537 26571
rect 4537 26537 4571 26571
rect 4571 26537 4580 26571
rect 4528 26528 4580 26537
rect 7104 26528 7156 26580
rect 8024 26571 8076 26580
rect 8024 26537 8033 26571
rect 8033 26537 8067 26571
rect 8067 26537 8076 26571
rect 8024 26528 8076 26537
rect 14280 26571 14332 26580
rect 14280 26537 14289 26571
rect 14289 26537 14323 26571
rect 14323 26537 14332 26571
rect 14280 26528 14332 26537
rect 16396 26571 16448 26580
rect 16396 26537 16405 26571
rect 16405 26537 16439 26571
rect 16439 26537 16448 26571
rect 16396 26528 16448 26537
rect 16672 26528 16724 26580
rect 9680 26503 9732 26512
rect 5080 26392 5132 26444
rect 9680 26469 9689 26503
rect 9689 26469 9723 26503
rect 9723 26469 9732 26503
rect 9680 26460 9732 26469
rect 16764 26460 16816 26512
rect 6460 26435 6512 26444
rect 6460 26401 6469 26435
rect 6469 26401 6503 26435
rect 6503 26401 6512 26435
rect 6460 26392 6512 26401
rect 6552 26392 6604 26444
rect 7472 26435 7524 26444
rect 4988 26299 5040 26308
rect 4988 26265 4997 26299
rect 4997 26265 5031 26299
rect 5031 26265 5040 26299
rect 4988 26256 5040 26265
rect 5264 26256 5316 26308
rect 6000 26324 6052 26376
rect 7472 26401 7481 26435
rect 7481 26401 7515 26435
rect 7515 26401 7524 26435
rect 7472 26392 7524 26401
rect 7656 26392 7708 26444
rect 10048 26392 10100 26444
rect 10508 26435 10560 26444
rect 10508 26401 10517 26435
rect 10517 26401 10551 26435
rect 10551 26401 10560 26435
rect 10508 26392 10560 26401
rect 10600 26435 10652 26444
rect 10600 26401 10609 26435
rect 10609 26401 10643 26435
rect 10643 26401 10652 26435
rect 10600 26392 10652 26401
rect 11428 26392 11480 26444
rect 12072 26392 12124 26444
rect 12440 26435 12492 26444
rect 12440 26401 12449 26435
rect 12449 26401 12483 26435
rect 12483 26401 12492 26435
rect 12716 26435 12768 26444
rect 12440 26392 12492 26401
rect 12716 26401 12725 26435
rect 12725 26401 12759 26435
rect 12759 26401 12768 26435
rect 12716 26392 12768 26401
rect 14096 26435 14148 26444
rect 14096 26401 14105 26435
rect 14105 26401 14139 26435
rect 14139 26401 14148 26435
rect 14096 26392 14148 26401
rect 15292 26435 15344 26444
rect 15292 26401 15301 26435
rect 15301 26401 15335 26435
rect 15335 26401 15344 26435
rect 15292 26392 15344 26401
rect 17684 26392 17736 26444
rect 23848 26528 23900 26580
rect 25964 26571 26016 26580
rect 25964 26537 25973 26571
rect 25973 26537 26007 26571
rect 26007 26537 26016 26571
rect 25964 26528 26016 26537
rect 27988 26571 28040 26580
rect 27988 26537 27997 26571
rect 27997 26537 28031 26571
rect 28031 26537 28040 26571
rect 27988 26528 28040 26537
rect 31024 26528 31076 26580
rect 32404 26528 32456 26580
rect 34704 26571 34756 26580
rect 34704 26537 34713 26571
rect 34713 26537 34747 26571
rect 34747 26537 34756 26571
rect 34704 26528 34756 26537
rect 35624 26528 35676 26580
rect 36084 26571 36136 26580
rect 36084 26537 36093 26571
rect 36093 26537 36127 26571
rect 36127 26537 36136 26571
rect 36084 26528 36136 26537
rect 19432 26460 19484 26512
rect 24860 26460 24912 26512
rect 26240 26503 26292 26512
rect 26240 26469 26249 26503
rect 26249 26469 26283 26503
rect 26283 26469 26292 26503
rect 26240 26460 26292 26469
rect 26608 26460 26660 26512
rect 27252 26460 27304 26512
rect 28816 26460 28868 26512
rect 29092 26503 29144 26512
rect 29092 26469 29101 26503
rect 29101 26469 29135 26503
rect 29135 26469 29144 26503
rect 29092 26460 29144 26469
rect 19524 26435 19576 26444
rect 9128 26367 9180 26376
rect 9128 26333 9137 26367
rect 9137 26333 9171 26367
rect 9171 26333 9180 26367
rect 9128 26324 9180 26333
rect 11796 26367 11848 26376
rect 11796 26333 11805 26367
rect 11805 26333 11839 26367
rect 11839 26333 11848 26367
rect 11796 26324 11848 26333
rect 12992 26367 13044 26376
rect 12992 26333 13001 26367
rect 13001 26333 13035 26367
rect 13035 26333 13044 26367
rect 12992 26324 13044 26333
rect 13176 26367 13228 26376
rect 13176 26333 13185 26367
rect 13185 26333 13219 26367
rect 13219 26333 13228 26367
rect 13176 26324 13228 26333
rect 17408 26367 17460 26376
rect 17408 26333 17417 26367
rect 17417 26333 17451 26367
rect 17451 26333 17460 26367
rect 17408 26324 17460 26333
rect 17500 26324 17552 26376
rect 19524 26401 19533 26435
rect 19533 26401 19567 26435
rect 19567 26401 19576 26435
rect 19524 26392 19576 26401
rect 21088 26435 21140 26444
rect 21088 26401 21097 26435
rect 21097 26401 21131 26435
rect 21131 26401 21140 26435
rect 21088 26392 21140 26401
rect 21456 26435 21508 26444
rect 21456 26401 21465 26435
rect 21465 26401 21499 26435
rect 21499 26401 21508 26435
rect 21456 26392 21508 26401
rect 22008 26392 22060 26444
rect 26792 26392 26844 26444
rect 20352 26324 20404 26376
rect 26240 26324 26292 26376
rect 6644 26256 6696 26308
rect 7748 26188 7800 26240
rect 8484 26256 8536 26308
rect 8852 26256 8904 26308
rect 11336 26299 11388 26308
rect 11336 26265 11345 26299
rect 11345 26265 11379 26299
rect 11379 26265 11388 26299
rect 11336 26256 11388 26265
rect 13452 26256 13504 26308
rect 15108 26256 15160 26308
rect 19892 26256 19944 26308
rect 21180 26256 21232 26308
rect 26884 26324 26936 26376
rect 27896 26392 27948 26444
rect 29552 26392 29604 26444
rect 29828 26435 29880 26444
rect 29828 26401 29837 26435
rect 29837 26401 29871 26435
rect 29871 26401 29880 26435
rect 29828 26392 29880 26401
rect 30012 26392 30064 26444
rect 30472 26392 30524 26444
rect 31208 26392 31260 26444
rect 34520 26435 34572 26444
rect 29092 26256 29144 26308
rect 34520 26401 34529 26435
rect 34529 26401 34563 26435
rect 34563 26401 34572 26435
rect 34520 26392 34572 26401
rect 33508 26256 33560 26308
rect 10968 26231 11020 26240
rect 10968 26197 10977 26231
rect 10977 26197 11011 26231
rect 11011 26197 11020 26231
rect 10968 26188 11020 26197
rect 11612 26188 11664 26240
rect 15752 26231 15804 26240
rect 15752 26197 15761 26231
rect 15761 26197 15795 26231
rect 15795 26197 15804 26231
rect 15752 26188 15804 26197
rect 18328 26188 18380 26240
rect 22836 26188 22888 26240
rect 27988 26188 28040 26240
rect 30840 26188 30892 26240
rect 35808 26188 35860 26240
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 2780 26027 2832 26036
rect 2780 25993 2789 26027
rect 2789 25993 2823 26027
rect 2823 25993 2832 26027
rect 2780 25984 2832 25993
rect 5080 25984 5132 26036
rect 8944 26027 8996 26036
rect 8944 25993 8953 26027
rect 8953 25993 8987 26027
rect 8987 25993 8996 26027
rect 8944 25984 8996 25993
rect 11796 26027 11848 26036
rect 11796 25993 11805 26027
rect 11805 25993 11839 26027
rect 11839 25993 11848 26027
rect 11796 25984 11848 25993
rect 13820 26027 13872 26036
rect 13820 25993 13829 26027
rect 13829 25993 13863 26027
rect 13863 25993 13872 26027
rect 13820 25984 13872 25993
rect 14648 25984 14700 26036
rect 15292 26027 15344 26036
rect 15292 25993 15301 26027
rect 15301 25993 15335 26027
rect 15335 25993 15344 26027
rect 15292 25984 15344 25993
rect 15936 25984 15988 26036
rect 16396 25984 16448 26036
rect 17500 25984 17552 26036
rect 17684 26027 17736 26036
rect 17684 25993 17693 26027
rect 17693 25993 17727 26027
rect 17727 25993 17736 26027
rect 17684 25984 17736 25993
rect 19524 25984 19576 26036
rect 21088 25984 21140 26036
rect 21456 25984 21508 26036
rect 22008 25984 22060 26036
rect 22468 26027 22520 26036
rect 22468 25993 22477 26027
rect 22477 25993 22511 26027
rect 22511 25993 22520 26027
rect 22468 25984 22520 25993
rect 25320 25984 25372 26036
rect 26148 25984 26200 26036
rect 26884 25984 26936 26036
rect 27804 26027 27856 26036
rect 27804 25993 27813 26027
rect 27813 25993 27847 26027
rect 27847 25993 27856 26027
rect 27804 25984 27856 25993
rect 29552 26027 29604 26036
rect 29552 25993 29561 26027
rect 29561 25993 29595 26027
rect 29595 25993 29604 26027
rect 29552 25984 29604 25993
rect 29828 25984 29880 26036
rect 30748 25984 30800 26036
rect 34520 26027 34572 26036
rect 34520 25993 34529 26027
rect 34529 25993 34563 26027
rect 34563 25993 34572 26027
rect 34520 25984 34572 25993
rect 37280 25984 37332 26036
rect 12440 25916 12492 25968
rect 12716 25916 12768 25968
rect 17408 25959 17460 25968
rect 17408 25925 17417 25959
rect 17417 25925 17451 25959
rect 17451 25925 17460 25959
rect 17408 25916 17460 25925
rect 27160 25916 27212 25968
rect 29184 25916 29236 25968
rect 30012 25916 30064 25968
rect 32312 25916 32364 25968
rect 1400 25891 1452 25900
rect 1400 25857 1409 25891
rect 1409 25857 1443 25891
rect 1443 25857 1452 25891
rect 1400 25848 1452 25857
rect 4620 25891 4672 25900
rect 4620 25857 4629 25891
rect 4629 25857 4663 25891
rect 4663 25857 4672 25891
rect 4620 25848 4672 25857
rect 7012 25848 7064 25900
rect 7104 25848 7156 25900
rect 8208 25848 8260 25900
rect 9128 25848 9180 25900
rect 10232 25891 10284 25900
rect 10232 25857 10241 25891
rect 10241 25857 10275 25891
rect 10275 25857 10284 25891
rect 10876 25891 10928 25900
rect 10232 25848 10284 25857
rect 10876 25857 10885 25891
rect 10885 25857 10919 25891
rect 10919 25857 10928 25891
rect 10876 25848 10928 25857
rect 1676 25823 1728 25832
rect 1676 25789 1685 25823
rect 1685 25789 1719 25823
rect 1719 25789 1728 25823
rect 1676 25780 1728 25789
rect 4528 25823 4580 25832
rect 4528 25789 4537 25823
rect 4537 25789 4571 25823
rect 4571 25789 4580 25823
rect 4528 25780 4580 25789
rect 5264 25687 5316 25696
rect 5264 25653 5273 25687
rect 5273 25653 5307 25687
rect 5307 25653 5316 25687
rect 5264 25644 5316 25653
rect 6000 25644 6052 25696
rect 6552 25687 6604 25696
rect 6552 25653 6561 25687
rect 6561 25653 6595 25687
rect 6595 25653 6604 25687
rect 6552 25644 6604 25653
rect 7472 25780 7524 25832
rect 7748 25780 7800 25832
rect 10968 25823 11020 25832
rect 8208 25687 8260 25696
rect 8208 25653 8217 25687
rect 8217 25653 8251 25687
rect 8251 25653 8260 25687
rect 8208 25644 8260 25653
rect 10968 25789 10977 25823
rect 10977 25789 11011 25823
rect 11011 25789 11020 25823
rect 10968 25780 11020 25789
rect 11060 25780 11112 25832
rect 12164 25780 12216 25832
rect 14096 25848 14148 25900
rect 15108 25848 15160 25900
rect 15752 25848 15804 25900
rect 18512 25891 18564 25900
rect 18512 25857 18521 25891
rect 18521 25857 18555 25891
rect 18555 25857 18564 25891
rect 18512 25848 18564 25857
rect 29644 25848 29696 25900
rect 30196 25848 30248 25900
rect 31852 25848 31904 25900
rect 13544 25780 13596 25832
rect 14372 25823 14424 25832
rect 14372 25789 14381 25823
rect 14381 25789 14415 25823
rect 14415 25789 14424 25823
rect 14372 25780 14424 25789
rect 15200 25780 15252 25832
rect 11612 25712 11664 25764
rect 13176 25712 13228 25764
rect 15384 25755 15436 25764
rect 15384 25721 15393 25755
rect 15393 25721 15427 25755
rect 15427 25721 15436 25755
rect 15384 25712 15436 25721
rect 15936 25823 15988 25832
rect 15936 25789 15945 25823
rect 15945 25789 15979 25823
rect 15979 25789 15988 25823
rect 15936 25780 15988 25789
rect 18236 25823 18288 25832
rect 18236 25789 18245 25823
rect 18245 25789 18279 25823
rect 18279 25789 18288 25823
rect 18236 25780 18288 25789
rect 22836 25780 22888 25832
rect 23664 25823 23716 25832
rect 23664 25789 23673 25823
rect 23673 25789 23707 25823
rect 23707 25789 23716 25823
rect 23664 25780 23716 25789
rect 23940 25823 23992 25832
rect 23940 25789 23949 25823
rect 23949 25789 23983 25823
rect 23983 25789 23992 25823
rect 23940 25780 23992 25789
rect 26884 25780 26936 25832
rect 8852 25644 8904 25696
rect 10048 25644 10100 25696
rect 10784 25644 10836 25696
rect 13084 25644 13136 25696
rect 14280 25644 14332 25696
rect 20352 25644 20404 25696
rect 25044 25687 25096 25696
rect 25044 25653 25053 25687
rect 25053 25653 25087 25687
rect 25087 25653 25096 25687
rect 25044 25644 25096 25653
rect 29092 25780 29144 25832
rect 29368 25823 29420 25832
rect 29368 25789 29377 25823
rect 29377 25789 29411 25823
rect 29411 25789 29420 25823
rect 29368 25780 29420 25789
rect 30196 25712 30248 25764
rect 32956 25780 33008 25832
rect 32404 25755 32456 25764
rect 32404 25721 32413 25755
rect 32413 25721 32447 25755
rect 32447 25721 32456 25755
rect 32404 25712 32456 25721
rect 28264 25644 28316 25696
rect 28724 25687 28776 25696
rect 28724 25653 28733 25687
rect 28733 25653 28767 25687
rect 28767 25653 28776 25687
rect 28724 25644 28776 25653
rect 32312 25687 32364 25696
rect 32312 25653 32321 25687
rect 32321 25653 32355 25687
rect 32355 25653 32364 25687
rect 33508 25780 33560 25832
rect 35808 25823 35860 25832
rect 35808 25789 35817 25823
rect 35817 25789 35851 25823
rect 35851 25789 35860 25823
rect 35808 25780 35860 25789
rect 36084 25823 36136 25832
rect 36084 25789 36093 25823
rect 36093 25789 36127 25823
rect 36127 25789 36136 25823
rect 36084 25780 36136 25789
rect 32312 25644 32364 25653
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 7104 25440 7156 25492
rect 7196 25415 7248 25424
rect 7196 25381 7205 25415
rect 7205 25381 7239 25415
rect 7239 25381 7248 25415
rect 7196 25372 7248 25381
rect 10600 25440 10652 25492
rect 12072 25483 12124 25492
rect 12072 25449 12081 25483
rect 12081 25449 12115 25483
rect 12115 25449 12124 25483
rect 12072 25440 12124 25449
rect 12624 25440 12676 25492
rect 14372 25483 14424 25492
rect 14372 25449 14381 25483
rect 14381 25449 14415 25483
rect 14415 25449 14424 25483
rect 14372 25440 14424 25449
rect 15016 25440 15068 25492
rect 15936 25440 15988 25492
rect 16764 25440 16816 25492
rect 18512 25440 18564 25492
rect 19432 25483 19484 25492
rect 19432 25449 19441 25483
rect 19441 25449 19475 25483
rect 19475 25449 19484 25483
rect 19432 25440 19484 25449
rect 21548 25440 21600 25492
rect 23204 25440 23256 25492
rect 23664 25483 23716 25492
rect 23664 25449 23673 25483
rect 23673 25449 23707 25483
rect 23707 25449 23716 25483
rect 23664 25440 23716 25449
rect 29552 25440 29604 25492
rect 30196 25483 30248 25492
rect 5080 25304 5132 25356
rect 5448 25304 5500 25356
rect 9496 25372 9548 25424
rect 16672 25415 16724 25424
rect 16672 25381 16681 25415
rect 16681 25381 16715 25415
rect 16715 25381 16724 25415
rect 16672 25372 16724 25381
rect 27436 25372 27488 25424
rect 30196 25449 30205 25483
rect 30205 25449 30239 25483
rect 30239 25449 30248 25483
rect 30196 25440 30248 25449
rect 30564 25440 30616 25492
rect 31852 25483 31904 25492
rect 31852 25449 31861 25483
rect 31861 25449 31895 25483
rect 31895 25449 31904 25483
rect 31852 25440 31904 25449
rect 32864 25440 32916 25492
rect 35808 25483 35860 25492
rect 35808 25449 35817 25483
rect 35817 25449 35851 25483
rect 35851 25449 35860 25483
rect 35808 25440 35860 25449
rect 32680 25415 32732 25424
rect 32680 25381 32689 25415
rect 32689 25381 32723 25415
rect 32723 25381 32732 25415
rect 32680 25372 32732 25381
rect 8116 25347 8168 25356
rect 8116 25313 8125 25347
rect 8125 25313 8159 25347
rect 8159 25313 8168 25347
rect 8116 25304 8168 25313
rect 8852 25304 8904 25356
rect 11244 25347 11296 25356
rect 11244 25313 11253 25347
rect 11253 25313 11287 25347
rect 11287 25313 11296 25347
rect 11244 25304 11296 25313
rect 11612 25347 11664 25356
rect 11612 25313 11621 25347
rect 11621 25313 11655 25347
rect 11655 25313 11664 25347
rect 11612 25304 11664 25313
rect 12900 25304 12952 25356
rect 13176 25347 13228 25356
rect 13176 25313 13185 25347
rect 13185 25313 13219 25347
rect 13219 25313 13228 25347
rect 13176 25304 13228 25313
rect 13360 25347 13412 25356
rect 13360 25313 13369 25347
rect 13369 25313 13403 25347
rect 13403 25313 13412 25347
rect 13360 25304 13412 25313
rect 13544 25347 13596 25356
rect 13544 25313 13553 25347
rect 13553 25313 13587 25347
rect 13587 25313 13596 25347
rect 13544 25304 13596 25313
rect 14096 25347 14148 25356
rect 14096 25313 14105 25347
rect 14105 25313 14139 25347
rect 14139 25313 14148 25347
rect 14096 25304 14148 25313
rect 16580 25304 16632 25356
rect 17408 25304 17460 25356
rect 17500 25347 17552 25356
rect 17500 25313 17509 25347
rect 17509 25313 17543 25347
rect 17543 25313 17552 25347
rect 17500 25304 17552 25313
rect 17868 25304 17920 25356
rect 21088 25304 21140 25356
rect 21916 25347 21968 25356
rect 21916 25313 21925 25347
rect 21925 25313 21959 25347
rect 21959 25313 21968 25347
rect 21916 25304 21968 25313
rect 25596 25304 25648 25356
rect 25964 25304 26016 25356
rect 29276 25347 29328 25356
rect 29276 25313 29285 25347
rect 29285 25313 29319 25347
rect 29319 25313 29328 25347
rect 29276 25304 29328 25313
rect 29460 25304 29512 25356
rect 30564 25304 30616 25356
rect 32220 25347 32272 25356
rect 4804 25236 4856 25288
rect 5264 25279 5316 25288
rect 5264 25245 5273 25279
rect 5273 25245 5307 25279
rect 5307 25245 5316 25279
rect 5264 25236 5316 25245
rect 7196 25236 7248 25288
rect 4988 25168 5040 25220
rect 7012 25168 7064 25220
rect 7840 25168 7892 25220
rect 8392 25236 8444 25288
rect 10876 25236 10928 25288
rect 11428 25236 11480 25288
rect 11520 25236 11572 25288
rect 11888 25236 11940 25288
rect 13728 25279 13780 25288
rect 13728 25245 13737 25279
rect 13737 25245 13771 25279
rect 13771 25245 13780 25279
rect 13728 25236 13780 25245
rect 15936 25279 15988 25288
rect 15936 25245 15945 25279
rect 15945 25245 15979 25279
rect 15979 25245 15988 25279
rect 15936 25236 15988 25245
rect 17224 25236 17276 25288
rect 21364 25279 21416 25288
rect 21364 25245 21373 25279
rect 21373 25245 21407 25279
rect 21407 25245 21416 25279
rect 21364 25236 21416 25245
rect 21732 25236 21784 25288
rect 27620 25236 27672 25288
rect 28264 25279 28316 25288
rect 28264 25245 28273 25279
rect 28273 25245 28307 25279
rect 28307 25245 28316 25279
rect 28264 25236 28316 25245
rect 32220 25313 32229 25347
rect 32229 25313 32263 25347
rect 32263 25313 32272 25347
rect 32220 25304 32272 25313
rect 32588 25304 32640 25356
rect 33508 25347 33560 25356
rect 33508 25313 33517 25347
rect 33517 25313 33551 25347
rect 33551 25313 33560 25347
rect 33508 25304 33560 25313
rect 13360 25168 13412 25220
rect 15384 25168 15436 25220
rect 16304 25168 16356 25220
rect 16672 25168 16724 25220
rect 17776 25168 17828 25220
rect 25688 25168 25740 25220
rect 26424 25168 26476 25220
rect 30472 25168 30524 25220
rect 32220 25168 32272 25220
rect 1676 25143 1728 25152
rect 1676 25109 1685 25143
rect 1685 25109 1719 25143
rect 1719 25109 1728 25143
rect 1676 25100 1728 25109
rect 2964 25100 3016 25152
rect 6460 25143 6512 25152
rect 6460 25109 6469 25143
rect 6469 25109 6503 25143
rect 6503 25109 6512 25143
rect 6460 25100 6512 25109
rect 6920 25143 6972 25152
rect 6920 25109 6929 25143
rect 6929 25109 6963 25143
rect 6963 25109 6972 25143
rect 6920 25100 6972 25109
rect 9588 25100 9640 25152
rect 11428 25100 11480 25152
rect 12624 25100 12676 25152
rect 16212 25143 16264 25152
rect 16212 25109 16221 25143
rect 16221 25109 16255 25143
rect 16255 25109 16264 25143
rect 16212 25100 16264 25109
rect 25872 25100 25924 25152
rect 26792 25143 26844 25152
rect 26792 25109 26801 25143
rect 26801 25109 26835 25143
rect 26835 25109 26844 25143
rect 26792 25100 26844 25109
rect 27068 25143 27120 25152
rect 27068 25109 27077 25143
rect 27077 25109 27111 25143
rect 27111 25109 27120 25143
rect 27068 25100 27120 25109
rect 31116 25100 31168 25152
rect 31576 25100 31628 25152
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 6920 24896 6972 24948
rect 10968 24896 11020 24948
rect 3332 24828 3384 24880
rect 3516 24828 3568 24880
rect 5448 24760 5500 24812
rect 6552 24760 6604 24812
rect 3516 24692 3568 24744
rect 5172 24692 5224 24744
rect 5632 24624 5684 24676
rect 8116 24828 8168 24880
rect 9496 24828 9548 24880
rect 10876 24828 10928 24880
rect 13728 24896 13780 24948
rect 17224 24939 17276 24948
rect 17224 24905 17233 24939
rect 17233 24905 17267 24939
rect 17267 24905 17276 24939
rect 17224 24896 17276 24905
rect 17408 24896 17460 24948
rect 27252 24896 27304 24948
rect 29276 24896 29328 24948
rect 13176 24828 13228 24880
rect 13360 24828 13412 24880
rect 7012 24692 7064 24744
rect 7288 24692 7340 24744
rect 8208 24692 8260 24744
rect 9404 24735 9456 24744
rect 9404 24701 9413 24735
rect 9413 24701 9447 24735
rect 9447 24701 9456 24735
rect 9404 24692 9456 24701
rect 7196 24667 7248 24676
rect 7196 24633 7205 24667
rect 7205 24633 7239 24667
rect 7239 24633 7248 24667
rect 7196 24624 7248 24633
rect 8944 24667 8996 24676
rect 8944 24633 8953 24667
rect 8953 24633 8987 24667
rect 8987 24633 8996 24667
rect 8944 24624 8996 24633
rect 9864 24760 9916 24812
rect 11796 24803 11848 24812
rect 11796 24769 11805 24803
rect 11805 24769 11839 24803
rect 11839 24769 11848 24803
rect 11796 24760 11848 24769
rect 12716 24760 12768 24812
rect 15292 24803 15344 24812
rect 15292 24769 15301 24803
rect 15301 24769 15335 24803
rect 15335 24769 15344 24803
rect 15292 24760 15344 24769
rect 16212 24803 16264 24812
rect 16212 24769 16221 24803
rect 16221 24769 16255 24803
rect 16255 24769 16264 24803
rect 16212 24760 16264 24769
rect 27068 24828 27120 24880
rect 27712 24871 27764 24880
rect 27712 24837 27721 24871
rect 27721 24837 27755 24871
rect 27755 24837 27764 24871
rect 27712 24828 27764 24837
rect 31576 24828 31628 24880
rect 9772 24735 9824 24744
rect 9772 24701 9781 24735
rect 9781 24701 9815 24735
rect 9815 24701 9824 24735
rect 10048 24735 10100 24744
rect 9772 24692 9824 24701
rect 10048 24701 10057 24735
rect 10057 24701 10091 24735
rect 10091 24701 10100 24735
rect 10048 24692 10100 24701
rect 10508 24692 10560 24744
rect 11428 24692 11480 24744
rect 11520 24692 11572 24744
rect 13084 24735 13136 24744
rect 13084 24701 13093 24735
rect 13093 24701 13127 24735
rect 13127 24701 13136 24735
rect 13084 24692 13136 24701
rect 11796 24624 11848 24676
rect 13268 24692 13320 24744
rect 13452 24735 13504 24744
rect 13452 24701 13461 24735
rect 13461 24701 13495 24735
rect 13495 24701 13504 24735
rect 13452 24692 13504 24701
rect 16304 24735 16356 24744
rect 16304 24701 16313 24735
rect 16313 24701 16347 24735
rect 16347 24701 16356 24735
rect 16304 24692 16356 24701
rect 20628 24760 20680 24812
rect 21916 24760 21968 24812
rect 16948 24692 17000 24744
rect 19892 24735 19944 24744
rect 19892 24701 19901 24735
rect 19901 24701 19935 24735
rect 19935 24701 19944 24735
rect 19892 24692 19944 24701
rect 25872 24760 25924 24812
rect 28264 24760 28316 24812
rect 31392 24760 31444 24812
rect 25596 24692 25648 24744
rect 25688 24735 25740 24744
rect 25688 24701 25697 24735
rect 25697 24701 25731 24735
rect 25731 24701 25740 24735
rect 26240 24735 26292 24744
rect 25688 24692 25740 24701
rect 26240 24701 26249 24735
rect 26249 24701 26283 24735
rect 26283 24701 26292 24735
rect 26240 24692 26292 24701
rect 27620 24735 27672 24744
rect 27620 24701 27629 24735
rect 27629 24701 27663 24735
rect 27663 24701 27672 24735
rect 27620 24692 27672 24701
rect 26424 24624 26476 24676
rect 29368 24692 29420 24744
rect 29460 24692 29512 24744
rect 31484 24735 31536 24744
rect 31484 24701 31493 24735
rect 31493 24701 31527 24735
rect 31527 24701 31536 24735
rect 31484 24692 31536 24701
rect 32128 24760 32180 24812
rect 37188 24760 37240 24812
rect 32956 24692 33008 24744
rect 35808 24735 35860 24744
rect 35808 24701 35817 24735
rect 35817 24701 35851 24735
rect 35851 24701 35860 24735
rect 35808 24692 35860 24701
rect 5080 24599 5132 24608
rect 5080 24565 5089 24599
rect 5089 24565 5123 24599
rect 5123 24565 5132 24599
rect 5080 24556 5132 24565
rect 6920 24556 6972 24608
rect 7840 24599 7892 24608
rect 7840 24565 7849 24599
rect 7849 24565 7883 24599
rect 7883 24565 7892 24599
rect 7840 24556 7892 24565
rect 11612 24556 11664 24608
rect 12256 24599 12308 24608
rect 12256 24565 12265 24599
rect 12265 24565 12299 24599
rect 12299 24565 12308 24599
rect 12256 24556 12308 24565
rect 15476 24556 15528 24608
rect 17040 24556 17092 24608
rect 20260 24556 20312 24608
rect 21732 24556 21784 24608
rect 24400 24599 24452 24608
rect 24400 24565 24409 24599
rect 24409 24565 24443 24599
rect 24443 24565 24452 24599
rect 24400 24556 24452 24565
rect 25964 24556 26016 24608
rect 28264 24624 28316 24676
rect 30012 24624 30064 24676
rect 31760 24624 31812 24676
rect 27620 24556 27672 24608
rect 29920 24556 29972 24608
rect 30472 24556 30524 24608
rect 32220 24599 32272 24608
rect 32220 24565 32229 24599
rect 32229 24565 32263 24599
rect 32263 24565 32272 24599
rect 32220 24556 32272 24565
rect 33508 24599 33560 24608
rect 33508 24565 33517 24599
rect 33517 24565 33551 24599
rect 33551 24565 33560 24599
rect 33508 24556 33560 24565
rect 36084 24556 36136 24608
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 3516 24395 3568 24404
rect 3516 24361 3525 24395
rect 3525 24361 3559 24395
rect 3559 24361 3568 24395
rect 3516 24352 3568 24361
rect 7748 24395 7800 24404
rect 7748 24361 7757 24395
rect 7757 24361 7791 24395
rect 7791 24361 7800 24395
rect 7748 24352 7800 24361
rect 4896 24284 4948 24336
rect 11244 24284 11296 24336
rect 12900 24284 12952 24336
rect 1400 24259 1452 24268
rect 1400 24225 1409 24259
rect 1409 24225 1443 24259
rect 1443 24225 1452 24259
rect 1400 24216 1452 24225
rect 5264 24216 5316 24268
rect 5540 24216 5592 24268
rect 6368 24259 6420 24268
rect 1584 24148 1636 24200
rect 4712 24148 4764 24200
rect 5172 24148 5224 24200
rect 6368 24225 6377 24259
rect 6377 24225 6411 24259
rect 6411 24225 6420 24259
rect 6368 24216 6420 24225
rect 7288 24216 7340 24268
rect 7472 24216 7524 24268
rect 7564 24259 7616 24268
rect 7564 24225 7573 24259
rect 7573 24225 7607 24259
rect 7607 24225 7616 24259
rect 7564 24216 7616 24225
rect 8852 24216 8904 24268
rect 10048 24216 10100 24268
rect 10232 24259 10284 24268
rect 10232 24225 10241 24259
rect 10241 24225 10275 24259
rect 10275 24225 10284 24259
rect 10232 24216 10284 24225
rect 9864 24148 9916 24200
rect 3424 24080 3476 24132
rect 7196 24080 7248 24132
rect 9772 24080 9824 24132
rect 13912 24259 13964 24268
rect 13912 24225 13921 24259
rect 13921 24225 13955 24259
rect 13955 24225 13964 24259
rect 13912 24216 13964 24225
rect 16212 24284 16264 24336
rect 16764 24352 16816 24404
rect 17500 24352 17552 24404
rect 21364 24352 21416 24404
rect 24032 24395 24084 24404
rect 24032 24361 24041 24395
rect 24041 24361 24075 24395
rect 24075 24361 24084 24395
rect 24032 24352 24084 24361
rect 26240 24352 26292 24404
rect 28264 24395 28316 24404
rect 28264 24361 28273 24395
rect 28273 24361 28307 24395
rect 28307 24361 28316 24395
rect 28264 24352 28316 24361
rect 16948 24284 17000 24336
rect 17408 24284 17460 24336
rect 25964 24327 26016 24336
rect 25964 24293 25973 24327
rect 25973 24293 26007 24327
rect 26007 24293 26016 24327
rect 25964 24284 26016 24293
rect 26884 24327 26936 24336
rect 26884 24293 26893 24327
rect 26893 24293 26927 24327
rect 26927 24293 26936 24327
rect 26884 24284 26936 24293
rect 16120 24259 16172 24268
rect 10876 24191 10928 24200
rect 10876 24157 10885 24191
rect 10885 24157 10919 24191
rect 10919 24157 10928 24191
rect 10876 24148 10928 24157
rect 11060 24191 11112 24200
rect 11060 24157 11069 24191
rect 11069 24157 11103 24191
rect 11103 24157 11112 24191
rect 11060 24148 11112 24157
rect 12440 24191 12492 24200
rect 12440 24157 12449 24191
rect 12449 24157 12483 24191
rect 12483 24157 12492 24191
rect 12992 24191 13044 24200
rect 12440 24148 12492 24157
rect 12992 24157 13001 24191
rect 13001 24157 13035 24191
rect 13035 24157 13044 24191
rect 12992 24148 13044 24157
rect 14096 24148 14148 24200
rect 16120 24225 16129 24259
rect 16129 24225 16163 24259
rect 16163 24225 16172 24259
rect 16120 24216 16172 24225
rect 17040 24216 17092 24268
rect 17684 24216 17736 24268
rect 23204 24216 23256 24268
rect 25504 24216 25556 24268
rect 27252 24259 27304 24268
rect 27252 24225 27261 24259
rect 27261 24225 27295 24259
rect 27295 24225 27304 24259
rect 27252 24216 27304 24225
rect 28448 24259 28500 24268
rect 28448 24225 28457 24259
rect 28457 24225 28491 24259
rect 28491 24225 28500 24259
rect 28448 24216 28500 24225
rect 30932 24352 30984 24404
rect 31392 24352 31444 24404
rect 32312 24395 32364 24404
rect 32312 24361 32321 24395
rect 32321 24361 32355 24395
rect 32355 24361 32364 24395
rect 32312 24352 32364 24361
rect 32588 24395 32640 24404
rect 32588 24361 32597 24395
rect 32597 24361 32631 24395
rect 32631 24361 32640 24395
rect 32588 24352 32640 24361
rect 32956 24395 33008 24404
rect 32956 24361 32965 24395
rect 32965 24361 32999 24395
rect 32999 24361 33008 24395
rect 32956 24352 33008 24361
rect 35808 24395 35860 24404
rect 35808 24361 35817 24395
rect 35817 24361 35851 24395
rect 35851 24361 35860 24395
rect 35808 24352 35860 24361
rect 29184 24284 29236 24336
rect 29644 24284 29696 24336
rect 30012 24259 30064 24268
rect 30012 24225 30021 24259
rect 30021 24225 30055 24259
rect 30055 24225 30064 24259
rect 30012 24216 30064 24225
rect 31024 24259 31076 24268
rect 31024 24225 31033 24259
rect 31033 24225 31067 24259
rect 31067 24225 31076 24259
rect 31024 24216 31076 24225
rect 31484 24216 31536 24268
rect 32220 24216 32272 24268
rect 32680 24216 32732 24268
rect 12348 24123 12400 24132
rect 12348 24089 12357 24123
rect 12357 24089 12391 24123
rect 12391 24089 12400 24123
rect 12348 24080 12400 24089
rect 13544 24080 13596 24132
rect 13728 24123 13780 24132
rect 13728 24089 13737 24123
rect 13737 24089 13771 24123
rect 13771 24089 13780 24123
rect 13728 24080 13780 24089
rect 15476 24148 15528 24200
rect 17960 24148 18012 24200
rect 18236 24148 18288 24200
rect 21088 24148 21140 24200
rect 22928 24191 22980 24200
rect 22928 24157 22937 24191
rect 22937 24157 22971 24191
rect 22971 24157 22980 24191
rect 22928 24148 22980 24157
rect 27712 24148 27764 24200
rect 29184 24191 29236 24200
rect 21548 24080 21600 24132
rect 26056 24080 26108 24132
rect 3884 24055 3936 24064
rect 3884 24021 3893 24055
rect 3893 24021 3927 24055
rect 3927 24021 3936 24055
rect 3884 24012 3936 24021
rect 6368 24012 6420 24064
rect 8668 24055 8720 24064
rect 8668 24021 8677 24055
rect 8677 24021 8711 24055
rect 8711 24021 8720 24055
rect 8668 24012 8720 24021
rect 11612 24012 11664 24064
rect 12164 24012 12216 24064
rect 12256 24012 12308 24064
rect 14372 24012 14424 24064
rect 18696 24012 18748 24064
rect 19892 24012 19944 24064
rect 20168 24012 20220 24064
rect 27620 24012 27672 24064
rect 29184 24157 29193 24191
rect 29193 24157 29227 24191
rect 29227 24157 29236 24191
rect 29184 24148 29236 24157
rect 29276 24080 29328 24132
rect 31576 24080 31628 24132
rect 29368 24012 29420 24064
rect 29552 24055 29604 24064
rect 29552 24021 29561 24055
rect 29561 24021 29595 24055
rect 29595 24021 29604 24055
rect 29552 24012 29604 24021
rect 30564 24012 30616 24064
rect 30840 24012 30892 24064
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 1584 23851 1636 23860
rect 1584 23817 1593 23851
rect 1593 23817 1627 23851
rect 1627 23817 1636 23851
rect 1584 23808 1636 23817
rect 3792 23851 3844 23860
rect 3792 23817 3801 23851
rect 3801 23817 3835 23851
rect 3835 23817 3844 23851
rect 3792 23808 3844 23817
rect 4712 23808 4764 23860
rect 9772 23851 9824 23860
rect 1400 23740 1452 23792
rect 5540 23740 5592 23792
rect 9772 23817 9781 23851
rect 9781 23817 9815 23851
rect 9815 23817 9824 23851
rect 9772 23808 9824 23817
rect 11060 23808 11112 23860
rect 11428 23808 11480 23860
rect 12440 23808 12492 23860
rect 12716 23851 12768 23860
rect 12716 23817 12725 23851
rect 12725 23817 12759 23851
rect 12759 23817 12768 23851
rect 12716 23808 12768 23817
rect 14004 23808 14056 23860
rect 15936 23808 15988 23860
rect 17408 23851 17460 23860
rect 17408 23817 17417 23851
rect 17417 23817 17451 23851
rect 17451 23817 17460 23851
rect 17408 23808 17460 23817
rect 18880 23851 18932 23860
rect 18880 23817 18889 23851
rect 18889 23817 18923 23851
rect 18923 23817 18932 23851
rect 18880 23808 18932 23817
rect 20260 23808 20312 23860
rect 3424 23715 3476 23724
rect 3424 23681 3433 23715
rect 3433 23681 3467 23715
rect 3467 23681 3476 23715
rect 3424 23672 3476 23681
rect 5908 23672 5960 23724
rect 13912 23740 13964 23792
rect 15384 23740 15436 23792
rect 6184 23647 6236 23656
rect 6184 23613 6193 23647
rect 6193 23613 6227 23647
rect 6227 23613 6236 23647
rect 6184 23604 6236 23613
rect 7564 23715 7616 23724
rect 7564 23681 7573 23715
rect 7573 23681 7607 23715
rect 7607 23681 7616 23715
rect 7564 23672 7616 23681
rect 10600 23672 10652 23724
rect 11520 23715 11572 23724
rect 7472 23604 7524 23656
rect 8668 23604 8720 23656
rect 9680 23604 9732 23656
rect 10784 23647 10836 23656
rect 10784 23613 10793 23647
rect 10793 23613 10827 23647
rect 10827 23613 10836 23647
rect 10784 23604 10836 23613
rect 11520 23681 11529 23715
rect 11529 23681 11563 23715
rect 11563 23681 11572 23715
rect 11520 23672 11572 23681
rect 11336 23604 11388 23656
rect 12348 23604 12400 23656
rect 3056 23579 3108 23588
rect 3056 23545 3065 23579
rect 3065 23545 3099 23579
rect 3099 23545 3108 23579
rect 3056 23536 3108 23545
rect 4804 23536 4856 23588
rect 7196 23579 7248 23588
rect 7196 23545 7205 23579
rect 7205 23545 7239 23579
rect 7239 23545 7248 23579
rect 7196 23536 7248 23545
rect 8944 23579 8996 23588
rect 8944 23545 8953 23579
rect 8953 23545 8987 23579
rect 8987 23545 8996 23579
rect 8944 23536 8996 23545
rect 9588 23536 9640 23588
rect 11244 23536 11296 23588
rect 13360 23536 13412 23588
rect 13820 23604 13872 23656
rect 14832 23672 14884 23724
rect 16580 23672 16632 23724
rect 23204 23808 23256 23860
rect 25872 23851 25924 23860
rect 25872 23817 25881 23851
rect 25881 23817 25915 23851
rect 25915 23817 25924 23851
rect 25872 23808 25924 23817
rect 24860 23783 24912 23792
rect 24860 23749 24869 23783
rect 24869 23749 24903 23783
rect 24903 23749 24912 23783
rect 24860 23740 24912 23749
rect 27252 23808 27304 23860
rect 28448 23808 28500 23860
rect 29460 23808 29512 23860
rect 30012 23808 30064 23860
rect 26884 23740 26936 23792
rect 27896 23740 27948 23792
rect 21732 23672 21784 23724
rect 14004 23647 14056 23656
rect 14004 23613 14013 23647
rect 14013 23613 14047 23647
rect 14047 23613 14056 23647
rect 14004 23604 14056 23613
rect 14372 23604 14424 23656
rect 16764 23604 16816 23656
rect 18604 23647 18656 23656
rect 13728 23536 13780 23588
rect 15476 23536 15528 23588
rect 16120 23579 16172 23588
rect 16120 23545 16129 23579
rect 16129 23545 16163 23579
rect 16163 23545 16172 23579
rect 16120 23536 16172 23545
rect 5264 23468 5316 23520
rect 6460 23468 6512 23520
rect 7104 23468 7156 23520
rect 8024 23511 8076 23520
rect 8024 23477 8033 23511
rect 8033 23477 8067 23511
rect 8067 23477 8076 23511
rect 8024 23468 8076 23477
rect 8392 23511 8444 23520
rect 8392 23477 8401 23511
rect 8401 23477 8435 23511
rect 8435 23477 8444 23511
rect 8392 23468 8444 23477
rect 11060 23468 11112 23520
rect 15108 23468 15160 23520
rect 18604 23613 18613 23647
rect 18613 23613 18647 23647
rect 18647 23613 18656 23647
rect 18604 23604 18656 23613
rect 18696 23647 18748 23656
rect 18696 23613 18705 23647
rect 18705 23613 18739 23647
rect 18739 23613 18748 23647
rect 18696 23604 18748 23613
rect 19892 23536 19944 23588
rect 21088 23604 21140 23656
rect 21548 23647 21600 23656
rect 21548 23613 21557 23647
rect 21557 23613 21591 23647
rect 21591 23613 21600 23647
rect 21548 23604 21600 23613
rect 29092 23715 29144 23724
rect 25872 23604 25924 23656
rect 27620 23647 27672 23656
rect 27620 23613 27629 23647
rect 27629 23613 27663 23647
rect 27663 23613 27672 23647
rect 27620 23604 27672 23613
rect 29092 23681 29101 23715
rect 29101 23681 29135 23715
rect 29135 23681 29144 23715
rect 29092 23672 29144 23681
rect 29552 23647 29604 23656
rect 29552 23613 29561 23647
rect 29561 23613 29595 23647
rect 29595 23613 29604 23647
rect 29552 23604 29604 23613
rect 30932 23672 30984 23724
rect 31116 23715 31168 23724
rect 31116 23681 31125 23715
rect 31125 23681 31159 23715
rect 31159 23681 31168 23715
rect 31116 23672 31168 23681
rect 36084 23715 36136 23724
rect 36084 23681 36093 23715
rect 36093 23681 36127 23715
rect 36127 23681 36136 23715
rect 36084 23672 36136 23681
rect 31576 23604 31628 23656
rect 31760 23647 31812 23656
rect 31760 23613 31769 23647
rect 31769 23613 31803 23647
rect 31803 23613 31812 23647
rect 35808 23647 35860 23656
rect 31760 23604 31812 23613
rect 35808 23613 35817 23647
rect 35817 23613 35851 23647
rect 35851 23613 35860 23647
rect 35808 23604 35860 23613
rect 22928 23536 22980 23588
rect 23388 23536 23440 23588
rect 26884 23536 26936 23588
rect 28816 23536 28868 23588
rect 32864 23536 32916 23588
rect 25320 23468 25372 23520
rect 25504 23511 25556 23520
rect 25504 23477 25513 23511
rect 25513 23477 25547 23511
rect 25547 23477 25556 23511
rect 25504 23468 25556 23477
rect 32680 23468 32732 23520
rect 37372 23511 37424 23520
rect 37372 23477 37381 23511
rect 37381 23477 37415 23511
rect 37415 23477 37424 23511
rect 37372 23468 37424 23477
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 3884 23307 3936 23316
rect 3884 23273 3893 23307
rect 3893 23273 3927 23307
rect 3927 23273 3936 23307
rect 3884 23264 3936 23273
rect 6460 23307 6512 23316
rect 6460 23273 6469 23307
rect 6469 23273 6503 23307
rect 6503 23273 6512 23307
rect 6460 23264 6512 23273
rect 8300 23264 8352 23316
rect 9864 23307 9916 23316
rect 9864 23273 9873 23307
rect 9873 23273 9907 23307
rect 9907 23273 9916 23307
rect 9864 23264 9916 23273
rect 10232 23264 10284 23316
rect 14648 23307 14700 23316
rect 14648 23273 14657 23307
rect 14657 23273 14691 23307
rect 14691 23273 14700 23307
rect 14648 23264 14700 23273
rect 15660 23307 15712 23316
rect 15660 23273 15669 23307
rect 15669 23273 15703 23307
rect 15703 23273 15712 23307
rect 15660 23264 15712 23273
rect 16764 23264 16816 23316
rect 17040 23264 17092 23316
rect 17684 23307 17736 23316
rect 17684 23273 17693 23307
rect 17693 23273 17727 23307
rect 17727 23273 17736 23307
rect 17684 23264 17736 23273
rect 6184 23196 6236 23248
rect 6644 23239 6696 23248
rect 6644 23205 6653 23239
rect 6653 23205 6687 23239
rect 6687 23205 6696 23239
rect 6644 23196 6696 23205
rect 7012 23239 7064 23248
rect 7012 23205 7021 23239
rect 7021 23205 7055 23239
rect 7055 23205 7064 23239
rect 7012 23196 7064 23205
rect 7564 23196 7616 23248
rect 1400 23128 1452 23180
rect 4620 23128 4672 23180
rect 5448 23128 5500 23180
rect 5632 23128 5684 23180
rect 6552 23171 6604 23180
rect 6552 23137 6561 23171
rect 6561 23137 6595 23171
rect 6595 23137 6604 23171
rect 6552 23128 6604 23137
rect 8208 23171 8260 23180
rect 8208 23137 8217 23171
rect 8217 23137 8251 23171
rect 8251 23137 8260 23171
rect 8208 23128 8260 23137
rect 8668 23196 8720 23248
rect 12348 23196 12400 23248
rect 12808 23196 12860 23248
rect 15936 23196 15988 23248
rect 17960 23239 18012 23248
rect 9772 23128 9824 23180
rect 11520 23171 11572 23180
rect 11520 23137 11529 23171
rect 11529 23137 11563 23171
rect 11563 23137 11572 23171
rect 11520 23128 11572 23137
rect 11612 23171 11664 23180
rect 11612 23137 11621 23171
rect 11621 23137 11655 23171
rect 11655 23137 11664 23171
rect 13360 23171 13412 23180
rect 11612 23128 11664 23137
rect 13360 23137 13369 23171
rect 13369 23137 13403 23171
rect 13403 23137 13412 23171
rect 13360 23128 13412 23137
rect 13544 23171 13596 23180
rect 13544 23137 13553 23171
rect 13553 23137 13587 23171
rect 13587 23137 13596 23171
rect 13544 23128 13596 23137
rect 14372 23128 14424 23180
rect 16120 23128 16172 23180
rect 17960 23205 17969 23239
rect 17969 23205 18003 23239
rect 18003 23205 18012 23239
rect 17960 23196 18012 23205
rect 21364 23264 21416 23316
rect 23480 23264 23532 23316
rect 25596 23307 25648 23316
rect 25596 23273 25605 23307
rect 25605 23273 25639 23307
rect 25639 23273 25648 23307
rect 25596 23264 25648 23273
rect 26240 23307 26292 23316
rect 26240 23273 26249 23307
rect 26249 23273 26283 23307
rect 26283 23273 26292 23307
rect 26240 23264 26292 23273
rect 27068 23264 27120 23316
rect 27620 23307 27672 23316
rect 27620 23273 27629 23307
rect 27629 23273 27663 23307
rect 27663 23273 27672 23307
rect 27620 23264 27672 23273
rect 27896 23264 27948 23316
rect 18880 23171 18932 23180
rect 18880 23137 18889 23171
rect 18889 23137 18923 23171
rect 18923 23137 18932 23171
rect 18880 23128 18932 23137
rect 19616 23196 19668 23248
rect 28264 23264 28316 23316
rect 29368 23264 29420 23316
rect 31024 23307 31076 23316
rect 31024 23273 31033 23307
rect 31033 23273 31067 23307
rect 31067 23273 31076 23307
rect 31024 23264 31076 23273
rect 31116 23264 31168 23316
rect 31760 23307 31812 23316
rect 31760 23273 31769 23307
rect 31769 23273 31803 23307
rect 31803 23273 31812 23307
rect 31760 23264 31812 23273
rect 35808 23307 35860 23316
rect 35808 23273 35817 23307
rect 35817 23273 35851 23307
rect 35851 23273 35860 23307
rect 35808 23264 35860 23273
rect 28724 23196 28776 23248
rect 1676 23060 1728 23112
rect 3516 23060 3568 23112
rect 7288 23060 7340 23112
rect 8024 23103 8076 23112
rect 8024 23069 8033 23103
rect 8033 23069 8067 23103
rect 8067 23069 8076 23103
rect 8024 23060 8076 23069
rect 10968 23060 11020 23112
rect 5172 23035 5224 23044
rect 5172 23001 5181 23035
rect 5181 23001 5215 23035
rect 5215 23001 5224 23035
rect 5172 22992 5224 23001
rect 10876 23035 10928 23044
rect 10876 23001 10885 23035
rect 10885 23001 10919 23035
rect 10919 23001 10928 23035
rect 10876 22992 10928 23001
rect 14280 23103 14332 23112
rect 14280 23069 14289 23103
rect 14289 23069 14323 23103
rect 14323 23069 14332 23103
rect 15844 23103 15896 23112
rect 14280 23060 14332 23069
rect 15844 23069 15853 23103
rect 15853 23069 15887 23103
rect 15887 23069 15896 23103
rect 15844 23060 15896 23069
rect 16304 23103 16356 23112
rect 16304 23069 16313 23103
rect 16313 23069 16347 23103
rect 16347 23069 16356 23103
rect 16304 23060 16356 23069
rect 16764 23060 16816 23112
rect 18420 23060 18472 23112
rect 20076 23128 20128 23180
rect 20720 23128 20772 23180
rect 22560 23128 22612 23180
rect 25964 23128 26016 23180
rect 29276 23128 29328 23180
rect 29460 23128 29512 23180
rect 32956 23128 33008 23180
rect 23204 23060 23256 23112
rect 26884 23103 26936 23112
rect 26884 23069 26893 23103
rect 26893 23069 26927 23103
rect 26927 23069 26936 23103
rect 26884 23060 26936 23069
rect 28540 23103 28592 23112
rect 28540 23069 28549 23103
rect 28549 23069 28583 23103
rect 28583 23069 28592 23103
rect 28540 23060 28592 23069
rect 31760 23060 31812 23112
rect 32128 23060 32180 23112
rect 32496 23060 32548 23112
rect 18696 23035 18748 23044
rect 3240 22924 3292 22976
rect 3332 22924 3384 22976
rect 3700 22924 3752 22976
rect 4896 22924 4948 22976
rect 5356 22924 5408 22976
rect 7104 22924 7156 22976
rect 9404 22967 9456 22976
rect 9404 22933 9413 22967
rect 9413 22933 9447 22967
rect 9447 22933 9456 22967
rect 9404 22924 9456 22933
rect 10784 22924 10836 22976
rect 11428 22924 11480 22976
rect 12440 22967 12492 22976
rect 12440 22933 12449 22967
rect 12449 22933 12483 22967
rect 12483 22933 12492 22967
rect 12808 22967 12860 22976
rect 12440 22924 12492 22933
rect 12808 22933 12817 22967
rect 12817 22933 12851 22967
rect 12851 22933 12860 22967
rect 12808 22924 12860 22933
rect 18696 23001 18705 23035
rect 18705 23001 18739 23035
rect 18739 23001 18748 23035
rect 18696 22992 18748 23001
rect 27252 22992 27304 23044
rect 14556 22924 14608 22976
rect 17408 22924 17460 22976
rect 18236 22924 18288 22976
rect 20996 22924 21048 22976
rect 25964 22967 26016 22976
rect 25964 22933 25973 22967
rect 25973 22933 26007 22967
rect 26007 22933 26016 22967
rect 25964 22924 26016 22933
rect 26056 22924 26108 22976
rect 26332 22924 26384 22976
rect 27160 22967 27212 22976
rect 27160 22933 27169 22967
rect 27169 22933 27203 22967
rect 27203 22933 27212 22967
rect 27160 22924 27212 22933
rect 30288 22967 30340 22976
rect 30288 22933 30297 22967
rect 30297 22933 30331 22967
rect 30331 22933 30340 22967
rect 30288 22924 30340 22933
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 1676 22763 1728 22772
rect 1676 22729 1685 22763
rect 1685 22729 1719 22763
rect 1719 22729 1728 22763
rect 1676 22720 1728 22729
rect 4620 22720 4672 22772
rect 5264 22720 5316 22772
rect 10968 22720 11020 22772
rect 11152 22720 11204 22772
rect 11612 22720 11664 22772
rect 12256 22763 12308 22772
rect 12256 22729 12265 22763
rect 12265 22729 12299 22763
rect 12299 22729 12308 22763
rect 12256 22720 12308 22729
rect 12532 22720 12584 22772
rect 13544 22720 13596 22772
rect 15200 22720 15252 22772
rect 16948 22720 17000 22772
rect 17408 22763 17460 22772
rect 17408 22729 17417 22763
rect 17417 22729 17451 22763
rect 17451 22729 17460 22763
rect 17408 22720 17460 22729
rect 18236 22763 18288 22772
rect 18236 22729 18245 22763
rect 18245 22729 18279 22763
rect 18279 22729 18288 22763
rect 18236 22720 18288 22729
rect 18604 22763 18656 22772
rect 18604 22729 18613 22763
rect 18613 22729 18647 22763
rect 18647 22729 18656 22763
rect 18604 22720 18656 22729
rect 18880 22720 18932 22772
rect 19616 22763 19668 22772
rect 19616 22729 19625 22763
rect 19625 22729 19659 22763
rect 19659 22729 19668 22763
rect 19616 22720 19668 22729
rect 19892 22720 19944 22772
rect 21548 22763 21600 22772
rect 3148 22652 3200 22704
rect 6920 22652 6972 22704
rect 8208 22652 8260 22704
rect 3516 22584 3568 22636
rect 3056 22516 3108 22568
rect 3240 22559 3292 22568
rect 3240 22525 3249 22559
rect 3249 22525 3283 22559
rect 3283 22525 3292 22559
rect 3240 22516 3292 22525
rect 5172 22584 5224 22636
rect 7104 22584 7156 22636
rect 3792 22559 3844 22568
rect 3792 22525 3801 22559
rect 3801 22525 3835 22559
rect 3835 22525 3844 22559
rect 3792 22516 3844 22525
rect 4068 22516 4120 22568
rect 4896 22559 4948 22568
rect 4896 22525 4905 22559
rect 4905 22525 4939 22559
rect 4939 22525 4948 22559
rect 4896 22516 4948 22525
rect 6644 22516 6696 22568
rect 8024 22584 8076 22636
rect 8760 22584 8812 22636
rect 9772 22652 9824 22704
rect 10692 22695 10744 22704
rect 10692 22661 10701 22695
rect 10701 22661 10735 22695
rect 10735 22661 10744 22695
rect 10692 22652 10744 22661
rect 11428 22695 11480 22704
rect 11428 22661 11437 22695
rect 11437 22661 11471 22695
rect 11471 22661 11480 22695
rect 11428 22652 11480 22661
rect 12624 22652 12676 22704
rect 9680 22584 9732 22636
rect 11060 22584 11112 22636
rect 13544 22627 13596 22636
rect 13544 22593 13553 22627
rect 13553 22593 13587 22627
rect 13587 22593 13596 22627
rect 13544 22584 13596 22593
rect 14280 22627 14332 22636
rect 14280 22593 14289 22627
rect 14289 22593 14323 22627
rect 14323 22593 14332 22627
rect 14280 22584 14332 22593
rect 14924 22584 14976 22636
rect 17040 22652 17092 22704
rect 17684 22652 17736 22704
rect 16764 22584 16816 22636
rect 18420 22584 18472 22636
rect 12992 22516 13044 22568
rect 13912 22516 13964 22568
rect 14004 22516 14056 22568
rect 15108 22516 15160 22568
rect 16948 22559 17000 22568
rect 16948 22525 16957 22559
rect 16957 22525 16991 22559
rect 16991 22525 17000 22559
rect 16948 22516 17000 22525
rect 18604 22516 18656 22568
rect 21548 22729 21557 22763
rect 21557 22729 21591 22763
rect 21591 22729 21600 22763
rect 21548 22720 21600 22729
rect 22560 22763 22612 22772
rect 22560 22729 22569 22763
rect 22569 22729 22603 22763
rect 22603 22729 22612 22763
rect 22560 22720 22612 22729
rect 20168 22627 20220 22636
rect 20168 22593 20184 22627
rect 20184 22593 20218 22627
rect 20218 22593 20220 22627
rect 23204 22720 23256 22772
rect 26884 22720 26936 22772
rect 25596 22652 25648 22704
rect 25504 22627 25556 22636
rect 20168 22584 20220 22593
rect 25504 22593 25513 22627
rect 25513 22593 25547 22627
rect 25547 22593 25556 22627
rect 25504 22584 25556 22593
rect 25964 22516 26016 22568
rect 27252 22720 27304 22772
rect 29276 22720 29328 22772
rect 32128 22763 32180 22772
rect 32128 22729 32137 22763
rect 32137 22729 32171 22763
rect 32171 22729 32180 22763
rect 32128 22720 32180 22729
rect 32496 22763 32548 22772
rect 32496 22729 32505 22763
rect 32505 22729 32539 22763
rect 32539 22729 32548 22763
rect 32496 22720 32548 22729
rect 28724 22652 28776 22704
rect 29552 22652 29604 22704
rect 32956 22695 33008 22704
rect 32956 22661 32965 22695
rect 32965 22661 32999 22695
rect 32999 22661 33008 22695
rect 32956 22652 33008 22661
rect 27068 22559 27120 22568
rect 27068 22525 27077 22559
rect 27077 22525 27111 22559
rect 27111 22525 27120 22559
rect 27068 22516 27120 22525
rect 30288 22584 30340 22636
rect 28448 22516 28500 22568
rect 29092 22516 29144 22568
rect 29184 22516 29236 22568
rect 37280 22627 37332 22636
rect 37280 22593 37289 22627
rect 37289 22593 37323 22627
rect 37323 22593 37332 22627
rect 37280 22584 37332 22593
rect 35808 22559 35860 22568
rect 35808 22525 35817 22559
rect 35817 22525 35851 22559
rect 35851 22525 35860 22559
rect 35808 22516 35860 22525
rect 36084 22559 36136 22568
rect 36084 22525 36093 22559
rect 36093 22525 36127 22559
rect 36127 22525 36136 22559
rect 36084 22516 36136 22525
rect 2596 22491 2648 22500
rect 2596 22457 2605 22491
rect 2605 22457 2639 22491
rect 2639 22457 2648 22491
rect 2596 22448 2648 22457
rect 7288 22491 7340 22500
rect 7288 22457 7297 22491
rect 7297 22457 7331 22491
rect 7331 22457 7340 22491
rect 7288 22448 7340 22457
rect 6552 22380 6604 22432
rect 7840 22448 7892 22500
rect 8300 22448 8352 22500
rect 9220 22491 9272 22500
rect 9220 22457 9229 22491
rect 9229 22457 9263 22491
rect 9263 22457 9272 22491
rect 9220 22448 9272 22457
rect 9588 22491 9640 22500
rect 9588 22457 9597 22491
rect 9597 22457 9631 22491
rect 9631 22457 9640 22491
rect 9588 22448 9640 22457
rect 10784 22448 10836 22500
rect 11520 22448 11572 22500
rect 12348 22448 12400 22500
rect 12808 22448 12860 22500
rect 16212 22448 16264 22500
rect 16304 22448 16356 22500
rect 27252 22448 27304 22500
rect 29460 22448 29512 22500
rect 30840 22448 30892 22500
rect 31576 22448 31628 22500
rect 7564 22423 7616 22432
rect 7564 22389 7573 22423
rect 7573 22389 7607 22423
rect 7607 22389 7616 22423
rect 7564 22380 7616 22389
rect 9404 22380 9456 22432
rect 10508 22380 10560 22432
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 3516 22176 3568 22228
rect 3792 22108 3844 22160
rect 2872 22040 2924 22092
rect 3976 22176 4028 22228
rect 5908 22176 5960 22228
rect 6184 22176 6236 22228
rect 4620 22108 4672 22160
rect 6092 22108 6144 22160
rect 7288 22176 7340 22228
rect 8760 22219 8812 22228
rect 8024 22151 8076 22160
rect 8024 22117 8033 22151
rect 8033 22117 8067 22151
rect 8067 22117 8076 22151
rect 8024 22108 8076 22117
rect 8760 22185 8769 22219
rect 8769 22185 8803 22219
rect 8803 22185 8812 22219
rect 8760 22176 8812 22185
rect 9404 22219 9456 22228
rect 9404 22185 9413 22219
rect 9413 22185 9447 22219
rect 9447 22185 9456 22219
rect 9404 22176 9456 22185
rect 13360 22176 13412 22228
rect 15844 22219 15896 22228
rect 10048 22151 10100 22160
rect 4712 22040 4764 22092
rect 5264 22040 5316 22092
rect 1860 21972 1912 22024
rect 5540 22040 5592 22092
rect 6460 22040 6512 22092
rect 6828 22040 6880 22092
rect 7012 22083 7064 22092
rect 7012 22049 7021 22083
rect 7021 22049 7055 22083
rect 7055 22049 7064 22083
rect 7012 22040 7064 22049
rect 8208 22040 8260 22092
rect 10048 22117 10057 22151
rect 10057 22117 10091 22151
rect 10091 22117 10100 22151
rect 10048 22108 10100 22117
rect 10508 22108 10560 22160
rect 12532 22151 12584 22160
rect 12532 22117 12541 22151
rect 12541 22117 12575 22151
rect 12575 22117 12584 22151
rect 12532 22108 12584 22117
rect 9220 22040 9272 22092
rect 11060 22083 11112 22092
rect 11060 22049 11069 22083
rect 11069 22049 11103 22083
rect 11103 22049 11112 22083
rect 11060 22040 11112 22049
rect 11336 22040 11388 22092
rect 11888 22040 11940 22092
rect 12256 22040 12308 22092
rect 12716 22040 12768 22092
rect 12808 22083 12860 22092
rect 12808 22049 12817 22083
rect 12817 22049 12851 22083
rect 12851 22049 12860 22083
rect 12808 22040 12860 22049
rect 6276 21972 6328 22024
rect 7380 22015 7432 22024
rect 7380 21981 7389 22015
rect 7389 21981 7423 22015
rect 7423 21981 7432 22015
rect 7380 21972 7432 21981
rect 7656 22015 7708 22024
rect 7656 21981 7665 22015
rect 7665 21981 7699 22015
rect 7699 21981 7708 22015
rect 7656 21972 7708 21981
rect 8392 21972 8444 22024
rect 9680 22015 9732 22024
rect 9680 21981 9689 22015
rect 9689 21981 9723 22015
rect 9723 21981 9732 22015
rect 9680 21972 9732 21981
rect 10692 21972 10744 22024
rect 15844 22185 15853 22219
rect 15853 22185 15887 22219
rect 15887 22185 15896 22219
rect 15844 22176 15896 22185
rect 16028 22176 16080 22228
rect 19432 22176 19484 22228
rect 20168 22219 20220 22228
rect 20168 22185 20177 22219
rect 20177 22185 20211 22219
rect 20211 22185 20220 22219
rect 20168 22176 20220 22185
rect 26332 22219 26384 22228
rect 26332 22185 26341 22219
rect 26341 22185 26375 22219
rect 26375 22185 26384 22219
rect 26332 22176 26384 22185
rect 29460 22176 29512 22228
rect 29828 22176 29880 22228
rect 35808 22219 35860 22228
rect 35808 22185 35817 22219
rect 35817 22185 35851 22219
rect 35851 22185 35860 22219
rect 35808 22176 35860 22185
rect 15936 22108 15988 22160
rect 13912 22083 13964 22092
rect 13912 22049 13921 22083
rect 13921 22049 13955 22083
rect 13955 22049 13964 22083
rect 13912 22040 13964 22049
rect 14648 22083 14700 22092
rect 14648 22049 14657 22083
rect 14657 22049 14691 22083
rect 14691 22049 14700 22083
rect 14648 22040 14700 22049
rect 16028 21972 16080 22024
rect 16212 21972 16264 22024
rect 17408 22040 17460 22092
rect 18604 22040 18656 22092
rect 21272 22083 21324 22092
rect 21272 22049 21281 22083
rect 21281 22049 21315 22083
rect 21315 22049 21324 22083
rect 21272 22040 21324 22049
rect 22284 22040 22336 22092
rect 16580 22015 16632 22024
rect 16580 21981 16589 22015
rect 16589 21981 16623 22015
rect 16623 21981 16632 22015
rect 16580 21972 16632 21981
rect 8668 21904 8720 21956
rect 16304 21904 16356 21956
rect 17224 21972 17276 22024
rect 17684 21904 17736 21956
rect 18788 21972 18840 22024
rect 21364 22015 21416 22024
rect 21364 21981 21373 22015
rect 21373 21981 21407 22015
rect 21407 21981 21416 22015
rect 21364 21972 21416 21981
rect 22376 21972 22428 22024
rect 23296 22015 23348 22024
rect 23296 21981 23305 22015
rect 23305 21981 23339 22015
rect 23339 21981 23348 22015
rect 23296 21972 23348 21981
rect 24492 22040 24544 22092
rect 27344 22083 27396 22092
rect 27344 22049 27353 22083
rect 27353 22049 27387 22083
rect 27387 22049 27396 22083
rect 27344 22040 27396 22049
rect 28816 22083 28868 22092
rect 28816 22049 28825 22083
rect 28825 22049 28859 22083
rect 28859 22049 28868 22083
rect 28816 22040 28868 22049
rect 30472 22083 30524 22092
rect 30472 22049 30481 22083
rect 30481 22049 30515 22083
rect 30515 22049 30524 22083
rect 30472 22040 30524 22049
rect 31300 22040 31352 22092
rect 33048 22040 33100 22092
rect 35256 22040 35308 22092
rect 23664 21904 23716 21956
rect 24032 21904 24084 21956
rect 27160 21972 27212 22024
rect 30288 22015 30340 22024
rect 30288 21981 30297 22015
rect 30297 21981 30331 22015
rect 30331 21981 30340 22015
rect 30288 21972 30340 21981
rect 30656 21972 30708 22024
rect 32956 22015 33008 22024
rect 32956 21981 32965 22015
rect 32965 21981 32999 22015
rect 32999 21981 33008 22015
rect 32956 21972 33008 21981
rect 27620 21904 27672 21956
rect 2044 21879 2096 21888
rect 2044 21845 2053 21879
rect 2053 21845 2087 21879
rect 2087 21845 2096 21879
rect 2044 21836 2096 21845
rect 3516 21879 3568 21888
rect 3516 21845 3525 21879
rect 3525 21845 3559 21879
rect 3559 21845 3568 21879
rect 3516 21836 3568 21845
rect 5080 21879 5132 21888
rect 5080 21845 5089 21879
rect 5089 21845 5123 21879
rect 5123 21845 5132 21879
rect 5080 21836 5132 21845
rect 5448 21836 5500 21888
rect 5632 21836 5684 21888
rect 7196 21836 7248 21888
rect 7564 21836 7616 21888
rect 8576 21836 8628 21888
rect 9128 21836 9180 21888
rect 9588 21836 9640 21888
rect 11244 21836 11296 21888
rect 12440 21836 12492 21888
rect 13268 21836 13320 21888
rect 15016 21879 15068 21888
rect 15016 21845 15025 21879
rect 15025 21845 15059 21879
rect 15059 21845 15068 21879
rect 15016 21836 15068 21845
rect 17960 21879 18012 21888
rect 17960 21845 17969 21879
rect 17969 21845 18003 21879
rect 18003 21845 18012 21879
rect 17960 21836 18012 21845
rect 25872 21836 25924 21888
rect 28632 21879 28684 21888
rect 28632 21845 28641 21879
rect 28641 21845 28675 21879
rect 28675 21845 28684 21879
rect 28632 21836 28684 21845
rect 31668 21836 31720 21888
rect 34060 21879 34112 21888
rect 34060 21845 34069 21879
rect 34069 21845 34103 21879
rect 34103 21845 34112 21879
rect 34060 21836 34112 21845
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 3884 21632 3936 21684
rect 5540 21675 5592 21684
rect 1952 21539 2004 21548
rect 1952 21505 1961 21539
rect 1961 21505 1995 21539
rect 1995 21505 2004 21539
rect 1952 21496 2004 21505
rect 2872 21496 2924 21548
rect 2044 21428 2096 21480
rect 3240 21428 3292 21480
rect 5540 21641 5549 21675
rect 5549 21641 5583 21675
rect 5583 21641 5592 21675
rect 5540 21632 5592 21641
rect 6460 21632 6512 21684
rect 9220 21632 9272 21684
rect 9956 21632 10008 21684
rect 10600 21632 10652 21684
rect 11152 21632 11204 21684
rect 8576 21564 8628 21616
rect 4712 21496 4764 21548
rect 7104 21496 7156 21548
rect 7196 21496 7248 21548
rect 6920 21428 6972 21480
rect 3148 21360 3200 21412
rect 7748 21496 7800 21548
rect 7380 21428 7432 21480
rect 7564 21403 7616 21412
rect 7564 21369 7573 21403
rect 7573 21369 7607 21403
rect 7607 21369 7616 21403
rect 7564 21360 7616 21369
rect 9588 21564 9640 21616
rect 10508 21564 10560 21616
rect 9956 21539 10008 21548
rect 9956 21505 9965 21539
rect 9965 21505 9999 21539
rect 9999 21505 10008 21539
rect 9956 21496 10008 21505
rect 10048 21496 10100 21548
rect 11796 21564 11848 21616
rect 14004 21632 14056 21684
rect 15936 21632 15988 21684
rect 17684 21632 17736 21684
rect 12716 21564 12768 21616
rect 12992 21496 13044 21548
rect 13452 21496 13504 21548
rect 15016 21496 15068 21548
rect 9772 21428 9824 21480
rect 11244 21428 11296 21480
rect 3056 21292 3108 21344
rect 6644 21292 6696 21344
rect 8024 21292 8076 21344
rect 8392 21335 8444 21344
rect 8392 21301 8401 21335
rect 8401 21301 8435 21335
rect 8435 21301 8444 21335
rect 8392 21292 8444 21301
rect 10048 21360 10100 21412
rect 8852 21292 8904 21344
rect 11336 21335 11388 21344
rect 11336 21301 11345 21335
rect 11345 21301 11379 21335
rect 11379 21301 11388 21335
rect 11336 21292 11388 21301
rect 11428 21292 11480 21344
rect 12716 21335 12768 21344
rect 12716 21301 12725 21335
rect 12725 21301 12759 21335
rect 12759 21301 12768 21335
rect 12716 21292 12768 21301
rect 13268 21428 13320 21480
rect 13912 21428 13964 21480
rect 15476 21471 15528 21480
rect 15476 21437 15485 21471
rect 15485 21437 15519 21471
rect 15519 21437 15528 21471
rect 15476 21428 15528 21437
rect 15660 21428 15712 21480
rect 19064 21471 19116 21480
rect 15844 21360 15896 21412
rect 13452 21292 13504 21344
rect 14096 21292 14148 21344
rect 15108 21292 15160 21344
rect 15936 21292 15988 21344
rect 16580 21292 16632 21344
rect 17316 21335 17368 21344
rect 17316 21301 17325 21335
rect 17325 21301 17359 21335
rect 17359 21301 17368 21335
rect 17316 21292 17368 21301
rect 18144 21292 18196 21344
rect 18604 21292 18656 21344
rect 19064 21437 19073 21471
rect 19073 21437 19107 21471
rect 19107 21437 19116 21471
rect 19064 21428 19116 21437
rect 19340 21428 19392 21480
rect 20260 21632 20312 21684
rect 21272 21632 21324 21684
rect 26056 21632 26108 21684
rect 27344 21632 27396 21684
rect 28816 21632 28868 21684
rect 32956 21632 33008 21684
rect 33048 21675 33100 21684
rect 33048 21641 33057 21675
rect 33057 21641 33091 21675
rect 33091 21641 33100 21675
rect 35256 21675 35308 21684
rect 33048 21632 33100 21641
rect 35256 21641 35265 21675
rect 35265 21641 35299 21675
rect 35299 21641 35308 21675
rect 35256 21632 35308 21641
rect 35348 21632 35400 21684
rect 22376 21564 22428 21616
rect 23572 21564 23624 21616
rect 26516 21607 26568 21616
rect 26516 21573 26525 21607
rect 26525 21573 26559 21607
rect 26559 21573 26568 21607
rect 26516 21564 26568 21573
rect 29184 21564 29236 21616
rect 29460 21564 29512 21616
rect 29644 21564 29696 21616
rect 29920 21564 29972 21616
rect 30288 21564 30340 21616
rect 23848 21539 23900 21548
rect 23848 21505 23857 21539
rect 23857 21505 23891 21539
rect 23891 21505 23900 21539
rect 23848 21496 23900 21505
rect 25872 21496 25924 21548
rect 21640 21471 21692 21480
rect 21640 21437 21649 21471
rect 21649 21437 21683 21471
rect 21683 21437 21692 21471
rect 21640 21428 21692 21437
rect 24032 21471 24084 21480
rect 24032 21437 24041 21471
rect 24041 21437 24075 21471
rect 24075 21437 24084 21471
rect 24032 21428 24084 21437
rect 24492 21471 24544 21480
rect 24492 21437 24501 21471
rect 24501 21437 24535 21471
rect 24535 21437 24544 21471
rect 24492 21428 24544 21437
rect 25504 21471 25556 21480
rect 25504 21437 25513 21471
rect 25513 21437 25547 21471
rect 25547 21437 25556 21471
rect 25504 21428 25556 21437
rect 25964 21471 26016 21480
rect 25964 21437 25973 21471
rect 25973 21437 26007 21471
rect 26007 21437 26016 21471
rect 25964 21428 26016 21437
rect 28264 21496 28316 21548
rect 28632 21496 28684 21548
rect 29552 21428 29604 21480
rect 21272 21403 21324 21412
rect 21272 21369 21281 21403
rect 21281 21369 21315 21403
rect 21315 21369 21324 21403
rect 21272 21360 21324 21369
rect 29920 21428 29972 21480
rect 30380 21428 30432 21480
rect 31300 21496 31352 21548
rect 31392 21471 31444 21480
rect 31392 21437 31401 21471
rect 31401 21437 31435 21471
rect 31435 21437 31444 21471
rect 31392 21428 31444 21437
rect 31668 21471 31720 21480
rect 31668 21437 31677 21471
rect 31677 21437 31711 21471
rect 31711 21437 31720 21471
rect 31668 21428 31720 21437
rect 32772 21496 32824 21548
rect 35716 21471 35768 21480
rect 35716 21437 35725 21471
rect 35725 21437 35759 21471
rect 35759 21437 35768 21471
rect 35716 21428 35768 21437
rect 35808 21471 35860 21480
rect 35808 21437 35817 21471
rect 35817 21437 35851 21471
rect 35851 21437 35860 21471
rect 35808 21428 35860 21437
rect 19156 21292 19208 21344
rect 19432 21292 19484 21344
rect 22376 21335 22428 21344
rect 22376 21301 22385 21335
rect 22385 21301 22419 21335
rect 22419 21301 22428 21335
rect 22376 21292 22428 21301
rect 22652 21335 22704 21344
rect 22652 21301 22661 21335
rect 22661 21301 22695 21335
rect 22695 21301 22704 21335
rect 22652 21292 22704 21301
rect 23296 21292 23348 21344
rect 27160 21292 27212 21344
rect 27620 21292 27672 21344
rect 29552 21292 29604 21344
rect 29828 21335 29880 21344
rect 29828 21301 29837 21335
rect 29837 21301 29871 21335
rect 29871 21301 29880 21335
rect 29828 21292 29880 21301
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 3884 21131 3936 21140
rect 3884 21097 3893 21131
rect 3893 21097 3927 21131
rect 3927 21097 3936 21131
rect 3884 21088 3936 21097
rect 4068 21088 4120 21140
rect 4528 21088 4580 21140
rect 6000 21131 6052 21140
rect 6000 21097 6009 21131
rect 6009 21097 6043 21131
rect 6043 21097 6052 21131
rect 6000 21088 6052 21097
rect 6920 21131 6972 21140
rect 6920 21097 6929 21131
rect 6929 21097 6963 21131
rect 6963 21097 6972 21131
rect 6920 21088 6972 21097
rect 7564 21088 7616 21140
rect 9404 21088 9456 21140
rect 12624 21131 12676 21140
rect 12624 21097 12633 21131
rect 12633 21097 12667 21131
rect 12667 21097 12676 21131
rect 12624 21088 12676 21097
rect 14832 21088 14884 21140
rect 15108 21088 15160 21140
rect 15384 21088 15436 21140
rect 16028 21088 16080 21140
rect 16764 21088 16816 21140
rect 22376 21088 22428 21140
rect 3148 21063 3200 21072
rect 3148 21029 3157 21063
rect 3157 21029 3191 21063
rect 3191 21029 3200 21063
rect 3148 21020 3200 21029
rect 1860 20952 1912 21004
rect 1952 20884 2004 20936
rect 4896 20952 4948 21004
rect 6276 21020 6328 21072
rect 8208 21020 8260 21072
rect 9220 21020 9272 21072
rect 9864 21063 9916 21072
rect 9864 21029 9873 21063
rect 9873 21029 9907 21063
rect 9907 21029 9916 21063
rect 9864 21020 9916 21029
rect 10324 21020 10376 21072
rect 10508 21020 10560 21072
rect 14648 21063 14700 21072
rect 14648 21029 14657 21063
rect 14657 21029 14691 21063
rect 14691 21029 14700 21063
rect 14648 21020 14700 21029
rect 24492 21088 24544 21140
rect 25964 21088 26016 21140
rect 26700 21131 26752 21140
rect 26700 21097 26709 21131
rect 26709 21097 26743 21131
rect 26743 21097 26752 21131
rect 26700 21088 26752 21097
rect 30472 21088 30524 21140
rect 28816 21020 28868 21072
rect 33324 21063 33376 21072
rect 33324 21029 33333 21063
rect 33333 21029 33367 21063
rect 33367 21029 33376 21063
rect 33324 21020 33376 21029
rect 5632 20995 5684 21004
rect 5632 20961 5641 20995
rect 5641 20961 5675 20995
rect 5675 20961 5684 20995
rect 6184 20995 6236 21004
rect 5632 20952 5684 20961
rect 6184 20961 6193 20995
rect 6193 20961 6227 20995
rect 6227 20961 6236 20995
rect 6184 20952 6236 20961
rect 7656 20952 7708 21004
rect 11060 20952 11112 21004
rect 11428 20995 11480 21004
rect 11428 20961 11437 20995
rect 11437 20961 11471 20995
rect 11471 20961 11480 20995
rect 11428 20952 11480 20961
rect 13912 20995 13964 21004
rect 13912 20961 13921 20995
rect 13921 20961 13955 20995
rect 13955 20961 13964 20995
rect 13912 20952 13964 20961
rect 14188 20995 14240 21004
rect 14188 20961 14197 20995
rect 14197 20961 14231 20995
rect 14231 20961 14240 20995
rect 14188 20952 14240 20961
rect 15384 20952 15436 21004
rect 17224 20995 17276 21004
rect 17224 20961 17233 20995
rect 17233 20961 17267 20995
rect 17267 20961 17276 20995
rect 17224 20952 17276 20961
rect 17592 20995 17644 21004
rect 17592 20961 17601 20995
rect 17601 20961 17635 20995
rect 17635 20961 17644 20995
rect 17592 20952 17644 20961
rect 18328 20952 18380 21004
rect 18604 20995 18656 21004
rect 18604 20961 18613 20995
rect 18613 20961 18647 20995
rect 18647 20961 18656 20995
rect 18604 20952 18656 20961
rect 20628 20952 20680 21004
rect 22652 20995 22704 21004
rect 22652 20961 22661 20995
rect 22661 20961 22695 20995
rect 22695 20961 22704 20995
rect 22652 20952 22704 20961
rect 23020 20952 23072 21004
rect 24676 20952 24728 21004
rect 26424 20952 26476 21004
rect 28448 20995 28500 21004
rect 28448 20961 28457 20995
rect 28457 20961 28491 20995
rect 28491 20961 28500 20995
rect 28448 20952 28500 20961
rect 28540 20952 28592 21004
rect 29092 20952 29144 21004
rect 29828 20952 29880 21004
rect 30656 20952 30708 21004
rect 32496 20952 32548 21004
rect 33048 20995 33100 21004
rect 33048 20961 33057 20995
rect 33057 20961 33091 20995
rect 33091 20961 33100 20995
rect 33048 20952 33100 20961
rect 35256 21088 35308 21140
rect 36268 21131 36320 21140
rect 36268 21097 36277 21131
rect 36277 21097 36311 21131
rect 36311 21097 36320 21131
rect 36268 21088 36320 21097
rect 5264 20884 5316 20936
rect 7104 20927 7156 20936
rect 7104 20893 7113 20927
rect 7113 20893 7147 20927
rect 7147 20893 7156 20927
rect 7104 20884 7156 20893
rect 7012 20816 7064 20868
rect 9128 20884 9180 20936
rect 9404 20884 9456 20936
rect 10508 20884 10560 20936
rect 13360 20927 13412 20936
rect 13360 20893 13369 20927
rect 13369 20893 13403 20927
rect 13403 20893 13412 20927
rect 13360 20884 13412 20893
rect 13820 20816 13872 20868
rect 14740 20884 14792 20936
rect 16948 20884 17000 20936
rect 21640 20927 21692 20936
rect 21640 20893 21649 20927
rect 21649 20893 21683 20927
rect 21683 20893 21692 20927
rect 21640 20884 21692 20893
rect 22376 20927 22428 20936
rect 22376 20893 22385 20927
rect 22385 20893 22419 20927
rect 22419 20893 22428 20927
rect 22376 20884 22428 20893
rect 24032 20884 24084 20936
rect 24768 20927 24820 20936
rect 24768 20893 24777 20927
rect 24777 20893 24811 20927
rect 24811 20893 24820 20927
rect 24768 20884 24820 20893
rect 25228 20927 25280 20936
rect 25228 20893 25237 20927
rect 25237 20893 25271 20927
rect 25271 20893 25280 20927
rect 25228 20884 25280 20893
rect 20260 20816 20312 20868
rect 23112 20859 23164 20868
rect 23112 20825 23121 20859
rect 23121 20825 23155 20859
rect 23155 20825 23164 20859
rect 23112 20816 23164 20825
rect 27620 20816 27672 20868
rect 5448 20748 5500 20800
rect 5816 20748 5868 20800
rect 7288 20748 7340 20800
rect 8392 20748 8444 20800
rect 9128 20748 9180 20800
rect 10324 20748 10376 20800
rect 12164 20748 12216 20800
rect 13360 20748 13412 20800
rect 13544 20748 13596 20800
rect 15844 20791 15896 20800
rect 15844 20757 15853 20791
rect 15853 20757 15887 20791
rect 15887 20757 15896 20791
rect 15844 20748 15896 20757
rect 18788 20748 18840 20800
rect 19064 20748 19116 20800
rect 20076 20791 20128 20800
rect 20076 20757 20085 20791
rect 20085 20757 20119 20791
rect 20119 20757 20128 20791
rect 20076 20748 20128 20757
rect 20444 20748 20496 20800
rect 22284 20748 22336 20800
rect 25688 20748 25740 20800
rect 27804 20748 27856 20800
rect 32312 20927 32364 20936
rect 32312 20893 32321 20927
rect 32321 20893 32355 20927
rect 32355 20893 32364 20927
rect 32312 20884 32364 20893
rect 35256 20884 35308 20936
rect 28724 20816 28776 20868
rect 30472 20791 30524 20800
rect 30472 20757 30481 20791
rect 30481 20757 30515 20791
rect 30515 20757 30524 20791
rect 30472 20748 30524 20757
rect 31300 20791 31352 20800
rect 31300 20757 31309 20791
rect 31309 20757 31343 20791
rect 31343 20757 31352 20791
rect 31300 20748 31352 20757
rect 32128 20748 32180 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 3516 20544 3568 20596
rect 4620 20587 4672 20596
rect 4620 20553 4629 20587
rect 4629 20553 4663 20587
rect 4663 20553 4672 20587
rect 4620 20544 4672 20553
rect 5264 20587 5316 20596
rect 5264 20553 5273 20587
rect 5273 20553 5307 20587
rect 5307 20553 5316 20587
rect 5264 20544 5316 20553
rect 4896 20476 4948 20528
rect 2412 20451 2464 20460
rect 2412 20417 2421 20451
rect 2421 20417 2455 20451
rect 2455 20417 2464 20451
rect 2412 20408 2464 20417
rect 3148 20451 3200 20460
rect 3148 20417 3157 20451
rect 3157 20417 3191 20451
rect 3191 20417 3200 20451
rect 3148 20408 3200 20417
rect 3240 20408 3292 20460
rect 3516 20408 3568 20460
rect 3056 20383 3108 20392
rect 3056 20349 3065 20383
rect 3065 20349 3099 20383
rect 3099 20349 3108 20383
rect 3056 20340 3108 20349
rect 3700 20272 3752 20324
rect 4896 20340 4948 20392
rect 6092 20544 6144 20596
rect 6920 20544 6972 20596
rect 7104 20587 7156 20596
rect 7104 20553 7113 20587
rect 7113 20553 7147 20587
rect 7147 20553 7156 20587
rect 7104 20544 7156 20553
rect 9404 20544 9456 20596
rect 9864 20587 9916 20596
rect 9864 20553 9873 20587
rect 9873 20553 9907 20587
rect 9907 20553 9916 20587
rect 9864 20544 9916 20553
rect 12440 20544 12492 20596
rect 12716 20544 12768 20596
rect 13820 20544 13872 20596
rect 16948 20544 17000 20596
rect 17224 20544 17276 20596
rect 18972 20587 19024 20596
rect 18972 20553 18981 20587
rect 18981 20553 19015 20587
rect 19015 20553 19024 20587
rect 18972 20544 19024 20553
rect 22376 20587 22428 20596
rect 22376 20553 22385 20587
rect 22385 20553 22419 20587
rect 22419 20553 22428 20587
rect 22376 20544 22428 20553
rect 22744 20544 22796 20596
rect 24676 20587 24728 20596
rect 24676 20553 24685 20587
rect 24685 20553 24719 20587
rect 24719 20553 24728 20587
rect 24676 20544 24728 20553
rect 26424 20544 26476 20596
rect 28448 20587 28500 20596
rect 28448 20553 28457 20587
rect 28457 20553 28491 20587
rect 28491 20553 28500 20587
rect 28448 20544 28500 20553
rect 30656 20587 30708 20596
rect 8668 20519 8720 20528
rect 8668 20485 8677 20519
rect 8677 20485 8711 20519
rect 8711 20485 8720 20519
rect 8668 20476 8720 20485
rect 7932 20451 7984 20460
rect 7932 20417 7941 20451
rect 7941 20417 7975 20451
rect 7975 20417 7984 20451
rect 7932 20408 7984 20417
rect 9588 20476 9640 20528
rect 10600 20519 10652 20528
rect 10600 20485 10609 20519
rect 10609 20485 10643 20519
rect 10643 20485 10652 20519
rect 10600 20476 10652 20485
rect 10784 20519 10836 20528
rect 10784 20485 10793 20519
rect 10793 20485 10827 20519
rect 10827 20485 10836 20519
rect 10784 20476 10836 20485
rect 11428 20519 11480 20528
rect 11428 20485 11437 20519
rect 11437 20485 11471 20519
rect 11471 20485 11480 20519
rect 11428 20476 11480 20485
rect 11888 20476 11940 20528
rect 14188 20476 14240 20528
rect 15660 20519 15712 20528
rect 15660 20485 15669 20519
rect 15669 20485 15703 20519
rect 15703 20485 15712 20519
rect 15660 20476 15712 20485
rect 17592 20476 17644 20528
rect 9680 20408 9732 20460
rect 11060 20408 11112 20460
rect 17224 20408 17276 20460
rect 25964 20519 26016 20528
rect 25964 20485 25973 20519
rect 25973 20485 26007 20519
rect 26007 20485 26016 20519
rect 25964 20476 26016 20485
rect 25596 20408 25648 20460
rect 30656 20553 30665 20587
rect 30665 20553 30699 20587
rect 30699 20553 30708 20587
rect 30656 20544 30708 20553
rect 35348 20544 35400 20596
rect 29828 20476 29880 20528
rect 31852 20476 31904 20528
rect 6920 20340 6972 20392
rect 7472 20383 7524 20392
rect 7472 20349 7481 20383
rect 7481 20349 7515 20383
rect 7515 20349 7524 20383
rect 7472 20340 7524 20349
rect 9036 20340 9088 20392
rect 10508 20340 10560 20392
rect 13084 20340 13136 20392
rect 13912 20340 13964 20392
rect 15844 20383 15896 20392
rect 3240 20204 3292 20256
rect 3976 20247 4028 20256
rect 3976 20213 3985 20247
rect 3985 20213 4019 20247
rect 4019 20213 4028 20247
rect 3976 20204 4028 20213
rect 4804 20204 4856 20256
rect 7104 20272 7156 20324
rect 7288 20272 7340 20324
rect 7840 20272 7892 20324
rect 9128 20315 9180 20324
rect 7380 20204 7432 20256
rect 7656 20204 7708 20256
rect 9128 20281 9137 20315
rect 9137 20281 9171 20315
rect 9171 20281 9180 20315
rect 9128 20272 9180 20281
rect 10600 20272 10652 20324
rect 13360 20272 13412 20324
rect 15844 20349 15853 20383
rect 15853 20349 15887 20383
rect 15887 20349 15896 20383
rect 15844 20340 15896 20349
rect 16028 20383 16080 20392
rect 16028 20349 16037 20383
rect 16037 20349 16071 20383
rect 16071 20349 16080 20383
rect 16028 20340 16080 20349
rect 17132 20340 17184 20392
rect 19156 20383 19208 20392
rect 19156 20349 19165 20383
rect 19165 20349 19199 20383
rect 19199 20349 19208 20383
rect 19156 20340 19208 20349
rect 25688 20383 25740 20392
rect 20812 20315 20864 20324
rect 20812 20281 20821 20315
rect 20821 20281 20855 20315
rect 20855 20281 20864 20315
rect 20812 20272 20864 20281
rect 22560 20272 22612 20324
rect 23020 20315 23072 20324
rect 23020 20281 23029 20315
rect 23029 20281 23063 20315
rect 23063 20281 23072 20315
rect 23020 20272 23072 20281
rect 24768 20272 24820 20324
rect 25688 20349 25697 20383
rect 25697 20349 25731 20383
rect 25731 20349 25740 20383
rect 25688 20340 25740 20349
rect 25964 20383 26016 20392
rect 25964 20349 25973 20383
rect 25973 20349 26007 20383
rect 26007 20349 26016 20383
rect 25964 20340 26016 20349
rect 27620 20383 27672 20392
rect 27620 20349 27629 20383
rect 27629 20349 27663 20383
rect 27663 20349 27672 20383
rect 27620 20340 27672 20349
rect 27896 20383 27948 20392
rect 27896 20349 27905 20383
rect 27905 20349 27939 20383
rect 27939 20349 27948 20383
rect 27896 20340 27948 20349
rect 28080 20383 28132 20392
rect 28080 20349 28089 20383
rect 28089 20349 28123 20383
rect 28123 20349 28132 20383
rect 28080 20340 28132 20349
rect 29368 20383 29420 20392
rect 29368 20349 29377 20383
rect 29377 20349 29411 20383
rect 29411 20349 29420 20383
rect 29368 20340 29420 20349
rect 26148 20272 26200 20324
rect 26332 20272 26384 20324
rect 27160 20272 27212 20324
rect 29092 20272 29144 20324
rect 9312 20204 9364 20256
rect 10968 20204 11020 20256
rect 11152 20204 11204 20256
rect 11888 20204 11940 20256
rect 15384 20204 15436 20256
rect 18328 20247 18380 20256
rect 18328 20213 18337 20247
rect 18337 20213 18371 20247
rect 18371 20213 18380 20247
rect 18328 20204 18380 20213
rect 18604 20247 18656 20256
rect 18604 20213 18613 20247
rect 18613 20213 18647 20247
rect 18647 20213 18656 20247
rect 18604 20204 18656 20213
rect 20720 20204 20772 20256
rect 22100 20204 22152 20256
rect 22652 20247 22704 20256
rect 22652 20213 22661 20247
rect 22661 20213 22695 20247
rect 22695 20213 22704 20247
rect 22652 20204 22704 20213
rect 24492 20204 24544 20256
rect 31116 20247 31168 20256
rect 31116 20213 31125 20247
rect 31125 20213 31159 20247
rect 31159 20213 31168 20247
rect 31484 20340 31536 20392
rect 32496 20408 32548 20460
rect 32128 20383 32180 20392
rect 32128 20349 32137 20383
rect 32137 20349 32171 20383
rect 32171 20349 32180 20383
rect 32128 20340 32180 20349
rect 32496 20272 32548 20324
rect 31116 20204 31168 20213
rect 32312 20204 32364 20256
rect 35164 20247 35216 20256
rect 35164 20213 35173 20247
rect 35173 20213 35207 20247
rect 35207 20213 35216 20247
rect 35164 20204 35216 20213
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 1952 20043 2004 20052
rect 1952 20009 1961 20043
rect 1961 20009 1995 20043
rect 1995 20009 2004 20043
rect 1952 20000 2004 20009
rect 2688 20000 2740 20052
rect 3056 20000 3108 20052
rect 3516 20043 3568 20052
rect 3516 20009 3525 20043
rect 3525 20009 3559 20043
rect 3559 20009 3568 20043
rect 3516 20000 3568 20009
rect 4620 20043 4672 20052
rect 4620 20009 4629 20043
rect 4629 20009 4663 20043
rect 4663 20009 4672 20043
rect 4620 20000 4672 20009
rect 5172 20000 5224 20052
rect 6184 20043 6236 20052
rect 6184 20009 6193 20043
rect 6193 20009 6227 20043
rect 6227 20009 6236 20043
rect 6184 20000 6236 20009
rect 6920 20000 6972 20052
rect 7840 20000 7892 20052
rect 8300 20043 8352 20052
rect 8300 20009 8309 20043
rect 8309 20009 8343 20043
rect 8343 20009 8352 20043
rect 8300 20000 8352 20009
rect 9404 20043 9456 20052
rect 9404 20009 9413 20043
rect 9413 20009 9447 20043
rect 9447 20009 9456 20043
rect 9404 20000 9456 20009
rect 10048 20000 10100 20052
rect 13544 20000 13596 20052
rect 13820 20000 13872 20052
rect 19156 20043 19208 20052
rect 19156 20009 19165 20043
rect 19165 20009 19199 20043
rect 19199 20009 19208 20043
rect 19156 20000 19208 20009
rect 24400 20000 24452 20052
rect 24676 20000 24728 20052
rect 25964 20000 26016 20052
rect 26332 20043 26384 20052
rect 26332 20009 26341 20043
rect 26341 20009 26375 20043
rect 26375 20009 26384 20043
rect 26332 20000 26384 20009
rect 27620 20043 27672 20052
rect 27620 20009 27629 20043
rect 27629 20009 27663 20043
rect 27663 20009 27672 20043
rect 27620 20000 27672 20009
rect 29092 20000 29144 20052
rect 31484 20043 31536 20052
rect 31484 20009 31493 20043
rect 31493 20009 31527 20043
rect 31527 20009 31536 20043
rect 31484 20000 31536 20009
rect 1860 19932 1912 19984
rect 3148 19932 3200 19984
rect 5264 19975 5316 19984
rect 5264 19941 5273 19975
rect 5273 19941 5307 19975
rect 5307 19941 5316 19975
rect 5264 19932 5316 19941
rect 5908 19932 5960 19984
rect 7380 19932 7432 19984
rect 7932 19932 7984 19984
rect 11612 19975 11664 19984
rect 11612 19941 11621 19975
rect 11621 19941 11655 19975
rect 11655 19941 11664 19975
rect 11612 19932 11664 19941
rect 15844 19975 15896 19984
rect 15844 19941 15853 19975
rect 15853 19941 15887 19975
rect 15887 19941 15896 19975
rect 15844 19932 15896 19941
rect 25688 19932 25740 19984
rect 5540 19864 5592 19916
rect 6184 19864 6236 19916
rect 7564 19907 7616 19916
rect 7288 19839 7340 19848
rect 7288 19805 7297 19839
rect 7297 19805 7331 19839
rect 7331 19805 7340 19839
rect 7288 19796 7340 19805
rect 7564 19873 7573 19907
rect 7573 19873 7607 19907
rect 7607 19873 7616 19907
rect 7564 19864 7616 19873
rect 10784 19864 10836 19916
rect 12348 19864 12400 19916
rect 12716 19864 12768 19916
rect 13912 19907 13964 19916
rect 13912 19873 13921 19907
rect 13921 19873 13955 19907
rect 13955 19873 13964 19907
rect 13912 19864 13964 19873
rect 15384 19907 15436 19916
rect 15384 19873 15393 19907
rect 15393 19873 15427 19907
rect 15427 19873 15436 19907
rect 15384 19864 15436 19873
rect 16948 19907 17000 19916
rect 16948 19873 16957 19907
rect 16957 19873 16991 19907
rect 16991 19873 17000 19907
rect 16948 19864 17000 19873
rect 17132 19864 17184 19916
rect 17408 19907 17460 19916
rect 17408 19873 17417 19907
rect 17417 19873 17451 19907
rect 17451 19873 17460 19907
rect 17408 19864 17460 19873
rect 17592 19864 17644 19916
rect 22100 19907 22152 19916
rect 22100 19873 22109 19907
rect 22109 19873 22143 19907
rect 22143 19873 22152 19907
rect 22100 19864 22152 19873
rect 22560 19864 22612 19916
rect 24032 19907 24084 19916
rect 24032 19873 24041 19907
rect 24041 19873 24075 19907
rect 24075 19873 24084 19907
rect 24032 19864 24084 19873
rect 24400 19907 24452 19916
rect 24400 19873 24409 19907
rect 24409 19873 24443 19907
rect 24443 19873 24452 19907
rect 24400 19864 24452 19873
rect 25228 19864 25280 19916
rect 27436 19864 27488 19916
rect 32496 19932 32548 19984
rect 10140 19796 10192 19848
rect 6460 19728 6512 19780
rect 10508 19796 10560 19848
rect 12164 19839 12216 19848
rect 12164 19805 12173 19839
rect 12173 19805 12207 19839
rect 12207 19805 12216 19839
rect 12164 19796 12216 19805
rect 12532 19796 12584 19848
rect 14556 19796 14608 19848
rect 15292 19839 15344 19848
rect 15292 19805 15301 19839
rect 15301 19805 15335 19839
rect 15335 19805 15344 19839
rect 21732 19839 21784 19848
rect 15292 19796 15344 19805
rect 12808 19728 12860 19780
rect 15660 19728 15712 19780
rect 3884 19703 3936 19712
rect 3884 19669 3893 19703
rect 3893 19669 3927 19703
rect 3927 19669 3936 19703
rect 3884 19660 3936 19669
rect 5264 19660 5316 19712
rect 7196 19660 7248 19712
rect 9036 19660 9088 19712
rect 9864 19660 9916 19712
rect 11060 19703 11112 19712
rect 11060 19669 11069 19703
rect 11069 19669 11103 19703
rect 11103 19669 11112 19703
rect 11060 19660 11112 19669
rect 13084 19660 13136 19712
rect 13636 19660 13688 19712
rect 14648 19703 14700 19712
rect 14648 19669 14657 19703
rect 14657 19669 14691 19703
rect 14691 19669 14700 19703
rect 14648 19660 14700 19669
rect 15476 19660 15528 19712
rect 16212 19703 16264 19712
rect 16212 19669 16221 19703
rect 16221 19669 16255 19703
rect 16255 19669 16264 19703
rect 16212 19660 16264 19669
rect 21732 19805 21741 19839
rect 21741 19805 21775 19839
rect 21775 19805 21784 19839
rect 21732 19796 21784 19805
rect 23940 19796 23992 19848
rect 28816 19864 28868 19916
rect 30012 19864 30064 19916
rect 30104 19907 30156 19916
rect 30104 19873 30113 19907
rect 30113 19873 30147 19907
rect 30147 19873 30156 19907
rect 30104 19864 30156 19873
rect 33140 19907 33192 19916
rect 28724 19796 28776 19848
rect 30196 19796 30248 19848
rect 33140 19873 33149 19907
rect 33149 19873 33183 19907
rect 33183 19873 33192 19907
rect 33140 19864 33192 19873
rect 34428 19932 34480 19984
rect 33968 19907 34020 19916
rect 33968 19873 33977 19907
rect 33977 19873 34011 19907
rect 34011 19873 34020 19907
rect 33968 19864 34020 19873
rect 35900 19907 35952 19916
rect 35900 19873 35909 19907
rect 35909 19873 35943 19907
rect 35943 19873 35952 19907
rect 35900 19864 35952 19873
rect 32128 19796 32180 19848
rect 33048 19796 33100 19848
rect 35624 19839 35676 19848
rect 35624 19805 35633 19839
rect 35633 19805 35667 19839
rect 35667 19805 35676 19839
rect 35624 19796 35676 19805
rect 36084 19839 36136 19848
rect 36084 19805 36093 19839
rect 36093 19805 36127 19839
rect 36127 19805 36136 19839
rect 36084 19796 36136 19805
rect 17316 19728 17368 19780
rect 22008 19728 22060 19780
rect 24308 19771 24360 19780
rect 24308 19737 24317 19771
rect 24317 19737 24351 19771
rect 24351 19737 24360 19771
rect 24308 19728 24360 19737
rect 26056 19728 26108 19780
rect 30288 19771 30340 19780
rect 30288 19737 30297 19771
rect 30297 19737 30331 19771
rect 30331 19737 30340 19771
rect 30288 19728 30340 19737
rect 17408 19660 17460 19712
rect 18420 19703 18472 19712
rect 18420 19669 18429 19703
rect 18429 19669 18463 19703
rect 18463 19669 18472 19703
rect 18420 19660 18472 19669
rect 19892 19660 19944 19712
rect 26792 19703 26844 19712
rect 26792 19669 26801 19703
rect 26801 19669 26835 19703
rect 26835 19669 26844 19703
rect 26792 19660 26844 19669
rect 27068 19703 27120 19712
rect 27068 19669 27077 19703
rect 27077 19669 27111 19703
rect 27111 19669 27120 19703
rect 27068 19660 27120 19669
rect 29368 19703 29420 19712
rect 29368 19669 29377 19703
rect 29377 19669 29411 19703
rect 29411 19669 29420 19703
rect 29368 19660 29420 19669
rect 31484 19660 31536 19712
rect 33048 19703 33100 19712
rect 33048 19669 33057 19703
rect 33057 19669 33091 19703
rect 33091 19669 33100 19703
rect 33048 19660 33100 19669
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 1952 19456 2004 19508
rect 3700 19499 3752 19508
rect 3700 19465 3709 19499
rect 3709 19465 3743 19499
rect 3743 19465 3752 19499
rect 3700 19456 3752 19465
rect 7840 19499 7892 19508
rect 7840 19465 7849 19499
rect 7849 19465 7883 19499
rect 7883 19465 7892 19499
rect 7840 19456 7892 19465
rect 8668 19456 8720 19508
rect 10140 19499 10192 19508
rect 3424 19320 3476 19372
rect 5264 19320 5316 19372
rect 5540 19320 5592 19372
rect 6460 19320 6512 19372
rect 10140 19465 10149 19499
rect 10149 19465 10183 19499
rect 10183 19465 10192 19499
rect 10140 19456 10192 19465
rect 12716 19456 12768 19508
rect 13084 19499 13136 19508
rect 13084 19465 13093 19499
rect 13093 19465 13127 19499
rect 13127 19465 13136 19499
rect 13084 19456 13136 19465
rect 16212 19456 16264 19508
rect 11428 19388 11480 19440
rect 12072 19388 12124 19440
rect 16028 19388 16080 19440
rect 16304 19388 16356 19440
rect 5080 19252 5132 19304
rect 4896 19184 4948 19236
rect 5172 19227 5224 19236
rect 5172 19193 5181 19227
rect 5181 19193 5215 19227
rect 5215 19193 5224 19227
rect 5172 19184 5224 19193
rect 5264 19184 5316 19236
rect 7288 19252 7340 19304
rect 12440 19320 12492 19372
rect 15936 19320 15988 19372
rect 9036 19252 9088 19304
rect 11336 19252 11388 19304
rect 12348 19252 12400 19304
rect 12624 19252 12676 19304
rect 12808 19295 12860 19304
rect 12808 19261 12817 19295
rect 12817 19261 12851 19295
rect 12851 19261 12860 19295
rect 12808 19252 12860 19261
rect 12900 19295 12952 19304
rect 12900 19261 12909 19295
rect 12909 19261 12943 19295
rect 12943 19261 12952 19295
rect 14188 19295 14240 19304
rect 12900 19252 12952 19261
rect 14188 19261 14197 19295
rect 14197 19261 14231 19295
rect 14231 19261 14240 19295
rect 14188 19252 14240 19261
rect 14740 19295 14792 19304
rect 7196 19227 7248 19236
rect 7196 19193 7205 19227
rect 7205 19193 7239 19227
rect 7239 19193 7248 19227
rect 7196 19184 7248 19193
rect 8300 19227 8352 19236
rect 8300 19193 8309 19227
rect 8309 19193 8343 19227
rect 8343 19193 8352 19227
rect 8300 19184 8352 19193
rect 9220 19184 9272 19236
rect 9864 19227 9916 19236
rect 9864 19193 9873 19227
rect 9873 19193 9907 19227
rect 9907 19193 9916 19227
rect 9864 19184 9916 19193
rect 11612 19184 11664 19236
rect 12532 19184 12584 19236
rect 4804 19116 4856 19168
rect 7012 19159 7064 19168
rect 7012 19125 7021 19159
rect 7021 19125 7055 19159
rect 7055 19125 7064 19159
rect 7012 19116 7064 19125
rect 7104 19159 7156 19168
rect 7104 19125 7113 19159
rect 7113 19125 7147 19159
rect 7147 19125 7156 19159
rect 7104 19116 7156 19125
rect 9404 19159 9456 19168
rect 9404 19125 9413 19159
rect 9413 19125 9447 19159
rect 9447 19125 9456 19159
rect 9404 19116 9456 19125
rect 10692 19159 10744 19168
rect 10692 19125 10701 19159
rect 10701 19125 10735 19159
rect 10735 19125 10744 19159
rect 10692 19116 10744 19125
rect 11060 19159 11112 19168
rect 11060 19125 11069 19159
rect 11069 19125 11103 19159
rect 11103 19125 11112 19159
rect 11060 19116 11112 19125
rect 12440 19116 12492 19168
rect 14096 19184 14148 19236
rect 14740 19261 14749 19295
rect 14749 19261 14783 19295
rect 14783 19261 14792 19295
rect 14740 19252 14792 19261
rect 17592 19499 17644 19508
rect 17592 19465 17601 19499
rect 17601 19465 17635 19499
rect 17635 19465 17644 19499
rect 17592 19456 17644 19465
rect 21732 19499 21784 19508
rect 21732 19465 21741 19499
rect 21741 19465 21775 19499
rect 21775 19465 21784 19499
rect 21732 19456 21784 19465
rect 23296 19456 23348 19508
rect 23940 19499 23992 19508
rect 23940 19465 23949 19499
rect 23949 19465 23983 19499
rect 23983 19465 23992 19499
rect 23940 19456 23992 19465
rect 16948 19388 17000 19440
rect 24032 19388 24084 19440
rect 25688 19388 25740 19440
rect 25780 19388 25832 19440
rect 31484 19388 31536 19440
rect 19892 19320 19944 19372
rect 16948 19295 17000 19304
rect 16948 19261 16957 19295
rect 16957 19261 16991 19295
rect 16991 19261 17000 19295
rect 16948 19252 17000 19261
rect 17408 19252 17460 19304
rect 19984 19295 20036 19304
rect 17316 19227 17368 19236
rect 17316 19193 17325 19227
rect 17325 19193 17359 19227
rect 17359 19193 17368 19227
rect 17316 19184 17368 19193
rect 18788 19184 18840 19236
rect 19984 19261 19993 19295
rect 19993 19261 20027 19295
rect 20027 19261 20036 19295
rect 19984 19252 20036 19261
rect 24308 19295 24360 19304
rect 24308 19261 24317 19295
rect 24317 19261 24351 19295
rect 24351 19261 24360 19295
rect 24308 19252 24360 19261
rect 25320 19295 25372 19304
rect 25320 19261 25329 19295
rect 25329 19261 25363 19295
rect 25363 19261 25372 19295
rect 25320 19252 25372 19261
rect 25688 19295 25740 19304
rect 25688 19261 25697 19295
rect 25697 19261 25731 19295
rect 25731 19261 25740 19295
rect 25688 19252 25740 19261
rect 26056 19252 26108 19304
rect 26332 19320 26384 19372
rect 26792 19363 26844 19372
rect 26792 19329 26801 19363
rect 26801 19329 26835 19363
rect 26835 19329 26844 19363
rect 26792 19320 26844 19329
rect 27436 19252 27488 19304
rect 28724 19320 28776 19372
rect 30012 19320 30064 19372
rect 21364 19227 21416 19236
rect 21364 19193 21373 19227
rect 21373 19193 21407 19227
rect 21407 19193 21416 19227
rect 21364 19184 21416 19193
rect 25228 19184 25280 19236
rect 28172 19252 28224 19304
rect 29276 19295 29328 19304
rect 29276 19261 29285 19295
rect 29285 19261 29319 19295
rect 29319 19261 29328 19295
rect 29276 19252 29328 19261
rect 29184 19184 29236 19236
rect 13820 19159 13872 19168
rect 13820 19125 13829 19159
rect 13829 19125 13863 19159
rect 13863 19125 13872 19159
rect 13820 19116 13872 19125
rect 15476 19159 15528 19168
rect 15476 19125 15485 19159
rect 15485 19125 15519 19159
rect 15519 19125 15528 19159
rect 15476 19116 15528 19125
rect 17132 19116 17184 19168
rect 17408 19116 17460 19168
rect 18144 19116 18196 19168
rect 18328 19116 18380 19168
rect 22100 19159 22152 19168
rect 22100 19125 22109 19159
rect 22109 19125 22143 19159
rect 22143 19125 22152 19159
rect 22100 19116 22152 19125
rect 22560 19116 22612 19168
rect 23112 19159 23164 19168
rect 23112 19125 23121 19159
rect 23121 19125 23155 19159
rect 23155 19125 23164 19159
rect 23112 19116 23164 19125
rect 25964 19116 26016 19168
rect 28080 19116 28132 19168
rect 28632 19159 28684 19168
rect 28632 19125 28641 19159
rect 28641 19125 28675 19159
rect 28675 19125 28684 19159
rect 28632 19116 28684 19125
rect 29276 19116 29328 19168
rect 30104 19184 30156 19236
rect 33968 19388 34020 19440
rect 32036 19363 32088 19372
rect 32036 19329 32045 19363
rect 32045 19329 32079 19363
rect 32079 19329 32088 19363
rect 32036 19320 32088 19329
rect 32956 19363 33008 19372
rect 32956 19329 32965 19363
rect 32965 19329 32999 19363
rect 32999 19329 33008 19363
rect 32956 19320 33008 19329
rect 31668 19184 31720 19236
rect 30288 19116 30340 19168
rect 30932 19159 30984 19168
rect 30932 19125 30941 19159
rect 30941 19125 30975 19159
rect 30975 19125 30984 19159
rect 30932 19116 30984 19125
rect 32496 19159 32548 19168
rect 32496 19125 32505 19159
rect 32505 19125 32539 19159
rect 32539 19125 32548 19159
rect 32496 19116 32548 19125
rect 32588 19116 32640 19168
rect 33140 19320 33192 19372
rect 33508 19295 33560 19304
rect 33508 19261 33517 19295
rect 33517 19261 33551 19295
rect 33551 19261 33560 19295
rect 33508 19252 33560 19261
rect 33784 19295 33836 19304
rect 33784 19261 33793 19295
rect 33793 19261 33827 19295
rect 33827 19261 33836 19295
rect 33784 19252 33836 19261
rect 33876 19252 33928 19304
rect 36084 19320 36136 19372
rect 35624 19184 35676 19236
rect 33140 19116 33192 19168
rect 33784 19116 33836 19168
rect 34428 19116 34480 19168
rect 35072 19159 35124 19168
rect 35072 19125 35081 19159
rect 35081 19125 35115 19159
rect 35115 19125 35124 19159
rect 35072 19116 35124 19125
rect 35900 19116 35952 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 3516 18955 3568 18964
rect 3516 18921 3525 18955
rect 3525 18921 3559 18955
rect 3559 18921 3568 18955
rect 3516 18912 3568 18921
rect 5448 18912 5500 18964
rect 6184 18955 6236 18964
rect 6184 18921 6193 18955
rect 6193 18921 6227 18955
rect 6227 18921 6236 18955
rect 6184 18912 6236 18921
rect 6460 18955 6512 18964
rect 6460 18921 6469 18955
rect 6469 18921 6503 18955
rect 6503 18921 6512 18955
rect 6460 18912 6512 18921
rect 6920 18912 6972 18964
rect 8760 18955 8812 18964
rect 8760 18921 8769 18955
rect 8769 18921 8803 18955
rect 8803 18921 8812 18955
rect 8760 18912 8812 18921
rect 5172 18887 5224 18896
rect 5172 18853 5181 18887
rect 5181 18853 5215 18887
rect 5215 18853 5224 18887
rect 5172 18844 5224 18853
rect 7472 18844 7524 18896
rect 10048 18844 10100 18896
rect 11060 18912 11112 18964
rect 11704 18955 11756 18964
rect 11704 18921 11713 18955
rect 11713 18921 11747 18955
rect 11747 18921 11756 18955
rect 11704 18912 11756 18921
rect 12164 18912 12216 18964
rect 13636 18912 13688 18964
rect 14648 18955 14700 18964
rect 14648 18921 14657 18955
rect 14657 18921 14691 18955
rect 14691 18921 14700 18955
rect 14648 18912 14700 18921
rect 16028 18912 16080 18964
rect 16212 18955 16264 18964
rect 16212 18921 16221 18955
rect 16221 18921 16255 18955
rect 16255 18921 16264 18955
rect 16212 18912 16264 18921
rect 17592 18912 17644 18964
rect 17684 18912 17736 18964
rect 18604 18912 18656 18964
rect 21364 18912 21416 18964
rect 23480 18912 23532 18964
rect 24308 18912 24360 18964
rect 26056 18912 26108 18964
rect 26240 18912 26292 18964
rect 26976 18955 27028 18964
rect 26976 18921 26985 18955
rect 26985 18921 27019 18955
rect 27019 18921 27028 18955
rect 26976 18912 27028 18921
rect 27712 18912 27764 18964
rect 30104 18912 30156 18964
rect 30196 18912 30248 18964
rect 31208 18912 31260 18964
rect 32956 18912 33008 18964
rect 10600 18844 10652 18896
rect 10784 18887 10836 18896
rect 10784 18853 10793 18887
rect 10793 18853 10827 18887
rect 10827 18853 10836 18887
rect 10784 18844 10836 18853
rect 15844 18844 15896 18896
rect 1676 18819 1728 18828
rect 1676 18785 1685 18819
rect 1685 18785 1719 18819
rect 1719 18785 1728 18819
rect 1676 18776 1728 18785
rect 1952 18776 2004 18828
rect 5632 18819 5684 18828
rect 5632 18785 5641 18819
rect 5641 18785 5675 18819
rect 5675 18785 5684 18819
rect 5632 18776 5684 18785
rect 7012 18776 7064 18828
rect 7380 18776 7432 18828
rect 7932 18819 7984 18828
rect 7932 18785 7941 18819
rect 7941 18785 7975 18819
rect 7975 18785 7984 18819
rect 7932 18776 7984 18785
rect 10692 18776 10744 18828
rect 8668 18708 8720 18760
rect 9220 18708 9272 18760
rect 9496 18708 9548 18760
rect 12440 18819 12492 18828
rect 12440 18785 12449 18819
rect 12449 18785 12483 18819
rect 12483 18785 12492 18819
rect 12440 18776 12492 18785
rect 12716 18776 12768 18828
rect 14280 18776 14332 18828
rect 16028 18776 16080 18828
rect 23112 18844 23164 18896
rect 4436 18683 4488 18692
rect 4436 18649 4445 18683
rect 4445 18649 4479 18683
rect 4479 18649 4488 18683
rect 4436 18640 4488 18649
rect 5448 18640 5500 18692
rect 6552 18640 6604 18692
rect 7196 18640 7248 18692
rect 8944 18640 8996 18692
rect 9404 18640 9456 18692
rect 9956 18640 10008 18692
rect 10600 18640 10652 18692
rect 10968 18640 11020 18692
rect 2596 18572 2648 18624
rect 3148 18572 3200 18624
rect 6460 18572 6512 18624
rect 7564 18572 7616 18624
rect 8116 18615 8168 18624
rect 8116 18581 8125 18615
rect 8125 18581 8159 18615
rect 8159 18581 8168 18615
rect 8116 18572 8168 18581
rect 9036 18572 9088 18624
rect 12532 18708 12584 18760
rect 17960 18776 18012 18828
rect 23940 18776 23992 18828
rect 25688 18844 25740 18896
rect 27436 18844 27488 18896
rect 27804 18887 27856 18896
rect 27804 18853 27813 18887
rect 27813 18853 27847 18887
rect 27847 18853 27856 18887
rect 27804 18844 27856 18853
rect 24400 18776 24452 18828
rect 18420 18708 18472 18760
rect 23204 18708 23256 18760
rect 24308 18708 24360 18760
rect 12808 18683 12860 18692
rect 12808 18649 12817 18683
rect 12817 18649 12851 18683
rect 12851 18649 12860 18683
rect 12808 18640 12860 18649
rect 14004 18640 14056 18692
rect 17500 18640 17552 18692
rect 23940 18683 23992 18692
rect 23940 18649 23949 18683
rect 23949 18649 23983 18683
rect 23983 18649 23992 18683
rect 23940 18640 23992 18649
rect 25596 18640 25648 18692
rect 26976 18776 27028 18828
rect 28172 18819 28224 18828
rect 28172 18785 28181 18819
rect 28181 18785 28215 18819
rect 28215 18785 28224 18819
rect 28172 18776 28224 18785
rect 28724 18776 28776 18828
rect 34060 18887 34112 18896
rect 34060 18853 34069 18887
rect 34069 18853 34103 18887
rect 34103 18853 34112 18887
rect 34060 18844 34112 18853
rect 33508 18819 33560 18828
rect 33508 18785 33517 18819
rect 33517 18785 33551 18819
rect 33551 18785 33560 18819
rect 33508 18776 33560 18785
rect 33784 18819 33836 18828
rect 33784 18785 33793 18819
rect 33793 18785 33827 18819
rect 33827 18785 33836 18819
rect 33784 18776 33836 18785
rect 29092 18751 29144 18760
rect 29092 18717 29101 18751
rect 29101 18717 29135 18751
rect 29135 18717 29144 18751
rect 29092 18708 29144 18717
rect 33048 18751 33100 18760
rect 33048 18717 33057 18751
rect 33057 18717 33091 18751
rect 33091 18717 33100 18751
rect 33048 18708 33100 18717
rect 26148 18640 26200 18692
rect 11336 18572 11388 18624
rect 13544 18572 13596 18624
rect 13912 18572 13964 18624
rect 14556 18572 14608 18624
rect 15384 18572 15436 18624
rect 16948 18572 17000 18624
rect 17132 18572 17184 18624
rect 17592 18615 17644 18624
rect 17592 18581 17601 18615
rect 17601 18581 17635 18615
rect 17635 18581 17644 18615
rect 17592 18572 17644 18581
rect 18788 18572 18840 18624
rect 19708 18615 19760 18624
rect 19708 18581 19717 18615
rect 19717 18581 19751 18615
rect 19751 18581 19760 18615
rect 19708 18572 19760 18581
rect 27620 18572 27672 18624
rect 30288 18572 30340 18624
rect 30656 18615 30708 18624
rect 30656 18581 30665 18615
rect 30665 18581 30699 18615
rect 30699 18581 30708 18615
rect 30656 18572 30708 18581
rect 30932 18572 30984 18624
rect 31668 18572 31720 18624
rect 32588 18572 32640 18624
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 1676 18411 1728 18420
rect 1676 18377 1685 18411
rect 1685 18377 1719 18411
rect 1719 18377 1728 18411
rect 1676 18368 1728 18377
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 4620 18368 4672 18420
rect 4896 18411 4948 18420
rect 4896 18377 4905 18411
rect 4905 18377 4939 18411
rect 4939 18377 4948 18411
rect 4896 18368 4948 18377
rect 5264 18411 5316 18420
rect 5264 18377 5273 18411
rect 5273 18377 5307 18411
rect 5307 18377 5316 18411
rect 5264 18368 5316 18377
rect 5632 18411 5684 18420
rect 5632 18377 5641 18411
rect 5641 18377 5675 18411
rect 5675 18377 5684 18411
rect 5632 18368 5684 18377
rect 5908 18411 5960 18420
rect 5908 18377 5917 18411
rect 5917 18377 5951 18411
rect 5951 18377 5960 18411
rect 5908 18368 5960 18377
rect 8576 18368 8628 18420
rect 10692 18411 10744 18420
rect 6920 18300 6972 18352
rect 7012 18232 7064 18284
rect 10692 18377 10701 18411
rect 10701 18377 10735 18411
rect 10735 18377 10744 18411
rect 10692 18368 10744 18377
rect 13820 18368 13872 18420
rect 9588 18275 9640 18284
rect 9588 18241 9597 18275
rect 9597 18241 9631 18275
rect 9631 18241 9640 18275
rect 9588 18232 9640 18241
rect 11336 18275 11388 18284
rect 11336 18241 11345 18275
rect 11345 18241 11379 18275
rect 11379 18241 11388 18275
rect 11336 18232 11388 18241
rect 12532 18300 12584 18352
rect 13636 18300 13688 18352
rect 15844 18368 15896 18420
rect 17316 18368 17368 18420
rect 18328 18368 18380 18420
rect 23204 18411 23256 18420
rect 23204 18377 23213 18411
rect 23213 18377 23247 18411
rect 23247 18377 23256 18411
rect 23204 18368 23256 18377
rect 24032 18368 24084 18420
rect 24308 18411 24360 18420
rect 24308 18377 24317 18411
rect 24317 18377 24351 18411
rect 24351 18377 24360 18411
rect 24308 18368 24360 18377
rect 28724 18411 28776 18420
rect 28724 18377 28733 18411
rect 28733 18377 28767 18411
rect 28767 18377 28776 18411
rect 28724 18368 28776 18377
rect 29920 18368 29972 18420
rect 30472 18368 30524 18420
rect 33048 18368 33100 18420
rect 7196 18207 7248 18216
rect 7196 18173 7205 18207
rect 7205 18173 7239 18207
rect 7239 18173 7248 18207
rect 7196 18164 7248 18173
rect 8760 18164 8812 18216
rect 8944 18164 8996 18216
rect 9772 18164 9824 18216
rect 10508 18207 10560 18216
rect 10508 18173 10517 18207
rect 10517 18173 10551 18207
rect 10551 18173 10560 18207
rect 10508 18164 10560 18173
rect 11980 18164 12032 18216
rect 13544 18207 13596 18216
rect 13544 18173 13553 18207
rect 13553 18173 13587 18207
rect 13587 18173 13596 18207
rect 13544 18164 13596 18173
rect 13912 18207 13964 18216
rect 13912 18173 13921 18207
rect 13921 18173 13955 18207
rect 13955 18173 13964 18207
rect 13912 18164 13964 18173
rect 17960 18300 18012 18352
rect 17684 18232 17736 18284
rect 19708 18275 19760 18284
rect 19708 18241 19717 18275
rect 19717 18241 19751 18275
rect 19751 18241 19760 18275
rect 19708 18232 19760 18241
rect 20444 18232 20496 18284
rect 21824 18232 21876 18284
rect 24216 18300 24268 18352
rect 31944 18300 31996 18352
rect 32956 18300 33008 18352
rect 14740 18207 14792 18216
rect 14740 18173 14749 18207
rect 14749 18173 14783 18207
rect 14783 18173 14792 18207
rect 14740 18164 14792 18173
rect 7932 18139 7984 18148
rect 4528 18071 4580 18080
rect 4528 18037 4537 18071
rect 4537 18037 4571 18071
rect 4571 18037 4580 18071
rect 4528 18028 4580 18037
rect 6000 18028 6052 18080
rect 6460 18028 6512 18080
rect 6920 18028 6972 18080
rect 7932 18105 7941 18139
rect 7941 18105 7975 18139
rect 7975 18105 7984 18139
rect 7932 18096 7984 18105
rect 9220 18139 9272 18148
rect 8208 18028 8260 18080
rect 8668 18028 8720 18080
rect 9220 18105 9229 18139
rect 9229 18105 9263 18139
rect 9263 18105 9272 18139
rect 9220 18096 9272 18105
rect 10784 18096 10836 18148
rect 13268 18139 13320 18148
rect 13268 18105 13277 18139
rect 13277 18105 13311 18139
rect 13311 18105 13320 18139
rect 13268 18096 13320 18105
rect 14188 18096 14240 18148
rect 16948 18164 17000 18216
rect 9036 18071 9088 18080
rect 9036 18037 9045 18071
rect 9045 18037 9079 18071
rect 9079 18037 9088 18071
rect 9036 18028 9088 18037
rect 9588 18028 9640 18080
rect 10232 18028 10284 18080
rect 10600 18028 10652 18080
rect 17408 18164 17460 18216
rect 16028 18071 16080 18080
rect 16028 18037 16037 18071
rect 16037 18037 16071 18071
rect 16071 18037 16080 18071
rect 16028 18028 16080 18037
rect 17776 18028 17828 18080
rect 19248 18028 19300 18080
rect 19432 18028 19484 18080
rect 20628 18164 20680 18216
rect 25780 18232 25832 18284
rect 28080 18275 28132 18284
rect 28080 18241 28089 18275
rect 28089 18241 28123 18275
rect 28123 18241 28132 18275
rect 28080 18232 28132 18241
rect 28172 18232 28224 18284
rect 30840 18232 30892 18284
rect 33508 18300 33560 18352
rect 21916 18096 21968 18148
rect 22008 18028 22060 18080
rect 22100 18028 22152 18080
rect 23664 18028 23716 18080
rect 24492 18028 24544 18080
rect 25136 18207 25188 18216
rect 25136 18173 25145 18207
rect 25145 18173 25179 18207
rect 25179 18173 25188 18207
rect 25136 18164 25188 18173
rect 25688 18207 25740 18216
rect 25688 18173 25697 18207
rect 25697 18173 25731 18207
rect 25731 18173 25740 18207
rect 25688 18164 25740 18173
rect 26056 18207 26108 18216
rect 26056 18173 26065 18207
rect 26065 18173 26099 18207
rect 26099 18173 26108 18207
rect 26056 18164 26108 18173
rect 27620 18164 27672 18216
rect 28632 18164 28684 18216
rect 29920 18164 29972 18216
rect 31208 18164 31260 18216
rect 31760 18164 31812 18216
rect 27804 18096 27856 18148
rect 32220 18096 32272 18148
rect 33048 18139 33100 18148
rect 33048 18105 33057 18139
rect 33057 18105 33091 18139
rect 33091 18105 33100 18139
rect 33048 18096 33100 18105
rect 24768 18028 24820 18080
rect 26976 18028 27028 18080
rect 27436 18028 27488 18080
rect 27896 18028 27948 18080
rect 29644 18028 29696 18080
rect 31484 18028 31536 18080
rect 32772 18028 32824 18080
rect 33784 18028 33836 18080
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 1860 17867 1912 17876
rect 1860 17833 1869 17867
rect 1869 17833 1903 17867
rect 1903 17833 1912 17867
rect 1860 17824 1912 17833
rect 1952 17799 2004 17808
rect 1952 17765 1961 17799
rect 1961 17765 1995 17799
rect 1995 17765 2004 17799
rect 1952 17756 2004 17765
rect 3332 17824 3384 17876
rect 4620 17867 4672 17876
rect 4620 17833 4629 17867
rect 4629 17833 4663 17867
rect 4663 17833 4672 17867
rect 4620 17824 4672 17833
rect 5172 17867 5224 17876
rect 5172 17833 5181 17867
rect 5181 17833 5215 17867
rect 5215 17833 5224 17867
rect 5172 17824 5224 17833
rect 7012 17824 7064 17876
rect 7380 17824 7432 17876
rect 8484 17824 8536 17876
rect 11520 17867 11572 17876
rect 11520 17833 11529 17867
rect 11529 17833 11563 17867
rect 11563 17833 11572 17867
rect 11520 17824 11572 17833
rect 11704 17824 11756 17876
rect 9128 17756 9180 17808
rect 9404 17756 9456 17808
rect 2412 17731 2464 17740
rect 2412 17697 2421 17731
rect 2421 17697 2455 17731
rect 2455 17697 2464 17731
rect 2412 17688 2464 17697
rect 2504 17688 2556 17740
rect 2688 17688 2740 17740
rect 3516 17688 3568 17740
rect 5540 17731 5592 17740
rect 3240 17620 3292 17672
rect 5540 17697 5549 17731
rect 5549 17697 5583 17731
rect 5583 17697 5592 17731
rect 5540 17688 5592 17697
rect 5908 17731 5960 17740
rect 5908 17697 5917 17731
rect 5917 17697 5951 17731
rect 5951 17697 5960 17731
rect 5908 17688 5960 17697
rect 6644 17688 6696 17740
rect 8024 17731 8076 17740
rect 8024 17697 8033 17731
rect 8033 17697 8067 17731
rect 8067 17697 8076 17731
rect 8024 17688 8076 17697
rect 8208 17688 8260 17740
rect 9680 17731 9732 17740
rect 9680 17697 9689 17731
rect 9689 17697 9723 17731
rect 9723 17697 9732 17731
rect 9680 17688 9732 17697
rect 10048 17756 10100 17808
rect 11612 17799 11664 17808
rect 11612 17765 11621 17799
rect 11621 17765 11655 17799
rect 11655 17765 11664 17799
rect 11612 17756 11664 17765
rect 11980 17799 12032 17808
rect 11980 17765 11989 17799
rect 11989 17765 12023 17799
rect 12023 17765 12032 17799
rect 11980 17756 12032 17765
rect 12440 17824 12492 17876
rect 12716 17867 12768 17876
rect 12716 17833 12725 17867
rect 12725 17833 12759 17867
rect 12759 17833 12768 17867
rect 12716 17824 12768 17833
rect 12532 17756 12584 17808
rect 15384 17824 15436 17876
rect 17408 17824 17460 17876
rect 17776 17824 17828 17876
rect 17960 17824 18012 17876
rect 18420 17867 18472 17876
rect 18420 17833 18429 17867
rect 18429 17833 18463 17867
rect 18463 17833 18472 17867
rect 18420 17824 18472 17833
rect 20260 17824 20312 17876
rect 20904 17824 20956 17876
rect 22008 17824 22060 17876
rect 25412 17824 25464 17876
rect 13544 17756 13596 17808
rect 11152 17688 11204 17740
rect 11336 17688 11388 17740
rect 13360 17688 13412 17740
rect 17592 17756 17644 17808
rect 22560 17799 22612 17808
rect 22560 17765 22569 17799
rect 22569 17765 22603 17799
rect 22603 17765 22612 17799
rect 22560 17756 22612 17765
rect 24400 17799 24452 17808
rect 24400 17765 24409 17799
rect 24409 17765 24443 17799
rect 24443 17765 24452 17799
rect 24400 17756 24452 17765
rect 16580 17688 16632 17740
rect 17776 17731 17828 17740
rect 5448 17620 5500 17672
rect 6920 17620 6972 17672
rect 8392 17663 8444 17672
rect 8392 17629 8401 17663
rect 8401 17629 8435 17663
rect 8435 17629 8444 17663
rect 8392 17620 8444 17629
rect 11060 17620 11112 17672
rect 13084 17663 13136 17672
rect 13084 17629 13093 17663
rect 13093 17629 13127 17663
rect 13127 17629 13136 17663
rect 13084 17620 13136 17629
rect 14740 17620 14792 17672
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 16028 17620 16080 17672
rect 8300 17595 8352 17604
rect 8300 17561 8309 17595
rect 8309 17561 8343 17595
rect 8343 17561 8352 17595
rect 8300 17552 8352 17561
rect 8576 17552 8628 17604
rect 3884 17527 3936 17536
rect 3884 17493 3893 17527
rect 3893 17493 3927 17527
rect 3927 17493 3936 17527
rect 3884 17484 3936 17493
rect 7472 17484 7524 17536
rect 8116 17484 8168 17536
rect 8944 17484 8996 17536
rect 9312 17552 9364 17604
rect 9772 17595 9824 17604
rect 9772 17561 9781 17595
rect 9781 17561 9815 17595
rect 9815 17561 9824 17595
rect 9772 17552 9824 17561
rect 17776 17697 17785 17731
rect 17785 17697 17819 17731
rect 17819 17697 17828 17731
rect 17776 17688 17828 17697
rect 18696 17620 18748 17672
rect 9588 17484 9640 17536
rect 14280 17527 14332 17536
rect 14280 17493 14289 17527
rect 14289 17493 14323 17527
rect 14323 17493 14332 17527
rect 14280 17484 14332 17493
rect 14832 17484 14884 17536
rect 15016 17527 15068 17536
rect 15016 17493 15025 17527
rect 15025 17493 15059 17527
rect 15059 17493 15068 17527
rect 15016 17484 15068 17493
rect 18788 17484 18840 17536
rect 23112 17731 23164 17740
rect 23112 17697 23121 17731
rect 23121 17697 23155 17731
rect 23155 17697 23164 17731
rect 23112 17688 23164 17697
rect 23204 17688 23256 17740
rect 22928 17620 22980 17672
rect 23664 17688 23716 17740
rect 23940 17688 23992 17740
rect 25964 17688 26016 17740
rect 26516 17731 26568 17740
rect 26516 17697 26525 17731
rect 26525 17697 26559 17731
rect 26559 17697 26568 17731
rect 26516 17688 26568 17697
rect 24216 17595 24268 17604
rect 19984 17484 20036 17536
rect 24216 17561 24225 17595
rect 24225 17561 24259 17595
rect 24259 17561 24268 17595
rect 24216 17552 24268 17561
rect 25412 17663 25464 17672
rect 25412 17629 25421 17663
rect 25421 17629 25455 17663
rect 25455 17629 25464 17663
rect 29184 17824 29236 17876
rect 29736 17824 29788 17876
rect 30840 17867 30892 17876
rect 30840 17833 30849 17867
rect 30849 17833 30883 17867
rect 30883 17833 30892 17867
rect 30840 17824 30892 17833
rect 27620 17688 27672 17740
rect 28080 17688 28132 17740
rect 29368 17756 29420 17808
rect 30380 17799 30432 17808
rect 30380 17765 30389 17799
rect 30389 17765 30423 17799
rect 30423 17765 30432 17799
rect 30380 17756 30432 17765
rect 28264 17731 28316 17740
rect 28264 17697 28273 17731
rect 28273 17697 28307 17731
rect 28307 17697 28316 17731
rect 29552 17731 29604 17740
rect 28264 17688 28316 17697
rect 29552 17697 29561 17731
rect 29561 17697 29595 17731
rect 29595 17697 29604 17731
rect 29552 17688 29604 17697
rect 30472 17688 30524 17740
rect 32496 17688 32548 17740
rect 33140 17688 33192 17740
rect 34520 17731 34572 17740
rect 34520 17697 34529 17731
rect 34529 17697 34563 17731
rect 34563 17697 34572 17731
rect 34520 17688 34572 17697
rect 34796 17731 34848 17740
rect 34796 17697 34805 17731
rect 34805 17697 34839 17731
rect 34839 17697 34848 17731
rect 34796 17688 34848 17697
rect 35256 17731 35308 17740
rect 35256 17697 35265 17731
rect 35265 17697 35299 17731
rect 35299 17697 35308 17731
rect 35256 17688 35308 17697
rect 35532 17731 35584 17740
rect 35532 17697 35541 17731
rect 35541 17697 35575 17731
rect 35575 17697 35584 17731
rect 35532 17688 35584 17697
rect 25412 17620 25464 17629
rect 27896 17620 27948 17672
rect 29736 17620 29788 17672
rect 32588 17620 32640 17672
rect 33508 17620 33560 17672
rect 33968 17620 34020 17672
rect 28172 17552 28224 17604
rect 25964 17527 26016 17536
rect 25964 17493 25973 17527
rect 25973 17493 26007 17527
rect 26007 17493 26016 17527
rect 25964 17484 26016 17493
rect 27068 17527 27120 17536
rect 27068 17493 27077 17527
rect 27077 17493 27111 17527
rect 27111 17493 27120 17527
rect 27068 17484 27120 17493
rect 27712 17527 27764 17536
rect 27712 17493 27721 17527
rect 27721 17493 27755 17527
rect 27755 17493 27764 17527
rect 27712 17484 27764 17493
rect 29368 17527 29420 17536
rect 29368 17493 29377 17527
rect 29377 17493 29411 17527
rect 29411 17493 29420 17527
rect 29368 17484 29420 17493
rect 29920 17484 29972 17536
rect 31208 17527 31260 17536
rect 31208 17493 31217 17527
rect 31217 17493 31251 17527
rect 31251 17493 31260 17527
rect 31208 17484 31260 17493
rect 31668 17484 31720 17536
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 3240 17280 3292 17332
rect 3516 17323 3568 17332
rect 3516 17289 3525 17323
rect 3525 17289 3559 17323
rect 3559 17289 3568 17323
rect 3516 17280 3568 17289
rect 5540 17280 5592 17332
rect 5724 17280 5776 17332
rect 8392 17280 8444 17332
rect 8668 17280 8720 17332
rect 5448 17212 5500 17264
rect 6000 17212 6052 17264
rect 6736 17212 6788 17264
rect 2412 17187 2464 17196
rect 2412 17153 2421 17187
rect 2421 17153 2455 17187
rect 2455 17153 2464 17187
rect 2412 17144 2464 17153
rect 6276 17187 6328 17196
rect 6276 17153 6285 17187
rect 6285 17153 6319 17187
rect 6319 17153 6328 17187
rect 6276 17144 6328 17153
rect 7104 17144 7156 17196
rect 9496 17280 9548 17332
rect 12440 17280 12492 17332
rect 14188 17323 14240 17332
rect 14188 17289 14197 17323
rect 14197 17289 14231 17323
rect 14231 17289 14240 17323
rect 14188 17280 14240 17289
rect 14280 17280 14332 17332
rect 16580 17280 16632 17332
rect 17592 17323 17644 17332
rect 17592 17289 17601 17323
rect 17601 17289 17635 17323
rect 17635 17289 17644 17323
rect 17592 17280 17644 17289
rect 17776 17280 17828 17332
rect 18788 17280 18840 17332
rect 19340 17280 19392 17332
rect 22928 17323 22980 17332
rect 22928 17289 22937 17323
rect 22937 17289 22971 17323
rect 22971 17289 22980 17323
rect 22928 17280 22980 17289
rect 25872 17280 25924 17332
rect 27436 17280 27488 17332
rect 28264 17280 28316 17332
rect 29552 17280 29604 17332
rect 30472 17280 30524 17332
rect 32588 17323 32640 17332
rect 32588 17289 32597 17323
rect 32597 17289 32631 17323
rect 32631 17289 32640 17323
rect 32588 17280 32640 17289
rect 34336 17280 34388 17332
rect 34520 17280 34572 17332
rect 11704 17212 11756 17264
rect 12256 17212 12308 17264
rect 14740 17212 14792 17264
rect 1860 17076 1912 17128
rect 2504 17076 2556 17128
rect 5448 17119 5500 17128
rect 5448 17085 5457 17119
rect 5457 17085 5491 17119
rect 5491 17085 5500 17119
rect 5448 17076 5500 17085
rect 7472 17076 7524 17128
rect 9404 17144 9456 17196
rect 11244 17144 11296 17196
rect 13360 17144 13412 17196
rect 14372 17144 14424 17196
rect 14648 17144 14700 17196
rect 8944 17076 8996 17128
rect 10232 17119 10284 17128
rect 10232 17085 10241 17119
rect 10241 17085 10275 17119
rect 10275 17085 10284 17119
rect 10232 17076 10284 17085
rect 10508 17119 10560 17128
rect 10508 17085 10517 17119
rect 10517 17085 10551 17119
rect 10551 17085 10560 17119
rect 10508 17076 10560 17085
rect 12440 17119 12492 17128
rect 12440 17085 12449 17119
rect 12449 17085 12483 17119
rect 12483 17085 12492 17119
rect 12440 17076 12492 17085
rect 7288 17051 7340 17060
rect 7288 17017 7297 17051
rect 7297 17017 7331 17051
rect 7331 17017 7340 17051
rect 7288 17008 7340 17017
rect 7656 17008 7708 17060
rect 8208 17008 8260 17060
rect 11980 17008 12032 17060
rect 14556 17076 14608 17128
rect 15016 17119 15068 17128
rect 15016 17085 15025 17119
rect 15025 17085 15059 17119
rect 15059 17085 15068 17119
rect 15016 17076 15068 17085
rect 15292 17076 15344 17128
rect 13360 17051 13412 17060
rect 13360 17017 13369 17051
rect 13369 17017 13403 17051
rect 13403 17017 13412 17051
rect 18052 17212 18104 17264
rect 18420 17212 18472 17264
rect 13360 17008 13412 17017
rect 2044 16940 2096 16992
rect 3516 16940 3568 16992
rect 6644 16983 6696 16992
rect 6644 16949 6653 16983
rect 6653 16949 6687 16983
rect 6687 16949 6696 16983
rect 6644 16940 6696 16949
rect 9772 16983 9824 16992
rect 9772 16949 9781 16983
rect 9781 16949 9815 16983
rect 9815 16949 9824 16983
rect 9772 16940 9824 16949
rect 11336 16983 11388 16992
rect 11336 16949 11345 16983
rect 11345 16949 11379 16983
rect 11379 16949 11388 16983
rect 11336 16940 11388 16949
rect 11612 16983 11664 16992
rect 11612 16949 11621 16983
rect 11621 16949 11655 16983
rect 11655 16949 11664 16983
rect 11612 16940 11664 16949
rect 13636 16983 13688 16992
rect 13636 16949 13645 16983
rect 13645 16949 13679 16983
rect 13679 16949 13688 16983
rect 13636 16940 13688 16949
rect 14924 16940 14976 16992
rect 16672 17144 16724 17196
rect 19432 17212 19484 17264
rect 19892 17255 19944 17264
rect 19892 17221 19901 17255
rect 19901 17221 19935 17255
rect 19935 17221 19944 17255
rect 19892 17212 19944 17221
rect 16856 17076 16908 17128
rect 17224 17076 17276 17128
rect 17316 17008 17368 17060
rect 17500 17008 17552 17060
rect 18696 17076 18748 17128
rect 19340 17076 19392 17128
rect 21364 17076 21416 17128
rect 22008 17212 22060 17264
rect 22192 17212 22244 17264
rect 26056 17212 26108 17264
rect 20720 17008 20772 17060
rect 23480 17076 23532 17128
rect 24032 17076 24084 17128
rect 22928 17008 22980 17060
rect 17224 16983 17276 16992
rect 17224 16949 17233 16983
rect 17233 16949 17267 16983
rect 17267 16949 17276 16983
rect 17224 16940 17276 16949
rect 18328 16940 18380 16992
rect 21364 16983 21416 16992
rect 21364 16949 21373 16983
rect 21373 16949 21407 16983
rect 21407 16949 21416 16983
rect 23204 16983 23256 16992
rect 21364 16940 21416 16949
rect 23204 16949 23213 16983
rect 23213 16949 23247 16983
rect 23247 16949 23256 16983
rect 23204 16940 23256 16949
rect 24124 16983 24176 16992
rect 24124 16949 24133 16983
rect 24133 16949 24167 16983
rect 24167 16949 24176 16983
rect 24124 16940 24176 16949
rect 24308 16940 24360 16992
rect 24952 16940 25004 16992
rect 26792 17144 26844 17196
rect 29092 17144 29144 17196
rect 30012 17187 30064 17196
rect 30012 17153 30021 17187
rect 30021 17153 30055 17187
rect 30055 17153 30064 17187
rect 30012 17144 30064 17153
rect 31300 17212 31352 17264
rect 31208 17144 31260 17196
rect 25964 17076 26016 17128
rect 27896 17119 27948 17128
rect 27896 17085 27905 17119
rect 27905 17085 27939 17119
rect 27939 17085 27948 17119
rect 27896 17076 27948 17085
rect 29368 17076 29420 17128
rect 31668 17119 31720 17128
rect 31668 17085 31677 17119
rect 31677 17085 31711 17119
rect 31711 17085 31720 17119
rect 31668 17076 31720 17085
rect 33324 17144 33376 17196
rect 27068 17008 27120 17060
rect 27620 17051 27672 17060
rect 27620 17017 27629 17051
rect 27629 17017 27663 17051
rect 27663 17017 27672 17051
rect 27620 17008 27672 17017
rect 27712 17008 27764 17060
rect 28540 17008 28592 17060
rect 29276 17051 29328 17060
rect 29276 17017 29285 17051
rect 29285 17017 29319 17051
rect 29319 17017 29328 17051
rect 29276 17008 29328 17017
rect 29736 17008 29788 17060
rect 31300 17008 31352 17060
rect 31760 17008 31812 17060
rect 32496 17076 32548 17128
rect 32864 17076 32916 17128
rect 33784 17119 33836 17128
rect 33784 17085 33793 17119
rect 33793 17085 33827 17119
rect 33827 17085 33836 17119
rect 33784 17076 33836 17085
rect 33600 17008 33652 17060
rect 26516 16940 26568 16992
rect 28080 16940 28132 16992
rect 29460 16983 29512 16992
rect 29460 16949 29469 16983
rect 29469 16949 29503 16983
rect 29503 16949 29512 16983
rect 29460 16940 29512 16949
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 1400 16736 1452 16788
rect 1860 16736 1912 16788
rect 2044 16779 2096 16788
rect 2044 16745 2053 16779
rect 2053 16745 2087 16779
rect 2087 16745 2096 16779
rect 2044 16736 2096 16745
rect 2412 16779 2464 16788
rect 2412 16745 2421 16779
rect 2421 16745 2455 16779
rect 2455 16745 2464 16779
rect 2412 16736 2464 16745
rect 3148 16779 3200 16788
rect 3148 16745 3157 16779
rect 3157 16745 3191 16779
rect 3191 16745 3200 16779
rect 3148 16736 3200 16745
rect 3976 16736 4028 16788
rect 5356 16736 5408 16788
rect 7104 16779 7156 16788
rect 7104 16745 7113 16779
rect 7113 16745 7147 16779
rect 7147 16745 7156 16779
rect 7104 16736 7156 16745
rect 9312 16736 9364 16788
rect 4068 16668 4120 16720
rect 7288 16668 7340 16720
rect 7472 16711 7524 16720
rect 7472 16677 7481 16711
rect 7481 16677 7515 16711
rect 7515 16677 7524 16711
rect 7472 16668 7524 16677
rect 4896 16643 4948 16652
rect 4896 16609 4905 16643
rect 4905 16609 4939 16643
rect 4939 16609 4948 16643
rect 4896 16600 4948 16609
rect 5172 16643 5224 16652
rect 5172 16609 5181 16643
rect 5181 16609 5215 16643
rect 5215 16609 5224 16643
rect 5172 16600 5224 16609
rect 5356 16643 5408 16652
rect 5356 16609 5365 16643
rect 5365 16609 5399 16643
rect 5399 16609 5408 16643
rect 5356 16600 5408 16609
rect 5632 16643 5684 16652
rect 5632 16609 5641 16643
rect 5641 16609 5675 16643
rect 5675 16609 5684 16643
rect 5632 16600 5684 16609
rect 6644 16643 6696 16652
rect 6644 16609 6653 16643
rect 6653 16609 6687 16643
rect 6687 16609 6696 16643
rect 7840 16668 7892 16720
rect 8024 16711 8076 16720
rect 8024 16677 8033 16711
rect 8033 16677 8067 16711
rect 8067 16677 8076 16711
rect 8024 16668 8076 16677
rect 7932 16643 7984 16652
rect 6644 16600 6696 16609
rect 7932 16609 7941 16643
rect 7941 16609 7975 16643
rect 7975 16609 7984 16643
rect 7932 16600 7984 16609
rect 4988 16464 5040 16516
rect 3148 16396 3200 16448
rect 8576 16668 8628 16720
rect 9680 16736 9732 16788
rect 11060 16736 11112 16788
rect 10232 16711 10284 16720
rect 10232 16677 10241 16711
rect 10241 16677 10275 16711
rect 10275 16677 10284 16711
rect 10232 16668 10284 16677
rect 11704 16668 11756 16720
rect 8392 16600 8444 16652
rect 9864 16600 9916 16652
rect 8944 16396 8996 16448
rect 10508 16396 10560 16448
rect 11060 16643 11112 16652
rect 11060 16609 11069 16643
rect 11069 16609 11103 16643
rect 11103 16609 11112 16643
rect 11060 16600 11112 16609
rect 11244 16600 11296 16652
rect 10876 16532 10928 16584
rect 11520 16575 11572 16584
rect 11520 16541 11529 16575
rect 11529 16541 11563 16575
rect 11563 16541 11572 16575
rect 11520 16532 11572 16541
rect 14096 16779 14148 16788
rect 14096 16745 14105 16779
rect 14105 16745 14139 16779
rect 14139 16745 14148 16779
rect 14096 16736 14148 16745
rect 14740 16779 14792 16788
rect 14740 16745 14749 16779
rect 14749 16745 14783 16779
rect 14783 16745 14792 16779
rect 14740 16736 14792 16745
rect 16028 16779 16080 16788
rect 16028 16745 16037 16779
rect 16037 16745 16071 16779
rect 16071 16745 16080 16779
rect 16028 16736 16080 16745
rect 16580 16736 16632 16788
rect 18144 16736 18196 16788
rect 20720 16779 20772 16788
rect 20720 16745 20729 16779
rect 20729 16745 20763 16779
rect 20763 16745 20772 16779
rect 20720 16736 20772 16745
rect 24860 16736 24912 16788
rect 26608 16736 26660 16788
rect 27896 16736 27948 16788
rect 28540 16736 28592 16788
rect 13176 16668 13228 16720
rect 14280 16668 14332 16720
rect 15016 16668 15068 16720
rect 17224 16668 17276 16720
rect 17316 16668 17368 16720
rect 12348 16600 12400 16652
rect 12532 16643 12584 16652
rect 12532 16609 12541 16643
rect 12541 16609 12575 16643
rect 12575 16609 12584 16643
rect 12532 16600 12584 16609
rect 12624 16643 12676 16652
rect 12624 16609 12633 16643
rect 12633 16609 12667 16643
rect 12667 16609 12676 16643
rect 12624 16600 12676 16609
rect 13636 16532 13688 16584
rect 14188 16600 14240 16652
rect 14372 16643 14424 16652
rect 14372 16609 14381 16643
rect 14381 16609 14415 16643
rect 14415 16609 14424 16643
rect 14372 16600 14424 16609
rect 15568 16643 15620 16652
rect 15568 16609 15577 16643
rect 15577 16609 15611 16643
rect 15611 16609 15620 16643
rect 15568 16600 15620 16609
rect 16672 16643 16724 16652
rect 16672 16609 16681 16643
rect 16681 16609 16715 16643
rect 16715 16609 16724 16643
rect 16672 16600 16724 16609
rect 16948 16600 17000 16652
rect 17500 16600 17552 16652
rect 18696 16600 18748 16652
rect 19156 16668 19208 16720
rect 19800 16711 19852 16720
rect 19800 16677 19809 16711
rect 19809 16677 19843 16711
rect 19843 16677 19852 16711
rect 19800 16668 19852 16677
rect 22928 16711 22980 16720
rect 22928 16677 22937 16711
rect 22937 16677 22971 16711
rect 22971 16677 22980 16711
rect 22928 16668 22980 16677
rect 25964 16668 26016 16720
rect 27252 16711 27304 16720
rect 27252 16677 27261 16711
rect 27261 16677 27295 16711
rect 27295 16677 27304 16711
rect 27252 16668 27304 16677
rect 29736 16736 29788 16788
rect 29828 16779 29880 16788
rect 29828 16745 29837 16779
rect 29837 16745 29871 16779
rect 29871 16745 29880 16779
rect 31300 16779 31352 16788
rect 29828 16736 29880 16745
rect 31300 16745 31309 16779
rect 31309 16745 31343 16779
rect 31343 16745 31352 16779
rect 31300 16736 31352 16745
rect 31392 16736 31444 16788
rect 32864 16779 32916 16788
rect 32864 16745 32873 16779
rect 32873 16745 32907 16779
rect 32907 16745 32916 16779
rect 32864 16736 32916 16745
rect 33600 16736 33652 16788
rect 34796 16779 34848 16788
rect 34796 16745 34805 16779
rect 34805 16745 34839 16779
rect 34839 16745 34848 16779
rect 34796 16736 34848 16745
rect 35256 16736 35308 16788
rect 29460 16668 29512 16720
rect 30288 16711 30340 16720
rect 30288 16677 30297 16711
rect 30297 16677 30331 16711
rect 30331 16677 30340 16711
rect 30288 16668 30340 16677
rect 31024 16668 31076 16720
rect 31668 16668 31720 16720
rect 19248 16600 19300 16652
rect 20996 16600 21048 16652
rect 21916 16643 21968 16652
rect 21916 16609 21925 16643
rect 21925 16609 21959 16643
rect 21959 16609 21968 16643
rect 21916 16600 21968 16609
rect 22100 16600 22152 16652
rect 24124 16600 24176 16652
rect 24676 16600 24728 16652
rect 24952 16600 25004 16652
rect 26056 16600 26108 16652
rect 17316 16532 17368 16584
rect 19340 16532 19392 16584
rect 21180 16532 21232 16584
rect 21364 16575 21416 16584
rect 21364 16541 21373 16575
rect 21373 16541 21407 16575
rect 21407 16541 21416 16575
rect 21364 16532 21416 16541
rect 21640 16532 21692 16584
rect 23112 16532 23164 16584
rect 23940 16575 23992 16584
rect 23940 16541 23949 16575
rect 23949 16541 23983 16575
rect 23983 16541 23992 16575
rect 23940 16532 23992 16541
rect 24400 16532 24452 16584
rect 26332 16532 26384 16584
rect 26700 16532 26752 16584
rect 29368 16600 29420 16652
rect 30196 16600 30248 16652
rect 30748 16643 30800 16652
rect 30748 16609 30757 16643
rect 30757 16609 30791 16643
rect 30791 16609 30800 16643
rect 30748 16600 30800 16609
rect 32496 16600 32548 16652
rect 33324 16668 33376 16720
rect 34704 16668 34756 16720
rect 33692 16600 33744 16652
rect 29276 16532 29328 16584
rect 16212 16396 16264 16448
rect 17776 16396 17828 16448
rect 18328 16396 18380 16448
rect 21548 16396 21600 16448
rect 24860 16396 24912 16448
rect 25044 16439 25096 16448
rect 25044 16405 25053 16439
rect 25053 16405 25087 16439
rect 25087 16405 25096 16439
rect 25872 16439 25924 16448
rect 25044 16396 25096 16405
rect 25872 16405 25881 16439
rect 25881 16405 25915 16439
rect 25915 16405 25924 16439
rect 25872 16396 25924 16405
rect 26608 16396 26660 16448
rect 28080 16439 28132 16448
rect 28080 16405 28089 16439
rect 28089 16405 28123 16439
rect 28123 16405 28132 16439
rect 28080 16396 28132 16405
rect 28540 16396 28592 16448
rect 28816 16396 28868 16448
rect 32864 16532 32916 16584
rect 33048 16575 33100 16584
rect 33048 16541 33057 16575
rect 33057 16541 33091 16575
rect 33091 16541 33100 16575
rect 33048 16532 33100 16541
rect 32220 16464 32272 16516
rect 33876 16532 33928 16584
rect 34060 16575 34112 16584
rect 34060 16541 34069 16575
rect 34069 16541 34103 16575
rect 34103 16541 34112 16575
rect 34060 16532 34112 16541
rect 30932 16439 30984 16448
rect 30932 16405 30941 16439
rect 30941 16405 30975 16439
rect 30975 16405 30984 16439
rect 30932 16396 30984 16405
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 4068 16192 4120 16244
rect 4804 16235 4856 16244
rect 4804 16201 4813 16235
rect 4813 16201 4847 16235
rect 4847 16201 4856 16235
rect 4804 16192 4856 16201
rect 5356 16192 5408 16244
rect 6644 16235 6696 16244
rect 6644 16201 6653 16235
rect 6653 16201 6687 16235
rect 6687 16201 6696 16235
rect 6644 16192 6696 16201
rect 7840 16192 7892 16244
rect 10876 16192 10928 16244
rect 13452 16192 13504 16244
rect 16672 16235 16724 16244
rect 16672 16201 16681 16235
rect 16681 16201 16715 16235
rect 16715 16201 16724 16235
rect 16672 16192 16724 16201
rect 4620 16167 4672 16176
rect 4620 16133 4629 16167
rect 4629 16133 4663 16167
rect 4663 16133 4672 16167
rect 4620 16124 4672 16133
rect 5080 16124 5132 16176
rect 5724 16124 5776 16176
rect 8024 16124 8076 16176
rect 9312 16124 9364 16176
rect 9956 16124 10008 16176
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 4712 16056 4764 16108
rect 5264 16099 5316 16108
rect 5264 16065 5273 16099
rect 5273 16065 5307 16099
rect 5307 16065 5316 16099
rect 5264 16056 5316 16065
rect 10232 16099 10284 16108
rect 10232 16065 10241 16099
rect 10241 16065 10275 16099
rect 10275 16065 10284 16099
rect 10232 16056 10284 16065
rect 5356 16031 5408 16040
rect 5356 15997 5365 16031
rect 5365 15997 5399 16031
rect 5399 15997 5408 16031
rect 5356 15988 5408 15997
rect 5724 16031 5776 16040
rect 5724 15997 5733 16031
rect 5733 15997 5767 16031
rect 5767 15997 5776 16031
rect 5724 15988 5776 15997
rect 6276 15988 6328 16040
rect 6644 15988 6696 16040
rect 6920 15988 6972 16040
rect 8852 16031 8904 16040
rect 8852 15997 8861 16031
rect 8861 15997 8895 16031
rect 8895 15997 8904 16031
rect 8852 15988 8904 15997
rect 9220 16031 9272 16040
rect 9220 15997 9229 16031
rect 9229 15997 9263 16031
rect 9263 15997 9272 16031
rect 9220 15988 9272 15997
rect 9956 15988 10008 16040
rect 10692 15988 10744 16040
rect 3884 15920 3936 15972
rect 5632 15920 5684 15972
rect 7196 15963 7248 15972
rect 6828 15852 6880 15904
rect 7196 15929 7205 15963
rect 7205 15929 7239 15963
rect 7239 15929 7248 15963
rect 7196 15920 7248 15929
rect 11152 15920 11204 15972
rect 13360 15988 13412 16040
rect 13636 16124 13688 16176
rect 14556 16124 14608 16176
rect 15108 16124 15160 16176
rect 15200 16124 15252 16176
rect 13912 16031 13964 16040
rect 13912 15997 13921 16031
rect 13921 15997 13955 16031
rect 13955 15997 13964 16031
rect 15568 16056 15620 16108
rect 13912 15988 13964 15997
rect 12440 15963 12492 15972
rect 7288 15852 7340 15904
rect 9864 15852 9916 15904
rect 11244 15852 11296 15904
rect 11612 15895 11664 15904
rect 11612 15861 11621 15895
rect 11621 15861 11655 15895
rect 11655 15861 11664 15895
rect 12440 15929 12449 15963
rect 12449 15929 12483 15963
rect 12483 15929 12492 15963
rect 12808 15963 12860 15972
rect 12440 15920 12492 15929
rect 12808 15929 12817 15963
rect 12817 15929 12851 15963
rect 12851 15929 12860 15963
rect 12808 15920 12860 15929
rect 13176 15963 13228 15972
rect 13176 15929 13185 15963
rect 13185 15929 13219 15963
rect 13219 15929 13228 15963
rect 13176 15920 13228 15929
rect 16120 15988 16172 16040
rect 17316 16192 17368 16244
rect 19156 16192 19208 16244
rect 21180 16192 21232 16244
rect 21640 16192 21692 16244
rect 23940 16192 23992 16244
rect 25228 16235 25280 16244
rect 25228 16201 25237 16235
rect 25237 16201 25271 16235
rect 25271 16201 25280 16235
rect 25228 16192 25280 16201
rect 26240 16192 26292 16244
rect 27804 16192 27856 16244
rect 17224 16124 17276 16176
rect 22376 16167 22428 16176
rect 22376 16133 22385 16167
rect 22385 16133 22419 16167
rect 22419 16133 22428 16167
rect 22376 16124 22428 16133
rect 25044 16167 25096 16176
rect 25044 16133 25053 16167
rect 25053 16133 25087 16167
rect 25087 16133 25096 16167
rect 25044 16124 25096 16133
rect 26056 16124 26108 16176
rect 26516 16167 26568 16176
rect 26516 16133 26540 16167
rect 26540 16133 26568 16167
rect 26516 16124 26568 16133
rect 17776 15988 17828 16040
rect 15568 15920 15620 15972
rect 18788 16056 18840 16108
rect 21364 16056 21416 16108
rect 22100 16056 22152 16108
rect 18512 15988 18564 16040
rect 18972 15988 19024 16040
rect 19248 15988 19300 16040
rect 11612 15852 11664 15861
rect 12348 15852 12400 15904
rect 12532 15852 12584 15904
rect 14188 15852 14240 15904
rect 15200 15895 15252 15904
rect 15200 15861 15209 15895
rect 15209 15861 15243 15895
rect 15243 15861 15252 15895
rect 15200 15852 15252 15861
rect 17684 15852 17736 15904
rect 18788 15963 18840 15972
rect 18788 15929 18797 15963
rect 18797 15929 18831 15963
rect 18831 15929 18840 15963
rect 18788 15920 18840 15929
rect 18144 15852 18196 15904
rect 18328 15852 18380 15904
rect 18696 15852 18748 15904
rect 19984 15988 20036 16040
rect 21824 15988 21876 16040
rect 22928 15988 22980 16040
rect 23756 15988 23808 16040
rect 20260 15852 20312 15904
rect 23480 15895 23532 15904
rect 23480 15861 23489 15895
rect 23489 15861 23523 15895
rect 23523 15861 23532 15895
rect 23480 15852 23532 15861
rect 24860 15988 24912 16040
rect 25320 15988 25372 16040
rect 26148 16056 26200 16108
rect 26700 16099 26752 16108
rect 26700 16065 26709 16099
rect 26709 16065 26743 16099
rect 26743 16065 26752 16099
rect 26700 16056 26752 16065
rect 28816 16192 28868 16244
rect 29276 16192 29328 16244
rect 30748 16192 30800 16244
rect 33876 16192 33928 16244
rect 31024 16124 31076 16176
rect 30196 16099 30248 16108
rect 30196 16065 30205 16099
rect 30205 16065 30239 16099
rect 30239 16065 30248 16099
rect 30196 16056 30248 16065
rect 30932 16056 30984 16108
rect 24676 15920 24728 15972
rect 27896 15920 27948 15972
rect 29092 15920 29144 15972
rect 29828 15988 29880 16040
rect 31852 16031 31904 16040
rect 31852 15997 31861 16031
rect 31861 15997 31895 16031
rect 31895 15997 31904 16031
rect 31852 15988 31904 15997
rect 33324 16031 33376 16040
rect 33324 15997 33333 16031
rect 33333 15997 33367 16031
rect 33367 15997 33376 16031
rect 33324 15988 33376 15997
rect 33508 15988 33560 16040
rect 34888 16031 34940 16040
rect 34888 15997 34897 16031
rect 34897 15997 34931 16031
rect 34931 15997 34940 16031
rect 34888 15988 34940 15997
rect 32220 15920 32272 15972
rect 23940 15852 23992 15904
rect 24308 15895 24360 15904
rect 24308 15861 24317 15895
rect 24317 15861 24351 15895
rect 24351 15861 24360 15895
rect 24308 15852 24360 15861
rect 26240 15895 26292 15904
rect 26240 15861 26249 15895
rect 26249 15861 26283 15895
rect 26283 15861 26292 15895
rect 26240 15852 26292 15861
rect 28080 15895 28132 15904
rect 28080 15861 28089 15895
rect 28089 15861 28123 15895
rect 28123 15861 28132 15895
rect 28080 15852 28132 15861
rect 28540 15852 28592 15904
rect 32864 15852 32916 15904
rect 33508 15852 33560 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 1676 15691 1728 15700
rect 1676 15657 1685 15691
rect 1685 15657 1719 15691
rect 1719 15657 1728 15691
rect 1676 15648 1728 15657
rect 4804 15648 4856 15700
rect 5356 15648 5408 15700
rect 6920 15648 6972 15700
rect 7932 15648 7984 15700
rect 8300 15648 8352 15700
rect 10876 15648 10928 15700
rect 11336 15648 11388 15700
rect 12992 15691 13044 15700
rect 12992 15657 13001 15691
rect 13001 15657 13035 15691
rect 13035 15657 13044 15691
rect 12992 15648 13044 15657
rect 16120 15691 16172 15700
rect 16120 15657 16129 15691
rect 16129 15657 16163 15691
rect 16163 15657 16172 15691
rect 16120 15648 16172 15657
rect 17132 15648 17184 15700
rect 17776 15648 17828 15700
rect 19156 15691 19208 15700
rect 19156 15657 19165 15691
rect 19165 15657 19199 15691
rect 19199 15657 19208 15691
rect 19156 15648 19208 15657
rect 20628 15648 20680 15700
rect 21824 15648 21876 15700
rect 5540 15580 5592 15632
rect 5908 15580 5960 15632
rect 4896 15512 4948 15564
rect 5816 15512 5868 15564
rect 6184 15512 6236 15564
rect 11612 15623 11664 15632
rect 7104 15555 7156 15564
rect 7104 15521 7113 15555
rect 7113 15521 7147 15555
rect 7147 15521 7156 15555
rect 7104 15512 7156 15521
rect 7840 15512 7892 15564
rect 9680 15555 9732 15564
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 10508 15512 10560 15564
rect 10692 15512 10744 15564
rect 11152 15555 11204 15564
rect 11152 15521 11161 15555
rect 11161 15521 11195 15555
rect 11195 15521 11204 15555
rect 11612 15589 11621 15623
rect 11621 15589 11655 15623
rect 11655 15589 11664 15623
rect 11612 15580 11664 15589
rect 12440 15580 12492 15632
rect 13084 15580 13136 15632
rect 16212 15580 16264 15632
rect 17224 15580 17276 15632
rect 18144 15580 18196 15632
rect 18972 15580 19024 15632
rect 19432 15580 19484 15632
rect 20996 15580 21048 15632
rect 21548 15580 21600 15632
rect 21732 15580 21784 15632
rect 22284 15648 22336 15700
rect 22744 15648 22796 15700
rect 23296 15648 23348 15700
rect 24308 15648 24360 15700
rect 25044 15648 25096 15700
rect 26976 15648 27028 15700
rect 27896 15691 27948 15700
rect 27896 15657 27905 15691
rect 27905 15657 27939 15691
rect 27939 15657 27948 15691
rect 27896 15648 27948 15657
rect 28448 15648 28500 15700
rect 23112 15580 23164 15632
rect 23480 15580 23532 15632
rect 24676 15580 24728 15632
rect 25964 15623 26016 15632
rect 25964 15589 25973 15623
rect 25973 15589 26007 15623
rect 26007 15589 26016 15623
rect 25964 15580 26016 15589
rect 28632 15623 28684 15632
rect 28632 15589 28641 15623
rect 28641 15589 28675 15623
rect 28675 15589 28684 15623
rect 28632 15580 28684 15589
rect 29092 15580 29144 15632
rect 29368 15623 29420 15632
rect 29368 15589 29377 15623
rect 29377 15589 29411 15623
rect 29411 15589 29420 15623
rect 29368 15580 29420 15589
rect 30472 15648 30524 15700
rect 31760 15648 31812 15700
rect 33692 15648 33744 15700
rect 30288 15580 30340 15632
rect 11152 15512 11204 15521
rect 11796 15512 11848 15564
rect 12256 15512 12308 15564
rect 13176 15555 13228 15564
rect 13176 15521 13185 15555
rect 13185 15521 13219 15555
rect 13219 15521 13228 15555
rect 13176 15512 13228 15521
rect 13636 15555 13688 15564
rect 13636 15521 13645 15555
rect 13645 15521 13679 15555
rect 13679 15521 13688 15555
rect 13636 15512 13688 15521
rect 3240 15444 3292 15496
rect 5080 15444 5132 15496
rect 5724 15444 5776 15496
rect 8300 15487 8352 15496
rect 8300 15453 8309 15487
rect 8309 15453 8343 15487
rect 8343 15453 8352 15487
rect 8300 15444 8352 15453
rect 10876 15487 10928 15496
rect 10876 15453 10885 15487
rect 10885 15453 10919 15487
rect 10919 15453 10928 15487
rect 10876 15444 10928 15453
rect 14740 15512 14792 15564
rect 15292 15555 15344 15564
rect 15292 15521 15301 15555
rect 15301 15521 15335 15555
rect 15335 15521 15344 15555
rect 15292 15512 15344 15521
rect 16764 15555 16816 15564
rect 16764 15521 16773 15555
rect 16773 15521 16807 15555
rect 16807 15521 16816 15555
rect 16764 15512 16816 15521
rect 18052 15512 18104 15564
rect 21824 15555 21876 15564
rect 21824 15521 21833 15555
rect 21833 15521 21867 15555
rect 21867 15521 21876 15555
rect 21824 15512 21876 15521
rect 4712 15376 4764 15428
rect 5448 15376 5500 15428
rect 6828 15376 6880 15428
rect 16672 15444 16724 15496
rect 18604 15444 18656 15496
rect 19340 15444 19392 15496
rect 15200 15376 15252 15428
rect 17960 15376 18012 15428
rect 22560 15376 22612 15428
rect 22744 15376 22796 15428
rect 23940 15512 23992 15564
rect 25504 15512 25556 15564
rect 26332 15512 26384 15564
rect 28356 15512 28408 15564
rect 29460 15512 29512 15564
rect 30012 15555 30064 15564
rect 30012 15521 30021 15555
rect 30021 15521 30055 15555
rect 30055 15521 30064 15555
rect 30012 15512 30064 15521
rect 23296 15444 23348 15496
rect 24400 15444 24452 15496
rect 25320 15487 25372 15496
rect 25320 15453 25329 15487
rect 25329 15453 25363 15487
rect 25363 15453 25372 15487
rect 25320 15444 25372 15453
rect 26056 15444 26108 15496
rect 26792 15444 26844 15496
rect 27344 15444 27396 15496
rect 27620 15444 27672 15496
rect 27896 15376 27948 15428
rect 29276 15444 29328 15496
rect 31944 15512 31996 15564
rect 32220 15512 32272 15564
rect 32404 15512 32456 15564
rect 32496 15512 32548 15564
rect 33140 15512 33192 15564
rect 34428 15555 34480 15564
rect 34428 15521 34437 15555
rect 34437 15521 34471 15555
rect 34471 15521 34480 15555
rect 34428 15512 34480 15521
rect 34796 15555 34848 15564
rect 34796 15521 34805 15555
rect 34805 15521 34839 15555
rect 34839 15521 34848 15555
rect 34796 15512 34848 15521
rect 30564 15487 30616 15496
rect 28448 15376 28500 15428
rect 29920 15376 29972 15428
rect 30564 15453 30573 15487
rect 30573 15453 30607 15487
rect 30607 15453 30616 15487
rect 30564 15444 30616 15453
rect 34336 15444 34388 15496
rect 34796 15419 34848 15428
rect 34796 15385 34805 15419
rect 34805 15385 34839 15419
rect 34839 15385 34848 15419
rect 34796 15376 34848 15385
rect 4988 15308 5040 15360
rect 6276 15308 6328 15360
rect 8024 15308 8076 15360
rect 8944 15351 8996 15360
rect 8944 15317 8953 15351
rect 8953 15317 8987 15351
rect 8987 15317 8996 15351
rect 8944 15308 8996 15317
rect 9220 15308 9272 15360
rect 9956 15308 10008 15360
rect 10508 15308 10560 15360
rect 12900 15308 12952 15360
rect 14740 15351 14792 15360
rect 14740 15317 14749 15351
rect 14749 15317 14783 15351
rect 14783 15317 14792 15351
rect 14740 15308 14792 15317
rect 15108 15351 15160 15360
rect 15108 15317 15117 15351
rect 15117 15317 15151 15351
rect 15151 15317 15160 15351
rect 15108 15308 15160 15317
rect 18052 15351 18104 15360
rect 18052 15317 18061 15351
rect 18061 15317 18095 15351
rect 18095 15317 18104 15351
rect 18052 15308 18104 15317
rect 19156 15308 19208 15360
rect 23848 15308 23900 15360
rect 24216 15308 24268 15360
rect 26792 15351 26844 15360
rect 26792 15317 26801 15351
rect 26801 15317 26835 15351
rect 26835 15317 26844 15351
rect 26792 15308 26844 15317
rect 27436 15308 27488 15360
rect 30196 15308 30248 15360
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 2872 15104 2924 15156
rect 5816 15104 5868 15156
rect 8484 15147 8536 15156
rect 8484 15113 8493 15147
rect 8493 15113 8527 15147
rect 8527 15113 8536 15147
rect 8484 15104 8536 15113
rect 10968 15147 11020 15156
rect 10968 15113 10992 15147
rect 10992 15113 11020 15147
rect 10968 15104 11020 15113
rect 11060 15147 11112 15156
rect 11060 15113 11069 15147
rect 11069 15113 11103 15147
rect 11103 15113 11112 15147
rect 11060 15104 11112 15113
rect 11336 15104 11388 15156
rect 7656 15079 7708 15088
rect 7656 15045 7665 15079
rect 7665 15045 7699 15079
rect 7699 15045 7708 15079
rect 7656 15036 7708 15045
rect 8392 15036 8444 15088
rect 9680 15036 9732 15088
rect 11244 15079 11296 15088
rect 1400 15011 1452 15020
rect 1400 14977 1409 15011
rect 1409 14977 1443 15011
rect 1443 14977 1452 15011
rect 1400 14968 1452 14977
rect 1584 14968 1636 15020
rect 2872 14968 2924 15020
rect 3424 14968 3476 15020
rect 4712 14968 4764 15020
rect 4344 14943 4396 14952
rect 4344 14909 4353 14943
rect 4353 14909 4387 14943
rect 4387 14909 4396 14943
rect 4344 14900 4396 14909
rect 4804 14900 4856 14952
rect 7196 14968 7248 15020
rect 7840 15011 7892 15020
rect 7840 14977 7849 15011
rect 7849 14977 7883 15011
rect 7883 14977 7892 15011
rect 7840 14968 7892 14977
rect 9404 14968 9456 15020
rect 11244 15045 11253 15079
rect 11253 15045 11287 15079
rect 11287 15045 11296 15079
rect 11244 15036 11296 15045
rect 5080 14943 5132 14952
rect 5080 14909 5089 14943
rect 5089 14909 5123 14943
rect 5123 14909 5132 14943
rect 5080 14900 5132 14909
rect 7104 14900 7156 14952
rect 7472 14900 7524 14952
rect 10784 14943 10836 14952
rect 10784 14909 10793 14943
rect 10793 14909 10827 14943
rect 10827 14909 10836 14943
rect 10784 14900 10836 14909
rect 11520 14968 11572 15020
rect 13176 15104 13228 15156
rect 13636 15104 13688 15156
rect 15292 15104 15344 15156
rect 16212 15104 16264 15156
rect 16764 15104 16816 15156
rect 17776 15104 17828 15156
rect 17960 15104 18012 15156
rect 19248 15104 19300 15156
rect 21824 15104 21876 15156
rect 23296 15104 23348 15156
rect 24308 15147 24360 15156
rect 24308 15113 24317 15147
rect 24317 15113 24351 15147
rect 24351 15113 24360 15147
rect 24308 15104 24360 15113
rect 24492 15147 24544 15156
rect 24492 15113 24501 15147
rect 24501 15113 24535 15147
rect 24535 15113 24544 15147
rect 24492 15104 24544 15113
rect 26056 15104 26108 15156
rect 26332 15104 26384 15156
rect 27068 15104 27120 15156
rect 28448 15104 28500 15156
rect 28632 15147 28684 15156
rect 28632 15113 28641 15147
rect 28641 15113 28675 15147
rect 28675 15113 28684 15147
rect 28632 15104 28684 15113
rect 29276 15104 29328 15156
rect 31852 15104 31904 15156
rect 31944 15147 31996 15156
rect 31944 15113 31953 15147
rect 31953 15113 31987 15147
rect 31987 15113 31996 15147
rect 31944 15104 31996 15113
rect 32588 15104 32640 15156
rect 33140 15104 33192 15156
rect 34336 15104 34388 15156
rect 34704 15104 34756 15156
rect 12348 15036 12400 15088
rect 16028 15036 16080 15088
rect 18328 15036 18380 15088
rect 12900 14968 12952 15020
rect 11796 14900 11848 14952
rect 14004 14900 14056 14952
rect 7380 14875 7432 14884
rect 7380 14841 7389 14875
rect 7389 14841 7423 14875
rect 7423 14841 7432 14875
rect 7380 14832 7432 14841
rect 7932 14832 7984 14884
rect 8944 14875 8996 14884
rect 8944 14841 8953 14875
rect 8953 14841 8987 14875
rect 8987 14841 8996 14875
rect 8944 14832 8996 14841
rect 9588 14832 9640 14884
rect 9864 14832 9916 14884
rect 12808 14875 12860 14884
rect 12808 14841 12817 14875
rect 12817 14841 12851 14875
rect 12851 14841 12860 14875
rect 12808 14832 12860 14841
rect 3424 14807 3476 14816
rect 3424 14773 3433 14807
rect 3433 14773 3467 14807
rect 3467 14773 3476 14807
rect 3424 14764 3476 14773
rect 3976 14807 4028 14816
rect 3976 14773 3985 14807
rect 3985 14773 4019 14807
rect 4019 14773 4028 14807
rect 3976 14764 4028 14773
rect 5908 14764 5960 14816
rect 6184 14764 6236 14816
rect 7012 14764 7064 14816
rect 7196 14807 7248 14816
rect 7196 14773 7205 14807
rect 7205 14773 7239 14807
rect 7239 14773 7248 14807
rect 7196 14764 7248 14773
rect 9128 14807 9180 14816
rect 9128 14773 9137 14807
rect 9137 14773 9171 14807
rect 9171 14773 9180 14807
rect 9128 14764 9180 14773
rect 9404 14764 9456 14816
rect 11152 14764 11204 14816
rect 12532 14764 12584 14816
rect 13820 14764 13872 14816
rect 16580 14968 16632 15020
rect 17500 14968 17552 15020
rect 19892 15036 19944 15088
rect 22468 15079 22520 15088
rect 22468 15045 22477 15079
rect 22477 15045 22511 15079
rect 22511 15045 22520 15079
rect 22468 15036 22520 15045
rect 25872 15036 25924 15088
rect 26792 15036 26844 15088
rect 27712 15079 27764 15088
rect 27712 15045 27721 15079
rect 27721 15045 27755 15079
rect 27755 15045 27764 15079
rect 27712 15036 27764 15045
rect 18788 14968 18840 15020
rect 19248 14968 19300 15020
rect 23848 14968 23900 15020
rect 24400 15011 24452 15020
rect 24400 14977 24409 15011
rect 24409 14977 24443 15011
rect 24443 14977 24452 15011
rect 24400 14968 24452 14977
rect 26332 15011 26384 15020
rect 26332 14977 26341 15011
rect 26341 14977 26375 15011
rect 26375 14977 26384 15011
rect 26332 14968 26384 14977
rect 26700 14968 26752 15020
rect 29828 14968 29880 15020
rect 30564 15011 30616 15020
rect 15384 14900 15436 14952
rect 15660 14943 15712 14952
rect 15660 14909 15669 14943
rect 15669 14909 15703 14943
rect 15703 14909 15712 14943
rect 15660 14900 15712 14909
rect 16304 14900 16356 14952
rect 18052 14900 18104 14952
rect 18328 14943 18380 14952
rect 18328 14909 18337 14943
rect 18337 14909 18371 14943
rect 18371 14909 18380 14943
rect 18328 14900 18380 14909
rect 19156 14900 19208 14952
rect 19340 14900 19392 14952
rect 20168 14943 20220 14952
rect 20168 14909 20177 14943
rect 20177 14909 20211 14943
rect 20211 14909 20220 14943
rect 20168 14900 20220 14909
rect 15568 14832 15620 14884
rect 19248 14832 19300 14884
rect 17132 14764 17184 14816
rect 18604 14764 18656 14816
rect 19156 14764 19208 14816
rect 22284 14900 22336 14952
rect 22560 14943 22612 14952
rect 22560 14909 22569 14943
rect 22569 14909 22603 14943
rect 22603 14909 22612 14943
rect 22560 14900 22612 14909
rect 23480 14900 23532 14952
rect 24124 14900 24176 14952
rect 25964 14943 26016 14952
rect 25964 14909 25973 14943
rect 25973 14909 26007 14943
rect 26007 14909 26016 14943
rect 25964 14900 26016 14909
rect 26608 14900 26660 14952
rect 27436 14900 27488 14952
rect 30196 14900 30248 14952
rect 30564 14977 30573 15011
rect 30573 14977 30607 15011
rect 30607 14977 30616 15011
rect 30564 14968 30616 14977
rect 34428 15036 34480 15088
rect 33048 15011 33100 15020
rect 33048 14977 33057 15011
rect 33057 14977 33091 15011
rect 33091 14977 33100 15011
rect 33048 14968 33100 14977
rect 32588 14900 32640 14952
rect 33508 14943 33560 14952
rect 33508 14909 33517 14943
rect 33517 14909 33551 14943
rect 33551 14909 33560 14943
rect 33508 14900 33560 14909
rect 26700 14875 26752 14884
rect 26700 14841 26709 14875
rect 26709 14841 26743 14875
rect 26743 14841 26752 14875
rect 26700 14832 26752 14841
rect 21824 14764 21876 14816
rect 24216 14764 24268 14816
rect 25504 14807 25556 14816
rect 25504 14773 25513 14807
rect 25513 14773 25547 14807
rect 25547 14773 25556 14807
rect 25504 14764 25556 14773
rect 25872 14807 25924 14816
rect 25872 14773 25881 14807
rect 25881 14773 25915 14807
rect 25915 14773 25924 14807
rect 25872 14764 25924 14773
rect 28080 14764 28132 14816
rect 30012 14832 30064 14884
rect 30380 14832 30432 14884
rect 33600 14832 33652 14884
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 1400 14560 1452 14612
rect 2688 14560 2740 14612
rect 3516 14603 3568 14612
rect 3516 14569 3525 14603
rect 3525 14569 3559 14603
rect 3559 14569 3568 14603
rect 3516 14560 3568 14569
rect 3884 14603 3936 14612
rect 3884 14569 3893 14603
rect 3893 14569 3927 14603
rect 3927 14569 3936 14603
rect 3884 14560 3936 14569
rect 4344 14603 4396 14612
rect 4344 14569 4353 14603
rect 4353 14569 4387 14603
rect 4387 14569 4396 14603
rect 4344 14560 4396 14569
rect 5356 14603 5408 14612
rect 5356 14569 5365 14603
rect 5365 14569 5399 14603
rect 5399 14569 5408 14603
rect 5356 14560 5408 14569
rect 6092 14603 6144 14612
rect 6092 14569 6101 14603
rect 6101 14569 6135 14603
rect 6135 14569 6144 14603
rect 6092 14560 6144 14569
rect 8116 14560 8168 14612
rect 8208 14560 8260 14612
rect 2504 14492 2556 14544
rect 4804 14492 4856 14544
rect 8484 14492 8536 14544
rect 9864 14492 9916 14544
rect 10876 14560 10928 14612
rect 11520 14560 11572 14612
rect 13360 14603 13412 14612
rect 13360 14569 13369 14603
rect 13369 14569 13403 14603
rect 13403 14569 13412 14603
rect 13360 14560 13412 14569
rect 14096 14560 14148 14612
rect 14924 14560 14976 14612
rect 15200 14560 15252 14612
rect 16212 14560 16264 14612
rect 17500 14603 17552 14612
rect 4068 14424 4120 14476
rect 6460 14467 6512 14476
rect 6460 14433 6469 14467
rect 6469 14433 6503 14467
rect 6503 14433 6512 14467
rect 6460 14424 6512 14433
rect 7932 14467 7984 14476
rect 7932 14433 7941 14467
rect 7941 14433 7975 14467
rect 7975 14433 7984 14467
rect 7932 14424 7984 14433
rect 8116 14467 8168 14476
rect 8116 14433 8125 14467
rect 8125 14433 8159 14467
rect 8159 14433 8168 14467
rect 8116 14424 8168 14433
rect 8208 14467 8260 14476
rect 8208 14433 8217 14467
rect 8217 14433 8251 14467
rect 8251 14433 8260 14467
rect 8208 14424 8260 14433
rect 9496 14424 9548 14476
rect 4896 14288 4948 14340
rect 5540 14288 5592 14340
rect 7196 14288 7248 14340
rect 7380 14288 7432 14340
rect 8576 14288 8628 14340
rect 9864 14288 9916 14340
rect 1584 14263 1636 14272
rect 1584 14229 1593 14263
rect 1593 14229 1627 14263
rect 1627 14229 1636 14263
rect 1584 14220 1636 14229
rect 5724 14263 5776 14272
rect 5724 14229 5733 14263
rect 5733 14229 5767 14263
rect 5767 14229 5776 14263
rect 5724 14220 5776 14229
rect 7932 14220 7984 14272
rect 8208 14220 8260 14272
rect 8668 14220 8720 14272
rect 9128 14220 9180 14272
rect 10232 14467 10284 14476
rect 10232 14433 10241 14467
rect 10241 14433 10275 14467
rect 10275 14433 10284 14467
rect 10232 14424 10284 14433
rect 10784 14492 10836 14544
rect 12256 14492 12308 14544
rect 12992 14492 13044 14544
rect 13636 14492 13688 14544
rect 15660 14492 15712 14544
rect 15936 14492 15988 14544
rect 12072 14424 12124 14476
rect 13268 14467 13320 14476
rect 13268 14433 13277 14467
rect 13277 14433 13311 14467
rect 13311 14433 13320 14467
rect 13268 14424 13320 14433
rect 15200 14424 15252 14476
rect 16580 14492 16632 14544
rect 17500 14569 17509 14603
rect 17509 14569 17543 14603
rect 17543 14569 17552 14603
rect 17500 14560 17552 14569
rect 17776 14603 17828 14612
rect 17776 14569 17785 14603
rect 17785 14569 17819 14603
rect 17819 14569 17828 14603
rect 17776 14560 17828 14569
rect 18144 14492 18196 14544
rect 18328 14535 18380 14544
rect 18328 14501 18337 14535
rect 18337 14501 18371 14535
rect 18371 14501 18380 14535
rect 18328 14492 18380 14501
rect 18788 14560 18840 14612
rect 19064 14603 19116 14612
rect 19064 14569 19073 14603
rect 19073 14569 19107 14603
rect 19107 14569 19116 14603
rect 19064 14560 19116 14569
rect 19248 14560 19300 14612
rect 19432 14560 19484 14612
rect 21732 14560 21784 14612
rect 22744 14603 22796 14612
rect 12348 14356 12400 14408
rect 13084 14399 13136 14408
rect 13084 14365 13093 14399
rect 13093 14365 13127 14399
rect 13127 14365 13136 14399
rect 13084 14356 13136 14365
rect 13912 14356 13964 14408
rect 15476 14356 15528 14408
rect 17500 14424 17552 14476
rect 18052 14424 18104 14476
rect 19340 14467 19392 14476
rect 19340 14433 19349 14467
rect 19349 14433 19383 14467
rect 19383 14433 19392 14467
rect 19340 14424 19392 14433
rect 19524 14535 19576 14544
rect 19524 14501 19533 14535
rect 19533 14501 19567 14535
rect 19567 14501 19576 14535
rect 19892 14535 19944 14544
rect 19524 14492 19576 14501
rect 19892 14501 19901 14535
rect 19901 14501 19935 14535
rect 19935 14501 19944 14535
rect 19892 14492 19944 14501
rect 22744 14569 22753 14603
rect 22753 14569 22787 14603
rect 22787 14569 22796 14603
rect 22744 14560 22796 14569
rect 25964 14560 26016 14612
rect 27344 14603 27396 14612
rect 27344 14569 27353 14603
rect 27353 14569 27387 14603
rect 27387 14569 27396 14603
rect 27344 14560 27396 14569
rect 27896 14603 27948 14612
rect 27896 14569 27905 14603
rect 27905 14569 27939 14603
rect 27939 14569 27948 14603
rect 27896 14560 27948 14569
rect 29920 14603 29972 14612
rect 29920 14569 29929 14603
rect 29929 14569 29963 14603
rect 29963 14569 29972 14603
rect 29920 14560 29972 14569
rect 30472 14560 30524 14612
rect 32588 14560 32640 14612
rect 33048 14603 33100 14612
rect 33048 14569 33057 14603
rect 33057 14569 33091 14603
rect 33091 14569 33100 14603
rect 33048 14560 33100 14569
rect 23480 14492 23532 14544
rect 26332 14492 26384 14544
rect 28264 14492 28316 14544
rect 20168 14424 20220 14476
rect 20996 14424 21048 14476
rect 21916 14467 21968 14476
rect 21916 14433 21925 14467
rect 21925 14433 21959 14467
rect 21959 14433 21968 14467
rect 21916 14424 21968 14433
rect 23940 14467 23992 14476
rect 10140 14288 10192 14340
rect 14004 14288 14056 14340
rect 10692 14220 10744 14272
rect 11336 14263 11388 14272
rect 11336 14229 11345 14263
rect 11345 14229 11379 14263
rect 11379 14229 11388 14263
rect 11336 14220 11388 14229
rect 11428 14220 11480 14272
rect 12072 14263 12124 14272
rect 12072 14229 12081 14263
rect 12081 14229 12115 14263
rect 12115 14229 12124 14263
rect 12072 14220 12124 14229
rect 12532 14263 12584 14272
rect 12532 14229 12541 14263
rect 12541 14229 12575 14263
rect 12575 14229 12584 14263
rect 12532 14220 12584 14229
rect 12900 14220 12952 14272
rect 19156 14399 19208 14408
rect 19156 14365 19165 14399
rect 19165 14365 19199 14399
rect 19199 14365 19208 14399
rect 19156 14356 19208 14365
rect 17776 14288 17828 14340
rect 18144 14288 18196 14340
rect 20260 14288 20312 14340
rect 23940 14433 23949 14467
rect 23949 14433 23983 14467
rect 23983 14433 23992 14467
rect 23940 14424 23992 14433
rect 24124 14467 24176 14476
rect 24124 14433 24130 14467
rect 24130 14433 24176 14467
rect 24124 14424 24176 14433
rect 23112 14356 23164 14408
rect 24308 14399 24360 14408
rect 24308 14365 24317 14399
rect 24317 14365 24351 14399
rect 24351 14365 24360 14399
rect 24308 14356 24360 14365
rect 25228 14356 25280 14408
rect 17132 14220 17184 14272
rect 22284 14220 22336 14272
rect 23848 14263 23900 14272
rect 23848 14229 23857 14263
rect 23857 14229 23891 14263
rect 23891 14229 23900 14263
rect 23848 14220 23900 14229
rect 24216 14263 24268 14272
rect 24216 14229 24225 14263
rect 24225 14229 24259 14263
rect 24259 14229 24268 14263
rect 24216 14220 24268 14229
rect 26792 14424 26844 14476
rect 31392 14492 31444 14544
rect 33600 14492 33652 14544
rect 26056 14356 26108 14408
rect 26516 14288 26568 14340
rect 29828 14424 29880 14476
rect 30380 14424 30432 14476
rect 31024 14424 31076 14476
rect 31668 14424 31720 14476
rect 32128 14467 32180 14476
rect 32128 14433 32137 14467
rect 32137 14433 32171 14467
rect 32171 14433 32180 14467
rect 32128 14424 32180 14433
rect 30196 14356 30248 14408
rect 31392 14356 31444 14408
rect 34152 14424 34204 14476
rect 33876 14356 33928 14408
rect 34336 14356 34388 14408
rect 29460 14331 29512 14340
rect 29460 14297 29469 14331
rect 29469 14297 29503 14331
rect 29503 14297 29512 14331
rect 29460 14288 29512 14297
rect 34244 14331 34296 14340
rect 34244 14297 34253 14331
rect 34253 14297 34287 14331
rect 34287 14297 34296 14331
rect 34244 14288 34296 14297
rect 26148 14220 26200 14272
rect 28448 14263 28500 14272
rect 28448 14229 28457 14263
rect 28457 14229 28491 14263
rect 28491 14229 28500 14263
rect 28448 14220 28500 14229
rect 31944 14263 31996 14272
rect 31944 14229 31953 14263
rect 31953 14229 31987 14263
rect 31987 14229 31996 14263
rect 31944 14220 31996 14229
rect 32588 14263 32640 14272
rect 32588 14229 32597 14263
rect 32597 14229 32631 14263
rect 32631 14229 32640 14263
rect 32588 14220 32640 14229
rect 33508 14220 33560 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 2688 14059 2740 14068
rect 2688 14025 2697 14059
rect 2697 14025 2731 14059
rect 2731 14025 2740 14059
rect 2688 14016 2740 14025
rect 4712 14016 4764 14068
rect 5448 14016 5500 14068
rect 6460 14016 6512 14068
rect 6920 13948 6972 14000
rect 2688 13812 2740 13864
rect 3976 13812 4028 13864
rect 6828 13855 6880 13864
rect 6828 13821 6837 13855
rect 6837 13821 6871 13855
rect 6871 13821 6880 13855
rect 6828 13812 6880 13821
rect 7012 13812 7064 13864
rect 9404 14016 9456 14068
rect 9220 13923 9272 13932
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 10232 14016 10284 14068
rect 10324 14016 10376 14068
rect 10876 14016 10928 14068
rect 13360 14016 13412 14068
rect 15384 14059 15436 14068
rect 15384 14025 15393 14059
rect 15393 14025 15427 14059
rect 15427 14025 15436 14059
rect 15384 14016 15436 14025
rect 15936 14059 15988 14068
rect 15936 14025 15945 14059
rect 15945 14025 15979 14059
rect 15979 14025 15988 14059
rect 15936 14016 15988 14025
rect 16580 14059 16632 14068
rect 16580 14025 16604 14059
rect 16604 14025 16632 14059
rect 16580 14016 16632 14025
rect 18052 14016 18104 14068
rect 18696 14016 18748 14068
rect 19340 14016 19392 14068
rect 20168 14016 20220 14068
rect 20996 14059 21048 14068
rect 20996 14025 21005 14059
rect 21005 14025 21039 14059
rect 21039 14025 21048 14059
rect 20996 14016 21048 14025
rect 23112 14059 23164 14068
rect 23112 14025 23121 14059
rect 23121 14025 23155 14059
rect 23155 14025 23164 14059
rect 23112 14016 23164 14025
rect 24308 14016 24360 14068
rect 25964 14016 26016 14068
rect 26148 14059 26200 14068
rect 26148 14025 26172 14059
rect 26172 14025 26200 14059
rect 26148 14016 26200 14025
rect 26608 14059 26660 14068
rect 26608 14025 26617 14059
rect 26617 14025 26651 14059
rect 26651 14025 26660 14059
rect 26608 14016 26660 14025
rect 26792 14016 26844 14068
rect 27804 14016 27856 14068
rect 28264 14016 28316 14068
rect 29828 14016 29880 14068
rect 30472 14016 30524 14068
rect 31760 14016 31812 14068
rect 32128 14016 32180 14068
rect 34152 14016 34204 14068
rect 12072 13948 12124 14000
rect 15108 13948 15160 14000
rect 16672 13991 16724 14000
rect 11060 13880 11112 13932
rect 11428 13880 11480 13932
rect 11704 13880 11756 13932
rect 13728 13880 13780 13932
rect 16672 13957 16681 13991
rect 16681 13957 16715 13991
rect 16715 13957 16724 13991
rect 16672 13948 16724 13957
rect 16856 13923 16908 13932
rect 16856 13889 16865 13923
rect 16865 13889 16899 13923
rect 16899 13889 16908 13923
rect 16856 13880 16908 13889
rect 10968 13812 11020 13864
rect 12532 13812 12584 13864
rect 8024 13744 8076 13796
rect 8576 13744 8628 13796
rect 9312 13744 9364 13796
rect 8668 13719 8720 13728
rect 8668 13685 8677 13719
rect 8677 13685 8711 13719
rect 8711 13685 8720 13719
rect 8668 13676 8720 13685
rect 9864 13719 9916 13728
rect 9864 13685 9873 13719
rect 9873 13685 9907 13719
rect 9907 13685 9916 13719
rect 10232 13719 10284 13728
rect 9864 13676 9916 13685
rect 10232 13685 10241 13719
rect 10241 13685 10275 13719
rect 10275 13685 10284 13719
rect 10232 13676 10284 13685
rect 11152 13719 11204 13728
rect 11152 13685 11161 13719
rect 11161 13685 11195 13719
rect 11195 13685 11204 13719
rect 11152 13676 11204 13685
rect 11336 13676 11388 13728
rect 11704 13676 11756 13728
rect 12900 13676 12952 13728
rect 14096 13812 14148 13864
rect 15200 13855 15252 13864
rect 15200 13821 15209 13855
rect 15209 13821 15243 13855
rect 15243 13821 15252 13855
rect 15200 13812 15252 13821
rect 16212 13812 16264 13864
rect 17684 13812 17736 13864
rect 19248 13880 19300 13932
rect 20260 13880 20312 13932
rect 18972 13855 19024 13864
rect 13728 13676 13780 13728
rect 14924 13744 14976 13796
rect 15476 13744 15528 13796
rect 17316 13744 17368 13796
rect 18972 13821 18981 13855
rect 18981 13821 19015 13855
rect 19015 13821 19024 13855
rect 18972 13812 19024 13821
rect 14188 13676 14240 13728
rect 15844 13676 15896 13728
rect 17776 13676 17828 13728
rect 18604 13744 18656 13796
rect 19064 13744 19116 13796
rect 21364 13948 21416 14000
rect 25872 13991 25924 14000
rect 25872 13957 25881 13991
rect 25881 13957 25915 13991
rect 25915 13957 25924 13991
rect 25872 13948 25924 13957
rect 26516 13948 26568 14000
rect 29920 13948 29972 14000
rect 31944 13948 31996 14000
rect 24032 13880 24084 13932
rect 20628 13812 20680 13864
rect 21732 13812 21784 13864
rect 22560 13812 22612 13864
rect 24400 13855 24452 13864
rect 24400 13821 24409 13855
rect 24409 13821 24443 13855
rect 24443 13821 24452 13855
rect 24400 13812 24452 13821
rect 25412 13880 25464 13932
rect 26332 13923 26384 13932
rect 26332 13889 26341 13923
rect 26341 13889 26375 13923
rect 26375 13889 26384 13923
rect 26332 13880 26384 13889
rect 25964 13855 26016 13864
rect 25964 13821 25973 13855
rect 25973 13821 26007 13855
rect 26007 13821 26016 13855
rect 25964 13812 26016 13821
rect 26700 13812 26752 13864
rect 27436 13855 27488 13864
rect 27436 13821 27445 13855
rect 27445 13821 27479 13855
rect 27479 13821 27488 13855
rect 27436 13812 27488 13821
rect 28448 13812 28500 13864
rect 29276 13855 29328 13864
rect 29276 13821 29285 13855
rect 29285 13821 29319 13855
rect 29319 13821 29328 13855
rect 29276 13812 29328 13821
rect 29460 13855 29512 13864
rect 29460 13821 29469 13855
rect 29469 13821 29503 13855
rect 29503 13821 29512 13855
rect 29460 13812 29512 13821
rect 30932 13855 30984 13864
rect 30932 13821 30941 13855
rect 30941 13821 30975 13855
rect 30975 13821 30984 13855
rect 30932 13812 30984 13821
rect 31392 13812 31444 13864
rect 25044 13744 25096 13796
rect 27896 13744 27948 13796
rect 28816 13744 28868 13796
rect 21824 13676 21876 13728
rect 23756 13676 23808 13728
rect 24216 13676 24268 13728
rect 30012 13787 30064 13796
rect 30012 13753 30021 13787
rect 30021 13753 30055 13787
rect 30055 13753 30064 13787
rect 30012 13744 30064 13753
rect 31576 13744 31628 13796
rect 32588 13812 32640 13864
rect 32864 13812 32916 13864
rect 33140 13855 33192 13864
rect 33140 13821 33149 13855
rect 33149 13821 33183 13855
rect 33183 13821 33192 13855
rect 33140 13812 33192 13821
rect 33600 13855 33652 13864
rect 33600 13821 33609 13855
rect 33609 13821 33643 13855
rect 33643 13821 33652 13855
rect 33600 13812 33652 13821
rect 34428 13812 34480 13864
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 5264 13515 5316 13524
rect 5264 13481 5273 13515
rect 5273 13481 5307 13515
rect 5307 13481 5316 13515
rect 5264 13472 5316 13481
rect 5632 13515 5684 13524
rect 5632 13481 5641 13515
rect 5641 13481 5675 13515
rect 5675 13481 5684 13515
rect 5632 13472 5684 13481
rect 6920 13472 6972 13524
rect 8116 13472 8168 13524
rect 8668 13472 8720 13524
rect 9772 13472 9824 13524
rect 9956 13472 10008 13524
rect 3056 13447 3108 13456
rect 3056 13413 3065 13447
rect 3065 13413 3099 13447
rect 3099 13413 3108 13447
rect 3056 13404 3108 13413
rect 1400 13379 1452 13388
rect 1400 13345 1409 13379
rect 1409 13345 1443 13379
rect 1443 13345 1452 13379
rect 1400 13336 1452 13345
rect 5724 13336 5776 13388
rect 5908 13336 5960 13388
rect 6184 13379 6236 13388
rect 6184 13345 6193 13379
rect 6193 13345 6227 13379
rect 6227 13345 6236 13379
rect 6184 13336 6236 13345
rect 6460 13336 6512 13388
rect 7012 13447 7064 13456
rect 7012 13413 7021 13447
rect 7021 13413 7055 13447
rect 7055 13413 7064 13447
rect 8392 13447 8444 13456
rect 7012 13404 7064 13413
rect 8392 13413 8401 13447
rect 8401 13413 8435 13447
rect 8435 13413 8444 13447
rect 8392 13404 8444 13413
rect 11704 13472 11756 13524
rect 12716 13472 12768 13524
rect 13452 13472 13504 13524
rect 13912 13515 13964 13524
rect 13912 13481 13921 13515
rect 13921 13481 13955 13515
rect 13955 13481 13964 13515
rect 13912 13472 13964 13481
rect 14372 13515 14424 13524
rect 14372 13481 14381 13515
rect 14381 13481 14415 13515
rect 14415 13481 14424 13515
rect 14372 13472 14424 13481
rect 15108 13472 15160 13524
rect 17132 13472 17184 13524
rect 10692 13404 10744 13456
rect 12348 13404 12400 13456
rect 14096 13404 14148 13456
rect 15936 13447 15988 13456
rect 15936 13413 15945 13447
rect 15945 13413 15979 13447
rect 15979 13413 15988 13447
rect 15936 13404 15988 13413
rect 16028 13404 16080 13456
rect 16580 13447 16632 13456
rect 16580 13413 16589 13447
rect 16589 13413 16623 13447
rect 16623 13413 16632 13447
rect 16580 13404 16632 13413
rect 16764 13404 16816 13456
rect 7932 13379 7984 13388
rect 7932 13345 7941 13379
rect 7941 13345 7975 13379
rect 7975 13345 7984 13379
rect 7932 13336 7984 13345
rect 1584 13268 1636 13320
rect 8024 13311 8076 13320
rect 8024 13277 8033 13311
rect 8033 13277 8067 13311
rect 8067 13277 8076 13311
rect 8024 13268 8076 13277
rect 8760 13311 8812 13320
rect 8760 13277 8769 13311
rect 8769 13277 8803 13311
rect 8803 13277 8812 13311
rect 8760 13268 8812 13277
rect 9864 13336 9916 13388
rect 10324 13336 10376 13388
rect 11152 13379 11204 13388
rect 11152 13345 11161 13379
rect 11161 13345 11195 13379
rect 11195 13345 11204 13379
rect 11152 13336 11204 13345
rect 11980 13336 12032 13388
rect 12716 13379 12768 13388
rect 12716 13345 12725 13379
rect 12725 13345 12759 13379
rect 12759 13345 12768 13379
rect 12716 13336 12768 13345
rect 12900 13379 12952 13388
rect 12900 13345 12909 13379
rect 12909 13345 12943 13379
rect 12943 13345 12952 13379
rect 12900 13336 12952 13345
rect 13084 13336 13136 13388
rect 13728 13336 13780 13388
rect 14188 13336 14240 13388
rect 14740 13336 14792 13388
rect 15384 13336 15436 13388
rect 17316 13336 17368 13388
rect 17500 13472 17552 13524
rect 19248 13472 19300 13524
rect 19340 13472 19392 13524
rect 20720 13515 20772 13524
rect 20720 13481 20729 13515
rect 20729 13481 20763 13515
rect 20763 13481 20772 13515
rect 20720 13472 20772 13481
rect 20996 13472 21048 13524
rect 22100 13472 22152 13524
rect 23848 13472 23900 13524
rect 25044 13515 25096 13524
rect 25044 13481 25053 13515
rect 25053 13481 25087 13515
rect 25087 13481 25096 13515
rect 25044 13472 25096 13481
rect 25412 13515 25464 13524
rect 25412 13481 25421 13515
rect 25421 13481 25455 13515
rect 25455 13481 25464 13515
rect 25412 13472 25464 13481
rect 26700 13515 26752 13524
rect 26700 13481 26709 13515
rect 26709 13481 26743 13515
rect 26743 13481 26752 13515
rect 26700 13472 26752 13481
rect 26792 13472 26844 13524
rect 27712 13472 27764 13524
rect 29276 13515 29328 13524
rect 29276 13481 29285 13515
rect 29285 13481 29319 13515
rect 29319 13481 29328 13515
rect 29276 13472 29328 13481
rect 31024 13472 31076 13524
rect 31576 13515 31628 13524
rect 31576 13481 31585 13515
rect 31585 13481 31619 13515
rect 31619 13481 31628 13515
rect 31576 13472 31628 13481
rect 31944 13472 31996 13524
rect 33140 13515 33192 13524
rect 33140 13481 33149 13515
rect 33149 13481 33183 13515
rect 33183 13481 33192 13515
rect 33140 13472 33192 13481
rect 33600 13515 33652 13524
rect 33600 13481 33609 13515
rect 33609 13481 33643 13515
rect 33643 13481 33652 13515
rect 33600 13472 33652 13481
rect 33876 13515 33928 13524
rect 33876 13481 33885 13515
rect 33885 13481 33919 13515
rect 33919 13481 33928 13515
rect 33876 13472 33928 13481
rect 17960 13404 18012 13456
rect 18604 13447 18656 13456
rect 18052 13379 18104 13388
rect 18052 13345 18061 13379
rect 18061 13345 18095 13379
rect 18095 13345 18104 13379
rect 18052 13336 18104 13345
rect 18604 13413 18613 13447
rect 18613 13413 18647 13447
rect 18647 13413 18656 13447
rect 18604 13404 18656 13413
rect 28264 13404 28316 13456
rect 18788 13336 18840 13388
rect 18972 13336 19024 13388
rect 19892 13336 19944 13388
rect 21456 13379 21508 13388
rect 21456 13345 21465 13379
rect 21465 13345 21499 13379
rect 21499 13345 21508 13379
rect 21456 13336 21508 13345
rect 22560 13336 22612 13388
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 16672 13268 16724 13320
rect 17776 13268 17828 13320
rect 4068 13200 4120 13252
rect 5080 13200 5132 13252
rect 8668 13200 8720 13252
rect 13268 13243 13320 13252
rect 13268 13209 13277 13243
rect 13277 13209 13311 13243
rect 13311 13209 13320 13243
rect 13268 13200 13320 13209
rect 14740 13200 14792 13252
rect 15476 13243 15528 13252
rect 15476 13209 15485 13243
rect 15485 13209 15519 13243
rect 15519 13209 15528 13243
rect 15476 13200 15528 13209
rect 19432 13200 19484 13252
rect 24124 13336 24176 13388
rect 25228 13379 25280 13388
rect 25228 13345 25237 13379
rect 25237 13345 25271 13379
rect 25271 13345 25280 13379
rect 25228 13336 25280 13345
rect 26056 13336 26108 13388
rect 27804 13336 27856 13388
rect 28356 13379 28408 13388
rect 28356 13345 28365 13379
rect 28365 13345 28399 13379
rect 28399 13345 28408 13379
rect 28356 13336 28408 13345
rect 29552 13404 29604 13456
rect 30104 13404 30156 13456
rect 29828 13336 29880 13388
rect 30196 13336 30248 13388
rect 31760 13336 31812 13388
rect 32496 13336 32548 13388
rect 24216 13268 24268 13320
rect 27252 13268 27304 13320
rect 31116 13311 31168 13320
rect 31116 13277 31125 13311
rect 31125 13277 31159 13311
rect 31159 13277 31168 13311
rect 31116 13268 31168 13277
rect 22928 13200 22980 13252
rect 27620 13200 27672 13252
rect 30012 13200 30064 13252
rect 30564 13200 30616 13252
rect 32864 13268 32916 13320
rect 4896 13175 4948 13184
rect 4896 13141 4905 13175
rect 4905 13141 4939 13175
rect 4939 13141 4948 13175
rect 4896 13132 4948 13141
rect 9864 13175 9916 13184
rect 9864 13141 9873 13175
rect 9873 13141 9907 13175
rect 9907 13141 9916 13175
rect 9864 13132 9916 13141
rect 10232 13175 10284 13184
rect 10232 13141 10241 13175
rect 10241 13141 10275 13175
rect 10275 13141 10284 13175
rect 10232 13132 10284 13141
rect 11336 13132 11388 13184
rect 12256 13175 12308 13184
rect 12256 13141 12265 13175
rect 12265 13141 12299 13175
rect 12299 13141 12308 13175
rect 12256 13132 12308 13141
rect 15108 13175 15160 13184
rect 15108 13141 15117 13175
rect 15117 13141 15151 13175
rect 15151 13141 15160 13175
rect 15108 13132 15160 13141
rect 17500 13132 17552 13184
rect 21916 13132 21968 13184
rect 23756 13132 23808 13184
rect 28816 13132 28868 13184
rect 29276 13132 29328 13184
rect 31852 13175 31904 13184
rect 31852 13141 31861 13175
rect 31861 13141 31895 13175
rect 31895 13141 31904 13175
rect 31852 13132 31904 13141
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 6184 12928 6236 12980
rect 5724 12860 5776 12912
rect 6460 12860 6512 12912
rect 1400 12792 1452 12844
rect 6920 12835 6972 12844
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 6920 12792 6972 12801
rect 8668 12928 8720 12980
rect 10692 12971 10744 12980
rect 10692 12937 10701 12971
rect 10701 12937 10735 12971
rect 10735 12937 10744 12971
rect 10692 12928 10744 12937
rect 11612 12928 11664 12980
rect 11796 12971 11848 12980
rect 11796 12937 11805 12971
rect 11805 12937 11839 12971
rect 11839 12937 11848 12971
rect 11796 12928 11848 12937
rect 12164 12928 12216 12980
rect 9588 12860 9640 12912
rect 10324 12903 10376 12912
rect 10324 12869 10333 12903
rect 10333 12869 10367 12903
rect 10367 12869 10376 12903
rect 10324 12860 10376 12869
rect 11060 12903 11112 12912
rect 11060 12869 11069 12903
rect 11069 12869 11103 12903
rect 11103 12869 11112 12903
rect 11060 12860 11112 12869
rect 11244 12903 11296 12912
rect 11244 12869 11253 12903
rect 11253 12869 11287 12903
rect 11287 12869 11296 12903
rect 11244 12860 11296 12869
rect 8852 12792 8904 12844
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 12716 12928 12768 12980
rect 13636 12928 13688 12980
rect 15108 12928 15160 12980
rect 16304 12928 16356 12980
rect 16580 12928 16632 12980
rect 18972 12971 19024 12980
rect 18972 12937 18981 12971
rect 18981 12937 19015 12971
rect 19015 12937 19024 12971
rect 18972 12928 19024 12937
rect 20996 12928 21048 12980
rect 24124 12971 24176 12980
rect 24124 12937 24133 12971
rect 24133 12937 24167 12971
rect 24167 12937 24176 12971
rect 24124 12928 24176 12937
rect 25228 12971 25280 12980
rect 25228 12937 25237 12971
rect 25237 12937 25271 12971
rect 25271 12937 25280 12971
rect 25228 12928 25280 12937
rect 26700 12928 26752 12980
rect 26976 12928 27028 12980
rect 27896 12928 27948 12980
rect 28632 12928 28684 12980
rect 30196 12971 30248 12980
rect 30196 12937 30205 12971
rect 30205 12937 30239 12971
rect 30239 12937 30248 12971
rect 30196 12928 30248 12937
rect 30564 12971 30616 12980
rect 30564 12937 30573 12971
rect 30573 12937 30607 12971
rect 30607 12937 30616 12971
rect 30564 12928 30616 12937
rect 32496 12971 32548 12980
rect 32496 12937 32505 12971
rect 32505 12937 32539 12971
rect 32539 12937 32548 12971
rect 32496 12928 32548 12937
rect 32864 12971 32916 12980
rect 32864 12937 32873 12971
rect 32873 12937 32907 12971
rect 32907 12937 32916 12971
rect 32864 12928 32916 12937
rect 8668 12724 8720 12776
rect 8760 12724 8812 12776
rect 9588 12724 9640 12776
rect 9772 12767 9824 12776
rect 9772 12733 9781 12767
rect 9781 12733 9815 12767
rect 9815 12733 9824 12767
rect 9772 12724 9824 12733
rect 10324 12724 10376 12776
rect 12256 12724 12308 12776
rect 12900 12792 12952 12844
rect 13912 12835 13964 12844
rect 13912 12801 13921 12835
rect 13921 12801 13955 12835
rect 13955 12801 13964 12835
rect 13912 12792 13964 12801
rect 15936 12860 15988 12912
rect 22468 12903 22520 12912
rect 22468 12869 22477 12903
rect 22477 12869 22511 12903
rect 22511 12869 22520 12903
rect 22468 12860 22520 12869
rect 24032 12903 24084 12912
rect 24032 12869 24056 12903
rect 24056 12869 24084 12903
rect 24032 12860 24084 12869
rect 24676 12860 24728 12912
rect 26332 12903 26384 12912
rect 26332 12869 26341 12903
rect 26341 12869 26375 12903
rect 26375 12869 26384 12903
rect 26332 12860 26384 12869
rect 13452 12724 13504 12776
rect 15108 12792 15160 12844
rect 15384 12792 15436 12844
rect 17776 12835 17828 12844
rect 17776 12801 17785 12835
rect 17785 12801 17819 12835
rect 17819 12801 17828 12835
rect 17776 12792 17828 12801
rect 19156 12792 19208 12844
rect 19340 12835 19392 12844
rect 19340 12801 19349 12835
rect 19349 12801 19383 12835
rect 19383 12801 19392 12835
rect 24216 12835 24268 12844
rect 19340 12792 19392 12801
rect 24216 12801 24225 12835
rect 24225 12801 24259 12835
rect 24259 12801 24268 12835
rect 24216 12792 24268 12801
rect 25504 12792 25556 12844
rect 25872 12792 25924 12844
rect 27620 12835 27672 12844
rect 27620 12801 27629 12835
rect 27629 12801 27663 12835
rect 27663 12801 27672 12835
rect 27620 12792 27672 12801
rect 32772 12860 32824 12912
rect 7472 12656 7524 12708
rect 9312 12656 9364 12708
rect 9864 12656 9916 12708
rect 10968 12656 11020 12708
rect 12532 12656 12584 12708
rect 12900 12656 12952 12708
rect 13084 12656 13136 12708
rect 5540 12588 5592 12640
rect 7012 12588 7064 12640
rect 11612 12588 11664 12640
rect 11980 12588 12032 12640
rect 14096 12724 14148 12776
rect 14556 12767 14608 12776
rect 14556 12733 14565 12767
rect 14565 12733 14599 12767
rect 14599 12733 14608 12767
rect 14556 12724 14608 12733
rect 14740 12724 14792 12776
rect 15844 12767 15896 12776
rect 15844 12733 15853 12767
rect 15853 12733 15887 12767
rect 15887 12733 15896 12767
rect 15844 12724 15896 12733
rect 17316 12724 17368 12776
rect 18604 12724 18656 12776
rect 15016 12656 15068 12708
rect 19432 12724 19484 12776
rect 20996 12724 21048 12776
rect 21824 12767 21876 12776
rect 21824 12733 21833 12767
rect 21833 12733 21867 12767
rect 21867 12733 21876 12767
rect 21824 12724 21876 12733
rect 22100 12767 22152 12776
rect 22100 12733 22109 12767
rect 22109 12733 22143 12767
rect 22143 12733 22152 12767
rect 22560 12767 22612 12776
rect 22100 12724 22152 12733
rect 22560 12733 22569 12767
rect 22569 12733 22603 12767
rect 22603 12733 22612 12767
rect 22560 12724 22612 12733
rect 23848 12767 23900 12776
rect 23848 12733 23857 12767
rect 23857 12733 23891 12767
rect 23891 12733 23900 12767
rect 23848 12724 23900 12733
rect 19984 12656 20036 12708
rect 20168 12656 20220 12708
rect 20812 12699 20864 12708
rect 20812 12665 20821 12699
rect 20821 12665 20855 12699
rect 20855 12665 20864 12699
rect 20812 12656 20864 12665
rect 23572 12656 23624 12708
rect 23940 12656 23992 12708
rect 26056 12767 26108 12776
rect 26056 12733 26065 12767
rect 26065 12733 26099 12767
rect 26099 12733 26108 12767
rect 26056 12724 26108 12733
rect 26332 12724 26384 12776
rect 27712 12724 27764 12776
rect 14372 12588 14424 12640
rect 15384 12631 15436 12640
rect 15384 12597 15393 12631
rect 15393 12597 15427 12631
rect 15427 12597 15436 12631
rect 15384 12588 15436 12597
rect 15476 12588 15528 12640
rect 16028 12588 16080 12640
rect 17960 12588 18012 12640
rect 19156 12588 19208 12640
rect 23296 12588 23348 12640
rect 26608 12656 26660 12708
rect 26792 12699 26844 12708
rect 26792 12665 26801 12699
rect 26801 12665 26835 12699
rect 26835 12665 26844 12699
rect 26792 12656 26844 12665
rect 27344 12656 27396 12708
rect 27804 12699 27856 12708
rect 24492 12631 24544 12640
rect 24492 12597 24501 12631
rect 24501 12597 24535 12631
rect 24535 12597 24544 12631
rect 24492 12588 24544 12597
rect 26240 12588 26292 12640
rect 26516 12588 26568 12640
rect 27804 12665 27813 12699
rect 27813 12665 27847 12699
rect 27847 12665 27856 12699
rect 27804 12656 27856 12665
rect 28264 12792 28316 12844
rect 30380 12792 30432 12844
rect 37280 12835 37332 12844
rect 29552 12767 29604 12776
rect 29552 12733 29561 12767
rect 29561 12733 29595 12767
rect 29595 12733 29604 12767
rect 29552 12724 29604 12733
rect 30656 12724 30708 12776
rect 31116 12767 31168 12776
rect 31116 12733 31125 12767
rect 31125 12733 31159 12767
rect 31159 12733 31168 12767
rect 31116 12724 31168 12733
rect 31668 12767 31720 12776
rect 31668 12733 31677 12767
rect 31677 12733 31711 12767
rect 31711 12733 31720 12767
rect 31668 12724 31720 12733
rect 31944 12767 31996 12776
rect 31944 12733 31953 12767
rect 31953 12733 31987 12767
rect 31987 12733 31996 12767
rect 31944 12724 31996 12733
rect 35808 12767 35860 12776
rect 35808 12733 35817 12767
rect 35817 12733 35851 12767
rect 35851 12733 35860 12767
rect 35808 12724 35860 12733
rect 37280 12801 37289 12835
rect 37289 12801 37323 12835
rect 37323 12801 37332 12835
rect 37280 12792 37332 12801
rect 37188 12724 37240 12776
rect 30564 12656 30616 12708
rect 28264 12588 28316 12640
rect 28448 12588 28500 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 5264 12427 5316 12436
rect 5264 12393 5273 12427
rect 5273 12393 5307 12427
rect 5307 12393 5316 12427
rect 5264 12384 5316 12393
rect 5540 12384 5592 12436
rect 6828 12384 6880 12436
rect 5816 12316 5868 12368
rect 6552 12316 6604 12368
rect 1584 12248 1636 12300
rect 3148 12291 3200 12300
rect 3148 12257 3157 12291
rect 3157 12257 3191 12291
rect 3191 12257 3200 12291
rect 3148 12248 3200 12257
rect 4620 12248 4672 12300
rect 6828 12291 6880 12300
rect 1952 12180 2004 12232
rect 4712 12112 4764 12164
rect 6828 12257 6837 12291
rect 6837 12257 6871 12291
rect 6871 12257 6880 12291
rect 6828 12248 6880 12257
rect 7932 12384 7984 12436
rect 8024 12427 8076 12436
rect 8024 12393 8033 12427
rect 8033 12393 8067 12427
rect 8067 12393 8076 12427
rect 8668 12427 8720 12436
rect 8024 12384 8076 12393
rect 8668 12393 8677 12427
rect 8677 12393 8711 12427
rect 8711 12393 8720 12427
rect 8668 12384 8720 12393
rect 8760 12384 8812 12436
rect 9956 12384 10008 12436
rect 11612 12427 11664 12436
rect 11612 12393 11621 12427
rect 11621 12393 11655 12427
rect 11655 12393 11664 12427
rect 11612 12384 11664 12393
rect 11796 12384 11848 12436
rect 12624 12427 12676 12436
rect 12624 12393 12633 12427
rect 12633 12393 12667 12427
rect 12667 12393 12676 12427
rect 12624 12384 12676 12393
rect 14188 12384 14240 12436
rect 15476 12384 15528 12436
rect 16580 12384 16632 12436
rect 16856 12384 16908 12436
rect 17408 12384 17460 12436
rect 11152 12316 11204 12368
rect 12440 12316 12492 12368
rect 13084 12316 13136 12368
rect 14096 12359 14148 12368
rect 14096 12325 14105 12359
rect 14105 12325 14139 12359
rect 14139 12325 14148 12359
rect 14096 12316 14148 12325
rect 14924 12316 14976 12368
rect 8208 12291 8260 12300
rect 8208 12257 8217 12291
rect 8217 12257 8251 12291
rect 8251 12257 8260 12291
rect 8208 12248 8260 12257
rect 9680 12291 9732 12300
rect 9680 12257 9689 12291
rect 9689 12257 9723 12291
rect 9723 12257 9732 12291
rect 10784 12291 10836 12300
rect 9680 12248 9732 12257
rect 10784 12257 10793 12291
rect 10793 12257 10827 12291
rect 10827 12257 10836 12291
rect 10784 12248 10836 12257
rect 11888 12248 11940 12300
rect 12164 12248 12216 12300
rect 14556 12248 14608 12300
rect 15384 12248 15436 12300
rect 16580 12291 16632 12300
rect 6276 12180 6328 12232
rect 7288 12223 7340 12232
rect 7288 12189 7297 12223
rect 7297 12189 7331 12223
rect 7331 12189 7340 12223
rect 7288 12180 7340 12189
rect 9956 12180 10008 12232
rect 11980 12180 12032 12232
rect 12900 12180 12952 12232
rect 13360 12180 13412 12232
rect 6460 12112 6512 12164
rect 9496 12112 9548 12164
rect 9772 12112 9824 12164
rect 10968 12112 11020 12164
rect 11336 12112 11388 12164
rect 14740 12180 14792 12232
rect 4620 12087 4672 12096
rect 4620 12053 4629 12087
rect 4629 12053 4663 12087
rect 4663 12053 4672 12087
rect 4620 12044 4672 12053
rect 5080 12044 5132 12096
rect 7472 12044 7524 12096
rect 9588 12044 9640 12096
rect 9680 12044 9732 12096
rect 13360 12044 13412 12096
rect 14740 12044 14792 12096
rect 16580 12257 16589 12291
rect 16589 12257 16623 12291
rect 16623 12257 16632 12291
rect 16580 12248 16632 12257
rect 16948 12248 17000 12300
rect 18052 12384 18104 12436
rect 18512 12384 18564 12436
rect 18696 12384 18748 12436
rect 18788 12384 18840 12436
rect 20168 12384 20220 12436
rect 16488 12180 16540 12232
rect 16672 12223 16724 12232
rect 16672 12189 16681 12223
rect 16681 12189 16715 12223
rect 16715 12189 16724 12223
rect 16672 12180 16724 12189
rect 17132 12223 17184 12232
rect 17132 12189 17141 12223
rect 17141 12189 17175 12223
rect 17175 12189 17184 12223
rect 17132 12180 17184 12189
rect 16948 12112 17000 12164
rect 17224 12112 17276 12164
rect 18052 12248 18104 12300
rect 22100 12427 22152 12436
rect 22100 12393 22109 12427
rect 22109 12393 22143 12427
rect 22143 12393 22152 12427
rect 22928 12427 22980 12436
rect 22100 12384 22152 12393
rect 22928 12393 22937 12427
rect 22937 12393 22971 12427
rect 22971 12393 22980 12427
rect 22928 12384 22980 12393
rect 23204 12384 23256 12436
rect 24676 12427 24728 12436
rect 24676 12393 24685 12427
rect 24685 12393 24719 12427
rect 24719 12393 24728 12427
rect 24676 12384 24728 12393
rect 26332 12384 26384 12436
rect 26700 12427 26752 12436
rect 26700 12393 26709 12427
rect 26709 12393 26743 12427
rect 26743 12393 26752 12427
rect 26700 12384 26752 12393
rect 27436 12384 27488 12436
rect 28356 12384 28408 12436
rect 28816 12427 28868 12436
rect 28816 12393 28825 12427
rect 28825 12393 28859 12427
rect 28859 12393 28868 12427
rect 28816 12384 28868 12393
rect 29552 12384 29604 12436
rect 30472 12427 30524 12436
rect 30472 12393 30481 12427
rect 30481 12393 30515 12427
rect 30515 12393 30524 12427
rect 30472 12384 30524 12393
rect 30564 12384 30616 12436
rect 32496 12384 32548 12436
rect 35900 12384 35952 12436
rect 36176 12384 36228 12436
rect 22560 12316 22612 12368
rect 19524 12291 19576 12300
rect 19524 12257 19533 12291
rect 19533 12257 19567 12291
rect 19567 12257 19576 12291
rect 19524 12248 19576 12257
rect 20904 12291 20956 12300
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 22100 12248 22152 12300
rect 22376 12291 22428 12300
rect 22376 12257 22385 12291
rect 22385 12257 22419 12291
rect 22419 12257 22428 12291
rect 22376 12248 22428 12257
rect 17592 12223 17644 12232
rect 17592 12189 17601 12223
rect 17601 12189 17635 12223
rect 17635 12189 17644 12223
rect 17592 12180 17644 12189
rect 18880 12180 18932 12232
rect 22008 12180 22060 12232
rect 23756 12316 23808 12368
rect 23480 12248 23532 12300
rect 24492 12248 24544 12300
rect 24860 12291 24912 12300
rect 24860 12257 24869 12291
rect 24869 12257 24903 12291
rect 24903 12257 24912 12291
rect 24860 12248 24912 12257
rect 24952 12180 25004 12232
rect 25596 12291 25648 12300
rect 25596 12257 25605 12291
rect 25605 12257 25639 12291
rect 25639 12257 25648 12291
rect 25596 12248 25648 12257
rect 26332 12248 26384 12300
rect 26976 12248 27028 12300
rect 28632 12291 28684 12300
rect 16120 12044 16172 12096
rect 16488 12044 16540 12096
rect 18328 12044 18380 12096
rect 20536 12044 20588 12096
rect 21456 12112 21508 12164
rect 23756 12112 23808 12164
rect 24124 12112 24176 12164
rect 25136 12155 25188 12164
rect 25136 12121 25145 12155
rect 25145 12121 25179 12155
rect 25179 12121 25188 12155
rect 25136 12112 25188 12121
rect 26608 12180 26660 12232
rect 27252 12180 27304 12232
rect 28632 12257 28641 12291
rect 28641 12257 28675 12291
rect 28675 12257 28684 12291
rect 28632 12248 28684 12257
rect 29644 12291 29696 12300
rect 29644 12257 29653 12291
rect 29653 12257 29687 12291
rect 29687 12257 29696 12291
rect 29644 12248 29696 12257
rect 30932 12248 30984 12300
rect 32496 12248 32548 12300
rect 32864 12248 32916 12300
rect 23296 12044 23348 12096
rect 25044 12087 25096 12096
rect 25044 12053 25068 12087
rect 25068 12053 25096 12087
rect 25044 12044 25096 12053
rect 25596 12044 25648 12096
rect 26148 12044 26200 12096
rect 27712 12112 27764 12164
rect 31024 12112 31076 12164
rect 27344 12087 27396 12096
rect 27344 12053 27353 12087
rect 27353 12053 27387 12087
rect 27387 12053 27396 12087
rect 27344 12044 27396 12053
rect 31484 12087 31536 12096
rect 31484 12053 31493 12087
rect 31493 12053 31527 12087
rect 31527 12053 31536 12087
rect 31484 12044 31536 12053
rect 31944 12044 31996 12096
rect 35808 12087 35860 12096
rect 35808 12053 35817 12087
rect 35817 12053 35851 12087
rect 35851 12053 35860 12087
rect 35808 12044 35860 12053
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 6276 11840 6328 11892
rect 7288 11883 7340 11892
rect 7288 11849 7297 11883
rect 7297 11849 7331 11883
rect 7331 11849 7340 11883
rect 7288 11840 7340 11849
rect 8208 11883 8260 11892
rect 8208 11849 8217 11883
rect 8217 11849 8251 11883
rect 8251 11849 8260 11883
rect 8208 11840 8260 11849
rect 9680 11840 9732 11892
rect 11888 11883 11940 11892
rect 11888 11849 11897 11883
rect 11897 11849 11931 11883
rect 11931 11849 11940 11883
rect 11888 11840 11940 11849
rect 14556 11840 14608 11892
rect 17408 11840 17460 11892
rect 4712 11772 4764 11824
rect 6552 11772 6604 11824
rect 11980 11772 12032 11824
rect 16120 11772 16172 11824
rect 3056 11704 3108 11756
rect 4620 11704 4672 11756
rect 7932 11704 7984 11756
rect 9772 11704 9824 11756
rect 12164 11704 12216 11756
rect 1952 11636 2004 11688
rect 3424 11679 3476 11688
rect 3424 11645 3433 11679
rect 3433 11645 3467 11679
rect 3467 11645 3476 11679
rect 3424 11636 3476 11645
rect 6644 11679 6696 11688
rect 6644 11645 6653 11679
rect 6653 11645 6687 11679
rect 6687 11645 6696 11679
rect 6644 11636 6696 11645
rect 5080 11611 5132 11620
rect 5080 11577 5089 11611
rect 5089 11577 5123 11611
rect 5123 11577 5132 11611
rect 5080 11568 5132 11577
rect 8300 11636 8352 11688
rect 8944 11636 8996 11688
rect 11336 11636 11388 11688
rect 13820 11704 13872 11756
rect 14740 11747 14792 11756
rect 14740 11713 14749 11747
rect 14749 11713 14783 11747
rect 14783 11713 14792 11747
rect 14740 11704 14792 11713
rect 16028 11704 16080 11756
rect 13084 11679 13136 11688
rect 13084 11645 13093 11679
rect 13093 11645 13127 11679
rect 13127 11645 13136 11679
rect 13084 11636 13136 11645
rect 13268 11679 13320 11688
rect 13268 11645 13277 11679
rect 13277 11645 13311 11679
rect 13311 11645 13320 11679
rect 13268 11636 13320 11645
rect 13360 11636 13412 11688
rect 14924 11679 14976 11688
rect 9404 11568 9456 11620
rect 14924 11645 14933 11679
rect 14933 11645 14967 11679
rect 14967 11645 14976 11679
rect 14924 11636 14976 11645
rect 15384 11679 15436 11688
rect 15384 11645 15393 11679
rect 15393 11645 15427 11679
rect 15427 11645 15436 11679
rect 15384 11636 15436 11645
rect 16764 11636 16816 11688
rect 17868 11840 17920 11892
rect 18880 11840 18932 11892
rect 19524 11883 19576 11892
rect 19524 11849 19533 11883
rect 19533 11849 19567 11883
rect 19567 11849 19576 11883
rect 19524 11840 19576 11849
rect 20904 11883 20956 11892
rect 20904 11849 20913 11883
rect 20913 11849 20947 11883
rect 20947 11849 20956 11883
rect 20904 11840 20956 11849
rect 23480 11883 23532 11892
rect 23480 11849 23489 11883
rect 23489 11849 23523 11883
rect 23523 11849 23532 11883
rect 23480 11840 23532 11849
rect 23848 11840 23900 11892
rect 24124 11840 24176 11892
rect 25136 11840 25188 11892
rect 27252 11883 27304 11892
rect 27252 11849 27261 11883
rect 27261 11849 27295 11883
rect 27295 11849 27304 11883
rect 27252 11840 27304 11849
rect 27712 11883 27764 11892
rect 27712 11849 27721 11883
rect 27721 11849 27755 11883
rect 27755 11849 27764 11883
rect 27712 11840 27764 11849
rect 28264 11840 28316 11892
rect 28632 11883 28684 11892
rect 28632 11849 28641 11883
rect 28641 11849 28675 11883
rect 28675 11849 28684 11883
rect 28632 11840 28684 11849
rect 29644 11883 29696 11892
rect 29644 11849 29653 11883
rect 29653 11849 29687 11883
rect 29687 11849 29696 11883
rect 29644 11840 29696 11849
rect 30748 11840 30800 11892
rect 32864 11883 32916 11892
rect 32864 11849 32873 11883
rect 32873 11849 32907 11883
rect 32907 11849 32916 11883
rect 32864 11840 32916 11849
rect 37280 11840 37332 11892
rect 22376 11772 22428 11824
rect 25228 11772 25280 11824
rect 19156 11704 19208 11756
rect 22560 11747 22612 11756
rect 22560 11713 22569 11747
rect 22569 11713 22603 11747
rect 22603 11713 22612 11747
rect 22560 11704 22612 11713
rect 26792 11704 26844 11756
rect 30932 11772 30984 11824
rect 31668 11747 31720 11756
rect 31668 11713 31677 11747
rect 31677 11713 31711 11747
rect 31711 11713 31720 11747
rect 31668 11704 31720 11713
rect 18328 11636 18380 11688
rect 20628 11636 20680 11688
rect 21824 11679 21876 11688
rect 21824 11645 21833 11679
rect 21833 11645 21867 11679
rect 21867 11645 21876 11679
rect 21824 11636 21876 11645
rect 22008 11679 22060 11688
rect 22008 11645 22017 11679
rect 22017 11645 22051 11679
rect 22051 11645 22060 11679
rect 22008 11636 22060 11645
rect 22100 11636 22152 11688
rect 24032 11636 24084 11688
rect 24860 11636 24912 11688
rect 25044 11636 25096 11688
rect 26700 11679 26752 11688
rect 26700 11645 26709 11679
rect 26709 11645 26743 11679
rect 26743 11645 26752 11679
rect 26700 11636 26752 11645
rect 27804 11679 27856 11688
rect 27804 11645 27813 11679
rect 27813 11645 27847 11679
rect 27847 11645 27856 11679
rect 27804 11636 27856 11645
rect 31024 11636 31076 11688
rect 18052 11611 18104 11620
rect 18052 11577 18061 11611
rect 18061 11577 18095 11611
rect 18095 11577 18104 11611
rect 18052 11568 18104 11577
rect 35808 11679 35860 11688
rect 35808 11645 35817 11679
rect 35817 11645 35851 11679
rect 35851 11645 35860 11679
rect 35808 11636 35860 11645
rect 36084 11679 36136 11688
rect 36084 11645 36093 11679
rect 36093 11645 36127 11679
rect 36127 11645 36136 11679
rect 36084 11636 36136 11645
rect 1492 11500 1544 11552
rect 1952 11543 2004 11552
rect 1952 11509 1961 11543
rect 1961 11509 1995 11543
rect 1995 11509 2004 11543
rect 1952 11500 2004 11509
rect 6460 11543 6512 11552
rect 6460 11509 6469 11543
rect 6469 11509 6503 11543
rect 6503 11509 6512 11543
rect 6460 11500 6512 11509
rect 10784 11500 10836 11552
rect 11060 11500 11112 11552
rect 11520 11500 11572 11552
rect 12532 11543 12584 11552
rect 12532 11509 12541 11543
rect 12541 11509 12575 11543
rect 12575 11509 12584 11543
rect 12532 11500 12584 11509
rect 16764 11500 16816 11552
rect 17132 11500 17184 11552
rect 24952 11500 25004 11552
rect 30380 11543 30432 11552
rect 30380 11509 30389 11543
rect 30389 11509 30423 11543
rect 30423 11509 30432 11543
rect 30380 11500 30432 11509
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 6644 11296 6696 11348
rect 8208 11296 8260 11348
rect 9404 11339 9456 11348
rect 9404 11305 9413 11339
rect 9413 11305 9447 11339
rect 9447 11305 9456 11339
rect 9404 11296 9456 11305
rect 10048 11296 10100 11348
rect 10232 11296 10284 11348
rect 10600 11296 10652 11348
rect 13268 11296 13320 11348
rect 14740 11339 14792 11348
rect 14740 11305 14749 11339
rect 14749 11305 14783 11339
rect 14783 11305 14792 11339
rect 14740 11296 14792 11305
rect 15200 11296 15252 11348
rect 17224 11296 17276 11348
rect 18328 11296 18380 11348
rect 18604 11296 18656 11348
rect 19156 11296 19208 11348
rect 20628 11339 20680 11348
rect 20628 11305 20637 11339
rect 20637 11305 20671 11339
rect 20671 11305 20680 11339
rect 20628 11296 20680 11305
rect 22008 11296 22060 11348
rect 22100 11339 22152 11348
rect 22100 11305 22109 11339
rect 22109 11305 22143 11339
rect 22143 11305 22152 11339
rect 22100 11296 22152 11305
rect 23756 11296 23808 11348
rect 24032 11339 24084 11348
rect 24032 11305 24041 11339
rect 24041 11305 24075 11339
rect 24075 11305 24084 11339
rect 24032 11296 24084 11305
rect 26240 11296 26292 11348
rect 3056 11271 3108 11280
rect 3056 11237 3065 11271
rect 3065 11237 3099 11271
rect 3099 11237 3108 11271
rect 3056 11228 3108 11237
rect 3608 11228 3660 11280
rect 8668 11271 8720 11280
rect 8668 11237 8677 11271
rect 8677 11237 8711 11271
rect 8711 11237 8720 11271
rect 8668 11228 8720 11237
rect 11336 11228 11388 11280
rect 12164 11271 12216 11280
rect 12164 11237 12173 11271
rect 12173 11237 12207 11271
rect 12207 11237 12216 11271
rect 12164 11228 12216 11237
rect 1952 11160 2004 11212
rect 4804 11160 4856 11212
rect 5080 11203 5132 11212
rect 5080 11169 5089 11203
rect 5089 11169 5123 11203
rect 5123 11169 5132 11203
rect 5080 11160 5132 11169
rect 1584 11092 1636 11144
rect 4160 11135 4212 11144
rect 4160 11101 4169 11135
rect 4169 11101 4203 11135
rect 4203 11101 4212 11135
rect 4160 11092 4212 11101
rect 4620 11135 4672 11144
rect 4620 11101 4629 11135
rect 4629 11101 4663 11135
rect 4663 11101 4672 11135
rect 4620 11092 4672 11101
rect 3424 11024 3476 11076
rect 3976 11024 4028 11076
rect 5448 11160 5500 11212
rect 6736 11203 6788 11212
rect 6736 11169 6745 11203
rect 6745 11169 6779 11203
rect 6779 11169 6788 11203
rect 6736 11160 6788 11169
rect 6920 11160 6972 11212
rect 8208 11203 8260 11212
rect 8208 11169 8217 11203
rect 8217 11169 8251 11203
rect 8251 11169 8260 11203
rect 8208 11160 8260 11169
rect 10324 11160 10376 11212
rect 11060 11203 11112 11212
rect 11060 11169 11069 11203
rect 11069 11169 11103 11203
rect 11103 11169 11112 11203
rect 11060 11160 11112 11169
rect 11796 11203 11848 11212
rect 11796 11169 11805 11203
rect 11805 11169 11839 11203
rect 11839 11169 11848 11203
rect 11796 11160 11848 11169
rect 13636 11203 13688 11212
rect 13636 11169 13645 11203
rect 13645 11169 13679 11203
rect 13679 11169 13688 11203
rect 13636 11160 13688 11169
rect 13820 11160 13872 11212
rect 15108 11160 15160 11212
rect 15844 11160 15896 11212
rect 16028 11203 16080 11212
rect 16028 11169 16037 11203
rect 16037 11169 16071 11203
rect 16071 11169 16080 11203
rect 16028 11160 16080 11169
rect 16120 11160 16172 11212
rect 17500 11271 17552 11280
rect 17500 11237 17509 11271
rect 17509 11237 17543 11271
rect 17543 11237 17552 11271
rect 17500 11228 17552 11237
rect 19432 11228 19484 11280
rect 20536 11228 20588 11280
rect 25228 11271 25280 11280
rect 25228 11237 25237 11271
rect 25237 11237 25271 11271
rect 25271 11237 25280 11271
rect 25228 11228 25280 11237
rect 6276 11092 6328 11144
rect 7932 11135 7984 11144
rect 3700 10956 3752 11008
rect 4712 10956 4764 11008
rect 6460 11024 6512 11076
rect 5632 10956 5684 11008
rect 6552 10956 6604 11008
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 8116 11135 8168 11144
rect 8116 11101 8125 11135
rect 8125 11101 8159 11135
rect 8159 11101 8168 11135
rect 8116 11092 8168 11101
rect 10784 11135 10836 11144
rect 10784 11101 10793 11135
rect 10793 11101 10827 11135
rect 10827 11101 10836 11135
rect 10784 11092 10836 11101
rect 13176 11135 13228 11144
rect 13176 11101 13185 11135
rect 13185 11101 13219 11135
rect 13219 11101 13228 11135
rect 13176 11092 13228 11101
rect 17408 11092 17460 11144
rect 19248 11160 19300 11212
rect 24124 11160 24176 11212
rect 24860 11203 24912 11212
rect 24860 11169 24869 11203
rect 24869 11169 24903 11203
rect 24903 11169 24912 11203
rect 24860 11160 24912 11169
rect 26240 11160 26292 11212
rect 27804 11160 27856 11212
rect 28540 11203 28592 11212
rect 28540 11169 28549 11203
rect 28549 11169 28583 11203
rect 28583 11169 28592 11203
rect 28540 11160 28592 11169
rect 30656 11203 30708 11212
rect 30656 11169 30665 11203
rect 30665 11169 30699 11203
rect 30699 11169 30708 11203
rect 30656 11160 30708 11169
rect 30748 11203 30800 11212
rect 30748 11169 30757 11203
rect 30757 11169 30791 11203
rect 30791 11169 30800 11203
rect 31024 11203 31076 11212
rect 30748 11160 30800 11169
rect 31024 11169 31033 11203
rect 31033 11169 31067 11203
rect 31067 11169 31076 11203
rect 31024 11160 31076 11169
rect 31484 11228 31536 11280
rect 23756 11092 23808 11144
rect 27344 11092 27396 11144
rect 27620 11092 27672 11144
rect 29920 11092 29972 11144
rect 13084 11024 13136 11076
rect 26976 11024 27028 11076
rect 8300 10956 8352 11008
rect 9496 10956 9548 11008
rect 10140 10956 10192 11008
rect 29000 11024 29052 11076
rect 27712 10956 27764 11008
rect 35348 10956 35400 11008
rect 35808 10999 35860 11008
rect 35808 10965 35817 10999
rect 35817 10965 35851 10999
rect 35851 10965 35860 10999
rect 35808 10956 35860 10965
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 3700 10795 3752 10804
rect 3700 10761 3709 10795
rect 3709 10761 3743 10795
rect 3743 10761 3752 10795
rect 3700 10752 3752 10761
rect 4804 10752 4856 10804
rect 8208 10795 8260 10804
rect 8208 10761 8217 10795
rect 8217 10761 8251 10795
rect 8251 10761 8260 10795
rect 8208 10752 8260 10761
rect 8484 10795 8536 10804
rect 8484 10761 8493 10795
rect 8493 10761 8527 10795
rect 8527 10761 8536 10795
rect 8484 10752 8536 10761
rect 10324 10752 10376 10804
rect 13176 10795 13228 10804
rect 4620 10684 4672 10736
rect 9680 10684 9732 10736
rect 13176 10761 13185 10795
rect 13185 10761 13219 10795
rect 13219 10761 13228 10795
rect 13912 10795 13964 10804
rect 13176 10752 13228 10761
rect 13912 10761 13921 10795
rect 13921 10761 13955 10795
rect 13955 10761 13964 10795
rect 13912 10752 13964 10761
rect 14648 10795 14700 10804
rect 14648 10761 14657 10795
rect 14657 10761 14691 10795
rect 14691 10761 14700 10795
rect 14648 10752 14700 10761
rect 15108 10752 15160 10804
rect 16028 10752 16080 10804
rect 16120 10795 16172 10804
rect 16120 10761 16129 10795
rect 16129 10761 16163 10795
rect 16163 10761 16172 10795
rect 16120 10752 16172 10761
rect 19340 10795 19392 10804
rect 19340 10761 19349 10795
rect 19349 10761 19383 10795
rect 19383 10761 19392 10795
rect 19340 10752 19392 10761
rect 20260 10752 20312 10804
rect 24124 10752 24176 10804
rect 25320 10795 25372 10804
rect 25320 10761 25329 10795
rect 25329 10761 25363 10795
rect 25363 10761 25372 10795
rect 25320 10752 25372 10761
rect 12532 10684 12584 10736
rect 12716 10684 12768 10736
rect 13636 10684 13688 10736
rect 13820 10684 13872 10736
rect 16672 10727 16724 10736
rect 16672 10693 16681 10727
rect 16681 10693 16715 10727
rect 16715 10693 16724 10727
rect 16672 10684 16724 10693
rect 15384 10616 15436 10668
rect 4712 10548 4764 10600
rect 6736 10548 6788 10600
rect 8668 10591 8720 10600
rect 8668 10557 8677 10591
rect 8677 10557 8711 10591
rect 8711 10557 8720 10591
rect 8668 10548 8720 10557
rect 8760 10591 8812 10600
rect 8760 10557 8769 10591
rect 8769 10557 8803 10591
rect 8803 10557 8812 10591
rect 8944 10591 8996 10600
rect 8760 10548 8812 10557
rect 8944 10557 8953 10591
rect 8953 10557 8987 10591
rect 8987 10557 8996 10591
rect 8944 10548 8996 10557
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 9496 10591 9548 10600
rect 9496 10557 9505 10591
rect 9505 10557 9539 10591
rect 9539 10557 9548 10591
rect 9496 10548 9548 10557
rect 12808 10548 12860 10600
rect 14464 10591 14516 10600
rect 14464 10557 14473 10591
rect 14473 10557 14507 10591
rect 14507 10557 14516 10591
rect 14464 10548 14516 10557
rect 15936 10548 15988 10600
rect 18420 10591 18472 10600
rect 18420 10557 18429 10591
rect 18429 10557 18463 10591
rect 18463 10557 18472 10591
rect 18420 10548 18472 10557
rect 24124 10591 24176 10600
rect 24124 10557 24133 10591
rect 24133 10557 24167 10591
rect 24167 10557 24176 10591
rect 24124 10548 24176 10557
rect 24860 10548 24912 10600
rect 25872 10752 25924 10804
rect 27712 10752 27764 10804
rect 28540 10752 28592 10804
rect 29000 10752 29052 10804
rect 30196 10752 30248 10804
rect 31024 10752 31076 10804
rect 30380 10684 30432 10736
rect 30748 10659 30800 10668
rect 30748 10625 30757 10659
rect 30757 10625 30791 10659
rect 30791 10625 30800 10659
rect 30748 10616 30800 10625
rect 26976 10591 27028 10600
rect 6828 10480 6880 10532
rect 11796 10480 11848 10532
rect 18328 10523 18380 10532
rect 18328 10489 18337 10523
rect 18337 10489 18371 10523
rect 18371 10489 18380 10523
rect 18328 10480 18380 10489
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 1952 10455 2004 10464
rect 1952 10421 1961 10455
rect 1961 10421 1995 10455
rect 1995 10421 2004 10455
rect 1952 10412 2004 10421
rect 3976 10412 4028 10464
rect 4620 10455 4672 10464
rect 4620 10421 4629 10455
rect 4629 10421 4663 10455
rect 4663 10421 4672 10455
rect 4620 10412 4672 10421
rect 6276 10412 6328 10464
rect 6552 10455 6604 10464
rect 6552 10421 6561 10455
rect 6561 10421 6595 10455
rect 6595 10421 6604 10455
rect 6552 10412 6604 10421
rect 8116 10412 8168 10464
rect 11336 10455 11388 10464
rect 11336 10421 11345 10455
rect 11345 10421 11379 10455
rect 11379 10421 11388 10455
rect 11336 10412 11388 10421
rect 11520 10412 11572 10464
rect 15108 10412 15160 10464
rect 17408 10455 17460 10464
rect 17408 10421 17417 10455
rect 17417 10421 17451 10455
rect 17451 10421 17460 10455
rect 17408 10412 17460 10421
rect 26148 10455 26200 10464
rect 26148 10421 26157 10455
rect 26157 10421 26191 10455
rect 26191 10421 26200 10455
rect 26148 10412 26200 10421
rect 26976 10557 26985 10591
rect 26985 10557 27019 10591
rect 27019 10557 27028 10591
rect 26976 10548 27028 10557
rect 30656 10548 30708 10600
rect 31392 10480 31444 10532
rect 27344 10412 27396 10464
rect 30656 10412 30708 10464
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 5080 10208 5132 10260
rect 6828 10251 6880 10260
rect 6828 10217 6837 10251
rect 6837 10217 6871 10251
rect 6871 10217 6880 10251
rect 6828 10208 6880 10217
rect 8668 10208 8720 10260
rect 9404 10208 9456 10260
rect 11704 10208 11756 10260
rect 12440 10251 12492 10260
rect 12440 10217 12449 10251
rect 12449 10217 12483 10251
rect 12483 10217 12492 10251
rect 12440 10208 12492 10217
rect 13728 10208 13780 10260
rect 16028 10208 16080 10260
rect 16580 10251 16632 10260
rect 16580 10217 16589 10251
rect 16589 10217 16623 10251
rect 16623 10217 16632 10251
rect 16580 10208 16632 10217
rect 17868 10208 17920 10260
rect 19156 10251 19208 10260
rect 19156 10217 19165 10251
rect 19165 10217 19199 10251
rect 19199 10217 19208 10251
rect 19156 10208 19208 10217
rect 20260 10208 20312 10260
rect 20352 10208 20404 10260
rect 25596 10251 25648 10260
rect 4712 10183 4764 10192
rect 4712 10149 4721 10183
rect 4721 10149 4755 10183
rect 4755 10149 4764 10183
rect 4712 10140 4764 10149
rect 13268 10140 13320 10192
rect 14372 10140 14424 10192
rect 15844 10183 15896 10192
rect 15844 10149 15853 10183
rect 15853 10149 15887 10183
rect 15887 10149 15896 10183
rect 15844 10140 15896 10149
rect 15936 10140 15988 10192
rect 16304 10140 16356 10192
rect 19892 10140 19944 10192
rect 5540 10115 5592 10124
rect 5540 10081 5549 10115
rect 5549 10081 5583 10115
rect 5583 10081 5592 10115
rect 5540 10072 5592 10081
rect 7104 10072 7156 10124
rect 4620 10004 4672 10056
rect 5448 10004 5500 10056
rect 6552 10004 6604 10056
rect 8208 10004 8260 10056
rect 8760 10072 8812 10124
rect 9496 10072 9548 10124
rect 11428 10115 11480 10124
rect 11428 10081 11437 10115
rect 11437 10081 11471 10115
rect 11471 10081 11480 10115
rect 11428 10072 11480 10081
rect 13452 10115 13504 10124
rect 13452 10081 13461 10115
rect 13461 10081 13495 10115
rect 13495 10081 13504 10115
rect 13452 10072 13504 10081
rect 14464 10072 14516 10124
rect 15292 10115 15344 10124
rect 15292 10081 15301 10115
rect 15301 10081 15335 10115
rect 15335 10081 15344 10115
rect 15292 10072 15344 10081
rect 18328 10072 18380 10124
rect 19064 10072 19116 10124
rect 21916 10115 21968 10124
rect 21916 10081 21925 10115
rect 21925 10081 21959 10115
rect 21959 10081 21968 10115
rect 21916 10072 21968 10081
rect 9588 10004 9640 10056
rect 9680 10004 9732 10056
rect 11796 10004 11848 10056
rect 12532 10004 12584 10056
rect 13820 10004 13872 10056
rect 25596 10217 25605 10251
rect 25605 10217 25639 10251
rect 25639 10217 25648 10251
rect 25596 10208 25648 10217
rect 27068 10208 27120 10260
rect 28080 10208 28132 10260
rect 30196 10251 30248 10260
rect 30196 10217 30205 10251
rect 30205 10217 30239 10251
rect 30239 10217 30248 10251
rect 30196 10208 30248 10217
rect 30748 10208 30800 10260
rect 36084 10208 36136 10260
rect 24124 10140 24176 10192
rect 22376 10072 22428 10124
rect 24400 10072 24452 10124
rect 25504 10072 25556 10124
rect 26148 10072 26200 10124
rect 26792 10115 26844 10124
rect 26792 10081 26801 10115
rect 26801 10081 26835 10115
rect 26835 10081 26844 10115
rect 26792 10072 26844 10081
rect 27620 10072 27672 10124
rect 30656 10072 30708 10124
rect 35256 10072 35308 10124
rect 22652 10004 22704 10056
rect 35348 10004 35400 10056
rect 8116 9936 8168 9988
rect 8760 9979 8812 9988
rect 8760 9945 8769 9979
rect 8769 9945 8803 9979
rect 8803 9945 8812 9979
rect 8760 9936 8812 9945
rect 17132 9979 17184 9988
rect 17132 9945 17141 9979
rect 17141 9945 17175 9979
rect 17175 9945 17184 9979
rect 17132 9936 17184 9945
rect 8300 9868 8352 9920
rect 9496 9911 9548 9920
rect 9496 9877 9505 9911
rect 9505 9877 9539 9911
rect 9539 9877 9548 9911
rect 9496 9868 9548 9877
rect 14280 9911 14332 9920
rect 14280 9877 14289 9911
rect 14289 9877 14323 9911
rect 14323 9877 14332 9911
rect 14280 9868 14332 9877
rect 15660 9868 15712 9920
rect 18144 9911 18196 9920
rect 18144 9877 18153 9911
rect 18153 9877 18187 9911
rect 18187 9877 18196 9911
rect 18144 9868 18196 9877
rect 18604 9868 18656 9920
rect 19524 9868 19576 9920
rect 27344 9911 27396 9920
rect 27344 9877 27353 9911
rect 27353 9877 27387 9911
rect 27387 9877 27396 9911
rect 27344 9868 27396 9877
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 2596 9664 2648 9716
rect 3884 9664 3936 9716
rect 11428 9664 11480 9716
rect 12532 9664 12584 9716
rect 13452 9707 13504 9716
rect 13452 9673 13461 9707
rect 13461 9673 13495 9707
rect 13495 9673 13504 9707
rect 13452 9664 13504 9673
rect 15292 9664 15344 9716
rect 18328 9707 18380 9716
rect 5540 9596 5592 9648
rect 1952 9503 2004 9512
rect 1952 9469 1961 9503
rect 1961 9469 1995 9503
rect 1995 9469 2004 9503
rect 1952 9460 2004 9469
rect 2872 9528 2924 9580
rect 6736 9528 6788 9580
rect 12072 9596 12124 9648
rect 8116 9528 8168 9580
rect 8208 9571 8260 9580
rect 8208 9537 8217 9571
rect 8217 9537 8251 9571
rect 8251 9537 8260 9571
rect 14372 9596 14424 9648
rect 18328 9673 18337 9707
rect 18337 9673 18371 9707
rect 18371 9673 18380 9707
rect 18328 9664 18380 9673
rect 19064 9664 19116 9716
rect 20904 9664 20956 9716
rect 21640 9664 21692 9716
rect 21916 9664 21968 9716
rect 26792 9707 26844 9716
rect 26792 9673 26801 9707
rect 26801 9673 26835 9707
rect 26835 9673 26844 9707
rect 26792 9664 26844 9673
rect 27620 9664 27672 9716
rect 8208 9528 8260 9537
rect 2320 9460 2372 9512
rect 5448 9460 5500 9512
rect 7104 9460 7156 9512
rect 7932 9503 7984 9512
rect 7932 9469 7941 9503
rect 7941 9469 7975 9503
rect 7975 9469 7984 9503
rect 7932 9460 7984 9469
rect 8300 9503 8352 9512
rect 8300 9469 8309 9503
rect 8309 9469 8343 9503
rect 8343 9469 8352 9503
rect 8300 9460 8352 9469
rect 8852 9503 8904 9512
rect 8852 9469 8861 9503
rect 8861 9469 8895 9503
rect 8895 9469 8904 9503
rect 8852 9460 8904 9469
rect 9496 9460 9548 9512
rect 7288 9435 7340 9444
rect 7288 9401 7297 9435
rect 7297 9401 7331 9435
rect 7331 9401 7340 9435
rect 7288 9392 7340 9401
rect 14096 9460 14148 9512
rect 19892 9596 19944 9648
rect 25780 9639 25832 9648
rect 25780 9605 25789 9639
rect 25789 9605 25823 9639
rect 25823 9605 25832 9639
rect 25780 9596 25832 9605
rect 35256 9639 35308 9648
rect 35256 9605 35265 9639
rect 35265 9605 35299 9639
rect 35299 9605 35308 9639
rect 35256 9596 35308 9605
rect 18604 9528 18656 9580
rect 12992 9367 13044 9376
rect 12992 9333 13001 9367
rect 13001 9333 13035 9367
rect 13035 9333 13044 9367
rect 14280 9392 14332 9444
rect 15016 9435 15068 9444
rect 15016 9401 15025 9435
rect 15025 9401 15059 9435
rect 15059 9401 15068 9435
rect 15016 9392 15068 9401
rect 16120 9367 16172 9376
rect 12992 9324 13044 9333
rect 16120 9333 16129 9367
rect 16129 9333 16163 9367
rect 16163 9333 16172 9367
rect 16120 9324 16172 9333
rect 19064 9392 19116 9444
rect 19524 9460 19576 9512
rect 35072 9528 35124 9580
rect 35348 9528 35400 9580
rect 24400 9503 24452 9512
rect 21916 9392 21968 9444
rect 24400 9469 24409 9503
rect 24409 9469 24443 9503
rect 24443 9469 24452 9503
rect 24400 9460 24452 9469
rect 24676 9503 24728 9512
rect 24676 9469 24685 9503
rect 24685 9469 24719 9503
rect 24719 9469 24728 9503
rect 24676 9460 24728 9469
rect 18236 9324 18288 9376
rect 19248 9367 19300 9376
rect 19248 9333 19257 9367
rect 19257 9333 19291 9367
rect 19291 9333 19300 9367
rect 19248 9324 19300 9333
rect 19984 9324 20036 9376
rect 22284 9367 22336 9376
rect 22284 9333 22293 9367
rect 22293 9333 22327 9367
rect 22327 9333 22336 9367
rect 22284 9324 22336 9333
rect 22652 9367 22704 9376
rect 22652 9333 22661 9367
rect 22661 9333 22695 9367
rect 22695 9333 22704 9367
rect 22652 9324 22704 9333
rect 23296 9367 23348 9376
rect 23296 9333 23305 9367
rect 23305 9333 23339 9367
rect 23339 9333 23348 9367
rect 23296 9324 23348 9333
rect 23480 9324 23532 9376
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 1952 9163 2004 9172
rect 1952 9129 1961 9163
rect 1961 9129 1995 9163
rect 1995 9129 2004 9163
rect 1952 9120 2004 9129
rect 8300 9120 8352 9172
rect 9680 9120 9732 9172
rect 9956 9120 10008 9172
rect 11152 9120 11204 9172
rect 12624 9163 12676 9172
rect 12624 9129 12633 9163
rect 12633 9129 12667 9163
rect 12667 9129 12676 9163
rect 13912 9163 13964 9172
rect 12624 9120 12676 9129
rect 12992 9052 13044 9104
rect 13912 9129 13921 9163
rect 13921 9129 13955 9163
rect 13955 9129 13964 9163
rect 13912 9120 13964 9129
rect 24400 9120 24452 9172
rect 25964 9163 26016 9172
rect 25964 9129 25973 9163
rect 25973 9129 26007 9163
rect 26007 9129 26016 9163
rect 25964 9120 26016 9129
rect 15384 9052 15436 9104
rect 19984 9095 20036 9104
rect 5540 8984 5592 9036
rect 6092 9027 6144 9036
rect 6092 8993 6101 9027
rect 6101 8993 6135 9027
rect 6135 8993 6144 9027
rect 6092 8984 6144 8993
rect 7196 8984 7248 9036
rect 8852 8984 8904 9036
rect 9864 9027 9916 9036
rect 9864 8993 9873 9027
rect 9873 8993 9907 9027
rect 9907 8993 9916 9027
rect 9864 8984 9916 8993
rect 10876 9027 10928 9036
rect 10876 8993 10885 9027
rect 10885 8993 10919 9027
rect 10919 8993 10928 9027
rect 10876 8984 10928 8993
rect 11612 9027 11664 9036
rect 11612 8993 11621 9027
rect 11621 8993 11655 9027
rect 11655 8993 11664 9027
rect 11612 8984 11664 8993
rect 11796 9027 11848 9036
rect 11796 8993 11805 9027
rect 11805 8993 11839 9027
rect 11839 8993 11848 9027
rect 11796 8984 11848 8993
rect 13176 9027 13228 9036
rect 13176 8993 13185 9027
rect 13185 8993 13219 9027
rect 13219 8993 13228 9027
rect 13176 8984 13228 8993
rect 13728 8984 13780 9036
rect 14832 8984 14884 9036
rect 15476 9027 15528 9036
rect 15476 8993 15485 9027
rect 15485 8993 15519 9027
rect 15519 8993 15528 9027
rect 15476 8984 15528 8993
rect 15660 8984 15712 9036
rect 19984 9061 19993 9095
rect 19993 9061 20027 9095
rect 20027 9061 20036 9095
rect 19984 9052 20036 9061
rect 25504 9095 25556 9104
rect 25504 9061 25513 9095
rect 25513 9061 25547 9095
rect 25547 9061 25556 9095
rect 25504 9052 25556 9061
rect 18420 8984 18472 9036
rect 18604 9027 18656 9036
rect 18604 8993 18613 9027
rect 18613 8993 18647 9027
rect 18647 8993 18656 9027
rect 18604 8984 18656 8993
rect 26148 9027 26200 9036
rect 26148 8993 26157 9027
rect 26157 8993 26191 9027
rect 26191 8993 26200 9027
rect 26148 8984 26200 8993
rect 7104 8959 7156 8968
rect 7104 8925 7113 8959
rect 7113 8925 7147 8959
rect 7147 8925 7156 8959
rect 7104 8916 7156 8925
rect 13084 8959 13136 8968
rect 13084 8925 13093 8959
rect 13093 8925 13127 8959
rect 13127 8925 13136 8959
rect 13084 8916 13136 8925
rect 13360 8916 13412 8968
rect 15200 8916 15252 8968
rect 6276 8891 6328 8900
rect 6276 8857 6285 8891
rect 6285 8857 6319 8891
rect 6319 8857 6328 8891
rect 6276 8848 6328 8857
rect 9956 8780 10008 8832
rect 12348 8780 12400 8832
rect 13360 8823 13412 8832
rect 13360 8789 13369 8823
rect 13369 8789 13403 8823
rect 13403 8789 13412 8823
rect 13360 8780 13412 8789
rect 14372 8823 14424 8832
rect 14372 8789 14381 8823
rect 14381 8789 14415 8823
rect 14415 8789 14424 8823
rect 14372 8780 14424 8789
rect 15200 8780 15252 8832
rect 16488 8823 16540 8832
rect 16488 8789 16497 8823
rect 16497 8789 16531 8823
rect 16531 8789 16540 8823
rect 16488 8780 16540 8789
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 6092 8619 6144 8628
rect 6092 8585 6101 8619
rect 6101 8585 6135 8619
rect 6135 8585 6144 8619
rect 6092 8576 6144 8585
rect 7104 8576 7156 8628
rect 11612 8619 11664 8628
rect 11612 8585 11621 8619
rect 11621 8585 11655 8619
rect 11655 8585 11664 8619
rect 11612 8576 11664 8585
rect 12900 8576 12952 8628
rect 13176 8619 13228 8628
rect 13176 8585 13185 8619
rect 13185 8585 13219 8619
rect 13219 8585 13228 8619
rect 13176 8576 13228 8585
rect 14280 8576 14332 8628
rect 15384 8619 15436 8628
rect 15384 8585 15393 8619
rect 15393 8585 15427 8619
rect 15427 8585 15436 8619
rect 15384 8576 15436 8585
rect 15476 8576 15528 8628
rect 18236 8619 18288 8628
rect 18236 8585 18245 8619
rect 18245 8585 18279 8619
rect 18279 8585 18288 8619
rect 18236 8576 18288 8585
rect 18328 8576 18380 8628
rect 18604 8576 18656 8628
rect 26148 8576 26200 8628
rect 7196 8551 7248 8560
rect 7196 8517 7205 8551
rect 7205 8517 7239 8551
rect 7239 8517 7248 8551
rect 7196 8508 7248 8517
rect 11796 8508 11848 8560
rect 7932 8440 7984 8492
rect 9680 8483 9732 8492
rect 9680 8449 9689 8483
rect 9689 8449 9723 8483
rect 9723 8449 9732 8483
rect 9680 8440 9732 8449
rect 10876 8440 10928 8492
rect 12900 8440 12952 8492
rect 9588 8415 9640 8424
rect 9588 8381 9597 8415
rect 9597 8381 9631 8415
rect 9631 8381 9640 8415
rect 9588 8372 9640 8381
rect 9956 8415 10008 8424
rect 9956 8381 9965 8415
rect 9965 8381 9999 8415
rect 9999 8381 10008 8415
rect 9956 8372 10008 8381
rect 10140 8415 10192 8424
rect 10140 8381 10149 8415
rect 10149 8381 10183 8415
rect 10183 8381 10192 8415
rect 10140 8372 10192 8381
rect 13728 8415 13780 8424
rect 13728 8381 13737 8415
rect 13737 8381 13771 8415
rect 13771 8381 13780 8415
rect 13728 8372 13780 8381
rect 1492 8304 1544 8356
rect 11060 8304 11112 8356
rect 13268 8347 13320 8356
rect 13268 8313 13277 8347
rect 13277 8313 13311 8347
rect 13311 8313 13320 8347
rect 13268 8304 13320 8313
rect 13636 8304 13688 8356
rect 14832 8440 14884 8492
rect 15752 8440 15804 8492
rect 16304 8440 16356 8492
rect 16948 8508 17000 8560
rect 18420 8508 18472 8560
rect 16856 8483 16908 8492
rect 16856 8449 16865 8483
rect 16865 8449 16899 8483
rect 16899 8449 16908 8483
rect 16856 8440 16908 8449
rect 14648 8347 14700 8356
rect 14648 8313 14657 8347
rect 14657 8313 14691 8347
rect 14691 8313 14700 8347
rect 14648 8304 14700 8313
rect 16672 8372 16724 8424
rect 18328 8372 18380 8424
rect 9956 8236 10008 8288
rect 13084 8236 13136 8288
rect 16028 8236 16080 8288
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 9036 8075 9088 8084
rect 9036 8041 9045 8075
rect 9045 8041 9079 8075
rect 9079 8041 9088 8075
rect 9036 8032 9088 8041
rect 11060 8075 11112 8084
rect 11060 8041 11069 8075
rect 11069 8041 11103 8075
rect 11103 8041 11112 8075
rect 11060 8032 11112 8041
rect 13360 7964 13412 8016
rect 12624 7939 12676 7948
rect 12624 7905 12633 7939
rect 12633 7905 12667 7939
rect 12667 7905 12676 7939
rect 12624 7896 12676 7905
rect 12716 7896 12768 7948
rect 13636 8032 13688 8084
rect 13820 8075 13872 8084
rect 13820 8041 13829 8075
rect 13829 8041 13863 8075
rect 13863 8041 13872 8075
rect 13820 8032 13872 8041
rect 15108 8075 15160 8084
rect 15108 8041 15117 8075
rect 15117 8041 15151 8075
rect 15151 8041 15160 8075
rect 15108 8032 15160 8041
rect 16672 8075 16724 8084
rect 16672 8041 16681 8075
rect 16681 8041 16715 8075
rect 16715 8041 16724 8075
rect 16672 8032 16724 8041
rect 20352 8032 20404 8084
rect 19708 7964 19760 8016
rect 21088 7964 21140 8016
rect 9680 7871 9732 7880
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 9680 7828 9732 7837
rect 9864 7828 9916 7880
rect 11336 7828 11388 7880
rect 12808 7828 12860 7880
rect 15200 7896 15252 7948
rect 16304 7896 16356 7948
rect 16580 7896 16632 7948
rect 17868 7896 17920 7948
rect 21180 7896 21232 7948
rect 15016 7828 15068 7880
rect 18420 7828 18472 7880
rect 20352 7828 20404 7880
rect 21548 7939 21600 7948
rect 21548 7905 21557 7939
rect 21557 7905 21591 7939
rect 21591 7905 21600 7939
rect 21916 7939 21968 7948
rect 21548 7896 21600 7905
rect 21916 7905 21925 7939
rect 21925 7905 21959 7939
rect 21959 7905 21968 7939
rect 21916 7896 21968 7905
rect 23112 7939 23164 7948
rect 23112 7905 23121 7939
rect 23121 7905 23155 7939
rect 23155 7905 23164 7939
rect 23112 7896 23164 7905
rect 19340 7735 19392 7744
rect 19340 7701 19349 7735
rect 19349 7701 19383 7735
rect 19383 7701 19392 7735
rect 19340 7692 19392 7701
rect 21180 7735 21232 7744
rect 21180 7701 21189 7735
rect 21189 7701 21223 7735
rect 21223 7701 21232 7735
rect 21180 7692 21232 7701
rect 23480 7692 23532 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 8484 7531 8536 7540
rect 8484 7497 8493 7531
rect 8493 7497 8527 7531
rect 8527 7497 8536 7531
rect 8484 7488 8536 7497
rect 9864 7488 9916 7540
rect 10048 7488 10100 7540
rect 10876 7395 10928 7404
rect 10876 7361 10885 7395
rect 10885 7361 10919 7395
rect 10919 7361 10928 7395
rect 10876 7352 10928 7361
rect 12624 7488 12676 7540
rect 15016 7531 15068 7540
rect 15016 7497 15025 7531
rect 15025 7497 15059 7531
rect 15059 7497 15068 7531
rect 15016 7488 15068 7497
rect 16304 7531 16356 7540
rect 16304 7497 16313 7531
rect 16313 7497 16347 7531
rect 16347 7497 16356 7531
rect 16304 7488 16356 7497
rect 17868 7531 17920 7540
rect 17868 7497 17877 7531
rect 17877 7497 17911 7531
rect 17911 7497 17920 7531
rect 17868 7488 17920 7497
rect 19432 7488 19484 7540
rect 21548 7488 21600 7540
rect 21916 7488 21968 7540
rect 23112 7488 23164 7540
rect 11152 7420 11204 7472
rect 12716 7420 12768 7472
rect 16028 7463 16080 7472
rect 16028 7429 16037 7463
rect 16037 7429 16071 7463
rect 16071 7429 16080 7463
rect 16028 7420 16080 7429
rect 11244 7395 11296 7404
rect 11244 7361 11253 7395
rect 11253 7361 11287 7395
rect 11287 7361 11296 7395
rect 11244 7352 11296 7361
rect 13268 7352 13320 7404
rect 20352 7352 20404 7404
rect 8484 7284 8536 7336
rect 10968 7327 11020 7336
rect 10968 7293 10977 7327
rect 10977 7293 11011 7327
rect 11011 7293 11020 7327
rect 10968 7284 11020 7293
rect 11336 7327 11388 7336
rect 11336 7293 11345 7327
rect 11345 7293 11379 7327
rect 11379 7293 11388 7327
rect 11336 7284 11388 7293
rect 12532 7284 12584 7336
rect 18420 7284 18472 7336
rect 20260 7284 20312 7336
rect 8668 7191 8720 7200
rect 8668 7157 8677 7191
rect 8677 7157 8711 7191
rect 8711 7157 8720 7191
rect 8668 7148 8720 7157
rect 10232 7148 10284 7200
rect 10968 7148 11020 7200
rect 12808 7216 12860 7268
rect 13636 7148 13688 7200
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 10876 6944 10928 6996
rect 12716 6944 12768 6996
rect 13268 6944 13320 6996
rect 20352 6944 20404 6996
rect 21088 6987 21140 6996
rect 21088 6953 21097 6987
rect 21097 6953 21131 6987
rect 21131 6953 21140 6987
rect 21088 6944 21140 6953
rect 21916 6944 21968 6996
rect 9680 6808 9732 6860
rect 11060 6808 11112 6860
rect 10968 6740 11020 6792
rect 13636 6808 13688 6860
rect 17868 6876 17920 6928
rect 18880 6876 18932 6928
rect 16856 6808 16908 6860
rect 16948 6808 17000 6860
rect 17224 6851 17276 6860
rect 17224 6817 17233 6851
rect 17233 6817 17267 6851
rect 17267 6817 17276 6851
rect 17224 6808 17276 6817
rect 19248 6808 19300 6860
rect 27160 6808 27212 6860
rect 28724 6851 28776 6860
rect 28724 6817 28733 6851
rect 28733 6817 28767 6851
rect 28767 6817 28776 6851
rect 28724 6808 28776 6817
rect 12440 6740 12492 6792
rect 13820 6783 13872 6792
rect 13820 6749 13829 6783
rect 13829 6749 13863 6783
rect 13863 6749 13872 6783
rect 13820 6740 13872 6749
rect 14004 6783 14056 6792
rect 14004 6749 14013 6783
rect 14013 6749 14047 6783
rect 14047 6749 14056 6783
rect 14004 6740 14056 6749
rect 16120 6783 16172 6792
rect 16120 6749 16129 6783
rect 16129 6749 16163 6783
rect 16163 6749 16172 6783
rect 16120 6740 16172 6749
rect 16672 6783 16724 6792
rect 16672 6749 16681 6783
rect 16681 6749 16715 6783
rect 16715 6749 16724 6783
rect 16672 6740 16724 6749
rect 19064 6783 19116 6792
rect 19064 6749 19073 6783
rect 19073 6749 19107 6783
rect 19107 6749 19116 6783
rect 19064 6740 19116 6749
rect 12348 6672 12400 6724
rect 15108 6672 15160 6724
rect 18512 6672 18564 6724
rect 19892 6740 19944 6792
rect 22192 6783 22244 6792
rect 22192 6749 22201 6783
rect 22201 6749 22235 6783
rect 22235 6749 22244 6783
rect 22192 6740 22244 6749
rect 22468 6783 22520 6792
rect 22468 6749 22477 6783
rect 22477 6749 22511 6783
rect 22511 6749 22520 6783
rect 22468 6740 22520 6749
rect 23572 6783 23624 6792
rect 23572 6749 23581 6783
rect 23581 6749 23615 6783
rect 23615 6749 23624 6783
rect 23572 6740 23624 6749
rect 27252 6740 27304 6792
rect 12532 6647 12584 6656
rect 12532 6613 12541 6647
rect 12541 6613 12575 6647
rect 12575 6613 12584 6647
rect 12532 6604 12584 6613
rect 14556 6647 14608 6656
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14556 6604 14608 6613
rect 18788 6647 18840 6656
rect 18788 6613 18797 6647
rect 18797 6613 18831 6647
rect 18831 6613 18840 6647
rect 18788 6604 18840 6613
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 9680 6400 9732 6452
rect 8208 6332 8260 6384
rect 10968 6400 11020 6452
rect 12716 6400 12768 6452
rect 13636 6400 13688 6452
rect 13912 6443 13964 6452
rect 13912 6409 13921 6443
rect 13921 6409 13955 6443
rect 13955 6409 13964 6443
rect 13912 6400 13964 6409
rect 17224 6400 17276 6452
rect 19248 6400 19300 6452
rect 20352 6400 20404 6452
rect 22192 6400 22244 6452
rect 22652 6400 22704 6452
rect 27252 6400 27304 6452
rect 12532 6332 12584 6384
rect 15936 6332 15988 6384
rect 16672 6332 16724 6384
rect 18512 6375 18564 6384
rect 18512 6341 18521 6375
rect 18521 6341 18555 6375
rect 18555 6341 18564 6375
rect 18512 6332 18564 6341
rect 16856 6264 16908 6316
rect 8668 6196 8720 6248
rect 13820 6196 13872 6248
rect 14556 6239 14608 6248
rect 14556 6205 14565 6239
rect 14565 6205 14599 6239
rect 14599 6205 14608 6239
rect 14556 6196 14608 6205
rect 14740 6239 14792 6248
rect 14740 6205 14749 6239
rect 14749 6205 14783 6239
rect 14783 6205 14792 6239
rect 14740 6196 14792 6205
rect 15108 6239 15160 6248
rect 15108 6205 15117 6239
rect 15117 6205 15151 6239
rect 15151 6205 15160 6239
rect 15108 6196 15160 6205
rect 19156 6196 19208 6248
rect 19340 6239 19392 6248
rect 19340 6205 19349 6239
rect 19349 6205 19383 6239
rect 19383 6205 19392 6239
rect 19340 6196 19392 6205
rect 14004 6128 14056 6180
rect 22468 6128 22520 6180
rect 23020 6128 23072 6180
rect 14372 6103 14424 6112
rect 14372 6069 14381 6103
rect 14381 6069 14415 6103
rect 14415 6069 14424 6103
rect 14372 6060 14424 6069
rect 16948 6103 17000 6112
rect 16948 6069 16957 6103
rect 16957 6069 16991 6103
rect 16991 6069 17000 6103
rect 16948 6060 17000 6069
rect 27068 6103 27120 6112
rect 27068 6069 27077 6103
rect 27077 6069 27111 6103
rect 27111 6069 27120 6103
rect 27068 6060 27120 6069
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 14740 5899 14792 5908
rect 14740 5865 14749 5899
rect 14749 5865 14783 5899
rect 14783 5865 14792 5899
rect 14740 5856 14792 5865
rect 16948 5856 17000 5908
rect 18880 5899 18932 5908
rect 18880 5865 18889 5899
rect 18889 5865 18923 5899
rect 18923 5865 18932 5899
rect 18880 5856 18932 5865
rect 19064 5788 19116 5840
rect 12348 5720 12400 5772
rect 12808 5720 12860 5772
rect 15936 5763 15988 5772
rect 15936 5729 15945 5763
rect 15945 5729 15979 5763
rect 15979 5729 15988 5763
rect 15936 5720 15988 5729
rect 23480 5720 23532 5772
rect 23848 5720 23900 5772
rect 12532 5652 12584 5704
rect 16028 5652 16080 5704
rect 18144 5516 18196 5568
rect 19156 5516 19208 5568
rect 23480 5559 23532 5568
rect 23480 5525 23489 5559
rect 23489 5525 23523 5559
rect 23523 5525 23532 5559
rect 23480 5516 23532 5525
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 10508 5312 10560 5364
rect 12808 5355 12860 5364
rect 12808 5321 12817 5355
rect 12817 5321 12851 5355
rect 12851 5321 12860 5355
rect 12808 5312 12860 5321
rect 16028 5355 16080 5364
rect 16028 5321 16037 5355
rect 16037 5321 16071 5355
rect 16071 5321 16080 5355
rect 16028 5312 16080 5321
rect 23848 5355 23900 5364
rect 23848 5321 23857 5355
rect 23857 5321 23891 5355
rect 23891 5321 23900 5355
rect 23848 5312 23900 5321
rect 12532 5244 12584 5296
rect 15936 5244 15988 5296
rect 8300 5108 8352 5160
rect 8852 5151 8904 5160
rect 8852 5117 8861 5151
rect 8861 5117 8895 5151
rect 8895 5117 8904 5151
rect 8852 5108 8904 5117
rect 9220 5108 9272 5160
rect 23480 5108 23532 5160
rect 21640 5015 21692 5024
rect 21640 4981 21649 5015
rect 21649 4981 21683 5015
rect 21683 4981 21692 5015
rect 21640 4972 21692 4981
rect 25412 5015 25464 5024
rect 25412 4981 25421 5015
rect 25421 4981 25455 5015
rect 25455 4981 25464 5015
rect 25412 4972 25464 4981
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 8852 4811 8904 4820
rect 8852 4777 8861 4811
rect 8861 4777 8895 4811
rect 8895 4777 8904 4811
rect 8852 4768 8904 4777
rect 12164 4811 12216 4820
rect 12164 4777 12173 4811
rect 12173 4777 12207 4811
rect 12207 4777 12216 4811
rect 12164 4768 12216 4777
rect 13820 4768 13872 4820
rect 17316 4768 17368 4820
rect 33508 4811 33560 4820
rect 33508 4777 33517 4811
rect 33517 4777 33551 4811
rect 33551 4777 33560 4811
rect 33508 4768 33560 4777
rect 19432 4743 19484 4752
rect 19432 4709 19441 4743
rect 19441 4709 19475 4743
rect 19475 4709 19484 4743
rect 19432 4700 19484 4709
rect 28908 4700 28960 4752
rect 11336 4632 11388 4684
rect 12532 4632 12584 4684
rect 16028 4632 16080 4684
rect 18144 4632 18196 4684
rect 32680 4632 32732 4684
rect 11060 4607 11112 4616
rect 11060 4573 11069 4607
rect 11069 4573 11103 4607
rect 11103 4573 11112 4607
rect 11060 4564 11112 4573
rect 17960 4564 18012 4616
rect 26516 4607 26568 4616
rect 26516 4573 26525 4607
rect 26525 4573 26559 4607
rect 26559 4573 26568 4607
rect 26516 4564 26568 4573
rect 26792 4607 26844 4616
rect 26792 4573 26801 4607
rect 26801 4573 26835 4607
rect 26835 4573 26844 4607
rect 26792 4564 26844 4573
rect 32128 4607 32180 4616
rect 32128 4573 32137 4607
rect 32137 4573 32171 4607
rect 32171 4573 32180 4607
rect 32128 4564 32180 4573
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 9956 4267 10008 4276
rect 9956 4233 9965 4267
rect 9965 4233 9999 4267
rect 9999 4233 10008 4267
rect 9956 4224 10008 4233
rect 11336 4224 11388 4276
rect 18144 4224 18196 4276
rect 8300 4088 8352 4140
rect 17868 4063 17920 4072
rect 17868 4029 17877 4063
rect 17877 4029 17911 4063
rect 17911 4029 17920 4063
rect 17868 4020 17920 4029
rect 26792 4224 26844 4276
rect 20536 4088 20588 4140
rect 21272 4088 21324 4140
rect 26884 4131 26936 4140
rect 19156 4063 19208 4072
rect 19156 4029 19165 4063
rect 19165 4029 19199 4063
rect 19199 4029 19208 4063
rect 19156 4020 19208 4029
rect 25412 4063 25464 4072
rect 25412 4029 25421 4063
rect 25421 4029 25455 4063
rect 25455 4029 25464 4063
rect 25412 4020 25464 4029
rect 26884 4097 26893 4131
rect 26893 4097 26927 4131
rect 26927 4097 26936 4131
rect 26884 4088 26936 4097
rect 25780 4020 25832 4072
rect 7840 3884 7892 3936
rect 9680 3952 9732 4004
rect 10968 3952 11020 4004
rect 32680 3952 32732 4004
rect 32128 3884 32180 3936
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 8300 3680 8352 3732
rect 11520 3723 11572 3732
rect 11520 3689 11529 3723
rect 11529 3689 11563 3723
rect 11563 3689 11572 3723
rect 11520 3680 11572 3689
rect 19156 3723 19208 3732
rect 19156 3689 19165 3723
rect 19165 3689 19199 3723
rect 19199 3689 19208 3723
rect 19156 3680 19208 3689
rect 19984 3680 20036 3732
rect 24676 3723 24728 3732
rect 24676 3689 24685 3723
rect 24685 3689 24719 3723
rect 24719 3689 24728 3723
rect 24676 3680 24728 3689
rect 33140 3680 33192 3732
rect 17040 3612 17092 3664
rect 1768 3587 1820 3596
rect 1768 3553 1777 3587
rect 1777 3553 1811 3587
rect 1811 3553 1820 3587
rect 1768 3544 1820 3553
rect 4620 3544 4672 3596
rect 10784 3544 10836 3596
rect 11336 3544 11388 3596
rect 15384 3544 15436 3596
rect 23204 3544 23256 3596
rect 1492 3519 1544 3528
rect 1492 3485 1501 3519
rect 1501 3485 1535 3519
rect 1535 3485 1544 3519
rect 1492 3476 1544 3485
rect 3148 3519 3200 3528
rect 3148 3485 3157 3519
rect 3157 3485 3191 3519
rect 3191 3485 3200 3519
rect 3148 3476 3200 3485
rect 3424 3476 3476 3528
rect 10508 3476 10560 3528
rect 15568 3519 15620 3528
rect 15568 3485 15577 3519
rect 15577 3485 15611 3519
rect 15611 3485 15620 3519
rect 15568 3476 15620 3485
rect 23112 3519 23164 3528
rect 23112 3485 23121 3519
rect 23121 3485 23155 3519
rect 23155 3485 23164 3519
rect 23112 3476 23164 3485
rect 32128 3519 32180 3528
rect 32128 3485 32137 3519
rect 32137 3485 32171 3519
rect 32171 3485 32180 3519
rect 32128 3476 32180 3485
rect 32404 3519 32456 3528
rect 32404 3485 32413 3519
rect 32413 3485 32447 3519
rect 32447 3485 32456 3519
rect 32404 3476 32456 3485
rect 4712 3340 4764 3392
rect 19984 3383 20036 3392
rect 19984 3349 19993 3383
rect 19993 3349 20027 3383
rect 20027 3349 20036 3383
rect 19984 3340 20036 3349
rect 25412 3340 25464 3392
rect 26516 3340 26568 3392
rect 27344 3340 27396 3392
rect 35808 3383 35860 3392
rect 35808 3349 35817 3383
rect 35817 3349 35851 3383
rect 35851 3349 35860 3383
rect 35808 3340 35860 3349
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 1492 3136 1544 3188
rect 3424 3136 3476 3188
rect 4620 3136 4672 3188
rect 10692 3136 10744 3188
rect 10784 3179 10836 3188
rect 10784 3145 10793 3179
rect 10793 3145 10827 3179
rect 10827 3145 10836 3179
rect 10784 3136 10836 3145
rect 14740 3136 14792 3188
rect 15568 3136 15620 3188
rect 17684 3136 17736 3188
rect 21272 3179 21324 3188
rect 21272 3145 21281 3179
rect 21281 3145 21315 3179
rect 21315 3145 21324 3179
rect 21272 3136 21324 3145
rect 23112 3136 23164 3188
rect 24584 3179 24636 3188
rect 24584 3145 24593 3179
rect 24593 3145 24627 3179
rect 24627 3145 24636 3179
rect 24584 3136 24636 3145
rect 26424 3136 26476 3188
rect 29552 3136 29604 3188
rect 32772 3136 32824 3188
rect 37372 3179 37424 3188
rect 37372 3145 37381 3179
rect 37381 3145 37415 3179
rect 37415 3145 37424 3179
rect 37372 3136 37424 3145
rect 1768 3068 1820 3120
rect 23204 3111 23256 3120
rect 23204 3077 23213 3111
rect 23213 3077 23247 3111
rect 23247 3077 23256 3111
rect 23204 3068 23256 3077
rect 4620 3000 4672 3052
rect 4804 3000 4856 3052
rect 8760 3043 8812 3052
rect 8760 3009 8769 3043
rect 8769 3009 8803 3043
rect 8803 3009 8812 3043
rect 8760 3000 8812 3009
rect 15384 3043 15436 3052
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 15660 3043 15712 3052
rect 15660 3009 15669 3043
rect 15669 3009 15703 3043
rect 15703 3009 15712 3043
rect 15660 3000 15712 3009
rect 8300 2932 8352 2984
rect 8484 2975 8536 2984
rect 8484 2941 8493 2975
rect 8493 2941 8527 2975
rect 8527 2941 8536 2975
rect 8484 2932 8536 2941
rect 10508 2975 10560 2984
rect 10508 2941 10517 2975
rect 10517 2941 10551 2975
rect 10551 2941 10560 2975
rect 10508 2932 10560 2941
rect 19984 2932 20036 2984
rect 20168 2975 20220 2984
rect 20168 2941 20177 2975
rect 20177 2941 20211 2975
rect 20211 2941 20220 2975
rect 20168 2932 20220 2941
rect 24860 2932 24912 2984
rect 29368 2932 29420 2984
rect 29552 2975 29604 2984
rect 29552 2941 29561 2975
rect 29561 2941 29595 2975
rect 29595 2941 29604 2975
rect 29552 2932 29604 2941
rect 32220 3000 32272 3052
rect 32128 2932 32180 2984
rect 35808 2975 35860 2984
rect 35808 2941 35817 2975
rect 35817 2941 35851 2975
rect 35851 2941 35860 2975
rect 35808 2932 35860 2941
rect 31300 2864 31352 2916
rect 3424 2796 3476 2848
rect 4344 2796 4396 2848
rect 19432 2796 19484 2848
rect 27528 2796 27580 2848
rect 35624 2839 35676 2848
rect 35624 2805 35633 2839
rect 35633 2805 35667 2839
rect 35667 2805 35676 2839
rect 35624 2796 35676 2805
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 3424 2635 3476 2644
rect 3424 2601 3433 2635
rect 3433 2601 3467 2635
rect 3467 2601 3476 2635
rect 3424 2592 3476 2601
rect 8484 2635 8536 2644
rect 8484 2601 8493 2635
rect 8493 2601 8527 2635
rect 8527 2601 8536 2635
rect 8484 2592 8536 2601
rect 11428 2635 11480 2644
rect 11428 2601 11437 2635
rect 11437 2601 11471 2635
rect 11471 2601 11480 2635
rect 11428 2592 11480 2601
rect 12532 2592 12584 2644
rect 15384 2592 15436 2644
rect 18328 2592 18380 2644
rect 19984 2592 20036 2644
rect 22836 2635 22888 2644
rect 22836 2601 22845 2635
rect 22845 2601 22879 2635
rect 22879 2601 22888 2635
rect 22836 2592 22888 2601
rect 29368 2635 29420 2644
rect 29368 2601 29377 2635
rect 29377 2601 29411 2635
rect 29411 2601 29420 2635
rect 29368 2592 29420 2601
rect 32128 2592 32180 2644
rect 35164 2635 35216 2644
rect 35164 2601 35173 2635
rect 35173 2601 35207 2635
rect 35207 2601 35216 2635
rect 35164 2592 35216 2601
rect 6184 2524 6236 2576
rect 11336 2524 11388 2576
rect 3700 2252 3752 2304
rect 10324 2499 10376 2508
rect 10324 2465 10333 2499
rect 10333 2465 10367 2499
rect 10367 2465 10376 2499
rect 10324 2456 10376 2465
rect 4344 2431 4396 2440
rect 4344 2397 4353 2431
rect 4353 2397 4387 2431
rect 4387 2397 4396 2431
rect 4344 2388 4396 2397
rect 29184 2524 29236 2576
rect 16120 2388 16172 2440
rect 21824 2456 21876 2508
rect 18328 2431 18380 2440
rect 18328 2397 18337 2431
rect 18337 2397 18371 2431
rect 18371 2397 18380 2431
rect 18328 2388 18380 2397
rect 19984 2388 20036 2440
rect 21640 2388 21692 2440
rect 23112 2388 23164 2440
rect 24860 2431 24912 2440
rect 24860 2397 24869 2431
rect 24869 2397 24903 2431
rect 24903 2397 24912 2431
rect 24860 2388 24912 2397
rect 27344 2388 27396 2440
rect 35808 2456 35860 2508
rect 27528 2388 27580 2440
rect 35164 2388 35216 2440
rect 18052 2363 18104 2372
rect 18052 2329 18061 2363
rect 18061 2329 18095 2363
rect 18095 2329 18104 2363
rect 18052 2320 18104 2329
rect 19800 2252 19852 2304
rect 32404 2252 32456 2304
rect 36360 2252 36412 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
rect 29092 2048 29144 2100
rect 37280 2048 37332 2100
rect 15660 1776 15712 1828
rect 16396 1776 16448 1828
rect 32404 1708 32456 1760
rect 33048 1708 33100 1760
rect 8300 1572 8352 1624
rect 17868 1572 17920 1624
rect 17040 1164 17092 1216
rect 17776 1164 17828 1216
<< metal2 >>
rect 478 40996 534 41796
rect 938 40996 994 41796
rect 1398 40996 1454 41796
rect 2318 40996 2374 41796
rect 2778 40996 2834 41796
rect 3238 41576 3294 41585
rect 3238 41511 3294 41520
rect 492 38486 520 40996
rect 952 38593 980 40996
rect 938 38584 994 38593
rect 938 38519 994 38528
rect 20 38480 72 38486
rect 20 38422 72 38428
rect 480 38480 532 38486
rect 480 38422 532 38428
rect 32 35193 60 38422
rect 1412 37777 1440 40996
rect 1492 38344 1544 38350
rect 1492 38286 1544 38292
rect 1676 38344 1728 38350
rect 1676 38286 1728 38292
rect 1504 38010 1532 38286
rect 1492 38004 1544 38010
rect 1492 37946 1544 37952
rect 1398 37768 1454 37777
rect 1398 37703 1454 37712
rect 1688 37670 1716 38286
rect 1676 37664 1728 37670
rect 1676 37606 1728 37612
rect 1584 37460 1636 37466
rect 1584 37402 1636 37408
rect 18 35184 74 35193
rect 18 35119 74 35128
rect 1596 34241 1624 37402
rect 1688 36922 1716 37606
rect 2332 37466 2360 40996
rect 2792 39098 2820 40996
rect 2962 40896 3018 40905
rect 2962 40831 3018 40840
rect 2976 40186 3004 40831
rect 2964 40180 3016 40186
rect 2964 40122 3016 40128
rect 3252 40118 3280 41511
rect 3698 40996 3754 41796
rect 4158 40996 4214 41796
rect 4618 40996 4674 41796
rect 5538 40996 5594 41796
rect 5998 40996 6054 41796
rect 6458 40996 6514 41796
rect 7378 40996 7434 41796
rect 7838 40996 7894 41796
rect 8758 40996 8814 41796
rect 9218 40996 9274 41796
rect 9678 40996 9734 41796
rect 10598 40996 10654 41796
rect 11058 40996 11114 41796
rect 11518 40996 11574 41796
rect 12438 40996 12494 41796
rect 12898 40996 12954 41796
rect 13818 40996 13874 41796
rect 14278 40996 14334 41796
rect 14738 40996 14794 41796
rect 15658 40996 15714 41796
rect 16118 40996 16174 41796
rect 16578 40996 16634 41796
rect 17498 40996 17554 41796
rect 17958 40996 18014 41796
rect 18418 40996 18474 41796
rect 19338 40996 19394 41796
rect 19798 40996 19854 41796
rect 20718 40996 20774 41796
rect 21178 40996 21234 41796
rect 21638 40996 21694 41796
rect 22558 40996 22614 41796
rect 23018 40996 23074 41796
rect 23478 40996 23534 41796
rect 24398 40996 24454 41796
rect 24858 40996 24914 41796
rect 25778 40996 25834 41796
rect 26238 40996 26294 41796
rect 26698 40996 26754 41796
rect 27618 40996 27674 41796
rect 28078 40996 28134 41796
rect 28538 40996 28594 41796
rect 29458 40996 29514 41796
rect 29918 40996 29974 41796
rect 30838 40996 30894 41796
rect 31298 40996 31354 41796
rect 31758 40996 31814 41796
rect 32678 40996 32734 41796
rect 33138 40996 33194 41796
rect 33598 40996 33654 41796
rect 34518 40996 34574 41796
rect 34978 40996 35034 41796
rect 35622 41576 35678 41585
rect 35622 41511 35678 41520
rect 3424 40248 3476 40254
rect 3422 40216 3424 40225
rect 3476 40216 3478 40225
rect 3422 40151 3478 40160
rect 3240 40112 3292 40118
rect 3240 40054 3292 40060
rect 2780 39092 2832 39098
rect 2780 39034 2832 39040
rect 2780 38752 2832 38758
rect 2700 38700 2780 38706
rect 2700 38694 2832 38700
rect 3422 38720 3478 38729
rect 2700 38678 2820 38694
rect 2700 38010 2728 38678
rect 3478 38678 3556 38706
rect 3422 38655 3478 38664
rect 2778 38176 2834 38185
rect 2778 38111 2834 38120
rect 2688 38004 2740 38010
rect 2688 37946 2740 37952
rect 2320 37460 2372 37466
rect 2320 37402 2372 37408
rect 1766 37360 1822 37369
rect 1766 37295 1822 37304
rect 1676 36916 1728 36922
rect 1676 36858 1728 36864
rect 1780 36802 1808 37295
rect 2318 37224 2374 37233
rect 2318 37159 2374 37168
rect 2332 36922 2360 37159
rect 2320 36916 2372 36922
rect 2320 36858 2372 36864
rect 1688 36774 1808 36802
rect 1582 34232 1638 34241
rect 1582 34167 1638 34176
rect 1688 29714 1716 36774
rect 1768 36712 1820 36718
rect 1768 36654 1820 36660
rect 1780 36038 1808 36654
rect 1768 36032 1820 36038
rect 1768 35974 1820 35980
rect 1676 29708 1728 29714
rect 1676 29650 1728 29656
rect 1398 29336 1454 29345
rect 1688 29306 1716 29650
rect 1398 29271 1454 29280
rect 1676 29300 1728 29306
rect 1412 28626 1440 29271
rect 1676 29242 1728 29248
rect 1400 28620 1452 28626
rect 1400 28562 1452 28568
rect 1412 28218 1440 28562
rect 1400 28212 1452 28218
rect 1400 28154 1452 28160
rect 1492 27532 1544 27538
rect 1492 27474 1544 27480
rect 1504 26790 1532 27474
rect 1492 26784 1544 26790
rect 1492 26726 1544 26732
rect 1400 26580 1452 26586
rect 1400 26522 1452 26528
rect 1412 25906 1440 26522
rect 1400 25900 1452 25906
rect 1400 25842 1452 25848
rect 1412 24274 1440 25842
rect 1400 24268 1452 24274
rect 1400 24210 1452 24216
rect 1412 23798 1440 24210
rect 1400 23792 1452 23798
rect 1400 23734 1452 23740
rect 1412 23186 1440 23734
rect 1400 23180 1452 23186
rect 1400 23122 1452 23128
rect 1400 16788 1452 16794
rect 1400 16730 1452 16736
rect 1412 16114 1440 16730
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1412 15026 1440 16050
rect 1400 15020 1452 15026
rect 1400 14962 1452 14968
rect 1412 14618 1440 14962
rect 1400 14612 1452 14618
rect 1400 14554 1452 14560
rect 1412 13394 1440 14554
rect 1400 13388 1452 13394
rect 1400 13330 1452 13336
rect 1412 12850 1440 13330
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1504 12322 1532 26726
rect 1676 25832 1728 25838
rect 1676 25774 1728 25780
rect 1688 25158 1716 25774
rect 1676 25152 1728 25158
rect 1676 25094 1728 25100
rect 1584 24200 1636 24206
rect 1584 24142 1636 24148
rect 1596 23905 1624 24142
rect 1582 23896 1638 23905
rect 1582 23831 1584 23840
rect 1636 23831 1638 23840
rect 1584 23802 1636 23808
rect 1676 23112 1728 23118
rect 1676 23054 1728 23060
rect 1688 22778 1716 23054
rect 1676 22772 1728 22778
rect 1676 22714 1728 22720
rect 1674 21176 1730 21185
rect 1674 21111 1730 21120
rect 1688 18834 1716 21111
rect 1780 19145 1808 35974
rect 2792 31346 2820 38111
rect 3422 34096 3478 34105
rect 3422 34031 3478 34040
rect 3436 33289 3464 34031
rect 3422 33280 3478 33289
rect 3422 33215 3478 33224
rect 3528 31906 3556 38678
rect 3712 38486 3740 40996
rect 4172 39370 4200 40996
rect 4160 39364 4212 39370
rect 4160 39306 4212 39312
rect 4220 39196 4516 39216
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4298 39142 4300 39194
rect 4362 39142 4374 39194
rect 4436 39142 4438 39194
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4220 39120 4516 39140
rect 3700 38480 3752 38486
rect 3700 38422 3752 38428
rect 4632 38418 4660 40996
rect 5172 39364 5224 39370
rect 5172 39306 5224 39312
rect 4620 38412 4672 38418
rect 4620 38354 4672 38360
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 4066 36816 4122 36825
rect 4066 36751 4122 36760
rect 4080 35465 4108 36751
rect 5184 36242 5212 39306
rect 5448 38888 5500 38894
rect 5448 38830 5500 38836
rect 5460 38350 5488 38830
rect 5552 38554 5580 40996
rect 5540 38548 5592 38554
rect 5540 38490 5592 38496
rect 5540 38412 5592 38418
rect 5540 38354 5592 38360
rect 5448 38344 5500 38350
rect 5448 38286 5500 38292
rect 5460 37874 5488 38286
rect 5552 38010 5580 38354
rect 5540 38004 5592 38010
rect 5540 37946 5592 37952
rect 5448 37868 5500 37874
rect 5448 37810 5500 37816
rect 5460 37330 5488 37810
rect 6012 37330 6040 40996
rect 6472 39030 6500 40996
rect 7012 40248 7064 40254
rect 7012 40190 7064 40196
rect 6460 39024 6512 39030
rect 6460 38966 6512 38972
rect 6736 38548 6788 38554
rect 6736 38490 6788 38496
rect 5448 37324 5500 37330
rect 5448 37266 5500 37272
rect 6000 37324 6052 37330
rect 6000 37266 6052 37272
rect 5460 36786 5488 37266
rect 6012 36922 6040 37266
rect 6000 36916 6052 36922
rect 6000 36858 6052 36864
rect 5448 36780 5500 36786
rect 5448 36722 5500 36728
rect 5460 36242 5488 36722
rect 5172 36236 5224 36242
rect 5172 36178 5224 36184
rect 5448 36236 5500 36242
rect 5448 36178 5500 36184
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 5184 35834 5212 36178
rect 5460 35834 5488 36178
rect 5172 35828 5224 35834
rect 5172 35770 5224 35776
rect 5448 35828 5500 35834
rect 5448 35770 5500 35776
rect 4066 35456 4122 35465
rect 4066 35391 4122 35400
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 6182 33416 6238 33425
rect 6182 33351 6238 33360
rect 6092 32972 6144 32978
rect 6092 32914 6144 32920
rect 5998 32872 6054 32881
rect 6104 32858 6132 32914
rect 6054 32830 6132 32858
rect 5998 32807 6054 32816
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 6012 32570 6040 32807
rect 6000 32564 6052 32570
rect 6000 32506 6052 32512
rect 3436 31878 3556 31906
rect 3436 31668 3464 31878
rect 3792 31680 3844 31686
rect 3436 31640 3556 31668
rect 3056 31408 3108 31414
rect 3056 31350 3108 31356
rect 2780 31340 2832 31346
rect 2780 31282 2832 31288
rect 2688 31136 2740 31142
rect 2688 31078 2740 31084
rect 2700 30580 2728 31078
rect 2700 30552 2820 30580
rect 2792 30258 2820 30552
rect 2780 30252 2832 30258
rect 2780 30194 2832 30200
rect 2044 29640 2096 29646
rect 2044 29582 2096 29588
rect 2056 29170 2084 29582
rect 2780 29504 2832 29510
rect 2780 29446 2832 29452
rect 2044 29164 2096 29170
rect 2044 29106 2096 29112
rect 2056 28626 2084 29106
rect 2044 28620 2096 28626
rect 2044 28562 2096 28568
rect 2056 28218 2084 28562
rect 2044 28212 2096 28218
rect 2044 28154 2096 28160
rect 2056 27470 2084 28154
rect 2792 27985 2820 29446
rect 2962 28520 3018 28529
rect 3068 28506 3096 31350
rect 3240 30184 3292 30190
rect 3422 30152 3478 30161
rect 3292 30132 3422 30138
rect 3240 30126 3422 30132
rect 3252 30110 3422 30126
rect 3422 30087 3478 30096
rect 3436 29850 3464 30087
rect 3424 29844 3476 29850
rect 3344 29804 3424 29832
rect 3344 29170 3372 29804
rect 3424 29786 3476 29792
rect 3332 29164 3384 29170
rect 3332 29106 3384 29112
rect 3148 29028 3200 29034
rect 3148 28970 3200 28976
rect 3160 28665 3188 28970
rect 3146 28656 3202 28665
rect 3146 28591 3202 28600
rect 3068 28478 3188 28506
rect 2962 28455 3018 28464
rect 2778 27976 2834 27985
rect 2778 27911 2834 27920
rect 2044 27464 2096 27470
rect 2044 27406 2096 27412
rect 2056 27130 2084 27406
rect 2044 27124 2096 27130
rect 2044 27066 2096 27072
rect 2056 26586 2084 27066
rect 2778 26616 2834 26625
rect 2044 26580 2096 26586
rect 2778 26551 2834 26560
rect 2044 26522 2096 26528
rect 2792 26042 2820 26551
rect 2780 26036 2832 26042
rect 2780 25978 2832 25984
rect 2976 25265 3004 28455
rect 3056 28416 3108 28422
rect 3056 28358 3108 28364
rect 3068 27577 3096 28358
rect 3054 27568 3110 27577
rect 3054 27503 3110 27512
rect 3056 27464 3108 27470
rect 3054 27432 3056 27441
rect 3108 27432 3110 27441
rect 3054 27367 3110 27376
rect 2962 25256 3018 25265
rect 2962 25191 3018 25200
rect 2964 25152 3016 25158
rect 2964 25094 3016 25100
rect 1950 23216 2006 23225
rect 1950 23151 2006 23160
rect 1860 22024 1912 22030
rect 1860 21966 1912 21972
rect 1872 21010 1900 21966
rect 1964 21554 1992 23151
rect 2596 22500 2648 22506
rect 2596 22442 2648 22448
rect 2044 21888 2096 21894
rect 2044 21830 2096 21836
rect 2410 21856 2466 21865
rect 1952 21548 2004 21554
rect 1952 21490 2004 21496
rect 2056 21486 2084 21830
rect 2410 21791 2466 21800
rect 2044 21480 2096 21486
rect 2044 21422 2096 21428
rect 1860 21004 1912 21010
rect 1860 20946 1912 20952
rect 1872 19990 1900 20946
rect 1952 20936 2004 20942
rect 1952 20878 2004 20884
rect 1964 20058 1992 20878
rect 2424 20466 2452 21791
rect 2608 20505 2636 22442
rect 2872 22092 2924 22098
rect 2872 22034 2924 22040
rect 2884 21554 2912 22034
rect 2872 21548 2924 21554
rect 2872 21490 2924 21496
rect 2594 20496 2650 20505
rect 2412 20460 2464 20466
rect 2594 20431 2650 20440
rect 2412 20402 2464 20408
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 2688 20052 2740 20058
rect 2688 19994 2740 20000
rect 1860 19984 1912 19990
rect 1860 19926 1912 19932
rect 1964 19514 1992 19994
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 1766 19136 1822 19145
rect 1766 19071 1822 19080
rect 1964 18834 1992 19450
rect 1676 18828 1728 18834
rect 1676 18770 1728 18776
rect 1952 18828 2004 18834
rect 1952 18770 2004 18776
rect 1688 18426 1716 18770
rect 1964 18426 1992 18770
rect 2596 18624 2648 18630
rect 2596 18566 2648 18572
rect 1676 18420 1728 18426
rect 1676 18362 1728 18368
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1964 17898 1992 18362
rect 1872 17882 1992 17898
rect 1860 17876 1992 17882
rect 1912 17870 1992 17876
rect 1860 17818 1912 17824
rect 1872 17134 1900 17818
rect 1952 17808 2004 17814
rect 1950 17776 1952 17785
rect 2004 17776 2006 17785
rect 1950 17711 2006 17720
rect 2412 17740 2464 17746
rect 2412 17682 2464 17688
rect 2504 17740 2556 17746
rect 2504 17682 2556 17688
rect 2424 17202 2452 17682
rect 2412 17196 2464 17202
rect 2412 17138 2464 17144
rect 1860 17128 1912 17134
rect 1860 17070 1912 17076
rect 1872 16794 1900 17070
rect 2044 16992 2096 16998
rect 2044 16934 2096 16940
rect 2056 16794 2084 16934
rect 2424 16794 2452 17138
rect 2516 17134 2544 17682
rect 2504 17128 2556 17134
rect 2504 17070 2556 17076
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 2044 16788 2096 16794
rect 2044 16730 2096 16736
rect 2412 16788 2464 16794
rect 2412 16730 2464 16736
rect 1674 16416 1730 16425
rect 1674 16351 1730 16360
rect 1688 16114 1716 16351
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1688 15706 1716 16050
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1596 14278 1624 14962
rect 2516 14550 2544 17070
rect 2504 14544 2556 14550
rect 2504 14486 2556 14492
rect 1584 14272 1636 14278
rect 1584 14214 1636 14220
rect 1596 13841 1624 14214
rect 1582 13832 1638 13841
rect 1582 13767 1638 13776
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 1596 13025 1624 13262
rect 1582 13016 1638 13025
rect 1582 12951 1584 12960
rect 1636 12951 1638 12960
rect 1584 12922 1636 12928
rect 1412 12294 1532 12322
rect 1584 12300 1636 12306
rect 18 5128 74 5137
rect 18 5063 74 5072
rect 32 800 60 5063
rect 938 3768 994 3777
rect 938 3703 994 3712
rect 478 3088 534 3097
rect 478 3023 534 3032
rect 492 800 520 3023
rect 952 800 980 3703
rect 18 0 74 800
rect 478 0 534 800
rect 938 0 994 800
rect 1412 785 1440 12294
rect 1584 12242 1636 12248
rect 1596 12186 1624 12242
rect 1504 12158 1624 12186
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1504 11558 1532 12158
rect 1964 11694 1992 12174
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 1964 11558 1992 11630
rect 1492 11552 1544 11558
rect 1492 11494 1544 11500
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 1504 11121 1532 11494
rect 1964 11218 1992 11494
rect 1952 11212 2004 11218
rect 1952 11154 2004 11160
rect 1584 11144 1636 11150
rect 1490 11112 1546 11121
rect 1584 11086 1636 11092
rect 1490 11047 1546 11056
rect 1596 10470 1624 11086
rect 1964 10470 1992 11154
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1596 10305 1624 10406
rect 1582 10296 1638 10305
rect 1582 10231 1638 10240
rect 1964 9518 1992 10406
rect 2608 9722 2636 18566
rect 2700 17746 2728 19994
rect 2688 17740 2740 17746
rect 2688 17682 2740 17688
rect 2884 15162 2912 21490
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2700 14074 2728 14554
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2700 13870 2728 14010
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2884 11121 2912 14962
rect 2870 11112 2926 11121
rect 2870 11047 2926 11056
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2410 9616 2466 9625
rect 2884 9586 2912 11047
rect 2410 9551 2466 9560
rect 2872 9580 2924 9586
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 1964 9178 1992 9454
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 7041 1532 8298
rect 1490 7032 1546 7041
rect 1490 6967 1546 6976
rect 1858 6760 1914 6769
rect 1858 6695 1914 6704
rect 1766 6216 1822 6225
rect 1766 6151 1822 6160
rect 1780 3602 1808 6151
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 1492 3528 1544 3534
rect 1492 3470 1544 3476
rect 1504 3194 1532 3470
rect 1492 3188 1544 3194
rect 1492 3130 1544 3136
rect 1780 3126 1808 3538
rect 1768 3120 1820 3126
rect 1768 3062 1820 3068
rect 1872 800 1900 6695
rect 2332 800 2360 9454
rect 2424 8945 2452 9551
rect 2872 9522 2924 9528
rect 2410 8936 2466 8945
rect 2410 8871 2466 8880
rect 2686 8256 2742 8265
rect 2742 8214 2820 8242
rect 2686 8191 2742 8200
rect 2792 7313 2820 8214
rect 2778 7304 2834 7313
rect 2778 7239 2834 7248
rect 2976 2802 3004 25094
rect 3054 23624 3110 23633
rect 3054 23559 3056 23568
rect 3108 23559 3110 23568
rect 3056 23530 3108 23536
rect 3160 22710 3188 28478
rect 3424 27328 3476 27334
rect 3424 27270 3476 27276
rect 3436 26994 3464 27270
rect 3424 26988 3476 26994
rect 3424 26930 3476 26936
rect 3332 26920 3384 26926
rect 3332 26862 3384 26868
rect 3344 26586 3372 26862
rect 3332 26580 3384 26586
rect 3332 26522 3384 26528
rect 3332 24880 3384 24886
rect 3332 24822 3384 24828
rect 3344 23066 3372 24822
rect 3436 24138 3464 26930
rect 3528 24886 3556 31640
rect 3792 31622 3844 31628
rect 3804 31278 3832 31622
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 4068 31340 4120 31346
rect 4068 31282 4120 31288
rect 3792 31272 3844 31278
rect 3792 31214 3844 31220
rect 3804 30394 3832 31214
rect 4080 30977 4108 31282
rect 4620 31204 4672 31210
rect 4620 31146 4672 31152
rect 4066 30968 4122 30977
rect 4066 30903 4068 30912
rect 4120 30903 4122 30912
rect 4068 30874 4120 30880
rect 4080 30843 4108 30874
rect 4068 30660 4120 30666
rect 4068 30602 4120 30608
rect 4080 30569 4108 30602
rect 4066 30560 4122 30569
rect 4066 30495 4122 30504
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 3792 30388 3844 30394
rect 3792 30330 3844 30336
rect 4632 30190 4660 31146
rect 4986 30968 5042 30977
rect 4986 30903 5042 30912
rect 4894 30288 4950 30297
rect 4894 30223 4950 30232
rect 4620 30184 4672 30190
rect 4620 30126 4672 30132
rect 4066 29744 4122 29753
rect 4066 29679 4122 29688
rect 3976 28756 4028 28762
rect 3976 28698 4028 28704
rect 3700 28212 3752 28218
rect 3700 28154 3752 28160
rect 3516 24880 3568 24886
rect 3516 24822 3568 24828
rect 3516 24744 3568 24750
rect 3516 24686 3568 24692
rect 3528 24410 3556 24686
rect 3516 24404 3568 24410
rect 3516 24346 3568 24352
rect 3424 24132 3476 24138
rect 3424 24074 3476 24080
rect 3422 23760 3478 23769
rect 3422 23695 3424 23704
rect 3476 23695 3478 23704
rect 3424 23666 3476 23672
rect 3516 23112 3568 23118
rect 3344 23038 3464 23066
rect 3516 23054 3568 23060
rect 3712 23066 3740 28154
rect 3882 27024 3938 27033
rect 3882 26959 3938 26968
rect 3896 26926 3924 26959
rect 3884 26920 3936 26926
rect 3884 26862 3936 26868
rect 3790 24168 3846 24177
rect 3790 24103 3846 24112
rect 3804 23866 3832 24103
rect 3884 24064 3936 24070
rect 3884 24006 3936 24012
rect 3792 23860 3844 23866
rect 3792 23802 3844 23808
rect 3896 23497 3924 24006
rect 3882 23488 3938 23497
rect 3882 23423 3938 23432
rect 3882 23352 3938 23361
rect 3988 23338 4016 28698
rect 4080 25945 4108 29679
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 4632 27130 4660 30126
rect 4908 29306 4936 30223
rect 4896 29300 4948 29306
rect 4896 29242 4948 29248
rect 4710 28928 4766 28937
rect 4710 28863 4766 28872
rect 4724 28626 4752 28863
rect 5000 28762 5028 30903
rect 4988 28756 5040 28762
rect 4988 28698 5040 28704
rect 4712 28620 4764 28626
rect 4712 28562 4764 28568
rect 5356 28620 5408 28626
rect 5356 28562 5408 28568
rect 4724 28218 4752 28562
rect 4712 28212 4764 28218
rect 4712 28154 4764 28160
rect 5368 27878 5396 28562
rect 6092 28416 6144 28422
rect 6092 28358 6144 28364
rect 5356 27872 5408 27878
rect 5356 27814 5408 27820
rect 4896 27328 4948 27334
rect 4896 27270 4948 27276
rect 4620 27124 4672 27130
rect 4620 27066 4672 27072
rect 4710 27024 4766 27033
rect 4710 26959 4766 26968
rect 4528 26852 4580 26858
rect 4528 26794 4580 26800
rect 4540 26586 4568 26794
rect 4528 26580 4580 26586
rect 4528 26522 4580 26528
rect 4540 26466 4568 26522
rect 4540 26438 4660 26466
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 4066 25936 4122 25945
rect 4632 25906 4660 26438
rect 4066 25871 4122 25880
rect 4620 25900 4672 25906
rect 4620 25842 4672 25848
rect 4528 25832 4580 25838
rect 4528 25774 4580 25780
rect 4540 25537 4568 25774
rect 4526 25528 4582 25537
rect 4526 25463 4582 25472
rect 4724 25106 4752 26959
rect 4804 25288 4856 25294
rect 4804 25230 4856 25236
rect 4632 25078 4752 25106
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 3988 23310 4108 23338
rect 3882 23287 3884 23296
rect 3936 23287 3938 23296
rect 3884 23258 3936 23264
rect 3974 23080 4030 23089
rect 3240 22976 3292 22982
rect 3240 22918 3292 22924
rect 3332 22976 3384 22982
rect 3332 22918 3384 22924
rect 3148 22704 3200 22710
rect 3068 22664 3148 22692
rect 3068 22574 3096 22664
rect 3148 22646 3200 22652
rect 3252 22574 3280 22918
rect 3056 22568 3108 22574
rect 3056 22510 3108 22516
rect 3240 22568 3292 22574
rect 3240 22510 3292 22516
rect 3240 21480 3292 21486
rect 3240 21422 3292 21428
rect 3148 21412 3200 21418
rect 3148 21354 3200 21360
rect 3056 21344 3108 21350
rect 3056 21286 3108 21292
rect 3068 20398 3096 21286
rect 3160 21078 3188 21354
rect 3148 21072 3200 21078
rect 3148 21014 3200 21020
rect 3252 20466 3280 21422
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 3240 20460 3292 20466
rect 3240 20402 3292 20408
rect 3056 20392 3108 20398
rect 3056 20334 3108 20340
rect 3068 20058 3096 20334
rect 3056 20052 3108 20058
rect 3056 19994 3108 20000
rect 3160 19990 3188 20402
rect 3252 20262 3280 20402
rect 3240 20256 3292 20262
rect 3240 20198 3292 20204
rect 3148 19984 3200 19990
rect 3148 19926 3200 19932
rect 3160 19417 3188 19926
rect 3146 19408 3202 19417
rect 3146 19343 3202 19352
rect 3054 18728 3110 18737
rect 3054 18663 3110 18672
rect 3068 13462 3096 18663
rect 3148 18624 3200 18630
rect 3148 18566 3200 18572
rect 3160 16794 3188 18566
rect 3252 17678 3280 20198
rect 3344 17882 3372 22918
rect 3436 19530 3464 23038
rect 3528 22642 3556 23054
rect 3712 23038 3924 23066
rect 3700 22976 3752 22982
rect 3700 22918 3752 22924
rect 3712 22681 3740 22918
rect 3698 22672 3754 22681
rect 3516 22636 3568 22642
rect 3698 22607 3754 22616
rect 3516 22578 3568 22584
rect 3528 22234 3556 22578
rect 3792 22568 3844 22574
rect 3792 22510 3844 22516
rect 3516 22228 3568 22234
rect 3516 22170 3568 22176
rect 3804 22166 3832 22510
rect 3792 22160 3844 22166
rect 3792 22102 3844 22108
rect 3516 21888 3568 21894
rect 3516 21830 3568 21836
rect 3528 21593 3556 21830
rect 3514 21584 3570 21593
rect 3514 21519 3570 21528
rect 3528 20602 3556 21519
rect 3516 20596 3568 20602
rect 3516 20538 3568 20544
rect 3516 20460 3568 20466
rect 3516 20402 3568 20408
rect 3528 20058 3556 20402
rect 3700 20324 3752 20330
rect 3700 20266 3752 20272
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3436 19502 3556 19530
rect 3712 19514 3740 20266
rect 3436 19417 3464 19443
rect 3422 19408 3478 19417
rect 3422 19343 3424 19352
rect 3476 19343 3478 19352
rect 3424 19314 3476 19320
rect 3332 17876 3384 17882
rect 3332 17818 3384 17824
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 3252 17338 3280 17614
rect 3240 17332 3292 17338
rect 3240 17274 3292 17280
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 3160 16454 3188 16730
rect 3148 16448 3200 16454
rect 3148 16390 3200 16396
rect 3252 15502 3280 17274
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 3436 15026 3464 19314
rect 3528 19224 3556 19502
rect 3700 19508 3752 19514
rect 3700 19450 3752 19456
rect 3528 19196 3648 19224
rect 3514 19136 3570 19145
rect 3514 19071 3570 19080
rect 3528 18970 3556 19071
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3516 17740 3568 17746
rect 3516 17682 3568 17688
rect 3528 17338 3556 17682
rect 3516 17332 3568 17338
rect 3516 17274 3568 17280
rect 3528 16998 3556 17274
rect 3516 16992 3568 16998
rect 3516 16934 3568 16940
rect 3514 15056 3570 15065
rect 3424 15020 3476 15026
rect 3514 14991 3570 15000
rect 3424 14962 3476 14968
rect 3424 14816 3476 14822
rect 3424 14758 3476 14764
rect 3436 14521 3464 14758
rect 3528 14618 3556 14991
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3422 14512 3478 14521
rect 3422 14447 3478 14456
rect 3056 13456 3108 13462
rect 3056 13398 3108 13404
rect 3146 12336 3202 12345
rect 3146 12271 3148 12280
rect 3200 12271 3202 12280
rect 3148 12242 3200 12248
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 3068 11286 3096 11698
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3056 11280 3108 11286
rect 3056 11222 3108 11228
rect 3436 11082 3464 11630
rect 3620 11286 3648 19196
rect 3804 18850 3832 22102
rect 3896 21690 3924 23038
rect 3974 23015 4030 23024
rect 3988 22234 4016 23015
rect 4080 22574 4108 23310
rect 4632 23186 4660 25078
rect 4710 24984 4766 24993
rect 4710 24919 4766 24928
rect 4724 24206 4752 24919
rect 4712 24200 4764 24206
rect 4712 24142 4764 24148
rect 4724 23866 4752 24142
rect 4712 23860 4764 23866
rect 4712 23802 4764 23808
rect 4816 23594 4844 25230
rect 4908 24342 4936 27270
rect 5078 26616 5134 26625
rect 5078 26551 5134 26560
rect 5092 26450 5120 26551
rect 5080 26444 5132 26450
rect 5080 26386 5132 26392
rect 4986 26344 5042 26353
rect 4986 26279 4988 26288
rect 5040 26279 5042 26288
rect 4988 26250 5040 26256
rect 5092 26042 5120 26386
rect 5264 26308 5316 26314
rect 5264 26250 5316 26256
rect 5080 26036 5132 26042
rect 5080 25978 5132 25984
rect 5092 25362 5120 25978
rect 5276 25702 5304 26250
rect 5264 25696 5316 25702
rect 5264 25638 5316 25644
rect 5080 25356 5132 25362
rect 5080 25298 5132 25304
rect 5276 25294 5304 25638
rect 5264 25288 5316 25294
rect 5264 25230 5316 25236
rect 4988 25220 5040 25226
rect 4988 25162 5040 25168
rect 4896 24336 4948 24342
rect 4896 24278 4948 24284
rect 4804 23588 4856 23594
rect 4804 23530 4856 23536
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 4632 22778 4660 23122
rect 4620 22772 4672 22778
rect 4620 22714 4672 22720
rect 4068 22568 4120 22574
rect 4068 22510 4120 22516
rect 4816 22420 4844 23530
rect 4896 22976 4948 22982
rect 4896 22918 4948 22924
rect 4908 22574 4936 22918
rect 4896 22568 4948 22574
rect 4896 22510 4948 22516
rect 4816 22392 4936 22420
rect 4802 22264 4858 22273
rect 3976 22228 4028 22234
rect 4802 22199 4858 22208
rect 3976 22170 4028 22176
rect 4620 22160 4672 22166
rect 4620 22102 4672 22108
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 3884 21684 3936 21690
rect 3884 21626 3936 21632
rect 4632 21400 4660 22102
rect 4712 22092 4764 22098
rect 4712 22034 4764 22040
rect 4724 21554 4752 22034
rect 4712 21548 4764 21554
rect 4712 21490 4764 21496
rect 4540 21372 4660 21400
rect 3882 21176 3938 21185
rect 4540 21146 4568 21372
rect 4816 21298 4844 22199
rect 4632 21270 4844 21298
rect 3882 21111 3884 21120
rect 3936 21111 3938 21120
rect 4068 21140 4120 21146
rect 3884 21082 3936 21088
rect 4068 21082 4120 21088
rect 4528 21140 4580 21146
rect 4528 21082 4580 21088
rect 3976 20256 4028 20262
rect 3976 20198 4028 20204
rect 3988 20097 4016 20198
rect 3974 20088 4030 20097
rect 3974 20023 4030 20032
rect 4080 19972 4108 21082
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 4632 20602 4660 21270
rect 4908 21162 4936 22392
rect 4724 21134 4936 21162
rect 4620 20596 4672 20602
rect 4620 20538 4672 20544
rect 4618 20496 4674 20505
rect 4618 20431 4674 20440
rect 4632 20058 4660 20431
rect 4620 20052 4672 20058
rect 4620 19994 4672 20000
rect 3988 19944 4108 19972
rect 3884 19712 3936 19718
rect 3884 19654 3936 19660
rect 3896 19281 3924 19654
rect 3882 19272 3938 19281
rect 3882 19207 3938 19216
rect 3712 18822 3832 18850
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3712 11098 3740 18822
rect 3884 17536 3936 17542
rect 3884 17478 3936 17484
rect 3896 16561 3924 17478
rect 3988 16969 4016 19944
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4066 19408 4122 19417
rect 4066 19343 4122 19352
rect 4080 18465 4108 19343
rect 4434 18728 4490 18737
rect 4434 18663 4436 18672
rect 4488 18663 4490 18672
rect 4436 18634 4488 18640
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4066 18456 4122 18465
rect 4220 18448 4516 18468
rect 4632 18426 4660 19994
rect 4066 18391 4122 18400
rect 4620 18420 4672 18426
rect 4620 18362 4672 18368
rect 4528 18080 4580 18086
rect 4528 18022 4580 18028
rect 4540 17649 4568 18022
rect 4618 17912 4674 17921
rect 4618 17847 4620 17856
rect 4672 17847 4674 17856
rect 4620 17818 4672 17824
rect 4526 17640 4582 17649
rect 4526 17575 4582 17584
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 3974 16960 4030 16969
rect 3974 16895 4030 16904
rect 3988 16794 4016 16895
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 4068 16720 4120 16726
rect 4068 16662 4120 16668
rect 3882 16552 3938 16561
rect 3882 16487 3938 16496
rect 4080 16250 4108 16662
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 4620 16176 4672 16182
rect 4620 16118 4672 16124
rect 3884 15972 3936 15978
rect 3884 15914 3936 15920
rect 3896 15473 3924 15914
rect 3882 15464 3938 15473
rect 3882 15399 3938 15408
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4632 15144 4660 16118
rect 4724 16114 4752 21134
rect 4896 21004 4948 21010
rect 4896 20946 4948 20952
rect 4908 20534 4936 20946
rect 4896 20528 4948 20534
rect 4896 20470 4948 20476
rect 4896 20392 4948 20398
rect 4896 20334 4948 20340
rect 4804 20256 4856 20262
rect 4804 20198 4856 20204
rect 4816 19174 4844 20198
rect 4908 19242 4936 20334
rect 4896 19236 4948 19242
rect 4896 19178 4948 19184
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4816 19009 4844 19110
rect 4802 19000 4858 19009
rect 4802 18935 4858 18944
rect 4894 18864 4950 18873
rect 4894 18799 4950 18808
rect 4908 18426 4936 18799
rect 4896 18420 4948 18426
rect 4896 18362 4948 18368
rect 4896 16652 4948 16658
rect 5000 16640 5028 25162
rect 5172 24744 5224 24750
rect 5172 24686 5224 24692
rect 5080 24608 5132 24614
rect 5080 24550 5132 24556
rect 5092 22001 5120 24550
rect 5184 24206 5212 24686
rect 5264 24268 5316 24274
rect 5264 24210 5316 24216
rect 5172 24200 5224 24206
rect 5172 24142 5224 24148
rect 5276 23526 5304 24210
rect 5264 23520 5316 23526
rect 5264 23462 5316 23468
rect 5172 23044 5224 23050
rect 5172 22986 5224 22992
rect 5184 22642 5212 22986
rect 5276 22778 5304 23462
rect 5368 23066 5396 27814
rect 6104 27606 6132 28358
rect 6092 27600 6144 27606
rect 6092 27542 6144 27548
rect 5724 27532 5776 27538
rect 5724 27474 5776 27480
rect 5816 27532 5868 27538
rect 5816 27474 5868 27480
rect 5736 27062 5764 27474
rect 5828 27130 5856 27474
rect 6104 27130 6132 27542
rect 5816 27124 5868 27130
rect 5816 27066 5868 27072
rect 6092 27124 6144 27130
rect 6092 27066 6144 27072
rect 5724 27056 5776 27062
rect 5724 26998 5776 27004
rect 5828 26489 5856 27066
rect 5814 26480 5870 26489
rect 5814 26415 5870 26424
rect 6000 26376 6052 26382
rect 6000 26318 6052 26324
rect 5722 26208 5778 26217
rect 5722 26143 5778 26152
rect 5448 25356 5500 25362
rect 5448 25298 5500 25304
rect 5460 24818 5488 25298
rect 5448 24812 5500 24818
rect 5448 24754 5500 24760
rect 5460 23186 5488 24754
rect 5632 24676 5684 24682
rect 5632 24618 5684 24624
rect 5540 24268 5592 24274
rect 5540 24210 5592 24216
rect 5552 23798 5580 24210
rect 5540 23792 5592 23798
rect 5540 23734 5592 23740
rect 5644 23610 5672 24618
rect 5552 23582 5672 23610
rect 5448 23180 5500 23186
rect 5448 23122 5500 23128
rect 5368 23038 5488 23066
rect 5356 22976 5408 22982
rect 5356 22918 5408 22924
rect 5264 22772 5316 22778
rect 5264 22714 5316 22720
rect 5368 22658 5396 22918
rect 5172 22636 5224 22642
rect 5172 22578 5224 22584
rect 5276 22630 5396 22658
rect 5170 22400 5226 22409
rect 5170 22335 5226 22344
rect 5078 21992 5134 22001
rect 5078 21927 5134 21936
rect 5080 21888 5132 21894
rect 5080 21830 5132 21836
rect 5092 19310 5120 21830
rect 5184 20058 5212 22335
rect 5276 22098 5304 22630
rect 5460 22556 5488 23038
rect 5368 22528 5488 22556
rect 5264 22092 5316 22098
rect 5264 22034 5316 22040
rect 5262 21992 5318 22001
rect 5262 21927 5318 21936
rect 5276 20942 5304 21927
rect 5264 20936 5316 20942
rect 5264 20878 5316 20884
rect 5276 20777 5304 20878
rect 5262 20768 5318 20777
rect 5262 20703 5318 20712
rect 5276 20602 5304 20703
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5172 20052 5224 20058
rect 5172 19994 5224 20000
rect 5264 19984 5316 19990
rect 5262 19952 5264 19961
rect 5316 19952 5318 19961
rect 5262 19887 5318 19896
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 5276 19378 5304 19654
rect 5264 19372 5316 19378
rect 5264 19314 5316 19320
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 4948 16612 5028 16640
rect 4896 16594 4948 16600
rect 4988 16516 5040 16522
rect 4988 16458 5040 16464
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4816 15706 4844 16186
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4896 15564 4948 15570
rect 4896 15506 4948 15512
rect 4712 15428 4764 15434
rect 4712 15370 4764 15376
rect 4356 15116 4660 15144
rect 4356 14958 4384 15116
rect 4724 15026 4752 15370
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4344 14952 4396 14958
rect 3882 14920 3938 14929
rect 4344 14894 4396 14900
rect 3882 14855 3938 14864
rect 3896 14618 3924 14855
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3988 14657 4016 14758
rect 3974 14648 4030 14657
rect 3884 14612 3936 14618
rect 4356 14618 4384 14894
rect 3974 14583 4030 14592
rect 4344 14612 4396 14618
rect 3884 14554 3936 14560
rect 4344 14554 4396 14560
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 3976 13864 4028 13870
rect 4080 13852 4108 14418
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4724 14074 4752 14962
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 4816 14550 4844 14894
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4028 13824 4108 13852
rect 3976 13806 4028 13812
rect 4080 13258 4108 13824
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4632 12102 4660 12242
rect 4712 12164 4764 12170
rect 4712 12106 4764 12112
rect 4620 12096 4672 12102
rect 4618 12064 4620 12073
rect 4672 12064 4674 12073
rect 4220 11996 4516 12016
rect 4618 11999 4674 12008
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4632 11762 4660 11999
rect 4724 11830 4752 12106
rect 4712 11824 4764 11830
rect 4712 11766 4764 11772
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 3790 11656 3846 11665
rect 3790 11591 3846 11600
rect 3424 11076 3476 11082
rect 3424 11018 3476 11024
rect 3620 11070 3740 11098
rect 3620 8401 3648 11070
rect 3700 11008 3752 11014
rect 3700 10950 3752 10956
rect 3712 10810 3740 10950
rect 3700 10804 3752 10810
rect 3700 10746 3752 10752
rect 3804 9489 3832 11591
rect 4160 11144 4212 11150
rect 4080 11092 4160 11098
rect 4080 11086 4212 11092
rect 4620 11144 4672 11150
rect 4724 11132 4752 11766
rect 4816 11218 4844 14486
rect 4908 14385 4936 15506
rect 5000 15366 5028 16458
rect 5092 16182 5120 19246
rect 5276 19242 5304 19314
rect 5172 19236 5224 19242
rect 5172 19178 5224 19184
rect 5264 19236 5316 19242
rect 5264 19178 5316 19184
rect 5184 18902 5212 19178
rect 5172 18896 5224 18902
rect 5172 18838 5224 18844
rect 5262 18456 5318 18465
rect 5262 18391 5264 18400
rect 5316 18391 5318 18400
rect 5264 18362 5316 18368
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 5184 16658 5212 17818
rect 5368 16794 5396 22528
rect 5552 22098 5580 23582
rect 5632 23180 5684 23186
rect 5632 23122 5684 23128
rect 5540 22092 5592 22098
rect 5540 22034 5592 22040
rect 5448 21888 5500 21894
rect 5448 21830 5500 21836
rect 5460 20806 5488 21830
rect 5552 21690 5580 22034
rect 5644 21894 5672 23122
rect 5632 21888 5684 21894
rect 5632 21830 5684 21836
rect 5540 21684 5592 21690
rect 5540 21626 5592 21632
rect 5632 21004 5684 21010
rect 5632 20946 5684 20952
rect 5448 20800 5500 20806
rect 5448 20742 5500 20748
rect 5644 19961 5672 20946
rect 5630 19952 5686 19961
rect 5540 19916 5592 19922
rect 5630 19887 5686 19896
rect 5540 19858 5592 19864
rect 5552 19378 5580 19858
rect 5540 19372 5592 19378
rect 5460 19332 5540 19360
rect 5460 18970 5488 19332
rect 5540 19314 5592 19320
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5448 18692 5500 18698
rect 5448 18634 5500 18640
rect 5460 17678 5488 18634
rect 5644 18426 5672 18770
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 5460 17270 5488 17614
rect 5552 17338 5580 17682
rect 5736 17338 5764 26143
rect 6012 25702 6040 26318
rect 6000 25696 6052 25702
rect 6000 25638 6052 25644
rect 5908 23724 5960 23730
rect 5908 23666 5960 23672
rect 5920 22234 5948 23666
rect 5908 22228 5960 22234
rect 5908 22170 5960 22176
rect 6012 21146 6040 25638
rect 6196 23746 6224 33351
rect 6368 32904 6420 32910
rect 6368 32846 6420 32852
rect 6380 32570 6408 32846
rect 6368 32564 6420 32570
rect 6368 32506 6420 32512
rect 6380 30161 6408 32506
rect 6366 30152 6422 30161
rect 6366 30087 6422 30096
rect 6644 27532 6696 27538
rect 6644 27474 6696 27480
rect 6276 27056 6328 27062
rect 6276 26998 6328 27004
rect 6288 25945 6316 26998
rect 6460 26920 6512 26926
rect 6460 26862 6512 26868
rect 6472 26450 6500 26862
rect 6656 26858 6684 27474
rect 6644 26852 6696 26858
rect 6644 26794 6696 26800
rect 6460 26444 6512 26450
rect 6460 26386 6512 26392
rect 6552 26444 6604 26450
rect 6552 26386 6604 26392
rect 6274 25936 6330 25945
rect 6274 25871 6330 25880
rect 6564 25702 6592 26386
rect 6656 26314 6684 26794
rect 6644 26308 6696 26314
rect 6644 26250 6696 26256
rect 6552 25696 6604 25702
rect 6552 25638 6604 25644
rect 6460 25152 6512 25158
rect 6460 25094 6512 25100
rect 6472 24596 6500 25094
rect 6564 24818 6592 25638
rect 6552 24812 6604 24818
rect 6552 24754 6604 24760
rect 6472 24568 6592 24596
rect 6368 24268 6420 24274
rect 6368 24210 6420 24216
rect 6380 24177 6408 24210
rect 6366 24168 6422 24177
rect 6366 24103 6422 24112
rect 6368 24064 6420 24070
rect 6368 24006 6420 24012
rect 6104 23718 6224 23746
rect 6104 22166 6132 23718
rect 6184 23656 6236 23662
rect 6184 23598 6236 23604
rect 6196 23254 6224 23598
rect 6184 23248 6236 23254
rect 6184 23190 6236 23196
rect 6196 22234 6224 23190
rect 6184 22228 6236 22234
rect 6184 22170 6236 22176
rect 6092 22160 6144 22166
rect 6092 22102 6144 22108
rect 6276 22024 6328 22030
rect 6276 21966 6328 21972
rect 6000 21140 6052 21146
rect 6000 21082 6052 21088
rect 6288 21078 6316 21966
rect 6276 21072 6328 21078
rect 6276 21014 6328 21020
rect 6184 21004 6236 21010
rect 6184 20946 6236 20952
rect 5816 20800 5868 20806
rect 5816 20742 5868 20748
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5448 17264 5500 17270
rect 5448 17206 5500 17212
rect 5448 17128 5500 17134
rect 5500 17088 5580 17116
rect 5448 17070 5500 17076
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5446 16688 5502 16697
rect 5172 16652 5224 16658
rect 5172 16594 5224 16600
rect 5356 16652 5408 16658
rect 5446 16623 5502 16632
rect 5356 16594 5408 16600
rect 5368 16250 5396 16594
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 5080 16176 5132 16182
rect 5080 16118 5132 16124
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5080 15496 5132 15502
rect 5080 15438 5132 15444
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 4894 14376 4950 14385
rect 4894 14311 4896 14320
rect 4948 14311 4950 14320
rect 4896 14282 4948 14288
rect 5000 13297 5028 15302
rect 5092 14958 5120 15438
rect 5276 15314 5304 16050
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5368 15706 5396 15982
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5460 15434 5488 16623
rect 5552 15638 5580 17088
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 5644 15978 5672 16594
rect 5724 16176 5776 16182
rect 5724 16118 5776 16124
rect 5736 16046 5764 16118
rect 5724 16040 5776 16046
rect 5724 15982 5776 15988
rect 5632 15972 5684 15978
rect 5632 15914 5684 15920
rect 5540 15632 5592 15638
rect 5540 15574 5592 15580
rect 5448 15428 5500 15434
rect 5448 15370 5500 15376
rect 5276 15286 5580 15314
rect 5446 15192 5502 15201
rect 5446 15127 5502 15136
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 5262 14784 5318 14793
rect 5262 14719 5318 14728
rect 5276 13530 5304 14719
rect 5354 14648 5410 14657
rect 5354 14583 5356 14592
rect 5408 14583 5410 14592
rect 5356 14554 5408 14560
rect 5460 14074 5488 15127
rect 5552 14346 5580 15286
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5644 13530 5672 15914
rect 5828 15570 5856 20742
rect 6090 20632 6146 20641
rect 6090 20567 6092 20576
rect 6144 20567 6146 20576
rect 6092 20538 6144 20544
rect 6196 20097 6224 20946
rect 6182 20088 6238 20097
rect 6182 20023 6184 20032
rect 6236 20023 6238 20032
rect 6184 19994 6236 20000
rect 5908 19984 5960 19990
rect 5908 19926 5960 19932
rect 5920 18426 5948 19926
rect 6184 19916 6236 19922
rect 6184 19858 6236 19864
rect 6196 18970 6224 19858
rect 6184 18964 6236 18970
rect 6184 18906 6236 18912
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 5906 17776 5962 17785
rect 5906 17711 5908 17720
rect 5960 17711 5962 17720
rect 5908 17682 5960 17688
rect 6012 17626 6040 18022
rect 5920 17598 6040 17626
rect 5920 15638 5948 17598
rect 6000 17264 6052 17270
rect 6000 17206 6052 17212
rect 6274 17232 6330 17241
rect 5908 15632 5960 15638
rect 5908 15574 5960 15580
rect 5816 15564 5868 15570
rect 5816 15506 5868 15512
rect 5724 15496 5776 15502
rect 5724 15438 5776 15444
rect 5736 14278 5764 15438
rect 5828 15162 5856 15506
rect 5816 15156 5868 15162
rect 5816 15098 5868 15104
rect 5920 14822 5948 15574
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 5814 14648 5870 14657
rect 5814 14583 5870 14592
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5736 13569 5764 14214
rect 5722 13560 5778 13569
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5632 13524 5684 13530
rect 5722 13495 5778 13504
rect 5632 13466 5684 13472
rect 5262 13424 5318 13433
rect 5262 13359 5318 13368
rect 5724 13388 5776 13394
rect 4986 13288 5042 13297
rect 4986 13223 5042 13232
rect 5080 13252 5132 13258
rect 5080 13194 5132 13200
rect 4896 13184 4948 13190
rect 4896 13126 4948 13132
rect 4908 13025 4936 13126
rect 4894 13016 4950 13025
rect 4894 12951 4950 12960
rect 5092 12102 5120 13194
rect 5276 12442 5304 13359
rect 5724 13330 5776 13336
rect 5736 13161 5764 13330
rect 5722 13152 5778 13161
rect 5722 13087 5778 13096
rect 5736 12918 5764 13087
rect 5724 12912 5776 12918
rect 5724 12854 5776 12860
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5552 12442 5580 12582
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5828 12374 5856 14583
rect 5920 13394 5948 14758
rect 5908 13388 5960 13394
rect 5908 13330 5960 13336
rect 5816 12368 5868 12374
rect 6012 12345 6040 17206
rect 6274 17167 6276 17176
rect 6328 17167 6330 17176
rect 6276 17138 6328 17144
rect 6276 16040 6328 16046
rect 6276 15982 6328 15988
rect 6090 15600 6146 15609
rect 6090 15535 6146 15544
rect 6184 15564 6236 15570
rect 6104 14618 6132 15535
rect 6184 15506 6236 15512
rect 6196 14822 6224 15506
rect 6288 15366 6316 15982
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6092 14612 6144 14618
rect 6092 14554 6144 14560
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 6196 12986 6224 13330
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 5816 12310 5868 12316
rect 5998 12336 6054 12345
rect 5998 12271 6054 12280
rect 5080 12096 5132 12102
rect 5080 12038 5132 12044
rect 5080 11620 5132 11626
rect 5080 11562 5132 11568
rect 5092 11218 5120 11562
rect 6196 11529 6224 12922
rect 6288 12238 6316 15302
rect 6380 12458 6408 24006
rect 6460 23520 6512 23526
rect 6460 23462 6512 23468
rect 6472 23322 6500 23462
rect 6460 23316 6512 23322
rect 6460 23258 6512 23264
rect 6564 23186 6592 24568
rect 6644 23248 6696 23254
rect 6644 23190 6696 23196
rect 6552 23180 6604 23186
rect 6552 23122 6604 23128
rect 6564 22438 6592 23122
rect 6656 23089 6684 23190
rect 6642 23080 6698 23089
rect 6642 23015 6698 23024
rect 6644 22568 6696 22574
rect 6644 22510 6696 22516
rect 6552 22432 6604 22438
rect 6552 22374 6604 22380
rect 6460 22092 6512 22098
rect 6460 22034 6512 22040
rect 6472 21690 6500 22034
rect 6460 21684 6512 21690
rect 6460 21626 6512 21632
rect 6460 19780 6512 19786
rect 6460 19722 6512 19728
rect 6472 19378 6500 19722
rect 6460 19372 6512 19378
rect 6460 19314 6512 19320
rect 6472 18970 6500 19314
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 6564 18698 6592 22374
rect 6656 21350 6684 22510
rect 6644 21344 6696 21350
rect 6644 21286 6696 21292
rect 6552 18692 6604 18698
rect 6552 18634 6604 18640
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 6472 18086 6500 18566
rect 6460 18080 6512 18086
rect 6460 18022 6512 18028
rect 6644 17740 6696 17746
rect 6644 17682 6696 17688
rect 6656 16998 6684 17682
rect 6748 17270 6776 38490
rect 7024 38010 7052 40190
rect 7392 38434 7420 40996
rect 7852 38457 7880 40996
rect 8772 40882 8800 40996
rect 8404 40854 8800 40882
rect 7116 38406 7420 38434
rect 7838 38448 7894 38457
rect 7012 38004 7064 38010
rect 7012 37946 7064 37952
rect 6826 37224 6882 37233
rect 6826 37159 6882 37168
rect 6840 36689 6868 37159
rect 7012 37120 7064 37126
rect 7012 37062 7064 37068
rect 6826 36680 6882 36689
rect 6826 36615 6882 36624
rect 6920 36032 6972 36038
rect 6920 35974 6972 35980
rect 6932 35154 6960 35974
rect 6920 35148 6972 35154
rect 6920 35090 6972 35096
rect 6932 34746 6960 35090
rect 6920 34740 6972 34746
rect 6920 34682 6972 34688
rect 6918 33552 6974 33561
rect 6918 33487 6974 33496
rect 6932 33289 6960 33487
rect 7024 33425 7052 37062
rect 7010 33416 7066 33425
rect 7010 33351 7066 33360
rect 7116 33289 7144 38406
rect 7838 38383 7894 38392
rect 7656 38344 7708 38350
rect 7656 38286 7708 38292
rect 7380 38208 7432 38214
rect 7380 38150 7432 38156
rect 7392 37806 7420 38150
rect 7380 37800 7432 37806
rect 7380 37742 7432 37748
rect 7392 37505 7420 37742
rect 7378 37496 7434 37505
rect 7378 37431 7434 37440
rect 7392 35086 7420 37431
rect 7380 35080 7432 35086
rect 7380 35022 7432 35028
rect 7392 34746 7420 35022
rect 7380 34740 7432 34746
rect 7380 34682 7432 34688
rect 6918 33280 6974 33289
rect 6918 33215 6974 33224
rect 7102 33280 7158 33289
rect 7102 33215 7158 33224
rect 7668 31260 7696 38286
rect 8404 35737 8432 40854
rect 8852 39364 8904 39370
rect 8852 39306 8904 39312
rect 8864 39098 8892 39306
rect 8852 39092 8904 39098
rect 8852 39034 8904 39040
rect 9036 37732 9088 37738
rect 9036 37674 9088 37680
rect 8390 35728 8446 35737
rect 8390 35663 8446 35672
rect 9048 34513 9076 37674
rect 9232 37369 9260 40996
rect 9692 39098 9720 40996
rect 9680 39092 9732 39098
rect 9680 39034 9732 39040
rect 9680 38888 9732 38894
rect 9680 38830 9732 38836
rect 9692 38214 9720 38830
rect 10612 38457 10640 40996
rect 10598 38448 10654 38457
rect 10598 38383 10654 38392
rect 9680 38208 9732 38214
rect 9680 38150 9732 38156
rect 9692 37505 9720 38150
rect 9954 38040 10010 38049
rect 9954 37975 10010 37984
rect 9678 37496 9734 37505
rect 9678 37431 9734 37440
rect 9218 37360 9274 37369
rect 9692 37330 9720 37431
rect 9968 37330 9996 37975
rect 10416 37664 10468 37670
rect 10416 37606 10468 37612
rect 10968 37664 11020 37670
rect 10968 37606 11020 37612
rect 10428 37369 10456 37606
rect 10414 37360 10470 37369
rect 9218 37295 9274 37304
rect 9680 37324 9732 37330
rect 9680 37266 9732 37272
rect 9956 37324 10008 37330
rect 10414 37295 10470 37304
rect 9956 37266 10008 37272
rect 9968 36922 9996 37266
rect 10048 37256 10100 37262
rect 10048 37198 10100 37204
rect 10060 36922 10088 37198
rect 9956 36916 10008 36922
rect 9956 36858 10008 36864
rect 10048 36916 10100 36922
rect 10048 36858 10100 36864
rect 10060 36378 10088 36858
rect 10980 36553 11008 37606
rect 11072 36922 11100 40996
rect 11428 39296 11480 39302
rect 11428 39238 11480 39244
rect 11440 39098 11468 39238
rect 11428 39092 11480 39098
rect 11428 39034 11480 39040
rect 11532 37913 11560 40996
rect 11704 38344 11756 38350
rect 11704 38286 11756 38292
rect 11888 38344 11940 38350
rect 11888 38286 11940 38292
rect 11518 37904 11574 37913
rect 11518 37839 11574 37848
rect 11716 37670 11744 38286
rect 11900 38010 11928 38286
rect 11888 38004 11940 38010
rect 11888 37946 11940 37952
rect 11704 37664 11756 37670
rect 11704 37606 11756 37612
rect 12164 37664 12216 37670
rect 12164 37606 12216 37612
rect 12176 37262 12204 37606
rect 12452 37482 12480 40996
rect 12912 38962 12940 40996
rect 12900 38956 12952 38962
rect 12900 38898 12952 38904
rect 13360 38888 13412 38894
rect 13360 38830 13412 38836
rect 13636 38888 13688 38894
rect 13636 38830 13688 38836
rect 13372 38554 13400 38830
rect 13648 38554 13676 38830
rect 13360 38548 13412 38554
rect 13360 38490 13412 38496
rect 13636 38548 13688 38554
rect 13636 38490 13688 38496
rect 13358 38448 13414 38457
rect 13358 38383 13360 38392
rect 13412 38383 13414 38392
rect 13360 38354 13412 38360
rect 13634 37768 13690 37777
rect 13634 37703 13690 37712
rect 12452 37454 12572 37482
rect 12360 37330 12480 37346
rect 12360 37324 12492 37330
rect 12360 37318 12440 37324
rect 12164 37256 12216 37262
rect 12164 37198 12216 37204
rect 11244 37120 11296 37126
rect 11244 37062 11296 37068
rect 11060 36916 11112 36922
rect 11060 36858 11112 36864
rect 10966 36544 11022 36553
rect 10966 36479 11022 36488
rect 10048 36372 10100 36378
rect 10048 36314 10100 36320
rect 9772 34944 9824 34950
rect 9772 34886 9824 34892
rect 9034 34504 9090 34513
rect 9034 34439 9090 34448
rect 7932 32768 7984 32774
rect 7932 32710 7984 32716
rect 7944 31929 7972 32710
rect 7930 31920 7986 31929
rect 7930 31855 7986 31864
rect 7748 31408 7800 31414
rect 7746 31376 7748 31385
rect 7800 31376 7802 31385
rect 7746 31311 7802 31320
rect 7668 31232 7788 31260
rect 6920 30592 6972 30598
rect 6920 30534 6972 30540
rect 6932 30297 6960 30534
rect 6918 30288 6974 30297
rect 6918 30223 6920 30232
rect 6972 30223 6974 30232
rect 7378 30288 7434 30297
rect 7378 30223 7434 30232
rect 6920 30194 6972 30200
rect 6932 30163 6960 30194
rect 7392 30190 7420 30223
rect 7380 30184 7432 30190
rect 7380 30126 7432 30132
rect 7104 30116 7156 30122
rect 7104 30058 7156 30064
rect 7012 28620 7064 28626
rect 7012 28562 7064 28568
rect 7024 28218 7052 28562
rect 7116 28558 7144 30058
rect 7392 29850 7420 30126
rect 7380 29844 7432 29850
rect 7380 29786 7432 29792
rect 7564 29708 7616 29714
rect 7564 29650 7616 29656
rect 7196 29640 7248 29646
rect 7196 29582 7248 29588
rect 7208 29034 7236 29582
rect 7576 29034 7604 29650
rect 7196 29028 7248 29034
rect 7196 28970 7248 28976
rect 7564 29028 7616 29034
rect 7564 28970 7616 28976
rect 7104 28552 7156 28558
rect 7104 28494 7156 28500
rect 7012 28212 7064 28218
rect 7012 28154 7064 28160
rect 7116 28150 7144 28494
rect 7104 28144 7156 28150
rect 7104 28086 7156 28092
rect 7104 27124 7156 27130
rect 7104 27066 7156 27072
rect 7010 26752 7066 26761
rect 7010 26687 7066 26696
rect 7024 25906 7052 26687
rect 7116 26586 7144 27066
rect 7104 26580 7156 26586
rect 7104 26522 7156 26528
rect 7116 25906 7144 26522
rect 7208 26217 7236 28970
rect 7472 28008 7524 28014
rect 7472 27950 7524 27956
rect 7484 27674 7512 27950
rect 7472 27668 7524 27674
rect 7472 27610 7524 27616
rect 7380 26784 7432 26790
rect 7380 26726 7432 26732
rect 7194 26208 7250 26217
rect 7194 26143 7250 26152
rect 7012 25900 7064 25906
rect 7012 25842 7064 25848
rect 7104 25900 7156 25906
rect 7104 25842 7156 25848
rect 7194 25800 7250 25809
rect 7194 25735 7250 25744
rect 7104 25492 7156 25498
rect 7104 25434 7156 25440
rect 7012 25220 7064 25226
rect 7012 25162 7064 25168
rect 6920 25152 6972 25158
rect 6920 25094 6972 25100
rect 6932 24954 6960 25094
rect 6920 24948 6972 24954
rect 6920 24890 6972 24896
rect 7024 24750 7052 25162
rect 7012 24744 7064 24750
rect 7012 24686 7064 24692
rect 6920 24608 6972 24614
rect 6920 24550 6972 24556
rect 6932 22964 6960 24550
rect 7010 24168 7066 24177
rect 7010 24103 7066 24112
rect 7024 23254 7052 24103
rect 7116 23526 7144 25434
rect 7208 25430 7236 25735
rect 7196 25424 7248 25430
rect 7196 25366 7248 25372
rect 7196 25288 7248 25294
rect 7196 25230 7248 25236
rect 7208 24682 7236 25230
rect 7288 24744 7340 24750
rect 7288 24686 7340 24692
rect 7196 24676 7248 24682
rect 7196 24618 7248 24624
rect 7208 24138 7236 24618
rect 7300 24274 7328 24686
rect 7288 24268 7340 24274
rect 7288 24210 7340 24216
rect 7196 24132 7248 24138
rect 7196 24074 7248 24080
rect 7196 23588 7248 23594
rect 7196 23530 7248 23536
rect 7104 23520 7156 23526
rect 7208 23497 7236 23530
rect 7104 23462 7156 23468
rect 7194 23488 7250 23497
rect 7194 23423 7250 23432
rect 7012 23248 7064 23254
rect 7012 23190 7064 23196
rect 7104 22976 7156 22982
rect 6932 22936 7104 22964
rect 7104 22918 7156 22924
rect 6920 22704 6972 22710
rect 6840 22652 6920 22658
rect 6840 22646 6972 22652
rect 6840 22630 6960 22646
rect 7116 22642 7144 22918
rect 7104 22636 7156 22642
rect 6840 22098 6868 22630
rect 7104 22578 7156 22584
rect 7116 22273 7144 22578
rect 7208 22545 7236 23423
rect 7288 23112 7340 23118
rect 7288 23054 7340 23060
rect 7194 22536 7250 22545
rect 7300 22506 7328 23054
rect 7194 22471 7250 22480
rect 7288 22500 7340 22506
rect 7288 22442 7340 22448
rect 7102 22264 7158 22273
rect 7300 22234 7328 22442
rect 7102 22199 7158 22208
rect 7288 22228 7340 22234
rect 7288 22170 7340 22176
rect 6828 22092 6880 22098
rect 6828 22034 6880 22040
rect 7012 22092 7064 22098
rect 7012 22034 7064 22040
rect 6920 21480 6972 21486
rect 6920 21422 6972 21428
rect 6932 21146 6960 21422
rect 6920 21140 6972 21146
rect 6920 21082 6972 21088
rect 6932 20602 6960 21082
rect 7024 20874 7052 22034
rect 7392 22030 7420 26726
rect 7472 26444 7524 26450
rect 7472 26386 7524 26392
rect 7484 25838 7512 26386
rect 7472 25832 7524 25838
rect 7472 25774 7524 25780
rect 7576 24449 7604 28970
rect 7760 28966 7788 31232
rect 7840 29572 7892 29578
rect 7840 29514 7892 29520
rect 7748 28960 7800 28966
rect 7748 28902 7800 28908
rect 7852 28626 7880 29514
rect 7840 28620 7892 28626
rect 7840 28562 7892 28568
rect 7656 27872 7708 27878
rect 7656 27814 7708 27820
rect 7668 26450 7696 27814
rect 7656 26444 7708 26450
rect 7656 26386 7708 26392
rect 7748 26240 7800 26246
rect 7748 26182 7800 26188
rect 7760 25838 7788 26182
rect 7748 25832 7800 25838
rect 7748 25774 7800 25780
rect 7562 24440 7618 24449
rect 7760 24410 7788 25774
rect 7840 25220 7892 25226
rect 7840 25162 7892 25168
rect 7852 24614 7880 25162
rect 7840 24608 7892 24614
rect 7840 24550 7892 24556
rect 7562 24375 7618 24384
rect 7748 24404 7800 24410
rect 7748 24346 7800 24352
rect 7472 24268 7524 24274
rect 7472 24210 7524 24216
rect 7564 24268 7616 24274
rect 7564 24210 7616 24216
rect 7484 23746 7512 24210
rect 7576 23848 7604 24210
rect 7576 23820 7696 23848
rect 7562 23760 7618 23769
rect 7484 23718 7562 23746
rect 7562 23695 7564 23704
rect 7616 23695 7618 23704
rect 7564 23666 7616 23672
rect 7472 23656 7524 23662
rect 7472 23598 7524 23604
rect 7380 22024 7432 22030
rect 7380 21966 7432 21972
rect 7196 21888 7248 21894
rect 7196 21830 7248 21836
rect 7208 21554 7236 21830
rect 7104 21548 7156 21554
rect 7104 21490 7156 21496
rect 7196 21548 7248 21554
rect 7196 21490 7248 21496
rect 7116 20942 7144 21490
rect 7104 20936 7156 20942
rect 7104 20878 7156 20884
rect 7012 20868 7064 20874
rect 7012 20810 7064 20816
rect 7116 20602 7144 20878
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 7104 20596 7156 20602
rect 7104 20538 7156 20544
rect 6932 20398 6960 20538
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 6932 20058 6960 20334
rect 7116 20330 7144 20538
rect 7104 20324 7156 20330
rect 7104 20266 7156 20272
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 6932 18970 6960 19994
rect 7208 19718 7236 21490
rect 7392 21486 7420 21966
rect 7380 21480 7432 21486
rect 7380 21422 7432 21428
rect 7288 20800 7340 20806
rect 7392 20777 7420 21422
rect 7288 20742 7340 20748
rect 7378 20768 7434 20777
rect 7300 20330 7328 20742
rect 7378 20703 7434 20712
rect 7484 20398 7512 23598
rect 7668 23361 7696 23820
rect 7654 23352 7710 23361
rect 7654 23287 7710 23296
rect 7564 23248 7616 23254
rect 7564 23190 7616 23196
rect 7576 22438 7604 23190
rect 7564 22432 7616 22438
rect 7562 22400 7564 22409
rect 7616 22400 7618 22409
rect 7562 22335 7618 22344
rect 7668 22030 7696 23287
rect 7852 22506 7880 24550
rect 7840 22500 7892 22506
rect 7840 22442 7892 22448
rect 7656 22024 7708 22030
rect 7656 21966 7708 21972
rect 7564 21888 7616 21894
rect 7564 21830 7616 21836
rect 7576 21418 7604 21830
rect 7748 21548 7800 21554
rect 7944 21536 7972 31855
rect 8024 30184 8076 30190
rect 8024 30126 8076 30132
rect 8574 30152 8630 30161
rect 8036 30025 8064 30126
rect 8574 30087 8630 30096
rect 8588 30054 8616 30087
rect 8576 30048 8628 30054
rect 8022 30016 8078 30025
rect 8576 29990 8628 29996
rect 8022 29951 8078 29960
rect 8036 29714 8064 29951
rect 8024 29708 8076 29714
rect 8024 29650 8076 29656
rect 8036 29306 8064 29650
rect 8588 29510 8616 29990
rect 8576 29504 8628 29510
rect 8576 29446 8628 29452
rect 8024 29300 8076 29306
rect 8024 29242 8076 29248
rect 8588 29102 8616 29446
rect 8576 29096 8628 29102
rect 8576 29038 8628 29044
rect 8944 29096 8996 29102
rect 8944 29038 8996 29044
rect 8666 28656 8722 28665
rect 8666 28591 8668 28600
rect 8720 28591 8722 28600
rect 8668 28562 8720 28568
rect 8024 28552 8076 28558
rect 8024 28494 8076 28500
rect 8036 28014 8064 28494
rect 8680 28218 8708 28562
rect 8668 28212 8720 28218
rect 8668 28154 8720 28160
rect 8956 28082 8984 29038
rect 9048 28422 9076 34439
rect 9784 34066 9812 34886
rect 9772 34060 9824 34066
rect 9772 34002 9824 34008
rect 9784 33658 9812 34002
rect 10060 33998 10088 36314
rect 10600 36236 10652 36242
rect 10600 36178 10652 36184
rect 10612 35834 10640 36178
rect 10600 35828 10652 35834
rect 10600 35770 10652 35776
rect 10612 35290 10640 35770
rect 10600 35284 10652 35290
rect 10600 35226 10652 35232
rect 11060 34740 11112 34746
rect 11060 34682 11112 34688
rect 10048 33992 10100 33998
rect 10048 33934 10100 33940
rect 10060 33658 10088 33934
rect 9772 33652 9824 33658
rect 9772 33594 9824 33600
rect 10048 33652 10100 33658
rect 10048 33594 10100 33600
rect 11072 33130 11100 34682
rect 10980 33114 11100 33130
rect 10968 33108 11100 33114
rect 11020 33102 11100 33108
rect 10968 33050 11020 33056
rect 10874 32192 10930 32201
rect 10874 32127 10930 32136
rect 10324 31136 10376 31142
rect 10324 31078 10376 31084
rect 9586 30696 9642 30705
rect 9586 30631 9588 30640
rect 9640 30631 9642 30640
rect 9588 30602 9640 30608
rect 9954 30424 10010 30433
rect 10336 30394 10364 31078
rect 10416 30592 10468 30598
rect 10416 30534 10468 30540
rect 9954 30359 10010 30368
rect 10324 30388 10376 30394
rect 9680 30320 9732 30326
rect 9678 30288 9680 30297
rect 9732 30288 9734 30297
rect 9678 30223 9734 30232
rect 9588 28960 9640 28966
rect 9588 28902 9640 28908
rect 9036 28416 9088 28422
rect 9036 28358 9088 28364
rect 9404 28416 9456 28422
rect 9404 28358 9456 28364
rect 8944 28076 8996 28082
rect 8944 28018 8996 28024
rect 8024 28008 8076 28014
rect 8024 27950 8076 27956
rect 8852 28008 8904 28014
rect 8852 27950 8904 27956
rect 8392 27872 8444 27878
rect 8392 27814 8444 27820
rect 8024 27532 8076 27538
rect 8024 27474 8076 27480
rect 8116 27532 8168 27538
rect 8116 27474 8168 27480
rect 8036 26586 8064 27474
rect 8128 27062 8156 27474
rect 8208 27328 8260 27334
rect 8208 27270 8260 27276
rect 8116 27056 8168 27062
rect 8114 27024 8116 27033
rect 8168 27024 8170 27033
rect 8114 26959 8170 26968
rect 8024 26580 8076 26586
rect 8024 26522 8076 26528
rect 8220 25906 8248 27270
rect 8404 26081 8432 27814
rect 8864 27674 8892 27950
rect 8852 27668 8904 27674
rect 8852 27610 8904 27616
rect 9312 27328 9364 27334
rect 9312 27270 9364 27276
rect 8852 26920 8904 26926
rect 8852 26862 8904 26868
rect 9128 26920 9180 26926
rect 9128 26862 9180 26868
rect 8864 26314 8892 26862
rect 9140 26382 9168 26862
rect 9128 26376 9180 26382
rect 9126 26344 9128 26353
rect 9180 26344 9182 26353
rect 8484 26308 8536 26314
rect 8484 26250 8536 26256
rect 8852 26308 8904 26314
rect 9126 26279 9182 26288
rect 8852 26250 8904 26256
rect 8390 26072 8446 26081
rect 8390 26007 8446 26016
rect 8208 25900 8260 25906
rect 8208 25842 8260 25848
rect 8208 25696 8260 25702
rect 8206 25664 8208 25673
rect 8260 25664 8262 25673
rect 8206 25599 8262 25608
rect 8116 25356 8168 25362
rect 8116 25298 8168 25304
rect 8128 24886 8156 25298
rect 8404 25294 8432 26007
rect 8392 25288 8444 25294
rect 8392 25230 8444 25236
rect 8116 24880 8168 24886
rect 8116 24822 8168 24828
rect 8208 24744 8260 24750
rect 8208 24686 8260 24692
rect 8220 24562 8248 24686
rect 8220 24534 8340 24562
rect 8024 23520 8076 23526
rect 8024 23462 8076 23468
rect 8036 23118 8064 23462
rect 8312 23322 8340 24534
rect 8392 23520 8444 23526
rect 8392 23462 8444 23468
rect 8300 23316 8352 23322
rect 8300 23258 8352 23264
rect 8404 23202 8432 23462
rect 8220 23186 8432 23202
rect 8208 23180 8432 23186
rect 8260 23174 8432 23180
rect 8208 23122 8260 23128
rect 8024 23112 8076 23118
rect 8024 23054 8076 23060
rect 8036 22642 8064 23054
rect 8220 22710 8248 23122
rect 8208 22704 8260 22710
rect 8208 22646 8260 22652
rect 8024 22636 8076 22642
rect 8024 22578 8076 22584
rect 8036 22166 8064 22578
rect 8300 22500 8352 22506
rect 8300 22442 8352 22448
rect 8024 22160 8076 22166
rect 8024 22102 8076 22108
rect 8208 22092 8260 22098
rect 8312 22080 8340 22442
rect 8260 22052 8340 22080
rect 8208 22034 8260 22040
rect 7748 21490 7800 21496
rect 7852 21508 7972 21536
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 7576 21146 7604 21354
rect 7564 21140 7616 21146
rect 7564 21082 7616 21088
rect 7656 21004 7708 21010
rect 7656 20946 7708 20952
rect 7472 20392 7524 20398
rect 7472 20334 7524 20340
rect 7288 20324 7340 20330
rect 7288 20266 7340 20272
rect 7300 19854 7328 20266
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7392 20097 7420 20198
rect 7378 20088 7434 20097
rect 7378 20023 7434 20032
rect 7380 19984 7432 19990
rect 7484 19972 7512 20334
rect 7668 20262 7696 20946
rect 7656 20256 7708 20262
rect 7656 20198 7708 20204
rect 7432 19944 7512 19972
rect 7380 19926 7432 19932
rect 7288 19848 7340 19854
rect 7288 19790 7340 19796
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7208 19360 7236 19654
rect 7116 19332 7236 19360
rect 7116 19174 7144 19332
rect 7300 19310 7328 19790
rect 7288 19304 7340 19310
rect 7194 19272 7250 19281
rect 7288 19246 7340 19252
rect 7194 19207 7196 19216
rect 7248 19207 7250 19216
rect 7196 19178 7248 19184
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 7104 19168 7156 19174
rect 7104 19110 7156 19116
rect 6920 18964 6972 18970
rect 6920 18906 6972 18912
rect 7024 18834 7052 19110
rect 7012 18828 7064 18834
rect 7012 18770 7064 18776
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 6932 18170 6960 18294
rect 7024 18290 7052 18770
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 6932 18142 7052 18170
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6932 17678 6960 18022
rect 7024 17882 7052 18142
rect 7012 17876 7064 17882
rect 7012 17818 7064 17824
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6736 17264 6788 17270
rect 6736 17206 6788 17212
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6826 16960 6882 16969
rect 6656 16658 6684 16934
rect 6826 16895 6882 16904
rect 6644 16652 6696 16658
rect 6644 16594 6696 16600
rect 6656 16250 6684 16594
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6656 16046 6684 16186
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 6734 16008 6790 16017
rect 6734 15943 6790 15952
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6472 14074 6500 14418
rect 6748 14249 6776 15943
rect 6840 15910 6868 16895
rect 6932 16046 6960 17614
rect 7116 17202 7144 19110
rect 7392 18834 7420 19926
rect 7564 19916 7616 19922
rect 7668 19904 7696 20198
rect 7616 19876 7696 19904
rect 7564 19858 7616 19864
rect 7472 18896 7524 18902
rect 7472 18838 7524 18844
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 7194 18728 7250 18737
rect 7194 18663 7196 18672
rect 7248 18663 7250 18672
rect 7196 18634 7248 18640
rect 7208 18222 7236 18634
rect 7196 18216 7248 18222
rect 7196 18158 7248 18164
rect 7392 17882 7420 18770
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7484 17542 7512 18838
rect 7576 18630 7604 19858
rect 7654 19136 7710 19145
rect 7654 19071 7710 19080
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7104 17196 7156 17202
rect 7104 17138 7156 17144
rect 7116 16794 7144 17138
rect 7484 17134 7512 17478
rect 7668 17184 7696 19071
rect 7760 18465 7788 21490
rect 7852 21185 7880 21508
rect 7930 21448 7986 21457
rect 7930 21383 7986 21392
rect 7838 21176 7894 21185
rect 7838 21111 7894 21120
rect 7852 20330 7880 21111
rect 7944 20466 7972 21383
rect 8024 21344 8076 21350
rect 8024 21286 8076 21292
rect 8036 21185 8064 21286
rect 8022 21176 8078 21185
rect 8022 21111 8078 21120
rect 7932 20460 7984 20466
rect 7932 20402 7984 20408
rect 7840 20324 7892 20330
rect 7840 20266 7892 20272
rect 7840 20052 7892 20058
rect 7840 19994 7892 20000
rect 7852 19514 7880 19994
rect 7932 19984 7984 19990
rect 7932 19926 7984 19932
rect 7840 19508 7892 19514
rect 7840 19450 7892 19456
rect 7944 19145 7972 19926
rect 7930 19136 7986 19145
rect 7930 19071 7986 19080
rect 7930 18864 7986 18873
rect 7930 18799 7932 18808
rect 7984 18799 7986 18808
rect 7932 18770 7984 18776
rect 7746 18456 7802 18465
rect 7746 18391 7802 18400
rect 7576 17156 7696 17184
rect 7472 17128 7524 17134
rect 7286 17096 7342 17105
rect 7472 17070 7524 17076
rect 7286 17031 7288 17040
rect 7340 17031 7342 17040
rect 7288 17002 7340 17008
rect 7104 16788 7156 16794
rect 7104 16730 7156 16736
rect 7300 16726 7328 17002
rect 7484 16726 7512 17070
rect 7288 16720 7340 16726
rect 7472 16720 7524 16726
rect 7288 16662 7340 16668
rect 7470 16688 7472 16697
rect 7524 16688 7526 16697
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6932 15706 6960 15982
rect 7196 15972 7248 15978
rect 7196 15914 7248 15920
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 6828 15428 6880 15434
rect 6828 15370 6880 15376
rect 6840 14657 6868 15370
rect 6826 14648 6882 14657
rect 6826 14583 6882 14592
rect 6734 14240 6790 14249
rect 6734 14175 6790 14184
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 6932 14006 6960 15642
rect 7102 15600 7158 15609
rect 7102 15535 7104 15544
rect 7156 15535 7158 15544
rect 7104 15506 7156 15512
rect 7208 15337 7236 15914
rect 7300 15910 7328 16662
rect 7470 16623 7526 16632
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7194 15328 7250 15337
rect 7194 15263 7250 15272
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6472 12918 6500 13330
rect 6460 12912 6512 12918
rect 6460 12854 6512 12860
rect 6380 12430 6592 12458
rect 6840 12442 6868 13806
rect 6932 13530 6960 13942
rect 7024 13870 7052 14758
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 7024 13462 7052 13806
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 6918 12880 6974 12889
rect 6918 12815 6920 12824
rect 6972 12815 6974 12824
rect 6920 12786 6972 12792
rect 7024 12646 7052 13398
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 6564 12374 6592 12430
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6288 11898 6316 12174
rect 6460 12164 6512 12170
rect 6460 12106 6512 12112
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6472 11558 6500 12106
rect 6564 11830 6592 12310
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6840 12209 6868 12242
rect 6826 12200 6882 12209
rect 6826 12135 6882 12144
rect 6552 11824 6604 11830
rect 6552 11766 6604 11772
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6460 11552 6512 11558
rect 6182 11520 6238 11529
rect 6460 11494 6512 11500
rect 6182 11455 6238 11464
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 4672 11104 4752 11132
rect 4620 11086 4672 11092
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 4080 11070 4200 11086
rect 3988 10470 4016 11018
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3790 9480 3846 9489
rect 3790 9415 3846 9424
rect 3606 8392 3662 8401
rect 3606 8327 3662 8336
rect 3514 7984 3570 7993
rect 3514 7919 3570 7928
rect 3528 4185 3556 7919
rect 3790 7168 3846 7177
rect 3790 7103 3846 7112
rect 3514 4176 3570 4185
rect 3514 4111 3570 4120
rect 3148 3528 3200 3534
rect 3146 3496 3148 3505
rect 3424 3528 3476 3534
rect 3200 3496 3202 3505
rect 3424 3470 3476 3476
rect 3146 3431 3202 3440
rect 3436 3194 3464 3470
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3436 2854 3464 3130
rect 2884 2774 3004 2802
rect 3424 2848 3476 2854
rect 3804 2825 3832 7103
rect 3424 2790 3476 2796
rect 3790 2816 3846 2825
rect 2884 2666 2912 2774
rect 2792 2638 2912 2666
rect 3436 2650 3464 2790
rect 3790 2751 3846 2760
rect 3424 2644 3476 2650
rect 2792 800 2820 2638
rect 3424 2586 3476 2592
rect 3700 2304 3752 2310
rect 3700 2246 3752 2252
rect 3712 800 3740 2246
rect 3896 1601 3924 9658
rect 4080 5692 4108 11070
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4632 10742 4660 11086
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 4724 10606 4752 10950
rect 4816 10810 4844 11154
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4632 10062 4660 10406
rect 4724 10198 4752 10542
rect 5092 10266 5120 11154
rect 5460 10962 5488 11154
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 5632 11008 5684 11014
rect 5460 10956 5632 10962
rect 5460 10950 5684 10956
rect 5460 10934 5672 10950
rect 6288 10470 6316 11086
rect 6472 11082 6500 11494
rect 6656 11354 6684 11630
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6564 10470 6592 10950
rect 6656 10849 6684 11290
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6642 10840 6698 10849
rect 6642 10775 6698 10784
rect 6748 10606 6776 11154
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 4712 10192 4764 10198
rect 4712 10134 4764 10140
rect 5538 10160 5594 10169
rect 5538 10095 5540 10104
rect 5592 10095 5594 10104
rect 5540 10066 5592 10072
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 5460 9518 5488 9998
rect 5552 9654 5580 10066
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5552 9042 5580 9590
rect 6182 9344 6238 9353
rect 6182 9279 6238 9288
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 6104 8634 6132 8978
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 5538 7712 5594 7721
rect 4220 7644 4516 7664
rect 5538 7647 5594 7656
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4802 7576 4858 7585
rect 4802 7511 4858 7520
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 3988 5664 4108 5692
rect 3988 3641 4016 5664
rect 4066 5536 4122 5545
rect 4066 5471 4122 5480
rect 4080 4593 4108 5471
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4618 4992 4674 5001
rect 4618 4927 4674 4936
rect 4066 4584 4122 4593
rect 4066 4519 4122 4528
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 3974 3632 4030 3641
rect 4632 3602 4660 4927
rect 3974 3567 4030 3576
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 4632 3194 4660 3538
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 4356 2553 4384 2790
rect 4342 2544 4398 2553
rect 4342 2479 4398 2488
rect 4356 2446 4384 2479
rect 4344 2440 4396 2446
rect 4066 2408 4122 2417
rect 4344 2382 4396 2388
rect 4066 2343 4122 2352
rect 3882 1592 3938 1601
rect 3882 1527 3938 1536
rect 4080 1465 4108 2343
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 4066 1456 4122 1465
rect 4632 1442 4660 2994
rect 4066 1391 4122 1400
rect 4172 1414 4660 1442
rect 4172 800 4200 1414
rect 4724 898 4752 3334
rect 4816 3058 4844 7511
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 4632 870 4752 898
rect 4632 800 4660 870
rect 5552 800 5580 7647
rect 5998 5944 6054 5953
rect 5998 5879 6054 5888
rect 6012 800 6040 5879
rect 6196 2582 6224 9279
rect 6288 8945 6316 10406
rect 6564 10062 6592 10406
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6748 9586 6776 10542
rect 6828 10532 6880 10538
rect 6828 10474 6880 10480
rect 6840 10266 6868 10474
rect 6828 10260 6880 10266
rect 6932 10248 6960 11154
rect 6880 10220 6960 10248
rect 6828 10202 6880 10208
rect 7116 10130 7144 14894
rect 7208 14822 7236 14962
rect 7472 14952 7524 14958
rect 7470 14920 7472 14929
rect 7524 14920 7526 14929
rect 7380 14884 7432 14890
rect 7470 14855 7526 14864
rect 7380 14826 7432 14832
rect 7196 14816 7248 14822
rect 7392 14793 7420 14826
rect 7196 14758 7248 14764
rect 7378 14784 7434 14793
rect 7208 14346 7236 14758
rect 7378 14719 7434 14728
rect 7392 14346 7420 14719
rect 7196 14340 7248 14346
rect 7196 14282 7248 14288
rect 7380 14340 7432 14346
rect 7380 14282 7432 14288
rect 7576 14249 7604 17156
rect 7760 17082 7788 18391
rect 8036 18306 8064 21111
rect 8208 21072 8260 21078
rect 8208 21014 8260 21020
rect 8220 20505 8248 21014
rect 8206 20496 8262 20505
rect 8206 20431 8262 20440
rect 8116 18624 8168 18630
rect 8116 18566 8168 18572
rect 7852 18278 8064 18306
rect 7852 17320 7880 18278
rect 7932 18148 7984 18154
rect 7932 18090 7984 18096
rect 7944 17921 7972 18090
rect 7930 17912 7986 17921
rect 7930 17847 7986 17856
rect 8024 17740 8076 17746
rect 8024 17682 8076 17688
rect 8036 17649 8064 17682
rect 8022 17640 8078 17649
rect 8022 17575 8078 17584
rect 8128 17542 8156 18566
rect 8220 18086 8248 20431
rect 8312 20058 8340 22052
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8404 21350 8432 21966
rect 8392 21344 8444 21350
rect 8392 21286 8444 21292
rect 8404 20806 8432 21286
rect 8392 20800 8444 20806
rect 8392 20742 8444 20748
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 8300 19236 8352 19242
rect 8300 19178 8352 19184
rect 8208 18080 8260 18086
rect 8312 18057 8340 19178
rect 8208 18022 8260 18028
rect 8298 18048 8354 18057
rect 8298 17983 8354 17992
rect 8298 17912 8354 17921
rect 8496 17882 8524 26250
rect 8944 26036 8996 26042
rect 8944 25978 8996 25984
rect 8852 25696 8904 25702
rect 8852 25638 8904 25644
rect 8864 25362 8892 25638
rect 8852 25356 8904 25362
rect 8852 25298 8904 25304
rect 8864 24313 8892 25298
rect 8956 24993 8984 25978
rect 9128 25900 9180 25906
rect 9128 25842 9180 25848
rect 8942 24984 8998 24993
rect 8942 24919 8998 24928
rect 8944 24676 8996 24682
rect 8944 24618 8996 24624
rect 8850 24304 8906 24313
rect 8850 24239 8852 24248
rect 8904 24239 8906 24248
rect 8852 24210 8904 24216
rect 8668 24064 8720 24070
rect 8668 24006 8720 24012
rect 8680 23662 8708 24006
rect 8668 23656 8720 23662
rect 8668 23598 8720 23604
rect 8668 23248 8720 23254
rect 8668 23190 8720 23196
rect 8680 21962 8708 23190
rect 8760 22636 8812 22642
rect 8760 22578 8812 22584
rect 8772 22234 8800 22578
rect 8760 22228 8812 22234
rect 8760 22170 8812 22176
rect 8864 22114 8892 24210
rect 8956 24177 8984 24618
rect 8942 24168 8998 24177
rect 8942 24103 8998 24112
rect 9140 23633 9168 25842
rect 9324 24857 9352 27270
rect 9310 24848 9366 24857
rect 9310 24783 9366 24792
rect 8942 23624 8998 23633
rect 8942 23559 8944 23568
rect 8996 23559 8998 23568
rect 9126 23624 9182 23633
rect 9126 23559 9182 23568
rect 8944 23530 8996 23536
rect 8956 22817 8984 23530
rect 8942 22808 8998 22817
rect 8942 22743 8998 22752
rect 9218 22672 9274 22681
rect 9218 22607 9274 22616
rect 9232 22506 9260 22607
rect 9220 22500 9272 22506
rect 9220 22442 9272 22448
rect 9232 22409 9260 22442
rect 9218 22400 9274 22409
rect 9218 22335 9274 22344
rect 9218 22264 9274 22273
rect 9218 22199 9274 22208
rect 8772 22086 8892 22114
rect 9232 22098 9260 22199
rect 9220 22092 9272 22098
rect 8668 21956 8720 21962
rect 8668 21898 8720 21904
rect 8576 21888 8628 21894
rect 8574 21856 8576 21865
rect 8628 21856 8630 21865
rect 8574 21791 8630 21800
rect 8588 21622 8616 21791
rect 8576 21616 8628 21622
rect 8680 21593 8708 21898
rect 8576 21558 8628 21564
rect 8666 21584 8722 21593
rect 8666 21519 8722 21528
rect 8666 20632 8722 20641
rect 8666 20567 8722 20576
rect 8680 20534 8708 20567
rect 8668 20528 8720 20534
rect 8668 20470 8720 20476
rect 8680 19514 8708 20470
rect 8668 19508 8720 19514
rect 8588 19468 8668 19496
rect 8588 18426 8616 19468
rect 8668 19450 8720 19456
rect 8772 18970 8800 22086
rect 9220 22034 9272 22040
rect 9232 22001 9260 22034
rect 9218 21992 9274 22001
rect 9218 21927 9274 21936
rect 9128 21888 9180 21894
rect 9128 21830 9180 21836
rect 8852 21344 8904 21350
rect 8850 21312 8852 21321
rect 8904 21312 8906 21321
rect 8850 21247 8906 21256
rect 9140 20942 9168 21830
rect 9232 21690 9260 21927
rect 9220 21684 9272 21690
rect 9220 21626 9272 21632
rect 9232 21078 9260 21626
rect 9220 21072 9272 21078
rect 9220 21014 9272 21020
rect 9128 20936 9180 20942
rect 9324 20924 9352 24783
rect 9416 24750 9444 28358
rect 9600 26353 9628 28902
rect 9772 28144 9824 28150
rect 9772 28086 9824 28092
rect 9784 28014 9812 28086
rect 9772 28008 9824 28014
rect 9772 27950 9824 27956
rect 9784 27169 9812 27950
rect 9770 27160 9826 27169
rect 9770 27095 9826 27104
rect 9680 26852 9732 26858
rect 9680 26794 9732 26800
rect 9692 26518 9720 26794
rect 9680 26512 9732 26518
rect 9680 26454 9732 26460
rect 9586 26344 9642 26353
rect 9586 26279 9642 26288
rect 9496 25424 9548 25430
rect 9496 25366 9548 25372
rect 9508 24886 9536 25366
rect 9588 25152 9640 25158
rect 9588 25094 9640 25100
rect 9496 24880 9548 24886
rect 9496 24822 9548 24828
rect 9404 24744 9456 24750
rect 9404 24686 9456 24692
rect 9600 23746 9628 25094
rect 9864 24812 9916 24818
rect 9864 24754 9916 24760
rect 9772 24744 9824 24750
rect 9772 24686 9824 24692
rect 9784 24138 9812 24686
rect 9876 24206 9904 24754
rect 9864 24200 9916 24206
rect 9864 24142 9916 24148
rect 9772 24132 9824 24138
rect 9772 24074 9824 24080
rect 9784 23866 9812 24074
rect 9772 23860 9824 23866
rect 9772 23802 9824 23808
rect 9600 23718 9720 23746
rect 9692 23662 9720 23718
rect 9680 23656 9732 23662
rect 9680 23598 9732 23604
rect 9588 23588 9640 23594
rect 9588 23530 9640 23536
rect 9404 22976 9456 22982
rect 9404 22918 9456 22924
rect 9416 22438 9444 22918
rect 9600 22658 9628 23530
rect 9876 23322 9904 24142
rect 9864 23316 9916 23322
rect 9864 23258 9916 23264
rect 9968 23202 9996 30359
rect 10324 30330 10376 30336
rect 10336 30297 10364 30330
rect 10322 30288 10378 30297
rect 10322 30223 10378 30232
rect 10428 30190 10456 30534
rect 10508 30320 10560 30326
rect 10508 30262 10560 30268
rect 10416 30184 10468 30190
rect 10416 30126 10468 30132
rect 10428 29714 10456 30126
rect 10324 29708 10376 29714
rect 10324 29650 10376 29656
rect 10416 29708 10468 29714
rect 10416 29650 10468 29656
rect 10336 29594 10364 29650
rect 10140 29572 10192 29578
rect 10336 29566 10456 29594
rect 10140 29514 10192 29520
rect 10152 29306 10180 29514
rect 10140 29300 10192 29306
rect 10140 29242 10192 29248
rect 10428 29034 10456 29566
rect 10416 29028 10468 29034
rect 10416 28970 10468 28976
rect 10428 28937 10456 28970
rect 10414 28928 10470 28937
rect 10336 28886 10414 28914
rect 10232 28008 10284 28014
rect 10336 27985 10364 28886
rect 10414 28863 10470 28872
rect 10416 28484 10468 28490
rect 10416 28426 10468 28432
rect 10232 27950 10284 27956
rect 10322 27976 10378 27985
rect 10140 26784 10192 26790
rect 10138 26752 10140 26761
rect 10192 26752 10194 26761
rect 10138 26687 10194 26696
rect 10244 26568 10272 27950
rect 10322 27911 10378 27920
rect 10324 27328 10376 27334
rect 10324 27270 10376 27276
rect 10336 27062 10364 27270
rect 10324 27056 10376 27062
rect 10324 26998 10376 27004
rect 10152 26540 10272 26568
rect 10048 26444 10100 26450
rect 10048 26386 10100 26392
rect 10060 25702 10088 26386
rect 10048 25696 10100 25702
rect 10046 25664 10048 25673
rect 10100 25664 10102 25673
rect 10046 25599 10102 25608
rect 10048 24744 10100 24750
rect 10048 24686 10100 24692
rect 10060 24274 10088 24686
rect 10048 24268 10100 24274
rect 10048 24210 10100 24216
rect 9772 23180 9824 23186
rect 9772 23122 9824 23128
rect 9876 23174 9996 23202
rect 9784 22710 9812 23122
rect 9772 22704 9824 22710
rect 9600 22642 9720 22658
rect 9772 22646 9824 22652
rect 9600 22636 9732 22642
rect 9600 22630 9680 22636
rect 9680 22578 9732 22584
rect 9588 22500 9640 22506
rect 9588 22442 9640 22448
rect 9404 22432 9456 22438
rect 9404 22374 9456 22380
rect 9416 22234 9444 22374
rect 9404 22228 9456 22234
rect 9404 22170 9456 22176
rect 9416 21146 9444 22170
rect 9600 22137 9628 22442
rect 9586 22128 9642 22137
rect 9586 22063 9642 22072
rect 9680 22024 9732 22030
rect 9680 21966 9732 21972
rect 9588 21888 9640 21894
rect 9692 21876 9720 21966
rect 9640 21848 9720 21876
rect 9588 21830 9640 21836
rect 9588 21616 9640 21622
rect 9508 21564 9588 21570
rect 9508 21558 9640 21564
rect 9692 21570 9720 21848
rect 9508 21542 9628 21558
rect 9692 21542 9812 21570
rect 9508 21434 9536 21542
rect 9784 21486 9812 21542
rect 9772 21480 9824 21486
rect 9508 21406 9720 21434
rect 9772 21422 9824 21428
rect 9404 21140 9456 21146
rect 9404 21082 9456 21088
rect 9128 20878 9180 20884
rect 9232 20896 9352 20924
rect 9404 20936 9456 20942
rect 9128 20800 9180 20806
rect 9128 20742 9180 20748
rect 9036 20392 9088 20398
rect 9036 20334 9088 20340
rect 9048 19718 9076 20334
rect 9140 20330 9168 20742
rect 9128 20324 9180 20330
rect 9128 20266 9180 20272
rect 9036 19712 9088 19718
rect 9036 19654 9088 19660
rect 8850 19544 8906 19553
rect 8850 19479 8906 19488
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 8576 18420 8628 18426
rect 8576 18362 8628 18368
rect 8680 18306 8708 18702
rect 8588 18278 8708 18306
rect 8298 17847 8354 17856
rect 8484 17876 8536 17882
rect 8208 17740 8260 17746
rect 8208 17682 8260 17688
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 7852 17292 8064 17320
rect 7668 17066 7788 17082
rect 7656 17060 7788 17066
rect 7708 17054 7788 17060
rect 7656 17002 7708 17008
rect 8036 16726 8064 17292
rect 7840 16720 7892 16726
rect 7840 16662 7892 16668
rect 8024 16720 8076 16726
rect 8024 16662 8076 16668
rect 7852 16250 7880 16662
rect 7932 16652 7984 16658
rect 7932 16594 7984 16600
rect 7944 16561 7972 16594
rect 7930 16552 7986 16561
rect 7930 16487 7986 16496
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 7944 15706 7972 16487
rect 8036 16182 8064 16662
rect 8024 16176 8076 16182
rect 8024 16118 8076 16124
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7840 15564 7892 15570
rect 7840 15506 7892 15512
rect 7656 15088 7708 15094
rect 7852 15065 7880 15506
rect 8024 15360 8076 15366
rect 8024 15302 8076 15308
rect 8036 15201 8064 15302
rect 8022 15192 8078 15201
rect 8022 15127 8078 15136
rect 7656 15030 7708 15036
rect 7838 15056 7894 15065
rect 7668 14521 7696 15030
rect 7838 14991 7840 15000
rect 7892 14991 7894 15000
rect 7840 14962 7892 14968
rect 7932 14884 7984 14890
rect 7932 14826 7984 14832
rect 7654 14512 7710 14521
rect 7944 14482 7972 14826
rect 8128 14618 8156 17478
rect 8220 17184 8248 17682
rect 8312 17610 8340 17847
rect 8484 17818 8536 17824
rect 8392 17672 8444 17678
rect 8390 17640 8392 17649
rect 8444 17640 8446 17649
rect 8300 17604 8352 17610
rect 8588 17610 8616 18278
rect 8772 18222 8800 18906
rect 8760 18216 8812 18222
rect 8760 18158 8812 18164
rect 8668 18080 8720 18086
rect 8720 18028 8800 18034
rect 8668 18022 8800 18028
rect 8680 18006 8800 18022
rect 8666 17912 8722 17921
rect 8666 17847 8722 17856
rect 8390 17575 8446 17584
rect 8576 17604 8628 17610
rect 8300 17546 8352 17552
rect 8404 17338 8432 17575
rect 8576 17546 8628 17552
rect 8392 17332 8444 17338
rect 8444 17292 8524 17320
rect 8392 17274 8444 17280
rect 8220 17156 8340 17184
rect 8208 17060 8260 17066
rect 8208 17002 8260 17008
rect 8220 15450 8248 17002
rect 8312 15706 8340 17156
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8300 15496 8352 15502
rect 8220 15444 8300 15450
rect 8220 15438 8352 15444
rect 8220 15422 8340 15438
rect 8220 14618 8248 15422
rect 8404 15094 8432 16594
rect 8496 15162 8524 17292
rect 8588 16726 8616 17546
rect 8680 17338 8708 17847
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8576 16720 8628 16726
rect 8576 16662 8628 16668
rect 8772 15858 8800 18006
rect 8864 17241 8892 19479
rect 9048 19310 9076 19654
rect 9036 19304 9088 19310
rect 9036 19246 9088 19252
rect 8944 18692 8996 18698
rect 8944 18634 8996 18640
rect 8956 18222 8984 18634
rect 9048 18630 9076 19246
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 8956 17542 8984 18158
rect 9048 18086 9076 18566
rect 9036 18080 9088 18086
rect 9036 18022 9088 18028
rect 9140 17814 9168 20266
rect 9232 19242 9260 20896
rect 9404 20878 9456 20884
rect 9416 20602 9444 20878
rect 9404 20596 9456 20602
rect 9404 20538 9456 20544
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 9220 19236 9272 19242
rect 9220 19178 9272 19184
rect 9232 18766 9260 19178
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 9218 18592 9274 18601
rect 9218 18527 9274 18536
rect 9232 18154 9260 18527
rect 9220 18148 9272 18154
rect 9220 18090 9272 18096
rect 9324 18034 9352 20198
rect 9416 20058 9444 20538
rect 9588 20528 9640 20534
rect 9588 20470 9640 20476
rect 9404 20052 9456 20058
rect 9404 19994 9456 20000
rect 9404 19168 9456 19174
rect 9404 19110 9456 19116
rect 9416 18698 9444 19110
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9404 18692 9456 18698
rect 9404 18634 9456 18640
rect 9232 18006 9352 18034
rect 9128 17808 9180 17814
rect 9128 17750 9180 17756
rect 9232 17660 9260 18006
rect 9404 17808 9456 17814
rect 9404 17750 9456 17756
rect 9048 17632 9260 17660
rect 8944 17536 8996 17542
rect 8944 17478 8996 17484
rect 8850 17232 8906 17241
rect 8850 17167 8906 17176
rect 8864 16046 8892 17167
rect 8956 17134 8984 17478
rect 8944 17128 8996 17134
rect 8944 17070 8996 17076
rect 8956 16454 8984 17070
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 8852 16040 8904 16046
rect 8852 15982 8904 15988
rect 8772 15830 8892 15858
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8392 15088 8444 15094
rect 8392 15030 8444 15036
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 8484 14544 8536 14550
rect 8484 14486 8536 14492
rect 7654 14447 7710 14456
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 7932 14272 7984 14278
rect 7562 14240 7618 14249
rect 7932 14214 7984 14220
rect 7562 14175 7618 14184
rect 7944 13394 7972 14214
rect 8024 13796 8076 13802
rect 8024 13738 8076 13744
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7300 11898 7328 12174
rect 7484 12102 7512 12650
rect 7944 12442 7972 13330
rect 8036 13326 8064 13738
rect 8128 13530 8156 14418
rect 8220 14278 8248 14418
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8496 13705 8524 14486
rect 8576 14340 8628 14346
rect 8576 14282 8628 14288
rect 8588 13802 8616 14282
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8576 13796 8628 13802
rect 8576 13738 8628 13744
rect 8680 13734 8708 14214
rect 8668 13728 8720 13734
rect 8482 13696 8538 13705
rect 8668 13670 8720 13676
rect 8482 13631 8538 13640
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 8392 13456 8444 13462
rect 8496 13433 8524 13631
rect 8680 13530 8708 13670
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8392 13398 8444 13404
rect 8482 13424 8538 13433
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 8036 12442 8064 13262
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 8206 12336 8262 12345
rect 8206 12271 8208 12280
rect 8260 12271 8262 12280
rect 8208 12242 8260 12248
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7484 11937 7512 12038
rect 7470 11928 7526 11937
rect 7288 11892 7340 11898
rect 8220 11898 8248 12242
rect 8404 12073 8432 13398
rect 8482 13359 8538 13368
rect 8680 13258 8708 13466
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8668 13252 8720 13258
rect 8668 13194 8720 13200
rect 8680 12986 8708 13194
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8772 12782 8800 13262
rect 8864 12850 8892 15830
rect 8956 15366 8984 16390
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8956 14890 8984 15302
rect 8944 14884 8996 14890
rect 8944 14826 8996 14832
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8680 12442 8708 12718
rect 8772 12442 8800 12718
rect 9048 12594 9076 17632
rect 9312 17604 9364 17610
rect 9312 17546 9364 17552
rect 9324 16794 9352 17546
rect 9416 17202 9444 17750
rect 9508 17338 9536 18702
rect 9600 18290 9628 20470
rect 9692 20466 9720 21406
rect 9876 21162 9904 23174
rect 10152 22964 10180 26540
rect 10230 26480 10286 26489
rect 10230 26415 10286 26424
rect 10244 25906 10272 26415
rect 10232 25900 10284 25906
rect 10232 25842 10284 25848
rect 10232 24268 10284 24274
rect 10232 24210 10284 24216
rect 10244 23322 10272 24210
rect 10232 23316 10284 23322
rect 10232 23258 10284 23264
rect 10244 23066 10272 23258
rect 10244 23038 10364 23066
rect 10152 22936 10272 22964
rect 10048 22160 10100 22166
rect 9954 22128 10010 22137
rect 10048 22102 10100 22108
rect 9954 22063 10010 22072
rect 9968 21690 9996 22063
rect 9956 21684 10008 21690
rect 9956 21626 10008 21632
rect 10060 21554 10088 22102
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 10048 21548 10100 21554
rect 10048 21490 10100 21496
rect 9968 21457 9996 21490
rect 9954 21448 10010 21457
rect 9954 21383 10010 21392
rect 10048 21412 10100 21418
rect 10048 21354 10100 21360
rect 9784 21134 9904 21162
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9784 18306 9812 21134
rect 9864 21072 9916 21078
rect 9864 21014 9916 21020
rect 9876 20602 9904 21014
rect 9864 20596 9916 20602
rect 9864 20538 9916 20544
rect 10060 20058 10088 21354
rect 10138 21312 10194 21321
rect 10138 21247 10194 21256
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 10152 19854 10180 21247
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 9876 19242 9904 19654
rect 10152 19514 10180 19790
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 9864 19236 9916 19242
rect 9864 19178 9916 19184
rect 9876 19145 9904 19178
rect 9862 19136 9918 19145
rect 9862 19071 9918 19080
rect 10048 18896 10100 18902
rect 10048 18838 10100 18844
rect 9956 18692 10008 18698
rect 9956 18634 10008 18640
rect 9588 18284 9640 18290
rect 9784 18278 9904 18306
rect 9588 18226 9640 18232
rect 9772 18216 9824 18222
rect 9772 18158 9824 18164
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 9678 18048 9734 18057
rect 9600 17626 9628 18022
rect 9678 17983 9734 17992
rect 9692 17746 9720 17983
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9600 17598 9720 17626
rect 9784 17610 9812 18158
rect 9588 17536 9640 17542
rect 9586 17504 9588 17513
rect 9640 17504 9642 17513
rect 9586 17439 9642 17448
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 9692 16794 9720 17598
rect 9772 17604 9824 17610
rect 9772 17546 9824 17552
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9678 16688 9734 16697
rect 9678 16623 9734 16632
rect 9312 16176 9364 16182
rect 9312 16118 9364 16124
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 9232 15366 9260 15982
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 9140 14278 9168 14758
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9232 13938 9260 15302
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9324 13802 9352 16118
rect 9692 15722 9720 16623
rect 9600 15694 9720 15722
rect 9404 15020 9456 15026
rect 9404 14962 9456 14968
rect 9416 14822 9444 14962
rect 9600 14890 9628 15694
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9692 15094 9720 15506
rect 9680 15088 9732 15094
rect 9680 15030 9732 15036
rect 9588 14884 9640 14890
rect 9588 14826 9640 14832
rect 9404 14816 9456 14822
rect 9402 14784 9404 14793
rect 9456 14784 9458 14793
rect 9402 14719 9458 14728
rect 9416 14074 9444 14719
rect 9496 14476 9548 14482
rect 9496 14418 9548 14424
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9312 13796 9364 13802
rect 9312 13738 9364 13744
rect 9324 13025 9352 13738
rect 9310 13016 9366 13025
rect 9310 12951 9366 12960
rect 9324 12714 9352 12951
rect 9312 12708 9364 12714
rect 9312 12650 9364 12656
rect 9048 12566 9352 12594
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8666 12200 8722 12209
rect 8666 12135 8722 12144
rect 8390 12064 8446 12073
rect 8390 11999 8446 12008
rect 7470 11863 7526 11872
rect 8208 11892 8260 11898
rect 7288 11834 7340 11840
rect 8208 11834 8260 11840
rect 8404 11778 8432 11999
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 8220 11750 8432 11778
rect 7944 11150 7972 11698
rect 8220 11354 8248 11750
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8206 11248 8262 11257
rect 8206 11183 8208 11192
rect 8260 11183 8262 11192
rect 8208 11154 8260 11160
rect 7932 11144 7984 11150
rect 7930 11112 7932 11121
rect 8116 11144 8168 11150
rect 7984 11112 7986 11121
rect 8116 11086 8168 11092
rect 7930 11047 7986 11056
rect 8128 10470 8156 11086
rect 8220 10810 8248 11154
rect 8312 11014 8340 11630
rect 8680 11286 8708 12135
rect 8944 11688 8996 11694
rect 8944 11630 8996 11636
rect 8668 11280 8720 11286
rect 8668 11222 8720 11228
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8666 10976 8722 10985
rect 8666 10911 8722 10920
rect 8482 10840 8538 10849
rect 8208 10804 8260 10810
rect 8482 10775 8484 10784
rect 8208 10746 8260 10752
rect 8536 10775 8538 10784
rect 8484 10746 8536 10752
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 8128 9994 8156 10406
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8128 9586 8156 9930
rect 8220 9586 8248 9998
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 7104 9512 7156 9518
rect 7932 9512 7984 9518
rect 7104 9454 7156 9460
rect 7286 9480 7342 9489
rect 7116 8974 7144 9454
rect 7932 9454 7984 9460
rect 7286 9415 7288 9424
rect 7340 9415 7342 9424
rect 7288 9386 7340 9392
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7104 8968 7156 8974
rect 6274 8936 6330 8945
rect 7104 8910 7156 8916
rect 6274 8871 6276 8880
rect 6328 8871 6330 8880
rect 6276 8842 6328 8848
rect 7116 8634 7144 8910
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7208 8566 7236 8978
rect 7196 8560 7248 8566
rect 7196 8502 7248 8508
rect 7944 8498 7972 9454
rect 8220 8537 8248 9522
rect 8312 9518 8340 9862
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8312 9178 8340 9454
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8206 8528 8262 8537
rect 7932 8492 7984 8498
rect 8206 8463 8262 8472
rect 7932 8434 7984 8440
rect 8496 7546 8524 10746
rect 8680 10606 8708 10911
rect 8956 10606 8984 11630
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8680 10266 8708 10542
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8772 10130 8800 10542
rect 9324 10305 9352 12566
rect 9508 12170 9536 14418
rect 9586 13016 9642 13025
rect 9586 12951 9642 12960
rect 9600 12918 9628 12951
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9496 12164 9548 12170
rect 9496 12106 9548 12112
rect 9600 12102 9628 12718
rect 9692 12306 9720 15030
rect 9784 13530 9812 16934
rect 9876 16776 9904 18278
rect 9968 17660 9996 18634
rect 10060 17814 10088 18838
rect 10244 18086 10272 22936
rect 10336 21078 10364 23038
rect 10324 21072 10376 21078
rect 10324 21014 10376 21020
rect 10336 20806 10364 21014
rect 10324 20800 10376 20806
rect 10324 20742 10376 20748
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 10048 17808 10100 17814
rect 10048 17750 10100 17756
rect 9968 17632 10088 17660
rect 9876 16748 9996 16776
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9876 15910 9904 16594
rect 9968 16182 9996 16748
rect 9956 16176 10008 16182
rect 9956 16118 10008 16124
rect 9956 16040 10008 16046
rect 9956 15982 10008 15988
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9968 15366 9996 15982
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 10060 14929 10088 17632
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10244 16726 10272 17070
rect 10232 16720 10284 16726
rect 10232 16662 10284 16668
rect 10230 16144 10286 16153
rect 10230 16079 10232 16088
rect 10284 16079 10286 16088
rect 10232 16050 10284 16056
rect 10046 14920 10102 14929
rect 9864 14884 9916 14890
rect 10046 14855 10102 14864
rect 9864 14826 9916 14832
rect 9876 14634 9904 14826
rect 9876 14606 10088 14634
rect 9864 14544 9916 14550
rect 9864 14486 9916 14492
rect 9876 14346 9904 14486
rect 9864 14340 9916 14346
rect 9916 14300 9996 14328
rect 9864 14282 9916 14288
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9784 12782 9812 13466
rect 9876 13394 9904 13670
rect 9968 13530 9996 14300
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9864 13184 9916 13190
rect 9862 13152 9864 13161
rect 9916 13152 9918 13161
rect 9862 13087 9918 13096
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9692 12102 9720 12242
rect 9772 12164 9824 12170
rect 9772 12106 9824 12112
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9600 11778 9628 12038
rect 9692 11898 9720 12038
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9600 11750 9720 11778
rect 9784 11762 9812 12106
rect 9404 11620 9456 11626
rect 9404 11562 9456 11568
rect 9416 11354 9444 11562
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9508 10849 9536 10950
rect 9494 10840 9550 10849
rect 9494 10775 9550 10784
rect 9402 10704 9458 10713
rect 9402 10639 9458 10648
rect 9416 10606 9444 10639
rect 9508 10606 9536 10775
rect 9692 10742 9720 11750
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9310 10296 9366 10305
rect 9416 10266 9444 10542
rect 9310 10231 9366 10240
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 8760 10124 8812 10130
rect 8760 10066 8812 10072
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 8758 10024 8814 10033
rect 8758 9959 8760 9968
rect 8812 9959 8814 9968
rect 8760 9930 8812 9936
rect 9508 9926 9536 10066
rect 9588 10056 9640 10062
rect 9680 10056 9732 10062
rect 9640 10016 9680 10044
rect 9588 9998 9640 10004
rect 9680 9998 9732 10004
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9508 9518 9536 9862
rect 8852 9512 8904 9518
rect 9496 9512 9548 9518
rect 8852 9454 8904 9460
rect 9494 9480 9496 9489
rect 9548 9480 9550 9489
rect 8864 9042 8892 9454
rect 9494 9415 9550 9424
rect 9508 9389 9536 9415
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 8852 9036 8904 9042
rect 8852 8978 8904 8984
rect 9586 8664 9642 8673
rect 9586 8599 9642 8608
rect 9034 8528 9090 8537
rect 9034 8463 9090 8472
rect 9048 8090 9076 8463
rect 9600 8430 9628 8599
rect 9692 8498 9720 9114
rect 9876 9042 9904 12650
rect 9968 12442 9996 13466
rect 9956 12436 10008 12442
rect 9956 12378 10008 12384
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9968 9178 9996 12174
rect 10060 11354 10088 14606
rect 10230 14512 10286 14521
rect 10230 14447 10232 14456
rect 10284 14447 10286 14456
rect 10232 14418 10284 14424
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10152 11014 10180 14282
rect 10244 14074 10272 14418
rect 10336 14074 10364 20742
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 10244 13190 10272 13670
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 10336 12918 10364 13330
rect 10324 12912 10376 12918
rect 10322 12880 10324 12889
rect 10376 12880 10378 12889
rect 10322 12815 10378 12824
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10152 9353 10180 10950
rect 10138 9344 10194 9353
rect 10138 9279 10194 9288
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 9876 7886 9904 8978
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9968 8430 9996 8774
rect 10138 8528 10194 8537
rect 10138 8463 10194 8472
rect 10152 8430 10180 8463
rect 9956 8424 10008 8430
rect 10140 8424 10192 8430
rect 9956 8366 10008 8372
rect 10046 8392 10102 8401
rect 10140 8366 10192 8372
rect 10046 8327 10102 8336
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8496 7342 8524 7482
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 6918 5536 6974 5545
rect 6918 5471 6974 5480
rect 6184 2576 6236 2582
rect 6184 2518 6236 2524
rect 6932 800 6960 5471
rect 8220 5250 8248 6326
rect 8680 6254 8708 7142
rect 9692 6866 9720 7822
rect 9876 7546 9904 7822
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9692 6458 9720 6802
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8220 5222 8340 5250
rect 8312 5166 8340 5222
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 7378 4720 7434 4729
rect 7378 4655 7434 4664
rect 7392 800 7420 4655
rect 8312 4146 8340 5102
rect 8864 4826 8892 5102
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7852 800 7880 3878
rect 8312 3738 8340 4082
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8312 2990 8340 3674
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8300 2984 8352 2990
rect 8300 2926 8352 2932
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8496 2650 8524 2926
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 8496 2553 8524 2586
rect 8482 2544 8538 2553
rect 8482 2479 8538 2488
rect 8300 1624 8352 1630
rect 8298 1592 8300 1601
rect 8352 1592 8354 1601
rect 8298 1527 8354 1536
rect 8772 800 8800 2994
rect 9232 800 9260 5102
rect 9968 4282 9996 8230
rect 10060 7546 10088 8327
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10244 7324 10272 11290
rect 10336 11218 10364 12718
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 10336 10810 10364 11154
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10152 7296 10272 7324
rect 10152 5545 10180 7296
rect 10232 7200 10284 7206
rect 10230 7168 10232 7177
rect 10284 7168 10286 7177
rect 10230 7103 10286 7112
rect 10138 5536 10194 5545
rect 10138 5471 10194 5480
rect 10428 4842 10456 28426
rect 10520 27554 10548 30262
rect 10600 29640 10652 29646
rect 10600 29582 10652 29588
rect 10612 28626 10640 29582
rect 10888 28626 10916 32127
rect 10980 31482 11008 33050
rect 11060 32972 11112 32978
rect 11060 32914 11112 32920
rect 11072 32230 11100 32914
rect 11060 32224 11112 32230
rect 11060 32166 11112 32172
rect 11072 32065 11100 32166
rect 11058 32056 11114 32065
rect 11058 31991 11114 32000
rect 10968 31476 11020 31482
rect 10968 31418 11020 31424
rect 11256 30433 11284 37062
rect 12360 36922 12388 37318
rect 12440 37266 12492 37272
rect 12348 36916 12400 36922
rect 12348 36858 12400 36864
rect 11888 35148 11940 35154
rect 11888 35090 11940 35096
rect 11900 34746 11928 35090
rect 11888 34740 11940 34746
rect 11888 34682 11940 34688
rect 11980 33856 12032 33862
rect 11980 33798 12032 33804
rect 11242 30424 11298 30433
rect 11242 30359 11298 30368
rect 11704 30184 11756 30190
rect 11704 30126 11756 30132
rect 11428 30048 11480 30054
rect 11428 29990 11480 29996
rect 11440 29714 11468 29990
rect 11716 29714 11744 30126
rect 11428 29708 11480 29714
rect 11428 29650 11480 29656
rect 11704 29708 11756 29714
rect 11704 29650 11756 29656
rect 11244 29640 11296 29646
rect 11244 29582 11296 29588
rect 11256 29306 11284 29582
rect 11716 29510 11744 29650
rect 11704 29504 11756 29510
rect 11704 29446 11756 29452
rect 11244 29300 11296 29306
rect 11244 29242 11296 29248
rect 11520 29232 11572 29238
rect 11520 29174 11572 29180
rect 11532 28665 11560 29174
rect 11716 28762 11744 29446
rect 11704 28756 11756 28762
rect 11704 28698 11756 28704
rect 11518 28656 11574 28665
rect 10600 28620 10652 28626
rect 10600 28562 10652 28568
rect 10876 28620 10928 28626
rect 11518 28591 11574 28600
rect 10876 28562 10928 28568
rect 10612 28218 10640 28562
rect 10600 28212 10652 28218
rect 10600 28154 10652 28160
rect 10888 28150 10916 28562
rect 11244 28552 11296 28558
rect 11244 28494 11296 28500
rect 11256 28218 11284 28494
rect 11244 28212 11296 28218
rect 11244 28154 11296 28160
rect 10876 28144 10928 28150
rect 10876 28086 10928 28092
rect 11256 28082 11284 28154
rect 11244 28076 11296 28082
rect 11244 28018 11296 28024
rect 10968 27872 11020 27878
rect 11532 27849 11560 28591
rect 11716 28218 11744 28698
rect 11704 28212 11756 28218
rect 11704 28154 11756 28160
rect 10968 27814 11020 27820
rect 11518 27840 11574 27849
rect 10520 27526 10640 27554
rect 10508 27396 10560 27402
rect 10508 27338 10560 27344
rect 10520 26450 10548 27338
rect 10612 26625 10640 27526
rect 10784 27328 10836 27334
rect 10784 27270 10836 27276
rect 10796 26926 10824 27270
rect 10784 26920 10836 26926
rect 10784 26862 10836 26868
rect 10598 26616 10654 26625
rect 10598 26551 10654 26560
rect 10612 26450 10640 26551
rect 10508 26444 10560 26450
rect 10508 26386 10560 26392
rect 10600 26444 10652 26450
rect 10600 26386 10652 26392
rect 10520 25265 10548 26386
rect 10612 25498 10640 26386
rect 10980 26330 11008 27814
rect 11518 27775 11574 27784
rect 11716 27577 11744 28154
rect 11058 27568 11114 27577
rect 11702 27568 11758 27577
rect 11058 27503 11060 27512
rect 11112 27503 11114 27512
rect 11520 27532 11572 27538
rect 11060 27474 11112 27480
rect 11702 27503 11758 27512
rect 11520 27474 11572 27480
rect 11428 26852 11480 26858
rect 11428 26794 11480 26800
rect 11440 26450 11468 26794
rect 11428 26444 11480 26450
rect 11428 26386 11480 26392
rect 10980 26302 11100 26330
rect 10968 26240 11020 26246
rect 10968 26182 11020 26188
rect 10876 25900 10928 25906
rect 10876 25842 10928 25848
rect 10784 25696 10836 25702
rect 10784 25638 10836 25644
rect 10600 25492 10652 25498
rect 10600 25434 10652 25440
rect 10506 25256 10562 25265
rect 10506 25191 10562 25200
rect 10506 24984 10562 24993
rect 10506 24919 10562 24928
rect 10520 24750 10548 24919
rect 10508 24744 10560 24750
rect 10508 24686 10560 24692
rect 10600 23724 10652 23730
rect 10600 23666 10652 23672
rect 10508 22432 10560 22438
rect 10508 22374 10560 22380
rect 10520 22166 10548 22374
rect 10508 22160 10560 22166
rect 10508 22102 10560 22108
rect 10612 21690 10640 23666
rect 10796 23662 10824 25638
rect 10888 25294 10916 25842
rect 10980 25838 11008 26182
rect 11072 25838 11100 26302
rect 11336 26308 11388 26314
rect 11336 26250 11388 26256
rect 10968 25832 11020 25838
rect 10966 25800 10968 25809
rect 11060 25832 11112 25838
rect 11020 25800 11022 25809
rect 11060 25774 11112 25780
rect 10966 25735 11022 25744
rect 11072 25537 11100 25774
rect 11058 25528 11114 25537
rect 11058 25463 11114 25472
rect 11244 25356 11296 25362
rect 11244 25298 11296 25304
rect 10876 25288 10928 25294
rect 10928 25248 11008 25276
rect 10876 25230 10928 25236
rect 10980 24954 11008 25248
rect 10968 24948 11020 24954
rect 10968 24890 11020 24896
rect 10876 24880 10928 24886
rect 10876 24822 10928 24828
rect 10888 24206 10916 24822
rect 11256 24342 11284 25298
rect 11244 24336 11296 24342
rect 11058 24304 11114 24313
rect 11244 24278 11296 24284
rect 11058 24239 11114 24248
rect 11072 24206 11100 24239
rect 10876 24200 10928 24206
rect 10876 24142 10928 24148
rect 11060 24200 11112 24206
rect 11060 24142 11112 24148
rect 10784 23656 10836 23662
rect 10784 23598 10836 23604
rect 10796 22982 10824 23598
rect 10888 23050 10916 24142
rect 11072 23866 11100 24142
rect 11060 23860 11112 23866
rect 11060 23802 11112 23808
rect 11348 23662 11376 26250
rect 11532 25294 11560 27474
rect 11716 27470 11744 27503
rect 11704 27464 11756 27470
rect 11704 27406 11756 27412
rect 11704 27328 11756 27334
rect 11704 27270 11756 27276
rect 11716 26790 11744 27270
rect 11704 26784 11756 26790
rect 11704 26726 11756 26732
rect 11610 26344 11666 26353
rect 11610 26279 11666 26288
rect 11624 26246 11652 26279
rect 11612 26240 11664 26246
rect 11612 26182 11664 26188
rect 11612 25764 11664 25770
rect 11612 25706 11664 25712
rect 11624 25362 11652 25706
rect 11612 25356 11664 25362
rect 11612 25298 11664 25304
rect 11428 25288 11480 25294
rect 11428 25230 11480 25236
rect 11520 25288 11572 25294
rect 11520 25230 11572 25236
rect 11440 25158 11468 25230
rect 11428 25152 11480 25158
rect 11428 25094 11480 25100
rect 11428 24744 11480 24750
rect 11428 24686 11480 24692
rect 11520 24744 11572 24750
rect 11520 24686 11572 24692
rect 11440 23866 11468 24686
rect 11428 23860 11480 23866
rect 11428 23802 11480 23808
rect 11532 23730 11560 24686
rect 11624 24614 11652 25298
rect 11612 24608 11664 24614
rect 11612 24550 11664 24556
rect 11624 24070 11652 24550
rect 11612 24064 11664 24070
rect 11612 24006 11664 24012
rect 11520 23724 11572 23730
rect 11520 23666 11572 23672
rect 11336 23656 11388 23662
rect 11336 23598 11388 23604
rect 11244 23588 11296 23594
rect 11244 23530 11296 23536
rect 11060 23520 11112 23526
rect 11060 23462 11112 23468
rect 10968 23112 11020 23118
rect 11072 23066 11100 23462
rect 11020 23060 11100 23066
rect 10968 23054 11100 23060
rect 10876 23044 10928 23050
rect 10980 23038 11100 23054
rect 10876 22986 10928 22992
rect 10784 22976 10836 22982
rect 10784 22918 10836 22924
rect 10692 22704 10744 22710
rect 10692 22646 10744 22652
rect 10782 22672 10838 22681
rect 10704 22030 10732 22646
rect 10782 22607 10838 22616
rect 10796 22506 10824 22607
rect 10784 22500 10836 22506
rect 10784 22442 10836 22448
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 10600 21684 10652 21690
rect 10600 21626 10652 21632
rect 10508 21616 10560 21622
rect 10508 21558 10560 21564
rect 10520 21078 10548 21558
rect 10508 21072 10560 21078
rect 10506 21040 10508 21049
rect 10560 21040 10562 21049
rect 10506 20975 10562 20984
rect 10508 20936 10560 20942
rect 10508 20878 10560 20884
rect 10520 20398 10548 20878
rect 10796 20534 10824 22442
rect 10888 21570 10916 22986
rect 10968 22772 11020 22778
rect 11072 22760 11100 23038
rect 11020 22732 11100 22760
rect 11152 22772 11204 22778
rect 10968 22714 11020 22720
rect 11152 22714 11204 22720
rect 11060 22636 11112 22642
rect 11060 22578 11112 22584
rect 11072 22098 11100 22578
rect 11060 22092 11112 22098
rect 11060 22034 11112 22040
rect 11164 21690 11192 22714
rect 11256 21894 11284 23530
rect 11520 23180 11572 23186
rect 11520 23122 11572 23128
rect 11612 23180 11664 23186
rect 11612 23122 11664 23128
rect 11428 22976 11480 22982
rect 11428 22918 11480 22924
rect 11440 22710 11468 22918
rect 11428 22704 11480 22710
rect 11428 22646 11480 22652
rect 11532 22506 11560 23122
rect 11624 22778 11652 23122
rect 11612 22772 11664 22778
rect 11612 22714 11664 22720
rect 11520 22500 11572 22506
rect 11520 22442 11572 22448
rect 11336 22092 11388 22098
rect 11388 22052 11468 22080
rect 11336 22034 11388 22040
rect 11244 21888 11296 21894
rect 11244 21830 11296 21836
rect 11242 21720 11298 21729
rect 11152 21684 11204 21690
rect 11242 21655 11298 21664
rect 11152 21626 11204 21632
rect 10888 21542 11192 21570
rect 11060 21004 11112 21010
rect 11060 20946 11112 20952
rect 10600 20528 10652 20534
rect 10600 20470 10652 20476
rect 10784 20528 10836 20534
rect 10784 20470 10836 20476
rect 10508 20392 10560 20398
rect 10508 20334 10560 20340
rect 10612 20330 10640 20470
rect 11072 20466 11100 20946
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 10600 20324 10652 20330
rect 10600 20266 10652 20272
rect 11164 20262 11192 21542
rect 11256 21486 11284 21655
rect 11244 21480 11296 21486
rect 11244 21422 11296 21428
rect 10968 20256 11020 20262
rect 10968 20198 11020 20204
rect 11152 20256 11204 20262
rect 11152 20198 11204 20204
rect 10784 19916 10836 19922
rect 10784 19858 10836 19864
rect 10508 19848 10560 19854
rect 10508 19790 10560 19796
rect 10520 18222 10548 19790
rect 10796 19417 10824 19858
rect 10782 19408 10838 19417
rect 10782 19343 10838 19352
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10704 19009 10732 19110
rect 10690 19000 10746 19009
rect 10690 18935 10746 18944
rect 10600 18896 10652 18902
rect 10600 18838 10652 18844
rect 10612 18698 10640 18838
rect 10704 18834 10732 18935
rect 10796 18902 10824 19343
rect 10784 18896 10836 18902
rect 10784 18838 10836 18844
rect 10692 18828 10744 18834
rect 10692 18770 10744 18776
rect 10704 18714 10732 18770
rect 10600 18692 10652 18698
rect 10704 18686 10824 18714
rect 10980 18698 11008 20198
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 11072 19174 11100 19654
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 11072 18970 11100 19110
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 10600 18634 10652 18640
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 10506 17232 10562 17241
rect 10506 17167 10562 17176
rect 10520 17134 10548 17167
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10506 16552 10562 16561
rect 10506 16487 10562 16496
rect 10520 16454 10548 16487
rect 10508 16448 10560 16454
rect 10508 16390 10560 16396
rect 10520 15570 10548 16390
rect 10508 15564 10560 15570
rect 10508 15506 10560 15512
rect 10508 15360 10560 15366
rect 10508 15302 10560 15308
rect 10520 13161 10548 15302
rect 10506 13152 10562 13161
rect 10506 13087 10562 13096
rect 10506 11792 10562 11801
rect 10506 11727 10562 11736
rect 10520 5370 10548 11727
rect 10612 11354 10640 18022
rect 10704 17649 10732 18362
rect 10796 18193 10824 18686
rect 10968 18692 11020 18698
rect 10968 18634 11020 18640
rect 11256 18306 11284 21422
rect 11440 21350 11468 22052
rect 11716 22001 11744 26726
rect 11796 26376 11848 26382
rect 11794 26344 11796 26353
rect 11848 26344 11850 26353
rect 11794 26279 11850 26288
rect 11794 26072 11850 26081
rect 11850 26030 11928 26058
rect 11794 26007 11796 26016
rect 11848 26007 11850 26016
rect 11796 25978 11848 25984
rect 11794 25936 11850 25945
rect 11794 25871 11850 25880
rect 11808 24818 11836 25871
rect 11900 25401 11928 26030
rect 11886 25392 11942 25401
rect 11886 25327 11942 25336
rect 11888 25288 11940 25294
rect 11888 25230 11940 25236
rect 11796 24812 11848 24818
rect 11796 24754 11848 24760
rect 11808 24682 11836 24754
rect 11796 24676 11848 24682
rect 11796 24618 11848 24624
rect 11900 22098 11928 25230
rect 11888 22092 11940 22098
rect 11888 22034 11940 22040
rect 11702 21992 11758 22001
rect 11702 21927 11758 21936
rect 11796 21616 11848 21622
rect 11796 21558 11848 21564
rect 11336 21344 11388 21350
rect 11336 21286 11388 21292
rect 11428 21344 11480 21350
rect 11428 21286 11480 21292
rect 11348 20641 11376 21286
rect 11440 21010 11468 21286
rect 11428 21004 11480 21010
rect 11428 20946 11480 20952
rect 11334 20632 11390 20641
rect 11334 20567 11390 20576
rect 11440 20534 11468 20946
rect 11428 20528 11480 20534
rect 11428 20470 11480 20476
rect 11808 20040 11836 21558
rect 11886 20632 11942 20641
rect 11886 20567 11942 20576
rect 11900 20534 11928 20567
rect 11888 20528 11940 20534
rect 11888 20470 11940 20476
rect 11900 20262 11928 20470
rect 11888 20256 11940 20262
rect 11888 20198 11940 20204
rect 11808 20012 11928 20040
rect 11612 19984 11664 19990
rect 11610 19952 11612 19961
rect 11664 19952 11666 19961
rect 11610 19887 11666 19896
rect 11794 19952 11850 19961
rect 11794 19887 11850 19896
rect 11428 19440 11480 19446
rect 11428 19382 11480 19388
rect 11336 19304 11388 19310
rect 11336 19246 11388 19252
rect 11348 18630 11376 19246
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11348 18329 11376 18566
rect 11164 18278 11284 18306
rect 11334 18320 11390 18329
rect 10782 18184 10838 18193
rect 10782 18119 10784 18128
rect 10836 18119 10838 18128
rect 10784 18090 10836 18096
rect 11164 17746 11192 18278
rect 11334 18255 11336 18264
rect 11388 18255 11390 18264
rect 11336 18226 11388 18232
rect 11152 17740 11204 17746
rect 11152 17682 11204 17688
rect 11336 17740 11388 17746
rect 11336 17682 11388 17688
rect 11060 17672 11112 17678
rect 10690 17640 10746 17649
rect 11060 17614 11112 17620
rect 10690 17575 10746 17584
rect 10704 16046 10732 17575
rect 10782 16824 10838 16833
rect 11072 16794 11100 17614
rect 11164 16969 11192 17682
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 11150 16960 11206 16969
rect 11150 16895 11206 16904
rect 10782 16759 10838 16768
rect 11060 16788 11112 16794
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10704 14278 10732 15506
rect 10796 14958 10824 16759
rect 11060 16730 11112 16736
rect 11256 16658 11284 17138
rect 11348 16998 11376 17682
rect 11336 16992 11388 16998
rect 11336 16934 11388 16940
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10888 16250 10916 16526
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 11072 15858 11100 16594
rect 11152 15972 11204 15978
rect 11152 15914 11204 15920
rect 10888 15830 11100 15858
rect 10888 15706 10916 15830
rect 10966 15736 11022 15745
rect 10876 15700 10928 15706
rect 10966 15671 11022 15680
rect 10876 15642 10928 15648
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10796 14550 10824 14894
rect 10888 14618 10916 15438
rect 10980 15162 11008 15671
rect 11164 15570 11192 15914
rect 11244 15904 11296 15910
rect 11348 15892 11376 16934
rect 11440 16425 11468 19382
rect 11612 19236 11664 19242
rect 11612 19178 11664 19184
rect 11624 18612 11652 19178
rect 11704 18964 11756 18970
rect 11704 18906 11756 18912
rect 11716 18737 11744 18906
rect 11702 18728 11758 18737
rect 11702 18663 11758 18672
rect 11624 18584 11744 18612
rect 11518 17912 11574 17921
rect 11716 17882 11744 18584
rect 11518 17847 11520 17856
rect 11572 17847 11574 17856
rect 11704 17876 11756 17882
rect 11520 17818 11572 17824
rect 11704 17818 11756 17824
rect 11612 17808 11664 17814
rect 11612 17750 11664 17756
rect 11624 16998 11652 17750
rect 11704 17264 11756 17270
rect 11704 17206 11756 17212
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 11426 16416 11482 16425
rect 11426 16351 11482 16360
rect 11296 15864 11376 15892
rect 11244 15846 11296 15852
rect 11348 15858 11376 15864
rect 11348 15830 11468 15858
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11152 15564 11204 15570
rect 11152 15506 11204 15512
rect 11058 15192 11114 15201
rect 10968 15156 11020 15162
rect 11058 15127 11060 15136
rect 10968 15098 11020 15104
rect 11112 15127 11114 15136
rect 11060 15098 11112 15104
rect 10966 14920 11022 14929
rect 10966 14855 11022 14864
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10782 14240 10838 14249
rect 10782 14175 10838 14184
rect 10692 13456 10744 13462
rect 10692 13398 10744 13404
rect 10704 12986 10732 13398
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10796 12866 10824 14175
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10704 12838 10824 12866
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10428 4814 10640 4842
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 9680 4004 9732 4010
rect 9680 3946 9732 3952
rect 9692 800 9720 3946
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 10520 2990 10548 3470
rect 10508 2984 10560 2990
rect 10506 2952 10508 2961
rect 10560 2952 10562 2961
rect 10506 2887 10562 2896
rect 10322 2544 10378 2553
rect 10322 2479 10324 2488
rect 10376 2479 10378 2488
rect 10324 2450 10376 2456
rect 10612 800 10640 4814
rect 10704 3194 10732 12838
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10796 11558 10824 12242
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10784 11144 10836 11150
rect 10782 11112 10784 11121
rect 10836 11112 10838 11121
rect 10782 11047 10838 11056
rect 10888 10033 10916 14010
rect 10980 13870 11008 14855
rect 11072 13938 11100 15098
rect 11164 14822 11192 15506
rect 11348 15162 11376 15642
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 11244 15088 11296 15094
rect 11242 15056 11244 15065
rect 11296 15056 11298 15065
rect 11242 14991 11298 15000
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11440 14278 11468 15830
rect 11532 15026 11560 16526
rect 11624 15910 11652 16934
rect 11716 16726 11744 17206
rect 11704 16720 11756 16726
rect 11704 16662 11756 16668
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11610 15736 11666 15745
rect 11610 15671 11666 15680
rect 11624 15638 11652 15671
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11610 15464 11666 15473
rect 11610 15399 11666 15408
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 11532 14618 11560 14962
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11428 14272 11480 14278
rect 11428 14214 11480 14220
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 11348 13734 11376 14214
rect 11428 13932 11480 13938
rect 11428 13874 11480 13880
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 10966 13560 11022 13569
rect 10966 13495 11022 13504
rect 10980 12714 11008 13495
rect 11164 13394 11192 13670
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 11242 13288 11298 13297
rect 11242 13223 11298 13232
rect 11256 12918 11284 13223
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 11244 12912 11296 12918
rect 11244 12854 11296 12860
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 11072 12186 11100 12854
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11164 12374 11192 12786
rect 11152 12368 11204 12374
rect 11152 12310 11204 12316
rect 10980 12170 11100 12186
rect 11348 12170 11376 13126
rect 10968 12164 11100 12170
rect 11020 12158 11100 12164
rect 11336 12164 11388 12170
rect 10968 12106 11020 12112
rect 11336 12106 11388 12112
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 11072 11257 11100 11494
rect 11348 11286 11376 11630
rect 11336 11280 11388 11286
rect 11058 11248 11114 11257
rect 11336 11222 11388 11228
rect 11058 11183 11060 11192
rect 11112 11183 11114 11192
rect 11060 11154 11112 11160
rect 11072 11123 11100 11154
rect 11348 10470 11376 11222
rect 11336 10464 11388 10470
rect 11334 10432 11336 10441
rect 11388 10432 11390 10441
rect 11334 10367 11390 10376
rect 11440 10130 11468 13874
rect 11624 13410 11652 15399
rect 11716 13938 11744 16662
rect 11808 15570 11836 19887
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11796 14952 11848 14958
rect 11796 14894 11848 14900
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11716 13530 11744 13670
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11532 13382 11652 13410
rect 11532 12764 11560 13382
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11624 12986 11652 13262
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11716 12866 11744 13466
rect 11808 12986 11836 14894
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11716 12838 11836 12866
rect 11532 12736 11744 12764
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11624 12442 11652 12582
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11532 10470 11560 11494
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11716 10266 11744 12736
rect 11808 12442 11836 12838
rect 11796 12436 11848 12442
rect 11900 12424 11928 20012
rect 11992 18306 12020 33798
rect 12544 31754 12572 37454
rect 12624 37256 12676 37262
rect 12624 37198 12676 37204
rect 12636 36922 12664 37198
rect 13544 37120 13596 37126
rect 13544 37062 13596 37068
rect 12624 36916 12676 36922
rect 12624 36858 12676 36864
rect 12624 32904 12676 32910
rect 12622 32872 12624 32881
rect 12808 32904 12860 32910
rect 12676 32872 12678 32881
rect 12808 32846 12860 32852
rect 12622 32807 12678 32816
rect 12636 32570 12664 32807
rect 12624 32564 12676 32570
rect 12624 32506 12676 32512
rect 12820 32230 12848 32846
rect 12808 32224 12860 32230
rect 13360 32224 13412 32230
rect 12808 32166 12860 32172
rect 13358 32192 13360 32201
rect 13412 32192 13414 32201
rect 12532 31748 12584 31754
rect 12532 31690 12584 31696
rect 12072 30728 12124 30734
rect 12072 30670 12124 30676
rect 12084 30258 12112 30670
rect 12716 30592 12768 30598
rect 12716 30534 12768 30540
rect 12532 30320 12584 30326
rect 12532 30262 12584 30268
rect 12072 30252 12124 30258
rect 12072 30194 12124 30200
rect 12084 29578 12112 30194
rect 12164 30048 12216 30054
rect 12164 29990 12216 29996
rect 12176 29782 12204 29990
rect 12544 29850 12572 30262
rect 12728 30190 12756 30534
rect 12716 30184 12768 30190
rect 12716 30126 12768 30132
rect 12728 29850 12756 30126
rect 12532 29844 12584 29850
rect 12532 29786 12584 29792
rect 12716 29844 12768 29850
rect 12716 29786 12768 29792
rect 12164 29776 12216 29782
rect 12164 29718 12216 29724
rect 12072 29572 12124 29578
rect 12072 29514 12124 29520
rect 12084 29034 12112 29514
rect 12176 29306 12204 29718
rect 12728 29510 12756 29786
rect 12716 29504 12768 29510
rect 12716 29446 12768 29452
rect 12164 29300 12216 29306
rect 12164 29242 12216 29248
rect 12072 29028 12124 29034
rect 12072 28970 12124 28976
rect 12348 29028 12400 29034
rect 12348 28970 12400 28976
rect 12084 27334 12112 28970
rect 12360 27606 12388 28970
rect 12622 27840 12678 27849
rect 12622 27775 12678 27784
rect 12348 27600 12400 27606
rect 12348 27542 12400 27548
rect 12072 27328 12124 27334
rect 12072 27270 12124 27276
rect 12084 27130 12112 27270
rect 12072 27124 12124 27130
rect 12072 27066 12124 27072
rect 12532 26784 12584 26790
rect 12532 26726 12584 26732
rect 12072 26444 12124 26450
rect 12072 26386 12124 26392
rect 12440 26444 12492 26450
rect 12440 26386 12492 26392
rect 12084 25498 12112 26386
rect 12452 25974 12480 26386
rect 12440 25968 12492 25974
rect 12440 25910 12492 25916
rect 12164 25832 12216 25838
rect 12164 25774 12216 25780
rect 12072 25492 12124 25498
rect 12072 25434 12124 25440
rect 12176 25378 12204 25774
rect 12084 25350 12204 25378
rect 12544 25378 12572 26726
rect 12636 25498 12664 27775
rect 12716 26444 12768 26450
rect 12716 26386 12768 26392
rect 12728 25974 12756 26386
rect 12716 25968 12768 25974
rect 12716 25910 12768 25916
rect 12624 25492 12676 25498
rect 12676 25452 12756 25480
rect 12624 25434 12676 25440
rect 12544 25350 12664 25378
rect 12084 19446 12112 25350
rect 12636 25158 12664 25350
rect 12624 25152 12676 25158
rect 12624 25094 12676 25100
rect 12256 24608 12308 24614
rect 12254 24576 12256 24585
rect 12308 24576 12310 24585
rect 12254 24511 12310 24520
rect 12440 24200 12492 24206
rect 12440 24142 12492 24148
rect 12348 24132 12400 24138
rect 12348 24074 12400 24080
rect 12164 24064 12216 24070
rect 12164 24006 12216 24012
rect 12256 24064 12308 24070
rect 12256 24006 12308 24012
rect 12176 20806 12204 24006
rect 12268 22778 12296 24006
rect 12360 23662 12388 24074
rect 12452 23866 12480 24142
rect 12440 23860 12492 23866
rect 12440 23802 12492 23808
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 12360 23254 12388 23598
rect 12348 23248 12400 23254
rect 12348 23190 12400 23196
rect 12440 22976 12492 22982
rect 12440 22918 12492 22924
rect 12256 22772 12308 22778
rect 12256 22714 12308 22720
rect 12452 22681 12480 22918
rect 12532 22772 12584 22778
rect 12532 22714 12584 22720
rect 12438 22672 12494 22681
rect 12438 22607 12494 22616
rect 12348 22500 12400 22506
rect 12348 22442 12400 22448
rect 12360 22386 12388 22442
rect 12360 22358 12480 22386
rect 12256 22092 12308 22098
rect 12256 22034 12308 22040
rect 12164 20800 12216 20806
rect 12164 20742 12216 20748
rect 12268 20097 12296 22034
rect 12452 21894 12480 22358
rect 12544 22166 12572 22714
rect 12636 22710 12664 25094
rect 12728 24818 12756 25452
rect 12716 24812 12768 24818
rect 12716 24754 12768 24760
rect 12728 23866 12756 24754
rect 12716 23860 12768 23866
rect 12716 23802 12768 23808
rect 12820 23254 12848 32166
rect 13358 32127 13414 32136
rect 12900 31680 12952 31686
rect 12900 31622 12952 31628
rect 12912 31346 12940 31622
rect 12900 31340 12952 31346
rect 12900 31282 12952 31288
rect 12912 30394 12940 31282
rect 12990 31240 13046 31249
rect 12990 31175 13046 31184
rect 13004 31142 13032 31175
rect 12992 31136 13044 31142
rect 12992 31078 13044 31084
rect 12900 30388 12952 30394
rect 12900 30330 12952 30336
rect 12900 28960 12952 28966
rect 12900 28902 12952 28908
rect 12912 28626 12940 28902
rect 12900 28620 12952 28626
rect 12900 28562 12952 28568
rect 12912 27946 12940 28562
rect 12900 27940 12952 27946
rect 12900 27882 12952 27888
rect 13004 27826 13032 31078
rect 13176 30796 13228 30802
rect 13176 30738 13228 30744
rect 13188 30258 13216 30738
rect 13360 30592 13412 30598
rect 13360 30534 13412 30540
rect 13176 30252 13228 30258
rect 13176 30194 13228 30200
rect 13188 29782 13216 30194
rect 13268 30116 13320 30122
rect 13268 30058 13320 30064
rect 13176 29776 13228 29782
rect 13176 29718 13228 29724
rect 13280 29306 13308 30058
rect 13372 30025 13400 30534
rect 13452 30388 13504 30394
rect 13452 30330 13504 30336
rect 13358 30016 13414 30025
rect 13358 29951 13414 29960
rect 13268 29300 13320 29306
rect 13268 29242 13320 29248
rect 13464 29102 13492 30330
rect 13452 29096 13504 29102
rect 13452 29038 13504 29044
rect 13268 28552 13320 28558
rect 13268 28494 13320 28500
rect 12912 27798 13032 27826
rect 12912 25362 12940 27798
rect 12992 26376 13044 26382
rect 12992 26318 13044 26324
rect 13176 26376 13228 26382
rect 13176 26318 13228 26324
rect 13004 25401 13032 26318
rect 13188 25770 13216 26318
rect 13176 25764 13228 25770
rect 13176 25706 13228 25712
rect 13084 25696 13136 25702
rect 13084 25638 13136 25644
rect 12990 25392 13046 25401
rect 12900 25356 12952 25362
rect 12990 25327 13046 25336
rect 12900 25298 12952 25304
rect 13096 24750 13124 25638
rect 13176 25356 13228 25362
rect 13176 25298 13228 25304
rect 13188 24886 13216 25298
rect 13176 24880 13228 24886
rect 13174 24848 13176 24857
rect 13228 24848 13230 24857
rect 13174 24783 13230 24792
rect 13188 24757 13216 24783
rect 13280 24750 13308 28494
rect 13556 28098 13584 37062
rect 13648 35057 13676 37703
rect 13832 37330 13860 40996
rect 13820 37324 13872 37330
rect 13820 37266 13872 37272
rect 14292 36009 14320 40996
rect 14372 38888 14424 38894
rect 14372 38830 14424 38836
rect 13726 36000 13782 36009
rect 13726 35935 13782 35944
rect 14278 36000 14334 36009
rect 14278 35935 14334 35944
rect 13634 35048 13690 35057
rect 13634 34983 13690 34992
rect 13740 32434 13768 35935
rect 14004 35216 14056 35222
rect 14004 35158 14056 35164
rect 14016 34746 14044 35158
rect 14004 34740 14056 34746
rect 14004 34682 14056 34688
rect 14094 33280 14150 33289
rect 14094 33215 14150 33224
rect 14004 32768 14056 32774
rect 14004 32710 14056 32716
rect 13728 32428 13780 32434
rect 13728 32370 13780 32376
rect 13636 32360 13688 32366
rect 13636 32302 13688 32308
rect 13648 32026 13676 32302
rect 13636 32020 13688 32026
rect 13636 31962 13688 31968
rect 14016 31890 14044 32710
rect 14004 31884 14056 31890
rect 14004 31826 14056 31832
rect 13820 31816 13872 31822
rect 13820 31758 13872 31764
rect 13832 30938 13860 31758
rect 14016 30938 14044 31826
rect 13820 30932 13872 30938
rect 13820 30874 13872 30880
rect 14004 30932 14056 30938
rect 14004 30874 14056 30880
rect 13728 30864 13780 30870
rect 13728 30806 13780 30812
rect 13740 30410 13768 30806
rect 13910 30424 13966 30433
rect 13740 30382 13910 30410
rect 13910 30359 13966 30368
rect 13924 30326 13952 30359
rect 13912 30320 13964 30326
rect 13912 30262 13964 30268
rect 13636 29708 13688 29714
rect 13636 29650 13688 29656
rect 13648 29617 13676 29650
rect 13634 29608 13690 29617
rect 13634 29543 13690 29552
rect 13648 29034 13676 29543
rect 14108 29345 14136 33215
rect 14384 32609 14412 38830
rect 14752 36961 14780 40996
rect 15292 38820 15344 38826
rect 15292 38762 15344 38768
rect 15304 38214 15332 38762
rect 15292 38208 15344 38214
rect 15292 38150 15344 38156
rect 15016 37324 15068 37330
rect 15016 37266 15068 37272
rect 14738 36952 14794 36961
rect 14738 36887 14794 36896
rect 14740 34944 14792 34950
rect 14740 34886 14792 34892
rect 14752 34610 14780 34886
rect 14740 34604 14792 34610
rect 14740 34546 14792 34552
rect 14554 34504 14610 34513
rect 14554 34439 14556 34448
rect 14608 34439 14610 34448
rect 14556 34410 14608 34416
rect 14568 33998 14596 34410
rect 14556 33992 14608 33998
rect 14556 33934 14608 33940
rect 14568 33658 14596 33934
rect 14556 33652 14608 33658
rect 14556 33594 14608 33600
rect 14462 33552 14518 33561
rect 14462 33487 14518 33496
rect 14370 32600 14426 32609
rect 14370 32535 14426 32544
rect 14186 30288 14242 30297
rect 14186 30223 14242 30232
rect 14200 30190 14228 30223
rect 14188 30184 14240 30190
rect 14188 30126 14240 30132
rect 14200 29850 14228 30126
rect 14188 29844 14240 29850
rect 14188 29786 14240 29792
rect 14094 29336 14150 29345
rect 14094 29271 14150 29280
rect 13912 29096 13964 29102
rect 14096 29096 14148 29102
rect 13912 29038 13964 29044
rect 14094 29064 14096 29073
rect 14148 29064 14150 29073
rect 13636 29028 13688 29034
rect 13636 28970 13688 28976
rect 13726 28656 13782 28665
rect 13726 28591 13782 28600
rect 13820 28620 13872 28626
rect 13556 28070 13676 28098
rect 13648 28014 13676 28070
rect 13452 28008 13504 28014
rect 13452 27950 13504 27956
rect 13636 28008 13688 28014
rect 13636 27950 13688 27956
rect 13360 27940 13412 27946
rect 13360 27882 13412 27888
rect 13372 27538 13400 27882
rect 13360 27532 13412 27538
rect 13360 27474 13412 27480
rect 13372 27130 13400 27474
rect 13464 27305 13492 27950
rect 13544 27328 13596 27334
rect 13450 27296 13506 27305
rect 13544 27270 13596 27276
rect 13450 27231 13506 27240
rect 13360 27124 13412 27130
rect 13360 27066 13412 27072
rect 13556 26790 13584 27270
rect 13740 26874 13768 28591
rect 13820 28562 13872 28568
rect 13832 27606 13860 28562
rect 13924 28558 13952 29038
rect 14094 28999 14150 29008
rect 14384 28762 14412 32535
rect 14476 29102 14504 33487
rect 14646 33416 14702 33425
rect 14646 33351 14702 33360
rect 14556 31204 14608 31210
rect 14556 31146 14608 31152
rect 14568 30394 14596 31146
rect 14556 30388 14608 30394
rect 14556 30330 14608 30336
rect 14464 29096 14516 29102
rect 14464 29038 14516 29044
rect 14372 28756 14424 28762
rect 14372 28698 14424 28704
rect 13912 28552 13964 28558
rect 13912 28494 13964 28500
rect 14004 28416 14056 28422
rect 14004 28358 14056 28364
rect 13820 27600 13872 27606
rect 13820 27542 13872 27548
rect 14016 26926 14044 28358
rect 14384 28082 14412 28698
rect 14372 28076 14424 28082
rect 14372 28018 14424 28024
rect 14188 28008 14240 28014
rect 14188 27950 14240 27956
rect 14200 27674 14228 27950
rect 14188 27668 14240 27674
rect 14188 27610 14240 27616
rect 14278 27160 14334 27169
rect 14278 27095 14334 27104
rect 13648 26846 13768 26874
rect 14004 26920 14056 26926
rect 14004 26862 14056 26868
rect 13544 26784 13596 26790
rect 13544 26726 13596 26732
rect 13452 26308 13504 26314
rect 13452 26250 13504 26256
rect 13360 25356 13412 25362
rect 13360 25298 13412 25304
rect 13372 25226 13400 25298
rect 13360 25220 13412 25226
rect 13360 25162 13412 25168
rect 13372 24886 13400 25162
rect 13360 24880 13412 24886
rect 13360 24822 13412 24828
rect 13464 24750 13492 26250
rect 13544 25832 13596 25838
rect 13544 25774 13596 25780
rect 13556 25362 13584 25774
rect 13544 25356 13596 25362
rect 13544 25298 13596 25304
rect 13084 24744 13136 24750
rect 13084 24686 13136 24692
rect 13268 24744 13320 24750
rect 13268 24686 13320 24692
rect 13452 24744 13504 24750
rect 13452 24686 13504 24692
rect 13174 24440 13230 24449
rect 13174 24375 13230 24384
rect 12900 24336 12952 24342
rect 12900 24278 12952 24284
rect 12808 23248 12860 23254
rect 12808 23190 12860 23196
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12624 22704 12676 22710
rect 12624 22646 12676 22652
rect 12820 22506 12848 22918
rect 12808 22500 12860 22506
rect 12808 22442 12860 22448
rect 12532 22160 12584 22166
rect 12532 22102 12584 22108
rect 12716 22092 12768 22098
rect 12716 22034 12768 22040
rect 12808 22092 12860 22098
rect 12912 22080 12940 24278
rect 12992 24200 13044 24206
rect 12992 24142 13044 24148
rect 13004 22574 13032 24142
rect 12992 22568 13044 22574
rect 12992 22510 13044 22516
rect 12860 22052 12940 22080
rect 12808 22034 12860 22040
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 12728 21622 12756 22034
rect 12716 21616 12768 21622
rect 12716 21558 12768 21564
rect 12622 21448 12678 21457
rect 12622 21383 12678 21392
rect 12636 21146 12664 21383
rect 12728 21350 12756 21558
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12624 21140 12676 21146
rect 12624 21082 12676 21088
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 12716 20596 12768 20602
rect 12716 20538 12768 20544
rect 12254 20088 12310 20097
rect 12254 20023 12310 20032
rect 12164 19848 12216 19854
rect 12164 19790 12216 19796
rect 12072 19440 12124 19446
rect 12072 19382 12124 19388
rect 12176 18970 12204 19790
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 11992 18278 12112 18306
rect 11980 18216 12032 18222
rect 11980 18158 12032 18164
rect 11992 17814 12020 18158
rect 11980 17808 12032 17814
rect 11980 17750 12032 17756
rect 11980 17060 12032 17066
rect 11980 17002 12032 17008
rect 11992 13394 12020 17002
rect 12084 14482 12112 18278
rect 12268 17270 12296 20023
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12360 19310 12388 19858
rect 12452 19378 12480 20538
rect 12728 19922 12756 20538
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 12544 19242 12572 19790
rect 12820 19786 12848 22034
rect 12992 21548 13044 21554
rect 12992 21490 13044 21496
rect 12808 19780 12860 19786
rect 12808 19722 12860 19728
rect 12716 19508 12768 19514
rect 12716 19450 12768 19456
rect 12624 19304 12676 19310
rect 12622 19272 12624 19281
rect 12676 19272 12678 19281
rect 12532 19236 12584 19242
rect 12622 19207 12678 19216
rect 12532 19178 12584 19184
rect 12440 19168 12492 19174
rect 12360 19128 12440 19156
rect 12256 17264 12308 17270
rect 12256 17206 12308 17212
rect 12360 17105 12388 19128
rect 12440 19110 12492 19116
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12452 17882 12480 18770
rect 12544 18766 12572 19178
rect 12728 18834 12756 19450
rect 12808 19304 12860 19310
rect 12900 19304 12952 19310
rect 12808 19246 12860 19252
rect 12898 19272 12900 19281
rect 12952 19272 12954 19281
rect 12716 18828 12768 18834
rect 12820 18816 12848 19246
rect 12898 19207 12954 19216
rect 12820 18788 12940 18816
rect 12716 18770 12768 18776
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12544 18358 12572 18702
rect 12532 18352 12584 18358
rect 12532 18294 12584 18300
rect 12728 17882 12756 18770
rect 12808 18692 12860 18698
rect 12808 18634 12860 18640
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 12452 17338 12480 17818
rect 12532 17808 12584 17814
rect 12820 17785 12848 18634
rect 12532 17750 12584 17756
rect 12806 17776 12862 17785
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12440 17128 12492 17134
rect 12346 17096 12402 17105
rect 12544 17116 12572 17750
rect 12806 17711 12862 17720
rect 12912 17513 12940 18788
rect 12714 17504 12770 17513
rect 12714 17439 12770 17448
rect 12898 17504 12954 17513
rect 12898 17439 12954 17448
rect 12492 17088 12572 17116
rect 12728 17105 12756 17439
rect 12714 17096 12770 17105
rect 12440 17070 12492 17076
rect 12346 17031 12402 17040
rect 12714 17031 12770 17040
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12162 16416 12218 16425
rect 12162 16351 12218 16360
rect 12176 15473 12204 16351
rect 12360 15910 12388 16594
rect 12544 15994 12572 16594
rect 12636 16153 12664 16594
rect 12622 16144 12678 16153
rect 12622 16079 12678 16088
rect 12440 15972 12492 15978
rect 12544 15966 12664 15994
rect 12440 15914 12492 15920
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 12452 15638 12480 15914
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 12440 15632 12492 15638
rect 12440 15574 12492 15580
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12162 15464 12218 15473
rect 12162 15399 12218 15408
rect 12268 14550 12296 15506
rect 12348 15088 12400 15094
rect 12348 15030 12400 15036
rect 12256 14544 12308 14550
rect 12256 14486 12308 14492
rect 12072 14476 12124 14482
rect 12124 14436 12204 14464
rect 12072 14418 12124 14424
rect 12072 14272 12124 14278
rect 12072 14214 12124 14220
rect 12084 14006 12112 14214
rect 12072 14000 12124 14006
rect 12072 13942 12124 13948
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11992 12646 12020 13330
rect 12176 13308 12204 14436
rect 12360 14414 12388 15030
rect 12544 14822 12572 15846
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12348 14408 12400 14414
rect 12544 14385 12572 14758
rect 12348 14350 12400 14356
rect 12530 14376 12586 14385
rect 12530 14311 12586 14320
rect 12544 14278 12572 14311
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12348 13456 12400 13462
rect 12254 13424 12310 13433
rect 12348 13398 12400 13404
rect 12254 13359 12310 13368
rect 12084 13280 12204 13308
rect 12084 12753 12112 13280
rect 12268 13190 12296 13359
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12070 12744 12126 12753
rect 12070 12679 12126 12688
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11900 12396 12020 12424
rect 11796 12378 11848 12384
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11900 11898 11928 12242
rect 11992 12238 12020 12396
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11992 11830 12020 12174
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 11808 10538 11836 11154
rect 11796 10532 11848 10538
rect 11796 10474 11848 10480
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11428 10124 11480 10130
rect 11428 10066 11480 10072
rect 10874 10024 10930 10033
rect 10874 9959 10930 9968
rect 10888 9042 10916 9959
rect 11440 9722 11468 10066
rect 11808 10062 11836 10474
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11426 9480 11482 9489
rect 11426 9415 11482 9424
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10888 8498 10916 8978
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 11072 8090 11100 8298
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11164 7478 11192 9114
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 10888 7002 10916 7346
rect 10968 7336 11020 7342
rect 11020 7296 11100 7324
rect 10968 7278 11020 7284
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 10888 6905 10916 6938
rect 10874 6896 10930 6905
rect 10874 6831 10930 6840
rect 10980 6798 11008 7142
rect 11072 6866 11100 7296
rect 11256 7177 11284 7346
rect 11348 7342 11376 7822
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11242 7168 11298 7177
rect 11242 7103 11298 7112
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10980 6458 11008 6734
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11072 4162 11100 4558
rect 11150 4312 11206 4321
rect 11348 4282 11376 4626
rect 11150 4247 11206 4256
rect 11336 4276 11388 4282
rect 10980 4134 11100 4162
rect 10980 4010 11008 4134
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10796 3194 10824 3538
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 11164 898 11192 4247
rect 11336 4218 11388 4224
rect 11348 3602 11376 4218
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11348 2582 11376 3538
rect 11440 2650 11468 9415
rect 11808 9042 11836 9998
rect 12084 9654 12112 12679
rect 12176 12306 12204 12922
rect 12268 12782 12296 13126
rect 12256 12776 12308 12782
rect 12256 12718 12308 12724
rect 12360 12594 12388 13398
rect 12544 12832 12572 13806
rect 12636 13025 12664 15966
rect 12728 15960 12756 17031
rect 12808 15972 12860 15978
rect 12728 15932 12808 15960
rect 12808 15914 12860 15920
rect 13004 15858 13032 21490
rect 13084 20392 13136 20398
rect 13084 20334 13136 20340
rect 13096 19718 13124 20334
rect 13084 19712 13136 19718
rect 13084 19654 13136 19660
rect 13096 19514 13124 19654
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 13096 16697 13124 17614
rect 13188 16726 13216 24375
rect 13360 23588 13412 23594
rect 13360 23530 13412 23536
rect 13372 23186 13400 23530
rect 13360 23180 13412 23186
rect 13360 23122 13412 23128
rect 13372 22234 13400 23122
rect 13360 22228 13412 22234
rect 13360 22170 13412 22176
rect 13268 21888 13320 21894
rect 13266 21856 13268 21865
rect 13320 21856 13322 21865
rect 13266 21791 13322 21800
rect 13280 21486 13308 21791
rect 13464 21554 13492 24686
rect 13556 24138 13584 25298
rect 13544 24132 13596 24138
rect 13544 24074 13596 24080
rect 13648 24018 13676 26846
rect 14292 26586 14320 27095
rect 14370 27024 14426 27033
rect 14370 26959 14426 26968
rect 14280 26580 14332 26586
rect 14280 26522 14332 26528
rect 14096 26444 14148 26450
rect 14096 26386 14148 26392
rect 13820 26036 13872 26042
rect 13820 25978 13872 25984
rect 13728 25288 13780 25294
rect 13728 25230 13780 25236
rect 13740 24954 13768 25230
rect 13728 24948 13780 24954
rect 13728 24890 13780 24896
rect 13728 24132 13780 24138
rect 13728 24074 13780 24080
rect 13556 23990 13676 24018
rect 13556 23338 13584 23990
rect 13740 23594 13768 24074
rect 13832 23662 13860 25978
rect 14108 25906 14136 26386
rect 14096 25900 14148 25906
rect 14096 25842 14148 25848
rect 14108 25362 14136 25842
rect 14384 25838 14412 26959
rect 14464 26920 14516 26926
rect 14464 26862 14516 26868
rect 14372 25832 14424 25838
rect 14372 25774 14424 25780
rect 14280 25696 14332 25702
rect 14280 25638 14332 25644
rect 14096 25356 14148 25362
rect 14096 25298 14148 25304
rect 14108 24585 14136 25298
rect 14094 24576 14150 24585
rect 14094 24511 14150 24520
rect 13910 24304 13966 24313
rect 13910 24239 13912 24248
rect 13964 24239 13966 24248
rect 13912 24210 13964 24216
rect 13924 23798 13952 24210
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 14004 23860 14056 23866
rect 14004 23802 14056 23808
rect 13912 23792 13964 23798
rect 13912 23734 13964 23740
rect 14016 23662 14044 23802
rect 13820 23656 13872 23662
rect 13820 23598 13872 23604
rect 14004 23656 14056 23662
rect 14004 23598 14056 23604
rect 13728 23588 13780 23594
rect 13728 23530 13780 23536
rect 13556 23310 13676 23338
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 13556 22778 13584 23122
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 13648 22658 13676 23310
rect 13544 22636 13596 22642
rect 13648 22630 13768 22658
rect 13544 22578 13596 22584
rect 13452 21548 13504 21554
rect 13452 21490 13504 21496
rect 13268 21480 13320 21486
rect 13268 21422 13320 21428
rect 13280 20210 13308 21422
rect 13452 21344 13504 21350
rect 13452 21286 13504 21292
rect 13360 20936 13412 20942
rect 13358 20904 13360 20913
rect 13412 20904 13414 20913
rect 13358 20839 13414 20848
rect 13360 20800 13412 20806
rect 13360 20742 13412 20748
rect 13372 20330 13400 20742
rect 13360 20324 13412 20330
rect 13360 20266 13412 20272
rect 13280 20182 13400 20210
rect 13268 18148 13320 18154
rect 13268 18090 13320 18096
rect 13280 18057 13308 18090
rect 13266 18048 13322 18057
rect 13266 17983 13322 17992
rect 13372 17898 13400 20182
rect 13280 17870 13400 17898
rect 13176 16720 13228 16726
rect 13082 16688 13138 16697
rect 13176 16662 13228 16668
rect 13082 16623 13138 16632
rect 13280 16130 13308 17870
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 13372 17202 13400 17682
rect 13360 17196 13412 17202
rect 13360 17138 13412 17144
rect 13372 17066 13400 17138
rect 13360 17060 13412 17066
rect 13360 17002 13412 17008
rect 13464 16250 13492 21286
rect 13556 21128 13584 22578
rect 13556 21100 13676 21128
rect 13544 20800 13596 20806
rect 13544 20742 13596 20748
rect 13556 20058 13584 20742
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13648 19718 13676 21100
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13648 18970 13676 19654
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13556 18222 13584 18566
rect 13648 18358 13676 18906
rect 13636 18352 13688 18358
rect 13636 18294 13688 18300
rect 13544 18216 13596 18222
rect 13544 18158 13596 18164
rect 13556 17814 13584 18158
rect 13544 17808 13596 17814
rect 13544 17750 13596 17756
rect 13740 17218 13768 22630
rect 13912 22568 13964 22574
rect 13912 22510 13964 22516
rect 14004 22568 14056 22574
rect 14004 22510 14056 22516
rect 13924 22098 13952 22510
rect 13912 22092 13964 22098
rect 13912 22034 13964 22040
rect 14016 21690 14044 22510
rect 14108 22409 14136 24142
rect 14292 23118 14320 25638
rect 14384 25498 14412 25774
rect 14372 25492 14424 25498
rect 14372 25434 14424 25440
rect 14372 24064 14424 24070
rect 14372 24006 14424 24012
rect 14384 23662 14412 24006
rect 14372 23656 14424 23662
rect 14372 23598 14424 23604
rect 14384 23186 14412 23598
rect 14372 23180 14424 23186
rect 14372 23122 14424 23128
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 14292 22642 14320 23054
rect 14280 22636 14332 22642
rect 14280 22578 14332 22584
rect 14094 22400 14150 22409
rect 14094 22335 14150 22344
rect 14004 21684 14056 21690
rect 14004 21626 14056 21632
rect 13912 21480 13964 21486
rect 13912 21422 13964 21428
rect 13924 21010 13952 21422
rect 14096 21344 14148 21350
rect 14094 21312 14096 21321
rect 14148 21312 14150 21321
rect 14094 21247 14150 21256
rect 13912 21004 13964 21010
rect 13912 20946 13964 20952
rect 13820 20868 13872 20874
rect 13820 20810 13872 20816
rect 13832 20602 13860 20810
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 13924 20482 13952 20946
rect 13832 20454 13952 20482
rect 13832 20058 13860 20454
rect 13912 20392 13964 20398
rect 13964 20352 14044 20380
rect 13912 20334 13964 20340
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 13912 19916 13964 19922
rect 13832 19876 13912 19904
rect 13832 19174 13860 19876
rect 13912 19858 13964 19864
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13832 18426 13860 19110
rect 14016 18698 14044 20352
rect 14108 19242 14136 21247
rect 14188 21004 14240 21010
rect 14188 20946 14240 20952
rect 14200 20534 14228 20946
rect 14188 20528 14240 20534
rect 14188 20470 14240 20476
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 14096 19236 14148 19242
rect 14096 19178 14148 19184
rect 14004 18692 14056 18698
rect 14004 18634 14056 18640
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13556 17190 13768 17218
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13280 16102 13492 16130
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 13176 15972 13228 15978
rect 13176 15914 13228 15920
rect 12728 15830 13032 15858
rect 12728 13705 12756 15830
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 13004 15609 13032 15642
rect 13084 15632 13136 15638
rect 12990 15600 13046 15609
rect 13084 15574 13136 15580
rect 12990 15535 13046 15544
rect 12806 15464 12862 15473
rect 12806 15399 12862 15408
rect 12820 14890 12848 15399
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12990 15328 13046 15337
rect 12912 15026 12940 15302
rect 12990 15263 13046 15272
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 12808 14884 12860 14890
rect 12808 14826 12860 14832
rect 13004 14770 13032 15263
rect 12820 14742 13032 14770
rect 12714 13696 12770 13705
rect 12714 13631 12770 13640
rect 12728 13530 12756 13631
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12622 13016 12678 13025
rect 12728 12986 12756 13330
rect 12622 12951 12678 12960
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12728 12889 12756 12922
rect 12714 12880 12770 12889
rect 12544 12804 12664 12832
rect 12714 12815 12770 12824
rect 12532 12708 12584 12714
rect 12636 12696 12664 12804
rect 12636 12668 12756 12696
rect 12532 12650 12584 12656
rect 12360 12566 12480 12594
rect 12452 12374 12480 12566
rect 12440 12368 12492 12374
rect 12440 12310 12492 12316
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12164 11756 12216 11762
rect 12164 11698 12216 11704
rect 12176 11286 12204 11698
rect 12544 11558 12572 12650
rect 12622 12608 12678 12617
rect 12622 12543 12678 12552
rect 12636 12442 12664 12543
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12728 12322 12756 12668
rect 12636 12294 12756 12322
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12164 11280 12216 11286
rect 12164 11222 12216 11228
rect 12438 11112 12494 11121
rect 12438 11047 12494 11056
rect 12452 10266 12480 11047
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12544 10062 12572 10678
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12544 9722 12572 9998
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12072 9648 12124 9654
rect 12072 9590 12124 9596
rect 12636 9178 12664 12294
rect 12714 10840 12770 10849
rect 12714 10775 12770 10784
rect 12728 10742 12756 10775
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12820 10606 12848 14742
rect 12992 14544 13044 14550
rect 12992 14486 13044 14492
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12912 13734 12940 14214
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12912 13394 12940 13670
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 12912 12850 12940 13330
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12900 12708 12952 12714
rect 12900 12650 12952 12656
rect 12912 12617 12940 12650
rect 12898 12608 12954 12617
rect 12898 12543 12954 12552
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11624 8634 11652 8978
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11808 8566 11836 8978
rect 12912 8945 12940 12174
rect 13004 11121 13032 14486
rect 13096 14414 13124 15574
rect 13188 15570 13216 15914
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 13188 15162 13216 15506
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 13372 14618 13400 15982
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13280 14113 13308 14418
rect 13266 14104 13322 14113
rect 13372 14074 13400 14554
rect 13266 14039 13322 14048
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13464 13954 13492 16102
rect 13372 13926 13492 13954
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 13096 12714 13124 13330
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13084 12708 13136 12714
rect 13084 12650 13136 12656
rect 13082 12608 13138 12617
rect 13082 12543 13138 12552
rect 13096 12374 13124 12543
rect 13084 12368 13136 12374
rect 13084 12310 13136 12316
rect 13280 11694 13308 13194
rect 13372 12238 13400 13926
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13464 12782 13492 13466
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13450 12472 13506 12481
rect 13450 12407 13506 12416
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13372 11694 13400 12038
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 12990 11112 13046 11121
rect 13096 11082 13124 11630
rect 13280 11354 13308 11630
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 12990 11047 13046 11056
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 13188 10810 13216 11086
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13464 10282 13492 12407
rect 13372 10254 13492 10282
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 13004 9110 13032 9318
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 13084 8968 13136 8974
rect 12898 8936 12954 8945
rect 13084 8910 13136 8916
rect 12898 8871 12954 8880
rect 12348 8832 12400 8838
rect 12162 8800 12218 8809
rect 12348 8774 12400 8780
rect 12162 8735 12218 8744
rect 11796 8560 11848 8566
rect 11796 8502 11848 8508
rect 11518 6624 11574 6633
rect 11518 6559 11574 6568
rect 11532 3738 11560 6559
rect 12176 4826 12204 8735
rect 12360 6730 12388 8774
rect 12912 8634 12940 8871
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12912 8498 12940 8570
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 13096 8294 13124 8910
rect 13188 8634 13216 8978
rect 13280 8945 13308 10134
rect 13372 8974 13400 10254
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13464 9722 13492 10066
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13360 8968 13412 8974
rect 13266 8936 13322 8945
rect 13360 8910 13412 8916
rect 13266 8871 13322 8880
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13268 8356 13320 8362
rect 13268 8298 13320 8304
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12636 7546 12664 7890
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12728 7478 12756 7890
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12716 7472 12768 7478
rect 12716 7414 12768 7420
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12348 6724 12400 6730
rect 12348 6666 12400 6672
rect 12360 5778 12388 6666
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 11978 4448 12034 4457
rect 11978 4383 12034 4392
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11428 2644 11480 2650
rect 11428 2586 11480 2592
rect 11336 2576 11388 2582
rect 11336 2518 11388 2524
rect 11072 870 11192 898
rect 11072 800 11100 870
rect 11992 800 12020 4383
rect 12452 800 12480 6734
rect 12544 6662 12572 7278
rect 12820 7274 12848 7822
rect 13280 7410 13308 8298
rect 13372 8022 13400 8774
rect 13360 8016 13412 8022
rect 13360 7958 13412 7964
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 12808 7268 12860 7274
rect 12808 7210 12860 7216
rect 13280 7002 13308 7346
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12544 6390 12572 6598
rect 12728 6458 12756 6938
rect 13556 6769 13584 17190
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 13648 16833 13676 16934
rect 13634 16824 13690 16833
rect 13634 16759 13690 16768
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13648 16182 13676 16526
rect 13636 16176 13688 16182
rect 13636 16118 13688 16124
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 13648 15162 13676 15506
rect 13636 15156 13688 15162
rect 13636 15098 13688 15104
rect 13648 14550 13676 15098
rect 13832 15065 13860 18362
rect 13924 18222 13952 18566
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 13818 15056 13874 15065
rect 13818 14991 13874 15000
rect 13924 14906 13952 15982
rect 14016 15337 14044 18634
rect 14108 16794 14136 19178
rect 14200 19009 14228 19246
rect 14186 19000 14242 19009
rect 14186 18935 14242 18944
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14188 18148 14240 18154
rect 14188 18090 14240 18096
rect 14200 17338 14228 18090
rect 14292 17542 14320 18770
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14292 17338 14320 17478
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 14280 17332 14332 17338
rect 14280 17274 14332 17280
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 14200 16658 14228 17274
rect 14384 17202 14412 23122
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14280 16720 14332 16726
rect 14280 16662 14332 16668
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14002 15328 14058 15337
rect 14002 15263 14058 15272
rect 13740 14878 13952 14906
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13634 14376 13690 14385
rect 13634 14311 13690 14320
rect 13648 13138 13676 14311
rect 13740 13938 13768 14878
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13726 13832 13782 13841
rect 13726 13767 13782 13776
rect 13740 13734 13768 13767
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13728 13388 13780 13394
rect 13832 13376 13860 14758
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 13924 13530 13952 14350
rect 14016 14346 14044 14894
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13780 13348 13860 13376
rect 13728 13330 13780 13336
rect 13648 13110 13768 13138
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13648 11778 13676 12922
rect 13740 12617 13768 13110
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 13726 12608 13782 12617
rect 13726 12543 13782 12552
rect 13648 11762 13860 11778
rect 13648 11756 13872 11762
rect 13648 11750 13820 11756
rect 13820 11698 13872 11704
rect 13634 11248 13690 11257
rect 13924 11234 13952 12786
rect 14016 12617 14044 14282
rect 14108 13870 14136 14554
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 14108 13462 14136 13806
rect 14200 13734 14228 15846
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 14096 13456 14148 13462
rect 14096 13398 14148 13404
rect 14188 13388 14240 13394
rect 14188 13330 14240 13336
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14002 12608 14058 12617
rect 14002 12543 14058 12552
rect 14108 12374 14136 12718
rect 14200 12442 14228 13330
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14096 12368 14148 12374
rect 14094 12336 14096 12345
rect 14148 12336 14150 12345
rect 14094 12271 14150 12280
rect 14108 12245 14136 12271
rect 14292 11801 14320 16662
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 14384 15201 14412 16594
rect 14370 15192 14426 15201
rect 14370 15127 14426 15136
rect 14370 13696 14426 13705
rect 14370 13631 14426 13640
rect 14384 13530 14412 13631
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14278 11792 14334 11801
rect 14278 11727 14334 11736
rect 13832 11218 13952 11234
rect 13634 11183 13636 11192
rect 13688 11183 13690 11192
rect 13820 11212 13952 11218
rect 13636 11154 13688 11160
rect 13872 11206 13952 11212
rect 13820 11154 13872 11160
rect 13648 10742 13676 11154
rect 13832 11098 13860 11154
rect 13740 11070 13860 11098
rect 13636 10736 13688 10742
rect 13636 10678 13688 10684
rect 13740 10266 13768 11070
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13832 10146 13860 10678
rect 13740 10118 13860 10146
rect 13740 9042 13768 10118
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13832 8650 13860 9998
rect 13924 9466 13952 10746
rect 14384 10198 14412 12582
rect 14476 10606 14504 26862
rect 14660 26042 14688 33351
rect 14740 30864 14792 30870
rect 14740 30806 14792 30812
rect 14752 30190 14780 30806
rect 14740 30184 14792 30190
rect 14740 30126 14792 30132
rect 15028 28121 15056 37266
rect 15304 37262 15332 38150
rect 15566 37904 15622 37913
rect 15566 37839 15622 37848
rect 15580 37330 15608 37839
rect 15672 37369 15700 40996
rect 15752 39432 15804 39438
rect 15752 39374 15804 39380
rect 15764 38962 15792 39374
rect 15752 38956 15804 38962
rect 15752 38898 15804 38904
rect 15658 37360 15714 37369
rect 15568 37324 15620 37330
rect 15658 37295 15714 37304
rect 15568 37266 15620 37272
rect 15292 37256 15344 37262
rect 15292 37198 15344 37204
rect 15304 36582 15332 37198
rect 15580 36922 15608 37266
rect 15750 37224 15806 37233
rect 15750 37159 15806 37168
rect 15568 36916 15620 36922
rect 15568 36858 15620 36864
rect 15292 36576 15344 36582
rect 15292 36518 15344 36524
rect 15292 34536 15344 34542
rect 15292 34478 15344 34484
rect 15108 34400 15160 34406
rect 15108 34342 15160 34348
rect 15120 34202 15148 34342
rect 15108 34196 15160 34202
rect 15108 34138 15160 34144
rect 15108 33992 15160 33998
rect 15108 33934 15160 33940
rect 15120 29034 15148 33934
rect 15304 32881 15332 34478
rect 15764 34202 15792 37159
rect 15936 35488 15988 35494
rect 15936 35430 15988 35436
rect 15752 34196 15804 34202
rect 15752 34138 15804 34144
rect 15660 34060 15712 34066
rect 15660 34002 15712 34008
rect 15672 33046 15700 34002
rect 15476 33040 15528 33046
rect 15476 32982 15528 32988
rect 15660 33040 15712 33046
rect 15660 32982 15712 32988
rect 15290 32872 15346 32881
rect 15290 32807 15346 32816
rect 15292 32360 15344 32366
rect 15292 32302 15344 32308
rect 15304 30258 15332 32302
rect 15384 32020 15436 32026
rect 15384 31962 15436 31968
rect 15396 31249 15424 31962
rect 15382 31240 15438 31249
rect 15382 31175 15438 31184
rect 15488 30977 15516 32982
rect 15844 32972 15896 32978
rect 15844 32914 15896 32920
rect 15660 32904 15712 32910
rect 15658 32872 15660 32881
rect 15712 32872 15714 32881
rect 15856 32858 15884 32914
rect 15658 32807 15714 32816
rect 15764 32830 15884 32858
rect 15764 31958 15792 32830
rect 15752 31952 15804 31958
rect 15750 31920 15752 31929
rect 15804 31920 15806 31929
rect 15750 31855 15806 31864
rect 15474 30968 15530 30977
rect 15474 30903 15530 30912
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 15568 30728 15620 30734
rect 15568 30670 15620 30676
rect 15292 30252 15344 30258
rect 15292 30194 15344 30200
rect 15488 29850 15516 30670
rect 15580 30394 15608 30670
rect 15568 30388 15620 30394
rect 15620 30348 15700 30376
rect 15568 30330 15620 30336
rect 15476 29844 15528 29850
rect 15476 29786 15528 29792
rect 15488 29646 15516 29786
rect 15476 29640 15528 29646
rect 15198 29608 15254 29617
rect 15476 29582 15528 29588
rect 15198 29543 15254 29552
rect 15212 29306 15240 29543
rect 15200 29300 15252 29306
rect 15200 29242 15252 29248
rect 15108 29028 15160 29034
rect 15108 28970 15160 28976
rect 15384 28620 15436 28626
rect 15384 28562 15436 28568
rect 15014 28112 15070 28121
rect 15014 28047 15070 28056
rect 15396 27878 15424 28562
rect 15488 28558 15516 29582
rect 15476 28552 15528 28558
rect 15476 28494 15528 28500
rect 15488 27878 15516 28494
rect 15384 27872 15436 27878
rect 15384 27814 15436 27820
rect 15476 27872 15528 27878
rect 15476 27814 15528 27820
rect 15292 27532 15344 27538
rect 15292 27474 15344 27480
rect 15016 27056 15068 27062
rect 15016 26998 15068 27004
rect 14648 26036 14700 26042
rect 14648 25978 14700 25984
rect 15028 25498 15056 26998
rect 15304 26858 15332 27474
rect 15292 26852 15344 26858
rect 15292 26794 15344 26800
rect 15304 26450 15332 26794
rect 15292 26444 15344 26450
rect 15292 26386 15344 26392
rect 15108 26308 15160 26314
rect 15108 26250 15160 26256
rect 15120 25906 15148 26250
rect 15304 26042 15332 26386
rect 15292 26036 15344 26042
rect 15292 25978 15344 25984
rect 15396 25922 15424 27814
rect 15476 27328 15528 27334
rect 15476 27270 15528 27276
rect 15488 27033 15516 27270
rect 15474 27024 15530 27033
rect 15474 26959 15476 26968
rect 15528 26959 15530 26968
rect 15476 26930 15528 26936
rect 15488 26899 15516 26930
rect 15568 26784 15620 26790
rect 15568 26726 15620 26732
rect 15108 25900 15160 25906
rect 15108 25842 15160 25848
rect 15304 25894 15424 25922
rect 15016 25492 15068 25498
rect 15016 25434 15068 25440
rect 14646 24168 14702 24177
rect 14646 24103 14702 24112
rect 14660 23322 14688 24103
rect 14832 23724 14884 23730
rect 14832 23666 14884 23672
rect 14738 23624 14794 23633
rect 14738 23559 14794 23568
rect 14648 23316 14700 23322
rect 14648 23258 14700 23264
rect 14556 22976 14608 22982
rect 14556 22918 14608 22924
rect 14568 19854 14596 22918
rect 14646 22128 14702 22137
rect 14646 22063 14648 22072
rect 14700 22063 14702 22072
rect 14648 22034 14700 22040
rect 14648 21072 14700 21078
rect 14646 21040 14648 21049
rect 14700 21040 14702 21049
rect 14752 21026 14780 23559
rect 14844 21146 14872 23666
rect 15120 23526 15148 25842
rect 15200 25832 15252 25838
rect 15200 25774 15252 25780
rect 15108 23520 15160 23526
rect 15108 23462 15160 23468
rect 15120 22658 15148 23462
rect 15212 22778 15240 25774
rect 15304 25106 15332 25894
rect 15384 25764 15436 25770
rect 15384 25706 15436 25712
rect 15396 25226 15424 25706
rect 15384 25220 15436 25226
rect 15384 25162 15436 25168
rect 15304 25078 15424 25106
rect 15290 24848 15346 24857
rect 15290 24783 15292 24792
rect 15344 24783 15346 24792
rect 15292 24754 15344 24760
rect 15396 23905 15424 25078
rect 15476 24608 15528 24614
rect 15476 24550 15528 24556
rect 15488 24206 15516 24550
rect 15476 24200 15528 24206
rect 15476 24142 15528 24148
rect 15382 23896 15438 23905
rect 15382 23831 15438 23840
rect 15384 23792 15436 23798
rect 15384 23734 15436 23740
rect 15290 23080 15346 23089
rect 15290 23015 15346 23024
rect 15200 22772 15252 22778
rect 15200 22714 15252 22720
rect 14924 22636 14976 22642
rect 15120 22630 15240 22658
rect 14924 22578 14976 22584
rect 14832 21140 14884 21146
rect 14832 21082 14884 21088
rect 14752 20998 14872 21026
rect 14646 20975 14702 20984
rect 14740 20936 14792 20942
rect 14740 20878 14792 20884
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14568 18630 14596 19790
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 14660 19417 14688 19654
rect 14646 19408 14702 19417
rect 14646 19343 14702 19352
rect 14752 19310 14780 20878
rect 14740 19304 14792 19310
rect 14740 19246 14792 19252
rect 14646 19136 14702 19145
rect 14646 19071 14702 19080
rect 14660 18970 14688 19071
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 14556 18624 14608 18630
rect 14556 18566 14608 18572
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 14752 18057 14780 18158
rect 14738 18048 14794 18057
rect 14738 17983 14794 17992
rect 14740 17672 14792 17678
rect 14738 17640 14740 17649
rect 14792 17640 14794 17649
rect 14738 17575 14794 17584
rect 14844 17542 14872 20998
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14740 17264 14792 17270
rect 14936 17218 14964 22578
rect 15108 22568 15160 22574
rect 15108 22510 15160 22516
rect 15016 21888 15068 21894
rect 15016 21830 15068 21836
rect 15028 21554 15056 21830
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 15120 21350 15148 22510
rect 15108 21344 15160 21350
rect 15212 21321 15240 22630
rect 15108 21286 15160 21292
rect 15198 21312 15254 21321
rect 15198 21247 15254 21256
rect 15108 21140 15160 21146
rect 15108 21082 15160 21088
rect 15016 17536 15068 17542
rect 15016 17478 15068 17484
rect 14740 17206 14792 17212
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 14556 17128 14608 17134
rect 14554 17096 14556 17105
rect 14608 17096 14610 17105
rect 14554 17031 14610 17040
rect 14556 16176 14608 16182
rect 14556 16118 14608 16124
rect 14568 14385 14596 16118
rect 14554 14376 14610 14385
rect 14554 14311 14610 14320
rect 14554 14104 14610 14113
rect 14554 14039 14610 14048
rect 14568 12782 14596 14039
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14554 12608 14610 12617
rect 14554 12543 14610 12552
rect 14568 12306 14596 12543
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14568 11898 14596 12242
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14660 10810 14688 17138
rect 14752 16794 14780 17206
rect 14844 17190 14964 17218
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 14740 15564 14792 15570
rect 14740 15506 14792 15512
rect 14752 15366 14780 15506
rect 14740 15360 14792 15366
rect 14738 15328 14740 15337
rect 14792 15328 14794 15337
rect 14738 15263 14794 15272
rect 14738 15056 14794 15065
rect 14738 14991 14794 15000
rect 14752 14521 14780 14991
rect 14738 14512 14794 14521
rect 14738 14447 14794 14456
rect 14752 13394 14780 14447
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14740 13252 14792 13258
rect 14740 13194 14792 13200
rect 14752 12782 14780 13194
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 14752 12238 14780 12718
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14752 11762 14780 12038
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14752 11354 14780 11698
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14372 10192 14424 10198
rect 14372 10134 14424 10140
rect 14476 10130 14504 10542
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14096 9512 14148 9518
rect 13924 9460 14096 9466
rect 13924 9454 14148 9460
rect 13924 9438 14136 9454
rect 14292 9450 14320 9862
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14280 9444 14332 9450
rect 13924 9178 13952 9438
rect 14280 9386 14332 9392
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 13740 8622 13860 8650
rect 14292 8634 14320 9386
rect 14384 8838 14412 9590
rect 14844 9042 14872 17190
rect 15028 17134 15056 17478
rect 15016 17128 15068 17134
rect 14922 17096 14978 17105
rect 15016 17070 15068 17076
rect 14922 17031 14978 17040
rect 14936 16998 14964 17031
rect 14924 16992 14976 16998
rect 14924 16934 14976 16940
rect 15028 16726 15056 17070
rect 15016 16720 15068 16726
rect 15016 16662 15068 16668
rect 15120 16182 15148 21082
rect 15212 18986 15240 21247
rect 15304 19854 15332 23015
rect 15396 21146 15424 23734
rect 15488 23594 15516 24142
rect 15476 23588 15528 23594
rect 15476 23530 15528 23536
rect 15488 21486 15516 23530
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15384 21140 15436 21146
rect 15384 21082 15436 21088
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 15396 20262 15424 20946
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15396 19922 15424 20198
rect 15384 19916 15436 19922
rect 15384 19858 15436 19864
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 15396 19156 15424 19858
rect 15488 19718 15516 21422
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15476 19168 15528 19174
rect 15396 19136 15476 19156
rect 15528 19136 15530 19145
rect 15396 19128 15474 19136
rect 15474 19071 15530 19080
rect 15212 18958 15516 18986
rect 15384 18624 15436 18630
rect 15384 18566 15436 18572
rect 15198 18320 15254 18329
rect 15198 18255 15254 18264
rect 15212 16182 15240 18255
rect 15396 17882 15424 18566
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15108 16176 15160 16182
rect 15108 16118 15160 16124
rect 15200 16176 15252 16182
rect 15200 16118 15252 16124
rect 15212 15994 15240 16118
rect 14936 15966 15240 15994
rect 14936 14618 14964 15966
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15212 15745 15240 15846
rect 15198 15736 15254 15745
rect 15198 15671 15254 15680
rect 15304 15570 15332 17070
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15028 15434 15240 15450
rect 15028 15428 15252 15434
rect 15028 15422 15200 15428
rect 15028 14793 15056 15422
rect 15200 15370 15252 15376
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 15014 14784 15070 14793
rect 15014 14719 15070 14728
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14924 13796 14976 13802
rect 14924 13738 14976 13744
rect 14936 12458 14964 13738
rect 15028 12714 15056 14719
rect 15120 14634 15148 15302
rect 15304 15162 15332 15506
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15304 14940 15332 15098
rect 15384 14952 15436 14958
rect 15304 14912 15384 14940
rect 15384 14894 15436 14900
rect 15488 14770 15516 18958
rect 15580 17921 15608 26726
rect 15672 23322 15700 30348
rect 15752 29096 15804 29102
rect 15752 29038 15804 29044
rect 15764 27062 15792 29038
rect 15844 29028 15896 29034
rect 15844 28970 15896 28976
rect 15752 27056 15804 27062
rect 15752 26998 15804 27004
rect 15856 26926 15884 28970
rect 15844 26920 15896 26926
rect 15844 26862 15896 26868
rect 15752 26240 15804 26246
rect 15752 26182 15804 26188
rect 15764 25906 15792 26182
rect 15948 26042 15976 35430
rect 16028 32360 16080 32366
rect 16132 32348 16160 40996
rect 16210 36680 16266 36689
rect 16210 36615 16266 36624
rect 16224 33658 16252 36615
rect 16488 36576 16540 36582
rect 16488 36518 16540 36524
rect 16302 36408 16358 36417
rect 16302 36343 16358 36352
rect 16212 33652 16264 33658
rect 16212 33594 16264 33600
rect 16316 32502 16344 36343
rect 16500 36242 16528 36518
rect 16592 36394 16620 40996
rect 17316 38412 17368 38418
rect 17316 38354 17368 38360
rect 17224 38344 17276 38350
rect 17224 38286 17276 38292
rect 17236 37670 17264 38286
rect 17328 37806 17356 38354
rect 17316 37800 17368 37806
rect 17314 37768 17316 37777
rect 17368 37768 17370 37777
rect 17314 37703 17370 37712
rect 17224 37664 17276 37670
rect 17224 37606 17276 37612
rect 16592 36366 16804 36394
rect 16488 36236 16540 36242
rect 16488 36178 16540 36184
rect 16500 35562 16528 36178
rect 16672 36168 16724 36174
rect 16672 36110 16724 36116
rect 16488 35556 16540 35562
rect 16488 35498 16540 35504
rect 16684 35494 16712 36110
rect 16672 35488 16724 35494
rect 16672 35430 16724 35436
rect 16488 34400 16540 34406
rect 16488 34342 16540 34348
rect 16500 34066 16528 34342
rect 16488 34060 16540 34066
rect 16488 34002 16540 34008
rect 16672 33856 16724 33862
rect 16672 33798 16724 33804
rect 16684 33522 16712 33798
rect 16672 33516 16724 33522
rect 16672 33458 16724 33464
rect 16684 32978 16712 33458
rect 16672 32972 16724 32978
rect 16672 32914 16724 32920
rect 16488 32904 16540 32910
rect 16488 32846 16540 32852
rect 16500 32570 16528 32846
rect 16488 32564 16540 32570
rect 16488 32506 16540 32512
rect 16304 32496 16356 32502
rect 16304 32438 16356 32444
rect 16132 32320 16528 32348
rect 16028 32302 16080 32308
rect 16040 32026 16068 32302
rect 16028 32020 16080 32026
rect 16028 31962 16080 31968
rect 16396 31816 16448 31822
rect 16396 31758 16448 31764
rect 16120 31748 16172 31754
rect 16120 31690 16172 31696
rect 16028 29028 16080 29034
rect 16028 28970 16080 28976
rect 15936 26036 15988 26042
rect 15936 25978 15988 25984
rect 15752 25900 15804 25906
rect 15752 25842 15804 25848
rect 15936 25832 15988 25838
rect 15936 25774 15988 25780
rect 15948 25498 15976 25774
rect 15936 25492 15988 25498
rect 15936 25434 15988 25440
rect 15936 25288 15988 25294
rect 15936 25230 15988 25236
rect 15750 24848 15806 24857
rect 15750 24783 15806 24792
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15660 21480 15712 21486
rect 15660 21422 15712 21428
rect 15672 20534 15700 21422
rect 15660 20528 15712 20534
rect 15660 20470 15712 20476
rect 15660 19780 15712 19786
rect 15660 19722 15712 19728
rect 15566 17912 15622 17921
rect 15566 17847 15622 17856
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15580 16114 15608 16594
rect 15672 16561 15700 19722
rect 15658 16552 15714 16561
rect 15658 16487 15714 16496
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15580 15978 15608 16050
rect 15568 15972 15620 15978
rect 15568 15914 15620 15920
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 15568 14884 15620 14890
rect 15568 14826 15620 14832
rect 15304 14742 15516 14770
rect 15120 14618 15240 14634
rect 15120 14612 15252 14618
rect 15120 14606 15200 14612
rect 15200 14554 15252 14560
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15108 14000 15160 14006
rect 15108 13942 15160 13948
rect 15120 13530 15148 13942
rect 15212 13870 15240 14418
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15198 13152 15254 13161
rect 15120 12986 15148 13126
rect 15198 13087 15254 13096
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15106 12880 15162 12889
rect 15106 12815 15108 12824
rect 15160 12815 15162 12824
rect 15108 12786 15160 12792
rect 15016 12708 15068 12714
rect 15016 12650 15068 12656
rect 14936 12430 15148 12458
rect 14924 12368 14976 12374
rect 14924 12310 14976 12316
rect 14936 11694 14964 12310
rect 14924 11688 14976 11694
rect 14924 11630 14976 11636
rect 15120 11218 15148 12430
rect 15212 11354 15240 13087
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15120 10810 15148 11154
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15120 10470 15148 10746
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 15198 10296 15254 10305
rect 15198 10231 15254 10240
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 15028 9081 15056 9386
rect 15014 9072 15070 9081
rect 14832 9036 14884 9042
rect 15014 9007 15070 9016
rect 14832 8978 14884 8984
rect 14372 8832 14424 8838
rect 14370 8800 14372 8809
rect 14424 8800 14426 8809
rect 14370 8735 14426 8744
rect 13740 8430 13768 8622
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13648 8090 13676 8298
rect 13832 8090 13860 8622
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14844 8498 14872 8978
rect 15212 8974 15240 10231
rect 15304 10130 15332 14742
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15382 14104 15438 14113
rect 15382 14039 15384 14048
rect 15436 14039 15438 14048
rect 15384 14010 15436 14016
rect 15488 13802 15516 14350
rect 15580 14249 15608 14826
rect 15672 14550 15700 14894
rect 15660 14544 15712 14550
rect 15660 14486 15712 14492
rect 15566 14240 15622 14249
rect 15566 14175 15622 14184
rect 15476 13796 15528 13802
rect 15476 13738 15528 13744
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15396 12850 15424 13330
rect 15488 13258 15516 13738
rect 15476 13252 15528 13258
rect 15476 13194 15528 13200
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15396 12646 15424 12786
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15396 12306 15424 12582
rect 15488 12442 15516 12582
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15384 11688 15436 11694
rect 15382 11656 15384 11665
rect 15436 11656 15438 11665
rect 15382 11591 15438 11600
rect 15396 10674 15424 11591
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 15304 9722 15332 10066
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15396 9110 15424 10610
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 15200 8968 15252 8974
rect 15120 8916 15200 8922
rect 15120 8910 15252 8916
rect 15120 8894 15240 8910
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 14646 8392 14702 8401
rect 14646 8327 14648 8336
rect 14700 8327 14702 8336
rect 14648 8298 14700 8304
rect 15120 8090 15148 8894
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15212 7954 15240 8774
rect 15396 8634 15424 9046
rect 15672 9042 15700 9862
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15488 8634 15516 8978
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15764 8498 15792 24783
rect 15948 23866 15976 25230
rect 15936 23860 15988 23866
rect 15936 23802 15988 23808
rect 15948 23254 15976 23802
rect 15936 23248 15988 23254
rect 15936 23190 15988 23196
rect 15844 23112 15896 23118
rect 15844 23054 15896 23060
rect 15856 22234 15884 23054
rect 15844 22228 15896 22234
rect 15844 22170 15896 22176
rect 15856 21418 15884 22170
rect 15948 22166 15976 23190
rect 16040 22234 16068 28970
rect 16132 25945 16160 31690
rect 16408 31414 16436 31758
rect 16396 31408 16448 31414
rect 16394 31376 16396 31385
rect 16448 31376 16450 31385
rect 16394 31311 16450 31320
rect 16396 31272 16448 31278
rect 16396 31214 16448 31220
rect 16408 30122 16436 31214
rect 16396 30116 16448 30122
rect 16396 30058 16448 30064
rect 16394 30016 16450 30025
rect 16394 29951 16450 29960
rect 16304 29708 16356 29714
rect 16304 29650 16356 29656
rect 16316 29306 16344 29650
rect 16304 29300 16356 29306
rect 16304 29242 16356 29248
rect 16316 29034 16344 29242
rect 16304 29028 16356 29034
rect 16304 28970 16356 28976
rect 16408 28529 16436 29951
rect 16394 28520 16450 28529
rect 16394 28455 16450 28464
rect 16304 27872 16356 27878
rect 16304 27814 16356 27820
rect 16316 27470 16344 27814
rect 16396 27532 16448 27538
rect 16396 27474 16448 27480
rect 16304 27464 16356 27470
rect 16304 27406 16356 27412
rect 16408 26586 16436 27474
rect 16396 26580 16448 26586
rect 16396 26522 16448 26528
rect 16396 26036 16448 26042
rect 16396 25978 16448 25984
rect 16118 25936 16174 25945
rect 16118 25871 16174 25880
rect 16304 25220 16356 25226
rect 16304 25162 16356 25168
rect 16212 25152 16264 25158
rect 16212 25094 16264 25100
rect 16224 24818 16252 25094
rect 16212 24812 16264 24818
rect 16212 24754 16264 24760
rect 16224 24342 16252 24754
rect 16316 24750 16344 25162
rect 16304 24744 16356 24750
rect 16304 24686 16356 24692
rect 16212 24336 16264 24342
rect 16212 24278 16264 24284
rect 16120 24268 16172 24274
rect 16120 24210 16172 24216
rect 16132 24177 16160 24210
rect 16118 24168 16174 24177
rect 16118 24103 16174 24112
rect 16120 23588 16172 23594
rect 16120 23530 16172 23536
rect 16132 23186 16160 23530
rect 16120 23180 16172 23186
rect 16120 23122 16172 23128
rect 16304 23112 16356 23118
rect 16302 23080 16304 23089
rect 16356 23080 16358 23089
rect 16302 23015 16358 23024
rect 16118 22536 16174 22545
rect 16316 22506 16344 23015
rect 16118 22471 16174 22480
rect 16212 22500 16264 22506
rect 16028 22228 16080 22234
rect 16028 22170 16080 22176
rect 15936 22160 15988 22166
rect 15936 22102 15988 22108
rect 15948 21690 15976 22102
rect 16028 22024 16080 22030
rect 16028 21966 16080 21972
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 15844 21412 15896 21418
rect 15844 21354 15896 21360
rect 15936 21344 15988 21350
rect 15936 21286 15988 21292
rect 15844 20800 15896 20806
rect 15844 20742 15896 20748
rect 15856 20398 15884 20742
rect 15844 20392 15896 20398
rect 15844 20334 15896 20340
rect 15856 19990 15884 20334
rect 15844 19984 15896 19990
rect 15844 19926 15896 19932
rect 15856 18902 15884 19926
rect 15948 19378 15976 21286
rect 16040 21146 16068 21966
rect 16028 21140 16080 21146
rect 16028 21082 16080 21088
rect 16026 20496 16082 20505
rect 16026 20431 16082 20440
rect 16040 20398 16068 20431
rect 16028 20392 16080 20398
rect 16028 20334 16080 20340
rect 16028 19440 16080 19446
rect 16028 19382 16080 19388
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 16040 18970 16068 19382
rect 16028 18964 16080 18970
rect 16028 18906 16080 18912
rect 15844 18896 15896 18902
rect 15844 18838 15896 18844
rect 15856 18426 15884 18838
rect 16028 18828 16080 18834
rect 16028 18770 16080 18776
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 16040 18086 16068 18770
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 16040 17678 16068 18022
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 16028 17672 16080 17678
rect 16028 17614 16080 17620
rect 15856 17241 15884 17614
rect 15842 17232 15898 17241
rect 15842 17167 15898 17176
rect 15934 17096 15990 17105
rect 15934 17031 15990 17040
rect 15948 14550 15976 17031
rect 16040 16794 16068 17614
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 16132 16130 16160 22471
rect 16212 22442 16264 22448
rect 16304 22500 16356 22506
rect 16304 22442 16356 22448
rect 16224 22030 16252 22442
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 16304 21956 16356 21962
rect 16304 21898 16356 21904
rect 16212 19712 16264 19718
rect 16212 19654 16264 19660
rect 16224 19514 16252 19654
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16316 19446 16344 21898
rect 16304 19440 16356 19446
rect 16304 19382 16356 19388
rect 16302 19000 16358 19009
rect 16212 18964 16264 18970
rect 16302 18935 16358 18944
rect 16212 18906 16264 18912
rect 16224 18873 16252 18906
rect 16210 18864 16266 18873
rect 16210 18799 16266 18808
rect 16212 16448 16264 16454
rect 16212 16390 16264 16396
rect 16040 16102 16160 16130
rect 16040 15094 16068 16102
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 16132 15706 16160 15982
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 16224 15638 16252 16390
rect 16212 15632 16264 15638
rect 16212 15574 16264 15580
rect 16224 15162 16252 15574
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 16028 15088 16080 15094
rect 16316 15042 16344 18935
rect 16028 15030 16080 15036
rect 16132 15014 16344 15042
rect 15936 14544 15988 14550
rect 15936 14486 15988 14492
rect 15948 14074 15976 14486
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 15844 13728 15896 13734
rect 15844 13670 15896 13676
rect 15856 12782 15884 13670
rect 15948 13546 15976 14010
rect 15948 13518 16068 13546
rect 16040 13462 16068 13518
rect 15936 13456 15988 13462
rect 15936 13398 15988 13404
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 15948 12918 15976 13398
rect 15936 12912 15988 12918
rect 16040 12889 16068 13398
rect 15936 12854 15988 12860
rect 16026 12880 16082 12889
rect 16026 12815 16082 12824
rect 15844 12776 15896 12782
rect 16132 12764 16160 15014
rect 16304 14952 16356 14958
rect 16304 14894 16356 14900
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16224 13870 16252 14554
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16210 13560 16266 13569
rect 16210 13495 16266 13504
rect 15844 12718 15896 12724
rect 15948 12736 16160 12764
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 15856 10198 15884 11154
rect 15948 10606 15976 12736
rect 16028 12640 16080 12646
rect 16028 12582 16080 12588
rect 16040 11762 16068 12582
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16132 11830 16160 12038
rect 16120 11824 16172 11830
rect 16120 11766 16172 11772
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 16040 11218 16068 11698
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 16040 10810 16068 11154
rect 16132 10810 16160 11154
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 15948 10198 15976 10542
rect 16040 10266 16068 10746
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 15844 10192 15896 10198
rect 15842 10160 15844 10169
rect 15936 10192 15988 10198
rect 15896 10160 15898 10169
rect 15936 10134 15988 10140
rect 15842 10095 15898 10104
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16026 8664 16082 8673
rect 16026 8599 16082 8608
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 16040 8294 16068 8599
rect 16132 8537 16160 9318
rect 16118 8528 16174 8537
rect 16118 8463 16174 8472
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 15200 7948 15252 7954
rect 15200 7890 15252 7896
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 15028 7546 15056 7822
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 16040 7478 16068 8230
rect 16028 7472 16080 7478
rect 16028 7414 16080 7420
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13910 7168 13966 7177
rect 13648 6866 13676 7142
rect 13910 7103 13966 7112
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13542 6760 13598 6769
rect 13542 6695 13598 6704
rect 12898 6624 12954 6633
rect 12898 6559 12954 6568
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12532 6384 12584 6390
rect 12532 6326 12584 6332
rect 12544 5710 12572 6326
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 12544 5302 12572 5646
rect 12820 5370 12848 5714
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 12544 4690 12572 5238
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 12530 2680 12586 2689
rect 12530 2615 12532 2624
rect 12584 2615 12586 2624
rect 12532 2586 12584 2592
rect 12912 800 12940 6559
rect 13648 6458 13676 6802
rect 13820 6792 13872 6798
rect 13818 6760 13820 6769
rect 13872 6760 13874 6769
rect 13818 6695 13874 6704
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13832 6254 13860 6695
rect 13924 6458 13952 7103
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 14016 6497 14044 6734
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14002 6488 14058 6497
rect 13912 6452 13964 6458
rect 14002 6423 14058 6432
rect 13912 6394 13964 6400
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 14016 6186 14044 6423
rect 14568 6361 14596 6598
rect 14554 6352 14610 6361
rect 14554 6287 14610 6296
rect 14568 6254 14596 6287
rect 15120 6254 15148 6666
rect 15936 6384 15988 6390
rect 15936 6326 15988 6332
rect 14556 6248 14608 6254
rect 14370 6216 14426 6225
rect 14004 6180 14056 6186
rect 14556 6190 14608 6196
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 14370 6151 14426 6160
rect 14004 6122 14056 6128
rect 14384 6118 14412 6151
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 14752 5914 14780 6190
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 15948 5778 15976 6326
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 15948 5302 15976 5714
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 16040 5370 16068 5646
rect 16028 5364 16080 5370
rect 16028 5306 16080 5312
rect 15936 5296 15988 5302
rect 15936 5238 15988 5244
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13832 800 13860 4762
rect 16040 4690 16068 5306
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 16132 4321 16160 6734
rect 16224 5273 16252 13495
rect 16316 12986 16344 14894
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16304 10192 16356 10198
rect 16304 10134 16356 10140
rect 16316 8498 16344 10134
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16316 7954 16344 8434
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16316 7546 16344 7890
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16210 5264 16266 5273
rect 16210 5199 16266 5208
rect 16118 4312 16174 4321
rect 16118 4247 16174 4256
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 14278 3360 14334 3369
rect 14278 3295 14334 3304
rect 14292 800 14320 3295
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 14752 800 14780 3130
rect 15396 3058 15424 3538
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15580 3194 15608 3470
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15658 3088 15714 3097
rect 15384 3052 15436 3058
rect 15658 3023 15660 3032
rect 15384 2994 15436 3000
rect 15712 3023 15714 3032
rect 15660 2994 15712 3000
rect 15396 2650 15424 2994
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 15660 1828 15712 1834
rect 15660 1770 15712 1776
rect 15672 800 15700 1770
rect 16132 800 16160 2382
rect 16408 1834 16436 25978
rect 16500 22681 16528 32320
rect 16578 32328 16634 32337
rect 16578 32263 16634 32272
rect 16592 31958 16620 32263
rect 16580 31952 16632 31958
rect 16580 31894 16632 31900
rect 16672 31272 16724 31278
rect 16672 31214 16724 31220
rect 16684 30938 16712 31214
rect 16672 30932 16724 30938
rect 16672 30874 16724 30880
rect 16670 29064 16726 29073
rect 16670 28999 16726 29008
rect 16684 28762 16712 28999
rect 16672 28756 16724 28762
rect 16672 28698 16724 28704
rect 16580 26852 16632 26858
rect 16580 26794 16632 26800
rect 16592 25362 16620 26794
rect 16672 26580 16724 26586
rect 16672 26522 16724 26528
rect 16684 25430 16712 26522
rect 16776 26518 16804 36366
rect 17132 34060 17184 34066
rect 17132 34002 17184 34008
rect 17144 33454 17172 34002
rect 16948 33448 17000 33454
rect 16948 33390 17000 33396
rect 17132 33448 17184 33454
rect 17132 33390 17184 33396
rect 16960 33114 16988 33390
rect 17144 33318 17172 33390
rect 17132 33312 17184 33318
rect 17130 33280 17132 33289
rect 17184 33280 17186 33289
rect 17130 33215 17186 33224
rect 17144 33189 17172 33215
rect 16948 33108 17000 33114
rect 16948 33050 17000 33056
rect 17512 32178 17540 40996
rect 17868 38752 17920 38758
rect 17868 38694 17920 38700
rect 17592 37324 17644 37330
rect 17592 37266 17644 37272
rect 17328 32150 17540 32178
rect 17040 31884 17092 31890
rect 17040 31826 17092 31832
rect 17224 31884 17276 31890
rect 17224 31826 17276 31832
rect 17052 31482 17080 31826
rect 17040 31476 17092 31482
rect 17040 31418 17092 31424
rect 16948 31272 17000 31278
rect 16948 31214 17000 31220
rect 16856 27940 16908 27946
rect 16856 27882 16908 27888
rect 16764 26512 16816 26518
rect 16764 26454 16816 26460
rect 16764 25492 16816 25498
rect 16764 25434 16816 25440
rect 16672 25424 16724 25430
rect 16672 25366 16724 25372
rect 16580 25356 16632 25362
rect 16580 25298 16632 25304
rect 16672 25220 16724 25226
rect 16672 25162 16724 25168
rect 16580 23724 16632 23730
rect 16580 23666 16632 23672
rect 16486 22672 16542 22681
rect 16486 22607 16542 22616
rect 16592 22545 16620 23666
rect 16578 22536 16634 22545
rect 16578 22471 16634 22480
rect 16486 22400 16542 22409
rect 16486 22335 16542 22344
rect 16500 12238 16528 22335
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 16592 21350 16620 21966
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16684 20505 16712 25162
rect 16776 24410 16804 25434
rect 16764 24404 16816 24410
rect 16764 24346 16816 24352
rect 16776 23662 16804 24346
rect 16764 23656 16816 23662
rect 16764 23598 16816 23604
rect 16776 23322 16804 23598
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 16764 23112 16816 23118
rect 16764 23054 16816 23060
rect 16776 22817 16804 23054
rect 16762 22808 16818 22817
rect 16762 22743 16818 22752
rect 16776 22642 16804 22743
rect 16764 22636 16816 22642
rect 16764 22578 16816 22584
rect 16868 22522 16896 27882
rect 16960 24750 16988 31214
rect 17236 30938 17264 31826
rect 17224 30932 17276 30938
rect 17224 30874 17276 30880
rect 17236 30394 17264 30874
rect 17224 30388 17276 30394
rect 17224 30330 17276 30336
rect 17040 27532 17092 27538
rect 17040 27474 17092 27480
rect 17052 27169 17080 27474
rect 17038 27160 17094 27169
rect 17038 27095 17094 27104
rect 17328 27010 17356 32150
rect 17604 32042 17632 37266
rect 17774 35592 17830 35601
rect 17774 35527 17776 35536
rect 17828 35527 17830 35536
rect 17776 35498 17828 35504
rect 17774 34096 17830 34105
rect 17774 34031 17830 34040
rect 17684 32564 17736 32570
rect 17684 32506 17736 32512
rect 17052 26982 17356 27010
rect 17420 32014 17632 32042
rect 17052 24857 17080 26982
rect 17420 26908 17448 32014
rect 17500 31952 17552 31958
rect 17500 31894 17552 31900
rect 17512 28966 17540 31894
rect 17592 31408 17644 31414
rect 17592 31350 17644 31356
rect 17604 30870 17632 31350
rect 17592 30864 17644 30870
rect 17592 30806 17644 30812
rect 17604 30394 17632 30806
rect 17592 30388 17644 30394
rect 17592 30330 17644 30336
rect 17592 30048 17644 30054
rect 17592 29990 17644 29996
rect 17604 29850 17632 29990
rect 17592 29844 17644 29850
rect 17592 29786 17644 29792
rect 17500 28960 17552 28966
rect 17500 28902 17552 28908
rect 17512 28558 17540 28902
rect 17500 28552 17552 28558
rect 17500 28494 17552 28500
rect 17512 27878 17540 28494
rect 17500 27872 17552 27878
rect 17500 27814 17552 27820
rect 17512 27470 17540 27814
rect 17696 27538 17724 32506
rect 17684 27532 17736 27538
rect 17684 27474 17736 27480
rect 17500 27464 17552 27470
rect 17500 27406 17552 27412
rect 17144 26880 17448 26908
rect 17038 24848 17094 24857
rect 17038 24783 17094 24792
rect 16948 24744 17000 24750
rect 16948 24686 17000 24692
rect 16960 24342 16988 24686
rect 17040 24608 17092 24614
rect 17040 24550 17092 24556
rect 16948 24336 17000 24342
rect 16948 24278 17000 24284
rect 17052 24274 17080 24550
rect 17040 24268 17092 24274
rect 17040 24210 17092 24216
rect 17040 23316 17092 23322
rect 17040 23258 17092 23264
rect 16948 22772 17000 22778
rect 16948 22714 17000 22720
rect 16960 22574 16988 22714
rect 17052 22710 17080 23258
rect 17040 22704 17092 22710
rect 17040 22646 17092 22652
rect 16776 22494 16896 22522
rect 16948 22568 17000 22574
rect 16948 22510 17000 22516
rect 16776 21146 16804 22494
rect 17038 21992 17094 22001
rect 17038 21927 17094 21936
rect 16764 21140 16816 21146
rect 16764 21082 16816 21088
rect 16948 20936 17000 20942
rect 16946 20904 16948 20913
rect 17000 20904 17002 20913
rect 16946 20839 17002 20848
rect 16960 20602 16988 20839
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 16670 20496 16726 20505
rect 16670 20431 16726 20440
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 16960 19446 16988 19858
rect 16948 19440 17000 19446
rect 16948 19382 17000 19388
rect 16948 19304 17000 19310
rect 16946 19272 16948 19281
rect 17000 19272 17002 19281
rect 16946 19207 17002 19216
rect 16946 18864 17002 18873
rect 16946 18799 17002 18808
rect 16960 18630 16988 18799
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16948 18216 17000 18222
rect 16670 18184 16726 18193
rect 16948 18158 17000 18164
rect 16670 18119 16726 18128
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16592 17338 16620 17682
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16592 16794 16620 17274
rect 16684 17202 16712 18119
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16580 16788 16632 16794
rect 16580 16730 16632 16736
rect 16684 16658 16712 17138
rect 16856 17128 16908 17134
rect 16960 17105 16988 18158
rect 16856 17070 16908 17076
rect 16946 17096 17002 17105
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16684 16250 16712 16594
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16764 15564 16816 15570
rect 16764 15506 16816 15512
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16578 15192 16634 15201
rect 16578 15127 16634 15136
rect 16592 15026 16620 15127
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16592 14550 16620 14962
rect 16580 14544 16632 14550
rect 16580 14486 16632 14492
rect 16684 14396 16712 15438
rect 16776 15162 16804 15506
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 16592 14368 16712 14396
rect 16592 14074 16620 14368
rect 16580 14068 16632 14074
rect 16868 14056 16896 17070
rect 16946 17031 17002 17040
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 16960 14249 16988 16594
rect 16946 14240 17002 14249
rect 16946 14175 17002 14184
rect 16580 14010 16632 14016
rect 16776 14028 16896 14056
rect 16592 13977 16620 14010
rect 16672 14000 16724 14006
rect 16578 13968 16634 13977
rect 16672 13942 16724 13948
rect 16578 13903 16634 13912
rect 16684 13705 16712 13942
rect 16670 13696 16726 13705
rect 16670 13631 16726 13640
rect 16580 13456 16632 13462
rect 16580 13398 16632 13404
rect 16592 12986 16620 13398
rect 16684 13326 16712 13631
rect 16776 13462 16804 14028
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16764 13456 16816 13462
rect 16868 13433 16896 13874
rect 16764 13398 16816 13404
rect 16854 13424 16910 13433
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16578 12880 16634 12889
rect 16578 12815 16634 12824
rect 16592 12442 16620 12815
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16500 10985 16528 12038
rect 16486 10976 16542 10985
rect 16486 10911 16542 10920
rect 16592 10266 16620 12242
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16684 11529 16712 12174
rect 16776 11694 16804 13398
rect 16854 13359 16910 13368
rect 16946 13016 17002 13025
rect 16946 12951 17002 12960
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16764 11552 16816 11558
rect 16670 11520 16726 11529
rect 16764 11494 16816 11500
rect 16670 11455 16726 11464
rect 16776 11370 16804 11494
rect 16684 11342 16804 11370
rect 16684 10742 16712 11342
rect 16672 10736 16724 10742
rect 16670 10704 16672 10713
rect 16724 10704 16726 10713
rect 16670 10639 16726 10648
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16500 7970 16528 8774
rect 16868 8650 16896 12378
rect 16960 12306 16988 12951
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16776 8622 16896 8650
rect 16684 8430 16712 8461
rect 16672 8424 16724 8430
rect 16670 8392 16672 8401
rect 16724 8392 16726 8401
rect 16670 8327 16726 8336
rect 16684 8090 16712 8327
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16500 7954 16620 7970
rect 16500 7948 16632 7954
rect 16500 7942 16580 7948
rect 16580 7890 16632 7896
rect 16672 6792 16724 6798
rect 16776 6780 16804 8622
rect 16960 8566 16988 12106
rect 16948 8560 17000 8566
rect 16854 8528 16910 8537
rect 16948 8502 17000 8508
rect 16854 8463 16856 8472
rect 16908 8463 16910 8472
rect 16856 8434 16908 8440
rect 16854 6896 16910 6905
rect 16854 6831 16856 6840
rect 16908 6831 16910 6840
rect 16948 6860 17000 6866
rect 16856 6802 16908 6808
rect 16948 6802 17000 6808
rect 16724 6752 16804 6780
rect 16672 6734 16724 6740
rect 16684 6390 16712 6734
rect 16672 6384 16724 6390
rect 16672 6326 16724 6332
rect 16684 5681 16712 6326
rect 16868 6322 16896 6802
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16960 6118 16988 6802
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 16960 5914 16988 6054
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 16670 5672 16726 5681
rect 16670 5607 16726 5616
rect 17052 3670 17080 21927
rect 17144 20482 17172 26880
rect 17512 26858 17540 27406
rect 17684 27328 17736 27334
rect 17684 27270 17736 27276
rect 17500 26852 17552 26858
rect 17500 26794 17552 26800
rect 17696 26450 17724 27270
rect 17684 26444 17736 26450
rect 17684 26386 17736 26392
rect 17408 26376 17460 26382
rect 17408 26318 17460 26324
rect 17500 26376 17552 26382
rect 17500 26318 17552 26324
rect 17420 25974 17448 26318
rect 17512 26042 17540 26318
rect 17696 26042 17724 26386
rect 17500 26036 17552 26042
rect 17500 25978 17552 25984
rect 17684 26036 17736 26042
rect 17684 25978 17736 25984
rect 17408 25968 17460 25974
rect 17408 25910 17460 25916
rect 17420 25809 17448 25910
rect 17406 25800 17462 25809
rect 17406 25735 17462 25744
rect 17408 25356 17460 25362
rect 17408 25298 17460 25304
rect 17500 25356 17552 25362
rect 17500 25298 17552 25304
rect 17224 25288 17276 25294
rect 17224 25230 17276 25236
rect 17236 24954 17264 25230
rect 17420 24954 17448 25298
rect 17512 24993 17540 25298
rect 17788 25226 17816 34031
rect 17880 31278 17908 38694
rect 17972 34921 18000 40996
rect 18432 38457 18460 40996
rect 19156 40180 19208 40186
rect 19156 40122 19208 40128
rect 18418 38448 18474 38457
rect 18418 38383 18474 38392
rect 18236 38208 18288 38214
rect 18236 38150 18288 38156
rect 18970 38176 19026 38185
rect 18144 37664 18196 37670
rect 18144 37606 18196 37612
rect 18156 37262 18184 37606
rect 18144 37256 18196 37262
rect 18144 37198 18196 37204
rect 18156 36718 18184 37198
rect 18144 36712 18196 36718
rect 18144 36654 18196 36660
rect 18052 36168 18104 36174
rect 18050 36136 18052 36145
rect 18104 36136 18106 36145
rect 18050 36071 18106 36080
rect 18156 36038 18184 36654
rect 18144 36032 18196 36038
rect 18144 35974 18196 35980
rect 18052 35624 18104 35630
rect 18156 35578 18184 35974
rect 18104 35572 18184 35578
rect 18052 35566 18184 35572
rect 18064 35550 18184 35566
rect 18156 35494 18184 35550
rect 18144 35488 18196 35494
rect 18144 35430 18196 35436
rect 18156 34950 18184 35430
rect 18144 34944 18196 34950
rect 17958 34912 18014 34921
rect 18144 34886 18196 34892
rect 17958 34847 18014 34856
rect 17958 34096 18014 34105
rect 17958 34031 17960 34040
rect 18012 34031 18014 34040
rect 17960 34002 18012 34008
rect 17972 33658 18000 34002
rect 18156 33998 18184 34886
rect 18144 33992 18196 33998
rect 18144 33934 18196 33940
rect 17960 33652 18012 33658
rect 17960 33594 18012 33600
rect 17960 33380 18012 33386
rect 17960 33322 18012 33328
rect 17972 32570 18000 33322
rect 18156 33318 18184 33934
rect 18144 33312 18196 33318
rect 18144 33254 18196 33260
rect 18156 32910 18184 33254
rect 18144 32904 18196 32910
rect 18144 32846 18196 32852
rect 17960 32564 18012 32570
rect 17960 32506 18012 32512
rect 18156 32502 18184 32846
rect 18144 32496 18196 32502
rect 18144 32438 18196 32444
rect 17960 32292 18012 32298
rect 17960 32234 18012 32240
rect 17868 31272 17920 31278
rect 17868 31214 17920 31220
rect 17866 30968 17922 30977
rect 17866 30903 17922 30912
rect 17880 25362 17908 30903
rect 17868 25356 17920 25362
rect 17868 25298 17920 25304
rect 17776 25220 17828 25226
rect 17776 25162 17828 25168
rect 17498 24984 17554 24993
rect 17224 24948 17276 24954
rect 17224 24890 17276 24896
rect 17408 24948 17460 24954
rect 17498 24919 17554 24928
rect 17408 24890 17460 24896
rect 17512 24410 17540 24919
rect 17500 24404 17552 24410
rect 17500 24346 17552 24352
rect 17408 24336 17460 24342
rect 17972 24290 18000 32234
rect 18144 32224 18196 32230
rect 18144 32166 18196 32172
rect 18156 31958 18184 32166
rect 18144 31952 18196 31958
rect 18144 31894 18196 31900
rect 18144 31272 18196 31278
rect 18144 31214 18196 31220
rect 18052 31136 18104 31142
rect 18052 31078 18104 31084
rect 18064 30258 18092 31078
rect 18052 30252 18104 30258
rect 18052 30194 18104 30200
rect 18052 28552 18104 28558
rect 18052 28494 18104 28500
rect 18064 27946 18092 28494
rect 18052 27940 18104 27946
rect 18052 27882 18104 27888
rect 18052 26784 18104 26790
rect 18052 26726 18104 26732
rect 17408 24278 17460 24284
rect 17420 23866 17448 24278
rect 17684 24268 17736 24274
rect 17684 24210 17736 24216
rect 17788 24262 18000 24290
rect 17408 23860 17460 23866
rect 17408 23802 17460 23808
rect 17420 23746 17448 23802
rect 17420 23718 17540 23746
rect 17408 22976 17460 22982
rect 17408 22918 17460 22924
rect 17420 22778 17448 22918
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 17408 22092 17460 22098
rect 17408 22034 17460 22040
rect 17224 22024 17276 22030
rect 17224 21966 17276 21972
rect 17236 21010 17264 21966
rect 17316 21344 17368 21350
rect 17316 21286 17368 21292
rect 17224 21004 17276 21010
rect 17224 20946 17276 20952
rect 17236 20602 17264 20946
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 17144 20466 17264 20482
rect 17144 20460 17276 20466
rect 17144 20454 17224 20460
rect 17224 20402 17276 20408
rect 17132 20392 17184 20398
rect 17132 20334 17184 20340
rect 17144 19922 17172 20334
rect 17328 20097 17356 21286
rect 17420 20992 17448 22034
rect 17512 21128 17540 23718
rect 17696 23322 17724 24210
rect 17684 23316 17736 23322
rect 17684 23258 17736 23264
rect 17684 22704 17736 22710
rect 17684 22646 17736 22652
rect 17696 21962 17724 22646
rect 17684 21956 17736 21962
rect 17684 21898 17736 21904
rect 17696 21690 17724 21898
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 17788 21298 17816 24262
rect 17960 24200 18012 24206
rect 17960 24142 18012 24148
rect 17972 23254 18000 24142
rect 17960 23248 18012 23254
rect 17960 23190 18012 23196
rect 17960 21888 18012 21894
rect 17960 21830 18012 21836
rect 17972 21729 18000 21830
rect 17958 21720 18014 21729
rect 17958 21655 18014 21664
rect 17788 21270 17908 21298
rect 17512 21100 17724 21128
rect 17592 21004 17644 21010
rect 17420 20964 17592 20992
rect 17592 20946 17644 20952
rect 17604 20534 17632 20946
rect 17592 20528 17644 20534
rect 17592 20470 17644 20476
rect 17314 20088 17370 20097
rect 17314 20023 17370 20032
rect 17132 19916 17184 19922
rect 17132 19858 17184 19864
rect 17408 19916 17460 19922
rect 17592 19916 17644 19922
rect 17460 19876 17540 19904
rect 17408 19858 17460 19864
rect 17144 19281 17172 19858
rect 17316 19780 17368 19786
rect 17236 19740 17316 19768
rect 17236 19689 17264 19740
rect 17316 19722 17368 19728
rect 17408 19712 17460 19718
rect 17222 19680 17278 19689
rect 17408 19654 17460 19660
rect 17222 19615 17278 19624
rect 17420 19310 17448 19654
rect 17408 19304 17460 19310
rect 17130 19272 17186 19281
rect 17408 19246 17460 19252
rect 17316 19236 17368 19242
rect 17130 19207 17186 19216
rect 17236 19196 17316 19224
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 17144 18630 17172 19110
rect 17132 18624 17184 18630
rect 17236 18601 17264 19196
rect 17316 19178 17368 19184
rect 17408 19168 17460 19174
rect 17408 19110 17460 19116
rect 17132 18566 17184 18572
rect 17222 18592 17278 18601
rect 17222 18527 17278 18536
rect 17236 17134 17264 18527
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 17328 17513 17356 18362
rect 17420 18222 17448 19110
rect 17512 18698 17540 19876
rect 17592 19858 17644 19864
rect 17604 19514 17632 19858
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 17590 19272 17646 19281
rect 17590 19207 17646 19216
rect 17604 18970 17632 19207
rect 17696 18970 17724 21100
rect 17774 20768 17830 20777
rect 17774 20703 17830 20712
rect 17592 18964 17644 18970
rect 17592 18906 17644 18912
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 17500 18692 17552 18698
rect 17500 18634 17552 18640
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17408 17876 17460 17882
rect 17408 17818 17460 17824
rect 17314 17504 17370 17513
rect 17314 17439 17370 17448
rect 17224 17128 17276 17134
rect 17224 17070 17276 17076
rect 17328 17066 17356 17439
rect 17316 17060 17368 17066
rect 17316 17002 17368 17008
rect 17224 16992 17276 16998
rect 17224 16934 17276 16940
rect 17236 16726 17264 16934
rect 17224 16720 17276 16726
rect 17224 16662 17276 16668
rect 17316 16720 17368 16726
rect 17316 16662 17368 16668
rect 17328 16590 17356 16662
rect 17316 16584 17368 16590
rect 17222 16552 17278 16561
rect 17316 16526 17368 16532
rect 17222 16487 17278 16496
rect 17236 16182 17264 16487
rect 17328 16250 17356 16526
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17224 16176 17276 16182
rect 17224 16118 17276 16124
rect 17132 15700 17184 15706
rect 17132 15642 17184 15648
rect 17144 14822 17172 15642
rect 17236 15638 17264 16118
rect 17224 15632 17276 15638
rect 17224 15574 17276 15580
rect 17132 14816 17184 14822
rect 17132 14758 17184 14764
rect 17144 14278 17172 14758
rect 17132 14272 17184 14278
rect 17132 14214 17184 14220
rect 17144 13530 17172 14214
rect 17316 13796 17368 13802
rect 17316 13738 17368 13744
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 17328 13394 17356 13738
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 17328 12782 17356 13330
rect 17316 12776 17368 12782
rect 17316 12718 17368 12724
rect 17420 12442 17448 17818
rect 17512 17184 17540 18634
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 17604 17814 17632 18566
rect 17696 18290 17724 18906
rect 17684 18284 17736 18290
rect 17684 18226 17736 18232
rect 17788 18193 17816 20703
rect 17774 18184 17830 18193
rect 17774 18119 17830 18128
rect 17776 18080 17828 18086
rect 17776 18022 17828 18028
rect 17788 17882 17816 18022
rect 17776 17876 17828 17882
rect 17776 17818 17828 17824
rect 17592 17808 17644 17814
rect 17592 17750 17644 17756
rect 17604 17338 17632 17750
rect 17776 17740 17828 17746
rect 17776 17682 17828 17688
rect 17788 17338 17816 17682
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 17512 17156 17632 17184
rect 17500 17060 17552 17066
rect 17500 17002 17552 17008
rect 17512 16658 17540 17002
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17498 16552 17554 16561
rect 17498 16487 17554 16496
rect 17512 16289 17540 16487
rect 17498 16280 17554 16289
rect 17498 16215 17554 16224
rect 17500 15020 17552 15026
rect 17500 14962 17552 14968
rect 17512 14618 17540 14962
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17512 13530 17540 14418
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17512 13190 17540 13466
rect 17500 13184 17552 13190
rect 17500 13126 17552 13132
rect 17512 12617 17540 13126
rect 17498 12608 17554 12617
rect 17498 12543 17554 12552
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 17314 12336 17370 12345
rect 17314 12271 17370 12280
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17144 11558 17172 12174
rect 17224 12164 17276 12170
rect 17224 12106 17276 12112
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17236 11354 17264 12106
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 17132 9988 17184 9994
rect 17132 9930 17184 9936
rect 17144 8242 17172 9930
rect 17144 8214 17264 8242
rect 17236 6866 17264 8214
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17236 6458 17264 6802
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 17130 4992 17186 5001
rect 17130 4927 17186 4936
rect 17144 4185 17172 4927
rect 17328 4826 17356 12271
rect 17420 11898 17448 12378
rect 17604 12238 17632 17156
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 17788 16046 17816 16390
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17684 15904 17736 15910
rect 17684 15846 17736 15852
rect 17696 13870 17724 15846
rect 17788 15706 17816 15982
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17788 15162 17816 15642
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17774 14920 17830 14929
rect 17774 14855 17830 14864
rect 17788 14618 17816 14855
rect 17776 14612 17828 14618
rect 17776 14554 17828 14560
rect 17776 14340 17828 14346
rect 17776 14282 17828 14288
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17788 13734 17816 14282
rect 17776 13728 17828 13734
rect 17776 13670 17828 13676
rect 17788 13326 17816 13670
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17682 12880 17738 12889
rect 17788 12850 17816 13262
rect 17682 12815 17738 12824
rect 17776 12844 17828 12850
rect 17592 12232 17644 12238
rect 17512 12192 17592 12220
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17512 11286 17540 12192
rect 17592 12174 17644 12180
rect 17696 12050 17724 12815
rect 17776 12786 17828 12792
rect 17880 12458 17908 21270
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 17972 18358 18000 18770
rect 17960 18352 18012 18358
rect 17960 18294 18012 18300
rect 17958 18048 18014 18057
rect 17958 17983 18014 17992
rect 17972 17882 18000 17983
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 18064 17270 18092 26726
rect 18156 22658 18184 31214
rect 18248 30977 18276 38150
rect 18970 38111 19026 38120
rect 18878 37632 18934 37641
rect 18878 37567 18934 37576
rect 18326 37360 18382 37369
rect 18326 37295 18382 37304
rect 18602 37360 18658 37369
rect 18602 37295 18604 37304
rect 18234 30968 18290 30977
rect 18234 30903 18290 30912
rect 18340 30818 18368 37295
rect 18656 37295 18658 37304
rect 18604 37266 18656 37272
rect 18616 36922 18644 37266
rect 18604 36916 18656 36922
rect 18604 36858 18656 36864
rect 18786 36544 18842 36553
rect 18786 36479 18842 36488
rect 18604 32904 18656 32910
rect 18604 32846 18656 32852
rect 18420 32360 18472 32366
rect 18420 32302 18472 32308
rect 18432 31890 18460 32302
rect 18616 32298 18644 32846
rect 18604 32292 18656 32298
rect 18604 32234 18656 32240
rect 18512 32020 18564 32026
rect 18512 31962 18564 31968
rect 18420 31884 18472 31890
rect 18420 31826 18472 31832
rect 18432 31142 18460 31826
rect 18524 31210 18552 31962
rect 18512 31204 18564 31210
rect 18512 31146 18564 31152
rect 18420 31136 18472 31142
rect 18420 31078 18472 31084
rect 18696 31136 18748 31142
rect 18696 31078 18748 31084
rect 18248 30790 18368 30818
rect 18420 30796 18472 30802
rect 18248 26081 18276 30790
rect 18604 30796 18656 30802
rect 18420 30738 18472 30744
rect 18524 30756 18604 30784
rect 18326 30696 18382 30705
rect 18326 30631 18328 30640
rect 18380 30631 18382 30640
rect 18328 30602 18380 30608
rect 18432 30546 18460 30738
rect 18340 30518 18460 30546
rect 18340 30394 18368 30518
rect 18328 30388 18380 30394
rect 18328 30330 18380 30336
rect 18340 29850 18368 30330
rect 18420 30320 18472 30326
rect 18420 30262 18472 30268
rect 18328 29844 18380 29850
rect 18328 29786 18380 29792
rect 18328 26852 18380 26858
rect 18328 26794 18380 26800
rect 18340 26246 18368 26794
rect 18328 26240 18380 26246
rect 18328 26182 18380 26188
rect 18234 26072 18290 26081
rect 18234 26007 18290 26016
rect 18236 25832 18288 25838
rect 18340 25820 18368 26182
rect 18288 25792 18368 25820
rect 18236 25774 18288 25780
rect 18248 24206 18276 25774
rect 18236 24200 18288 24206
rect 18236 24142 18288 24148
rect 18432 23118 18460 30262
rect 18524 29850 18552 30756
rect 18604 30738 18656 30744
rect 18604 30252 18656 30258
rect 18604 30194 18656 30200
rect 18512 29844 18564 29850
rect 18512 29786 18564 29792
rect 18616 29170 18644 30194
rect 18604 29164 18656 29170
rect 18604 29106 18656 29112
rect 18708 27538 18736 31078
rect 18696 27532 18748 27538
rect 18696 27474 18748 27480
rect 18604 27396 18656 27402
rect 18604 27338 18656 27344
rect 18510 26344 18566 26353
rect 18510 26279 18566 26288
rect 18524 25906 18552 26279
rect 18512 25900 18564 25906
rect 18512 25842 18564 25848
rect 18524 25498 18552 25842
rect 18512 25492 18564 25498
rect 18512 25434 18564 25440
rect 18510 25256 18566 25265
rect 18510 25191 18566 25200
rect 18420 23112 18472 23118
rect 18420 23054 18472 23060
rect 18236 22976 18288 22982
rect 18236 22918 18288 22924
rect 18248 22778 18276 22918
rect 18236 22772 18288 22778
rect 18236 22714 18288 22720
rect 18156 22630 18276 22658
rect 18432 22642 18460 23054
rect 18144 21344 18196 21350
rect 18142 21312 18144 21321
rect 18196 21312 18198 21321
rect 18142 21247 18198 21256
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 18156 18873 18184 19110
rect 18142 18864 18198 18873
rect 18142 18799 18198 18808
rect 18142 17776 18198 17785
rect 18142 17711 18198 17720
rect 18052 17264 18104 17270
rect 18052 17206 18104 17212
rect 18156 16794 18184 17711
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18144 15904 18196 15910
rect 18064 15864 18144 15892
rect 18064 15570 18092 15864
rect 18144 15846 18196 15852
rect 18144 15632 18196 15638
rect 18144 15574 18196 15580
rect 18052 15564 18104 15570
rect 18052 15506 18104 15512
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17972 15162 18000 15370
rect 18064 15366 18092 15506
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 18064 14958 18092 15302
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 18064 14482 18092 14894
rect 18156 14550 18184 15574
rect 18144 14544 18196 14550
rect 18144 14486 18196 14492
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 17958 14104 18014 14113
rect 18064 14074 18092 14418
rect 18156 14346 18184 14486
rect 18144 14340 18196 14346
rect 18144 14282 18196 14288
rect 17958 14039 18014 14048
rect 18052 14068 18104 14074
rect 17972 13462 18000 14039
rect 18052 14010 18104 14016
rect 17960 13456 18012 13462
rect 17960 13398 18012 13404
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 17604 12022 17724 12050
rect 17788 12430 17908 12458
rect 17500 11280 17552 11286
rect 17500 11222 17552 11228
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17420 10470 17448 11086
rect 17604 10826 17632 12022
rect 17682 11928 17738 11937
rect 17682 11863 17738 11872
rect 17512 10798 17632 10826
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17420 10305 17448 10406
rect 17406 10296 17462 10305
rect 17406 10231 17462 10240
rect 17512 5953 17540 10798
rect 17590 10704 17646 10713
rect 17590 10639 17646 10648
rect 17498 5944 17554 5953
rect 17498 5879 17554 5888
rect 17316 4820 17368 4826
rect 17316 4762 17368 4768
rect 17222 4720 17278 4729
rect 17222 4655 17278 4664
rect 17236 4321 17264 4655
rect 17222 4312 17278 4321
rect 17222 4247 17278 4256
rect 17130 4176 17186 4185
rect 17130 4111 17186 4120
rect 17040 3664 17092 3670
rect 17040 3606 17092 3612
rect 16396 1828 16448 1834
rect 16396 1770 16448 1776
rect 17040 1216 17092 1222
rect 17040 1158 17092 1164
rect 17052 800 17080 1158
rect 17604 898 17632 10639
rect 17696 3194 17724 11863
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17788 1222 17816 12430
rect 17868 11892 17920 11898
rect 17972 11880 18000 12582
rect 18064 12442 18092 13330
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17920 11852 18000 11880
rect 17868 11834 17920 11840
rect 18064 11778 18092 12242
rect 17972 11750 18092 11778
rect 17866 10296 17922 10305
rect 17866 10231 17868 10240
rect 17920 10231 17922 10240
rect 17868 10202 17920 10208
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17880 7546 17908 7890
rect 17972 7585 18000 11750
rect 18050 11656 18106 11665
rect 18050 11591 18052 11600
rect 18104 11591 18106 11600
rect 18052 11562 18104 11568
rect 18144 9920 18196 9926
rect 18142 9888 18144 9897
rect 18196 9888 18198 9897
rect 18142 9823 18198 9832
rect 18248 9382 18276 22630
rect 18420 22636 18472 22642
rect 18420 22578 18472 22584
rect 18328 21004 18380 21010
rect 18328 20946 18380 20952
rect 18340 20262 18368 20946
rect 18328 20256 18380 20262
rect 18328 20198 18380 20204
rect 18340 19174 18368 20198
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18340 18426 18368 19110
rect 18432 19009 18460 19654
rect 18418 19000 18474 19009
rect 18418 18935 18474 18944
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18432 17882 18460 18702
rect 18420 17876 18472 17882
rect 18420 17818 18472 17824
rect 18420 17264 18472 17270
rect 18420 17206 18472 17212
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 18340 16454 18368 16934
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 18328 15904 18380 15910
rect 18328 15846 18380 15852
rect 18340 15094 18368 15846
rect 18328 15088 18380 15094
rect 18328 15030 18380 15036
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18340 14550 18368 14894
rect 18328 14544 18380 14550
rect 18328 14486 18380 14492
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18340 11694 18368 12038
rect 18328 11688 18380 11694
rect 18328 11630 18380 11636
rect 18340 11354 18368 11630
rect 18328 11348 18380 11354
rect 18328 11290 18380 11296
rect 18432 10606 18460 17206
rect 18524 16046 18552 25191
rect 18616 23662 18644 27338
rect 18708 26790 18736 27474
rect 18696 26784 18748 26790
rect 18696 26726 18748 26732
rect 18696 24064 18748 24070
rect 18696 24006 18748 24012
rect 18708 23662 18736 24006
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 18696 23656 18748 23662
rect 18696 23598 18748 23604
rect 18616 22778 18644 23598
rect 18694 23080 18750 23089
rect 18694 23015 18696 23024
rect 18748 23015 18750 23024
rect 18696 22986 18748 22992
rect 18604 22772 18656 22778
rect 18604 22714 18656 22720
rect 18616 22574 18644 22714
rect 18800 22658 18828 36479
rect 18892 31414 18920 37567
rect 18984 32570 19012 38111
rect 19064 33856 19116 33862
rect 19064 33798 19116 33804
rect 19076 33425 19104 33798
rect 19062 33416 19118 33425
rect 19062 33351 19118 33360
rect 19064 33312 19116 33318
rect 19064 33254 19116 33260
rect 18972 32564 19024 32570
rect 18972 32506 19024 32512
rect 18984 32366 19012 32506
rect 19076 32366 19104 33254
rect 18972 32360 19024 32366
rect 18972 32302 19024 32308
rect 19064 32360 19116 32366
rect 19064 32302 19116 32308
rect 19168 32178 19196 40122
rect 19352 37097 19380 40996
rect 19812 38842 19840 40996
rect 20076 40112 20128 40118
rect 20076 40054 20128 40060
rect 19984 39024 20036 39030
rect 19984 38966 20036 38972
rect 19812 38814 19932 38842
rect 19580 38652 19876 38672
rect 19636 38650 19660 38652
rect 19716 38650 19740 38652
rect 19796 38650 19820 38652
rect 19658 38598 19660 38650
rect 19722 38598 19734 38650
rect 19796 38598 19798 38650
rect 19636 38596 19660 38598
rect 19716 38596 19740 38598
rect 19796 38596 19820 38598
rect 19430 38584 19486 38593
rect 19580 38576 19876 38596
rect 19430 38519 19432 38528
rect 19484 38519 19486 38528
rect 19432 38490 19484 38496
rect 19432 38208 19484 38214
rect 19432 38150 19484 38156
rect 19444 37806 19472 38150
rect 19432 37800 19484 37806
rect 19432 37742 19484 37748
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 19432 37120 19484 37126
rect 19338 37088 19394 37097
rect 19432 37062 19484 37068
rect 19338 37023 19394 37032
rect 19444 36786 19472 37062
rect 19432 36780 19484 36786
rect 19432 36722 19484 36728
rect 19904 36689 19932 38814
rect 19996 37874 20024 38966
rect 19984 37868 20036 37874
rect 19984 37810 20036 37816
rect 20088 37754 20116 40054
rect 19996 37726 20116 37754
rect 20732 37754 20760 40996
rect 20732 37726 21036 37754
rect 19890 36680 19946 36689
rect 19890 36615 19946 36624
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 19892 35556 19944 35562
rect 19892 35498 19944 35504
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 19432 34536 19484 34542
rect 19432 34478 19484 34484
rect 19444 33998 19472 34478
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 19432 33992 19484 33998
rect 19432 33934 19484 33940
rect 19338 33280 19394 33289
rect 19338 33215 19394 33224
rect 19352 32586 19380 33215
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 18984 32150 19196 32178
rect 19260 32558 19380 32586
rect 18880 31408 18932 31414
rect 18880 31350 18932 31356
rect 18880 31272 18932 31278
rect 18880 31214 18932 31220
rect 18892 30938 18920 31214
rect 18880 30932 18932 30938
rect 18880 30874 18932 30880
rect 18878 27976 18934 27985
rect 18878 27911 18934 27920
rect 18892 27402 18920 27911
rect 18880 27396 18932 27402
rect 18880 27338 18932 27344
rect 18880 27056 18932 27062
rect 18880 26998 18932 27004
rect 18892 24721 18920 26998
rect 18878 24712 18934 24721
rect 18878 24647 18934 24656
rect 18880 23860 18932 23866
rect 18880 23802 18932 23808
rect 18892 23186 18920 23802
rect 18880 23180 18932 23186
rect 18880 23122 18932 23128
rect 18892 22778 18920 23122
rect 18880 22772 18932 22778
rect 18880 22714 18932 22720
rect 18800 22630 18920 22658
rect 18604 22568 18656 22574
rect 18604 22510 18656 22516
rect 18604 22092 18656 22098
rect 18604 22034 18656 22040
rect 18616 21350 18644 22034
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18604 21344 18656 21350
rect 18604 21286 18656 21292
rect 18604 21004 18656 21010
rect 18604 20946 18656 20952
rect 18616 20262 18644 20946
rect 18800 20806 18828 21966
rect 18788 20800 18840 20806
rect 18788 20742 18840 20748
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 18616 19417 18644 20198
rect 18602 19408 18658 19417
rect 18602 19343 18658 19352
rect 18788 19236 18840 19242
rect 18788 19178 18840 19184
rect 18602 19136 18658 19145
rect 18602 19071 18658 19080
rect 18616 18970 18644 19071
rect 18604 18964 18656 18970
rect 18604 18906 18656 18912
rect 18800 18630 18828 19178
rect 18788 18624 18840 18630
rect 18788 18566 18840 18572
rect 18602 18184 18658 18193
rect 18602 18119 18658 18128
rect 18512 16040 18564 16046
rect 18512 15982 18564 15988
rect 18616 15586 18644 18119
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18708 17134 18736 17614
rect 18800 17542 18828 18566
rect 18788 17536 18840 17542
rect 18788 17478 18840 17484
rect 18800 17338 18828 17478
rect 18788 17332 18840 17338
rect 18788 17274 18840 17280
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 18708 16658 18736 17070
rect 18786 16688 18842 16697
rect 18696 16652 18748 16658
rect 18786 16623 18842 16632
rect 18696 16594 18748 16600
rect 18708 15910 18736 16594
rect 18800 16114 18828 16623
rect 18788 16108 18840 16114
rect 18788 16050 18840 16056
rect 18788 15972 18840 15978
rect 18788 15914 18840 15920
rect 18696 15904 18748 15910
rect 18696 15846 18748 15852
rect 18524 15558 18644 15586
rect 18524 13954 18552 15558
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 18616 14822 18644 15438
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 18708 14074 18736 15846
rect 18800 15026 18828 15914
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18800 14618 18828 14962
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 18696 14068 18748 14074
rect 18696 14010 18748 14016
rect 18524 13926 18736 13954
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 18616 13462 18644 13738
rect 18604 13456 18656 13462
rect 18604 13398 18656 13404
rect 18604 12776 18656 12782
rect 18602 12744 18604 12753
rect 18656 12744 18658 12753
rect 18602 12679 18658 12688
rect 18510 12608 18566 12617
rect 18510 12543 18566 12552
rect 18524 12442 18552 12543
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18510 12336 18566 12345
rect 18510 12271 18566 12280
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18328 10532 18380 10538
rect 18328 10474 18380 10480
rect 18340 10130 18368 10474
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 18340 9722 18368 10066
rect 18328 9716 18380 9722
rect 18328 9658 18380 9664
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18248 8634 18276 9318
rect 18340 8634 18368 9658
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18340 8430 18368 8570
rect 18432 8566 18460 8978
rect 18420 8560 18472 8566
rect 18420 8502 18472 8508
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 18432 7886 18460 8502
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 17958 7576 18014 7585
rect 17868 7540 17920 7546
rect 17958 7511 18014 7520
rect 17868 7482 17920 7488
rect 17880 6934 17908 7482
rect 18432 7342 18460 7822
rect 18524 7449 18552 12271
rect 18616 11354 18644 12679
rect 18708 12442 18736 13926
rect 18788 13388 18840 13394
rect 18788 13330 18840 13336
rect 18800 12442 18828 13330
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18892 12322 18920 22630
rect 18984 20602 19012 32150
rect 19062 32056 19118 32065
rect 19062 31991 19118 32000
rect 19076 31142 19104 31991
rect 19260 31906 19288 32558
rect 19340 32428 19392 32434
rect 19340 32370 19392 32376
rect 19352 32026 19380 32370
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19340 32020 19392 32026
rect 19340 31962 19392 31968
rect 19432 32020 19484 32026
rect 19432 31962 19484 31968
rect 19260 31890 19380 31906
rect 19260 31884 19392 31890
rect 19260 31878 19340 31884
rect 19340 31826 19392 31832
rect 19248 31748 19300 31754
rect 19248 31690 19300 31696
rect 19156 31408 19208 31414
rect 19156 31350 19208 31356
rect 19064 31136 19116 31142
rect 19064 31078 19116 31084
rect 19168 31090 19196 31350
rect 19260 31278 19288 31690
rect 19248 31272 19300 31278
rect 19248 31214 19300 31220
rect 19076 30297 19104 31078
rect 19168 31062 19288 31090
rect 19062 30288 19118 30297
rect 19062 30223 19118 30232
rect 19156 30252 19208 30258
rect 19156 30194 19208 30200
rect 19168 29850 19196 30194
rect 19156 29844 19208 29850
rect 19156 29786 19208 29792
rect 19260 29730 19288 31062
rect 19352 30938 19380 31826
rect 19340 30932 19392 30938
rect 19340 30874 19392 30880
rect 19338 30832 19394 30841
rect 19338 30767 19394 30776
rect 19352 30705 19380 30767
rect 19338 30696 19394 30705
rect 19338 30631 19394 30640
rect 19340 30048 19392 30054
rect 19338 30016 19340 30025
rect 19392 30016 19394 30025
rect 19338 29951 19394 29960
rect 19168 29702 19288 29730
rect 19064 28144 19116 28150
rect 19064 28086 19116 28092
rect 19076 27985 19104 28086
rect 19062 27976 19118 27985
rect 19062 27911 19118 27920
rect 19168 24993 19196 29702
rect 19248 29096 19300 29102
rect 19300 29044 19380 29050
rect 19248 29038 19380 29044
rect 19260 29022 19380 29038
rect 19248 28960 19300 28966
rect 19248 28902 19300 28908
rect 19260 28014 19288 28902
rect 19352 28762 19380 29022
rect 19340 28756 19392 28762
rect 19340 28698 19392 28704
rect 19444 28150 19472 31962
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 19904 29714 19932 35498
rect 19892 29708 19944 29714
rect 19892 29650 19944 29656
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 19800 28416 19852 28422
rect 19904 28404 19932 29650
rect 19852 28376 19932 28404
rect 19800 28358 19852 28364
rect 19812 28257 19840 28358
rect 19798 28248 19854 28257
rect 19798 28183 19854 28192
rect 19432 28144 19484 28150
rect 19432 28086 19484 28092
rect 19248 28008 19300 28014
rect 19248 27950 19300 27956
rect 19892 28008 19944 28014
rect 19892 27950 19944 27956
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19352 26994 19380 27270
rect 19340 26988 19392 26994
rect 19340 26930 19392 26936
rect 19248 26852 19300 26858
rect 19248 26794 19300 26800
rect 19154 24984 19210 24993
rect 19154 24919 19210 24928
rect 19064 21480 19116 21486
rect 19062 21448 19064 21457
rect 19116 21448 19118 21457
rect 19062 21383 19118 21392
rect 19156 21344 19208 21350
rect 19156 21286 19208 21292
rect 19064 20800 19116 20806
rect 19064 20742 19116 20748
rect 18972 20596 19024 20602
rect 18972 20538 19024 20544
rect 19076 20482 19104 20742
rect 18984 20454 19104 20482
rect 18984 16674 19012 20454
rect 19168 20398 19196 21286
rect 19156 20392 19208 20398
rect 19156 20334 19208 20340
rect 19168 20058 19196 20334
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 19260 19961 19288 26794
rect 19352 26353 19380 26930
rect 19904 26926 19932 27950
rect 19432 26920 19484 26926
rect 19432 26862 19484 26868
rect 19892 26920 19944 26926
rect 19892 26862 19944 26868
rect 19444 26518 19472 26862
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19432 26512 19484 26518
rect 19432 26454 19484 26460
rect 19524 26444 19576 26450
rect 19524 26386 19576 26392
rect 19338 26344 19394 26353
rect 19338 26279 19394 26288
rect 19536 26042 19564 26386
rect 19904 26314 19932 26862
rect 19892 26308 19944 26314
rect 19892 26250 19944 26256
rect 19524 26036 19576 26042
rect 19524 25978 19576 25984
rect 19536 25786 19564 25978
rect 19444 25758 19564 25786
rect 19444 25498 19472 25758
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19432 25492 19484 25498
rect 19432 25434 19484 25440
rect 19892 24744 19944 24750
rect 19892 24686 19944 24692
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 19904 24070 19932 24686
rect 19892 24064 19944 24070
rect 19892 24006 19944 24012
rect 19890 23624 19946 23633
rect 19890 23559 19892 23568
rect 19944 23559 19946 23568
rect 19892 23530 19944 23536
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19616 23248 19668 23254
rect 19616 23190 19668 23196
rect 19628 22778 19656 23190
rect 19904 22778 19932 23530
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19892 22772 19944 22778
rect 19892 22714 19944 22720
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19432 22228 19484 22234
rect 19432 22170 19484 22176
rect 19340 21480 19392 21486
rect 19340 21422 19392 21428
rect 19246 19952 19302 19961
rect 19246 19887 19302 19896
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19260 17354 19288 18022
rect 19352 17490 19380 21422
rect 19444 21350 19472 22170
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19904 19378 19932 19654
rect 19892 19372 19944 19378
rect 19892 19314 19944 19320
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19904 18952 19932 19314
rect 19996 19310 20024 37726
rect 20720 37664 20772 37670
rect 20720 37606 20772 37612
rect 20534 35728 20590 35737
rect 20534 35663 20590 35672
rect 20074 35456 20130 35465
rect 20074 35391 20130 35400
rect 20088 34610 20116 35391
rect 20076 34604 20128 34610
rect 20076 34546 20128 34552
rect 20352 33856 20404 33862
rect 20352 33798 20404 33804
rect 20364 33454 20392 33798
rect 20442 33552 20498 33561
rect 20548 33522 20576 35663
rect 20442 33487 20444 33496
rect 20496 33487 20498 33496
rect 20536 33516 20588 33522
rect 20444 33458 20496 33464
rect 20536 33458 20588 33464
rect 20352 33448 20404 33454
rect 20352 33390 20404 33396
rect 20364 33046 20392 33390
rect 20352 33040 20404 33046
rect 20352 32982 20404 32988
rect 20076 32224 20128 32230
rect 20076 32166 20128 32172
rect 20088 31346 20116 32166
rect 20444 31816 20496 31822
rect 20444 31758 20496 31764
rect 20076 31340 20128 31346
rect 20076 31282 20128 31288
rect 20088 30938 20116 31282
rect 20260 31272 20312 31278
rect 20260 31214 20312 31220
rect 20076 30932 20128 30938
rect 20076 30874 20128 30880
rect 20272 30802 20300 31214
rect 20260 30796 20312 30802
rect 20260 30738 20312 30744
rect 20272 30274 20300 30738
rect 20180 30258 20300 30274
rect 20168 30252 20300 30258
rect 20220 30246 20300 30252
rect 20168 30194 20220 30200
rect 20352 29640 20404 29646
rect 20352 29582 20404 29588
rect 20364 29102 20392 29582
rect 20352 29096 20404 29102
rect 20352 29038 20404 29044
rect 20364 28762 20392 29038
rect 20352 28756 20404 28762
rect 20352 28698 20404 28704
rect 20364 27674 20392 28698
rect 20352 27668 20404 27674
rect 20352 27610 20404 27616
rect 20352 26376 20404 26382
rect 20352 26318 20404 26324
rect 20258 25800 20314 25809
rect 20258 25735 20314 25744
rect 20272 24614 20300 25735
rect 20364 25702 20392 26318
rect 20352 25696 20404 25702
rect 20352 25638 20404 25644
rect 20260 24608 20312 24614
rect 20260 24550 20312 24556
rect 20168 24064 20220 24070
rect 20168 24006 20220 24012
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 20088 22114 20116 23122
rect 20180 22642 20208 24006
rect 20272 23866 20300 24550
rect 20260 23860 20312 23866
rect 20260 23802 20312 23808
rect 20258 22808 20314 22817
rect 20258 22743 20314 22752
rect 20168 22636 20220 22642
rect 20168 22578 20220 22584
rect 20180 22234 20208 22578
rect 20168 22228 20220 22234
rect 20168 22170 20220 22176
rect 20088 22086 20208 22114
rect 20076 20800 20128 20806
rect 20076 20742 20128 20748
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 19720 18924 19932 18952
rect 19720 18630 19748 18924
rect 19708 18624 19760 18630
rect 19708 18566 19760 18572
rect 19720 18290 19748 18566
rect 19708 18284 19760 18290
rect 19708 18226 19760 18232
rect 19432 18080 19484 18086
rect 19430 18048 19432 18057
rect 19484 18048 19486 18057
rect 19430 17983 19486 17992
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19984 17536 20036 17542
rect 19352 17462 19472 17490
rect 19984 17478 20036 17484
rect 19260 17338 19380 17354
rect 19260 17332 19392 17338
rect 19260 17326 19340 17332
rect 19340 17274 19392 17280
rect 19444 17270 19472 17462
rect 19432 17264 19484 17270
rect 19432 17206 19484 17212
rect 19892 17264 19944 17270
rect 19892 17206 19944 17212
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19156 16720 19208 16726
rect 18984 16668 19156 16674
rect 18984 16662 19208 16668
rect 18984 16646 19196 16662
rect 19248 16652 19300 16658
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 18984 15638 19012 15982
rect 18972 15632 19024 15638
rect 18972 15574 19024 15580
rect 19076 15484 19104 16646
rect 19248 16594 19300 16600
rect 19156 16244 19208 16250
rect 19156 16186 19208 16192
rect 19168 15706 19196 16186
rect 19260 16046 19288 16594
rect 19352 16590 19380 17070
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19800 16720 19852 16726
rect 19798 16688 19800 16697
rect 19852 16688 19854 16697
rect 19798 16623 19854 16632
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 19156 15700 19208 15706
rect 19156 15642 19208 15648
rect 19432 15632 19484 15638
rect 19432 15574 19484 15580
rect 19340 15496 19392 15502
rect 18984 15456 19104 15484
rect 19260 15456 19340 15484
rect 18984 14113 19012 15456
rect 19156 15360 19208 15366
rect 19156 15302 19208 15308
rect 19168 14958 19196 15302
rect 19260 15162 19288 15456
rect 19340 15438 19392 15444
rect 19338 15328 19394 15337
rect 19338 15263 19394 15272
rect 19248 15156 19300 15162
rect 19248 15098 19300 15104
rect 19352 15042 19380 15263
rect 19260 15026 19380 15042
rect 19248 15020 19380 15026
rect 19300 15014 19380 15020
rect 19248 14962 19300 14968
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 19156 14816 19208 14822
rect 19156 14758 19208 14764
rect 19064 14612 19116 14618
rect 19064 14554 19116 14560
rect 18970 14104 19026 14113
rect 18970 14039 19026 14048
rect 19076 13954 19104 14554
rect 19168 14414 19196 14758
rect 19260 14618 19288 14826
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19352 14482 19380 14894
rect 19444 14618 19472 15574
rect 19904 15201 19932 17206
rect 19996 16046 20024 17478
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 19890 15192 19946 15201
rect 19890 15127 19946 15136
rect 19892 15088 19944 15094
rect 19892 15030 19944 15036
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19904 14550 19932 15030
rect 19524 14544 19576 14550
rect 19524 14486 19576 14492
rect 19892 14544 19944 14550
rect 19892 14486 19944 14492
rect 19340 14476 19392 14482
rect 19392 14436 19472 14464
rect 19340 14418 19392 14424
rect 19156 14408 19208 14414
rect 19156 14350 19208 14356
rect 18984 13926 19104 13954
rect 19168 14090 19196 14350
rect 19168 14074 19380 14090
rect 19168 14068 19392 14074
rect 19168 14062 19340 14068
rect 18984 13870 19012 13926
rect 18972 13864 19024 13870
rect 18972 13806 19024 13812
rect 18984 13394 19012 13806
rect 19064 13796 19116 13802
rect 19064 13738 19116 13744
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18984 12986 19012 13330
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 18800 12294 18920 12322
rect 18604 11348 18656 11354
rect 18604 11290 18656 11296
rect 18604 9920 18656 9926
rect 18604 9862 18656 9868
rect 18616 9586 18644 9862
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 18616 9081 18644 9522
rect 18602 9072 18658 9081
rect 18602 9007 18604 9016
rect 18656 9007 18658 9016
rect 18604 8978 18656 8984
rect 18616 8634 18644 8978
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18694 7848 18750 7857
rect 18694 7783 18750 7792
rect 18510 7440 18566 7449
rect 18510 7375 18566 7384
rect 18420 7336 18472 7342
rect 18420 7278 18472 7284
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 18512 6724 18564 6730
rect 18512 6666 18564 6672
rect 18524 6497 18552 6666
rect 18510 6488 18566 6497
rect 18510 6423 18566 6432
rect 18524 6390 18552 6423
rect 18512 6384 18564 6390
rect 18512 6326 18564 6332
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18156 4690 18184 5510
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 17868 4072 17920 4078
rect 17866 4040 17868 4049
rect 17920 4040 17922 4049
rect 17972 4026 18000 4558
rect 18156 4282 18184 4626
rect 18144 4276 18196 4282
rect 18144 4218 18196 4224
rect 17922 3998 18000 4026
rect 17866 3975 17922 3984
rect 18328 2644 18380 2650
rect 18328 2586 18380 2592
rect 18340 2446 18368 2586
rect 18328 2440 18380 2446
rect 18050 2408 18106 2417
rect 18328 2382 18380 2388
rect 18050 2343 18052 2352
rect 18104 2343 18106 2352
rect 18052 2314 18104 2320
rect 17868 1624 17920 1630
rect 17866 1592 17868 1601
rect 17920 1592 17922 1601
rect 17866 1527 17922 1536
rect 17776 1216 17828 1222
rect 17776 1158 17828 1164
rect 18708 921 18736 7783
rect 18800 7585 18828 12294
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18892 11898 18920 12174
rect 18880 11892 18932 11898
rect 18880 11834 18932 11840
rect 19076 10130 19104 13738
rect 19168 12850 19196 14062
rect 19340 14010 19392 14016
rect 19338 13968 19394 13977
rect 19248 13932 19300 13938
rect 19338 13903 19394 13912
rect 19248 13874 19300 13880
rect 19260 13530 19288 13874
rect 19352 13530 19380 13903
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19444 13258 19472 14436
rect 19536 14385 19564 14486
rect 19522 14376 19578 14385
rect 19522 14311 19578 14320
rect 19890 14376 19946 14385
rect 19890 14311 19946 14320
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 19904 13394 19932 14311
rect 19892 13388 19944 13394
rect 19892 13330 19944 13336
rect 19432 13252 19484 13258
rect 19432 13194 19484 13200
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 19168 12646 19196 12786
rect 19352 12753 19380 12786
rect 19432 12776 19484 12782
rect 19338 12744 19394 12753
rect 19432 12718 19484 12724
rect 19338 12679 19394 12688
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19168 11762 19196 12582
rect 19260 12396 19380 12424
rect 19156 11756 19208 11762
rect 19156 11698 19208 11704
rect 19156 11348 19208 11354
rect 19156 11290 19208 11296
rect 19168 11257 19196 11290
rect 19154 11248 19210 11257
rect 19260 11218 19288 12396
rect 19352 12345 19380 12396
rect 19338 12336 19394 12345
rect 19338 12271 19394 12280
rect 19444 11286 19472 12718
rect 19996 12714 20024 15982
rect 20088 13025 20116 20742
rect 20180 17649 20208 22086
rect 20272 21690 20300 22743
rect 20260 21684 20312 21690
rect 20260 21626 20312 21632
rect 20260 20868 20312 20874
rect 20260 20810 20312 20816
rect 20272 20641 20300 20810
rect 20258 20632 20314 20641
rect 20258 20567 20314 20576
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 20166 17640 20222 17649
rect 20166 17575 20222 17584
rect 20272 15994 20300 17818
rect 20180 15966 20300 15994
rect 20180 14958 20208 15966
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20168 14952 20220 14958
rect 20166 14920 20168 14929
rect 20220 14920 20222 14929
rect 20166 14855 20222 14864
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 20180 14074 20208 14418
rect 20272 14346 20300 15846
rect 20260 14340 20312 14346
rect 20260 14282 20312 14288
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20272 13938 20300 14282
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 20074 13016 20130 13025
rect 20074 12951 20130 12960
rect 19984 12708 20036 12714
rect 19984 12650 20036 12656
rect 20168 12708 20220 12714
rect 20168 12650 20220 12656
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 20180 12442 20208 12650
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 20364 12356 20392 25638
rect 20456 20806 20484 31758
rect 20534 27976 20590 27985
rect 20534 27911 20590 27920
rect 20444 20800 20496 20806
rect 20444 20742 20496 20748
rect 20444 18284 20496 18290
rect 20444 18226 20496 18232
rect 20272 12328 20392 12356
rect 19524 12300 19576 12306
rect 19524 12242 19576 12248
rect 19536 11898 19564 12242
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 19432 11280 19484 11286
rect 19432 11222 19484 11228
rect 19154 11183 19210 11192
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 19260 11098 19288 11154
rect 19260 11070 19380 11098
rect 19352 10810 19380 11070
rect 20272 10810 20300 12328
rect 20456 12288 20484 18226
rect 20364 12260 20484 12288
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 20260 10804 20312 10810
rect 20260 10746 20312 10752
rect 19154 10432 19210 10441
rect 19154 10367 19210 10376
rect 19168 10266 19196 10367
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 20272 10266 20300 10746
rect 20364 10266 20392 12260
rect 20548 12186 20576 27911
rect 20628 24812 20680 24818
rect 20732 24800 20760 37606
rect 20812 36644 20864 36650
rect 20812 36586 20864 36592
rect 20680 24772 20760 24800
rect 20628 24754 20680 24760
rect 20732 23186 20760 24772
rect 20720 23180 20772 23186
rect 20720 23122 20772 23128
rect 20628 21004 20680 21010
rect 20628 20946 20680 20952
rect 20640 20369 20668 20946
rect 20824 20482 20852 36586
rect 20904 34604 20956 34610
rect 20904 34546 20956 34552
rect 20916 21729 20944 34546
rect 21008 33697 21036 37726
rect 20994 33688 21050 33697
rect 20994 33623 21050 33632
rect 21192 33289 21220 40996
rect 21652 34184 21680 40996
rect 22572 37913 22600 40996
rect 22928 39364 22980 39370
rect 22928 39306 22980 39312
rect 22742 38448 22798 38457
rect 22742 38383 22798 38392
rect 22558 37904 22614 37913
rect 22558 37839 22614 37848
rect 22756 35329 22784 38383
rect 22836 36372 22888 36378
rect 22836 36314 22888 36320
rect 22742 35320 22798 35329
rect 22742 35255 22798 35264
rect 22374 34912 22430 34921
rect 22374 34847 22430 34856
rect 21652 34156 22048 34184
rect 21824 34060 21876 34066
rect 21824 34002 21876 34008
rect 21732 33992 21784 33998
rect 21732 33934 21784 33940
rect 21744 33658 21772 33934
rect 21732 33652 21784 33658
rect 21732 33594 21784 33600
rect 21364 33448 21416 33454
rect 21836 33425 21864 34002
rect 21914 33824 21970 33833
rect 21914 33759 21970 33768
rect 21364 33390 21416 33396
rect 21822 33416 21878 33425
rect 21178 33280 21234 33289
rect 21178 33215 21234 33224
rect 21376 33114 21404 33390
rect 21822 33351 21878 33360
rect 21836 33318 21864 33351
rect 21824 33312 21876 33318
rect 21824 33254 21876 33260
rect 21364 33108 21416 33114
rect 21364 33050 21416 33056
rect 21364 32904 21416 32910
rect 21364 32846 21416 32852
rect 21376 32230 21404 32846
rect 21364 32224 21416 32230
rect 21364 32166 21416 32172
rect 21086 31648 21142 31657
rect 21086 31583 21142 31592
rect 20996 31136 21048 31142
rect 20996 31078 21048 31084
rect 21008 30433 21036 31078
rect 20994 30424 21050 30433
rect 20994 30359 21050 30368
rect 21100 30258 21128 31583
rect 21376 30802 21404 32166
rect 21546 31784 21602 31793
rect 21546 31719 21602 31728
rect 21364 30796 21416 30802
rect 21364 30738 21416 30744
rect 21272 30728 21324 30734
rect 21272 30670 21324 30676
rect 21284 30569 21312 30670
rect 21270 30560 21326 30569
rect 21270 30495 21326 30504
rect 21284 30394 21312 30495
rect 21272 30388 21324 30394
rect 21272 30330 21324 30336
rect 21088 30252 21140 30258
rect 21088 30194 21140 30200
rect 21376 29850 21404 30738
rect 21364 29844 21416 29850
rect 21364 29786 21416 29792
rect 21272 29504 21324 29510
rect 21272 29446 21324 29452
rect 21178 29336 21234 29345
rect 21178 29271 21234 29280
rect 21192 29238 21220 29271
rect 21180 29232 21232 29238
rect 21180 29174 21232 29180
rect 21284 29102 21312 29446
rect 21456 29164 21508 29170
rect 21456 29106 21508 29112
rect 21272 29096 21324 29102
rect 21272 29038 21324 29044
rect 21088 28008 21140 28014
rect 21088 27950 21140 27956
rect 21100 27130 21128 27950
rect 21284 27946 21312 29038
rect 21272 27940 21324 27946
rect 21272 27882 21324 27888
rect 21364 27940 21416 27946
rect 21364 27882 21416 27888
rect 21088 27124 21140 27130
rect 21088 27066 21140 27072
rect 21088 26852 21140 26858
rect 21088 26794 21140 26800
rect 21100 26450 21128 26794
rect 21088 26444 21140 26450
rect 21088 26386 21140 26392
rect 21100 26042 21128 26386
rect 21180 26308 21232 26314
rect 21180 26250 21232 26256
rect 21088 26036 21140 26042
rect 21088 25978 21140 25984
rect 21088 25356 21140 25362
rect 21088 25298 21140 25304
rect 21100 24206 21128 25298
rect 21088 24200 21140 24206
rect 21088 24142 21140 24148
rect 21100 23662 21128 24142
rect 21088 23656 21140 23662
rect 21008 23604 21088 23610
rect 21008 23598 21140 23604
rect 21008 23582 21128 23598
rect 21008 22982 21036 23582
rect 20996 22976 21048 22982
rect 20996 22918 21048 22924
rect 20902 21720 20958 21729
rect 20902 21655 20958 21664
rect 20824 20454 20944 20482
rect 20626 20360 20682 20369
rect 20626 20295 20682 20304
rect 20812 20324 20864 20330
rect 20640 20244 20668 20295
rect 20812 20266 20864 20272
rect 20720 20256 20772 20262
rect 20640 20216 20720 20244
rect 20640 18222 20668 20216
rect 20720 20198 20772 20204
rect 20628 18216 20680 18222
rect 20628 18158 20680 18164
rect 20720 17060 20772 17066
rect 20720 17002 20772 17008
rect 20732 16794 20760 17002
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20824 15881 20852 20266
rect 20916 17882 20944 20454
rect 20904 17876 20956 17882
rect 20904 17818 20956 17824
rect 21008 16658 21036 22918
rect 21192 22794 21220 26250
rect 21100 22766 21220 22794
rect 20996 16652 21048 16658
rect 20996 16594 21048 16600
rect 20810 15872 20866 15881
rect 20810 15807 20866 15816
rect 20824 15722 20852 15807
rect 20640 15706 20852 15722
rect 20628 15700 20852 15706
rect 20680 15694 20852 15700
rect 20628 15642 20680 15648
rect 21008 15638 21036 16594
rect 20996 15632 21048 15638
rect 20996 15574 21048 15580
rect 20718 15192 20774 15201
rect 20718 15127 20774 15136
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20456 12158 20576 12186
rect 20640 12730 20668 13806
rect 20732 13530 20760 15127
rect 20996 14476 21048 14482
rect 20996 14418 21048 14424
rect 21008 14074 21036 14418
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 21008 13530 21036 14010
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 21008 12986 21036 13466
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 21008 12782 21036 12922
rect 20996 12776 21048 12782
rect 20718 12744 20774 12753
rect 20640 12702 20718 12730
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 19892 10192 19944 10198
rect 19892 10134 19944 10140
rect 19064 10124 19116 10130
rect 19064 10066 19116 10072
rect 19076 9722 19104 10066
rect 19524 9920 19576 9926
rect 19524 9862 19576 9868
rect 19064 9716 19116 9722
rect 19064 9658 19116 9664
rect 19536 9518 19564 9862
rect 19904 9654 19932 10134
rect 19892 9648 19944 9654
rect 19892 9590 19944 9596
rect 19524 9512 19576 9518
rect 19246 9480 19302 9489
rect 19064 9444 19116 9450
rect 19524 9454 19576 9460
rect 19246 9415 19302 9424
rect 19064 9386 19116 9392
rect 18970 9072 19026 9081
rect 18970 9007 19026 9016
rect 18786 7576 18842 7585
rect 18786 7511 18842 7520
rect 18880 6928 18932 6934
rect 18880 6870 18932 6876
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 18800 5817 18828 6598
rect 18892 5914 18920 6870
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 18786 5808 18842 5817
rect 18786 5743 18842 5752
rect 18984 2802 19012 9007
rect 19076 6798 19104 9386
rect 19260 9382 19288 9415
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 19708 8016 19760 8022
rect 19708 7958 19760 7964
rect 19340 7744 19392 7750
rect 19720 7721 19748 7958
rect 19340 7686 19392 7692
rect 19706 7712 19762 7721
rect 19352 6882 19380 7686
rect 19706 7647 19762 7656
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19444 6905 19472 7482
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19260 6866 19380 6882
rect 19248 6860 19380 6866
rect 19300 6854 19380 6860
rect 19430 6896 19486 6905
rect 19430 6831 19486 6840
rect 19248 6802 19300 6808
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 19076 6361 19104 6734
rect 19260 6458 19288 6802
rect 19904 6798 19932 9590
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19996 9110 20024 9318
rect 19984 9104 20036 9110
rect 19984 9046 20036 9052
rect 20364 8090 20392 10202
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 20364 7970 20392 8026
rect 20272 7942 20392 7970
rect 20272 7342 20300 7942
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 20364 7449 20392 7822
rect 20350 7440 20406 7449
rect 20350 7375 20352 7384
rect 20404 7375 20406 7384
rect 20352 7346 20404 7352
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 20364 7002 20392 7346
rect 20352 6996 20404 7002
rect 20352 6938 20404 6944
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 20364 6458 20392 6938
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 19062 6352 19118 6361
rect 19062 6287 19118 6296
rect 19076 5846 19104 6287
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19340 6248 19392 6254
rect 19340 6190 19392 6196
rect 19064 5840 19116 5846
rect 19064 5782 19116 5788
rect 19168 5574 19196 6190
rect 19156 5568 19208 5574
rect 19156 5510 19208 5516
rect 19156 4072 19208 4078
rect 19156 4014 19208 4020
rect 19168 3738 19196 4014
rect 19156 3732 19208 3738
rect 19156 3674 19208 3680
rect 18800 2774 19012 2802
rect 18800 2666 18828 2774
rect 18800 2638 18920 2666
rect 17512 870 17632 898
rect 17958 912 18014 921
rect 17512 800 17540 870
rect 17958 847 18014 856
rect 18694 912 18750 921
rect 18694 847 18750 856
rect 17972 800 18000 847
rect 18892 800 18920 2638
rect 19352 800 19380 6190
rect 19982 6080 20038 6089
rect 19580 6012 19876 6032
rect 19982 6015 20038 6024
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 19430 5672 19486 5681
rect 19430 5607 19486 5616
rect 19444 4758 19472 5607
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 19432 4752 19484 4758
rect 19432 4694 19484 4700
rect 19996 4593 20024 6015
rect 20456 5953 20484 12158
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20548 11286 20576 12038
rect 20640 11694 20668 12702
rect 20996 12718 21048 12724
rect 20718 12679 20774 12688
rect 20812 12708 20864 12714
rect 20812 12650 20864 12656
rect 20824 12288 20852 12650
rect 20904 12300 20956 12306
rect 20824 12260 20904 12288
rect 20904 12242 20956 12248
rect 20916 11898 20944 12242
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 20628 11688 20680 11694
rect 20628 11630 20680 11636
rect 20640 11354 20668 11630
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20536 11280 20588 11286
rect 20536 11222 20588 11228
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 20810 9616 20866 9625
rect 20810 9551 20866 9560
rect 20824 8945 20852 9551
rect 20810 8936 20866 8945
rect 20810 8871 20866 8880
rect 20916 6361 20944 9658
rect 21100 8022 21128 22766
rect 21284 22098 21312 27882
rect 21376 27674 21404 27882
rect 21364 27668 21416 27674
rect 21364 27610 21416 27616
rect 21468 26450 21496 29106
rect 21456 26444 21508 26450
rect 21456 26386 21508 26392
rect 21468 26042 21496 26386
rect 21456 26036 21508 26042
rect 21456 25978 21508 25984
rect 21560 25498 21588 31719
rect 21836 29170 21864 33254
rect 21928 32910 21956 33759
rect 21916 32904 21968 32910
rect 21916 32846 21968 32852
rect 21928 32570 21956 32846
rect 21916 32564 21968 32570
rect 21916 32506 21968 32512
rect 22020 32450 22048 34156
rect 22388 33930 22416 34847
rect 22468 34060 22520 34066
rect 22468 34002 22520 34008
rect 22376 33924 22428 33930
rect 22376 33866 22428 33872
rect 22480 33590 22508 34002
rect 22848 33844 22876 36314
rect 22940 36258 22968 39306
rect 23032 36378 23060 40996
rect 23492 38593 23520 40996
rect 23478 38584 23534 38593
rect 23478 38519 23534 38528
rect 24412 38457 24440 40996
rect 24584 38548 24636 38554
rect 24584 38490 24636 38496
rect 24596 38457 24624 38490
rect 23202 38448 23258 38457
rect 23202 38383 23204 38392
rect 23256 38383 23258 38392
rect 24398 38448 24454 38457
rect 24398 38383 24454 38392
rect 24582 38448 24638 38457
rect 24582 38383 24638 38392
rect 23204 38354 23256 38360
rect 23216 38010 23244 38354
rect 23388 38344 23440 38350
rect 23388 38286 23440 38292
rect 23204 38004 23256 38010
rect 23204 37946 23256 37952
rect 23400 37670 23428 38286
rect 24308 38208 24360 38214
rect 24308 38150 24360 38156
rect 23388 37664 23440 37670
rect 23388 37606 23440 37612
rect 23570 37496 23626 37505
rect 23570 37431 23626 37440
rect 23020 36372 23072 36378
rect 23020 36314 23072 36320
rect 22940 36230 23244 36258
rect 22848 33816 22968 33844
rect 22468 33584 22520 33590
rect 22466 33552 22468 33561
rect 22520 33552 22522 33561
rect 22466 33487 22522 33496
rect 22376 33448 22428 33454
rect 22376 33390 22428 33396
rect 22098 33144 22154 33153
rect 22098 33079 22154 33088
rect 21928 32422 22048 32450
rect 21824 29164 21876 29170
rect 21824 29106 21876 29112
rect 21638 28112 21694 28121
rect 21638 28047 21694 28056
rect 21548 25492 21600 25498
rect 21548 25434 21600 25440
rect 21362 25392 21418 25401
rect 21652 25378 21680 28047
rect 21732 27668 21784 27674
rect 21732 27610 21784 27616
rect 21744 26994 21772 27610
rect 21732 26988 21784 26994
rect 21732 26930 21784 26936
rect 21928 25922 21956 32422
rect 22112 28744 22140 33079
rect 22284 30184 22336 30190
rect 22282 30152 22284 30161
rect 22336 30152 22338 30161
rect 22192 30116 22244 30122
rect 22282 30087 22338 30096
rect 22192 30058 22244 30064
rect 22204 29850 22232 30058
rect 22284 30048 22336 30054
rect 22388 30025 22416 33390
rect 22284 29990 22336 29996
rect 22374 30016 22430 30025
rect 22192 29844 22244 29850
rect 22192 29786 22244 29792
rect 22296 29646 22324 29990
rect 22374 29951 22430 29960
rect 22284 29640 22336 29646
rect 22284 29582 22336 29588
rect 22020 28716 22140 28744
rect 22020 28150 22048 28716
rect 22190 28656 22246 28665
rect 22190 28591 22192 28600
rect 22244 28591 22246 28600
rect 22192 28562 22244 28568
rect 22100 28552 22152 28558
rect 22100 28494 22152 28500
rect 22008 28144 22060 28150
rect 22008 28086 22060 28092
rect 22020 27674 22048 28086
rect 22112 27878 22140 28494
rect 22100 27872 22152 27878
rect 22100 27814 22152 27820
rect 22008 27668 22060 27674
rect 22008 27610 22060 27616
rect 22112 27146 22140 27814
rect 22192 27464 22244 27470
rect 22192 27406 22244 27412
rect 22020 27118 22140 27146
rect 22020 27062 22048 27118
rect 22008 27056 22060 27062
rect 22008 26998 22060 27004
rect 22020 26450 22048 26998
rect 22204 26926 22232 27406
rect 22192 26920 22244 26926
rect 22192 26862 22244 26868
rect 22008 26444 22060 26450
rect 22008 26386 22060 26392
rect 22020 26042 22048 26386
rect 22008 26036 22060 26042
rect 22008 25978 22060 25984
rect 21928 25894 22048 25922
rect 21362 25327 21418 25336
rect 21468 25350 21680 25378
rect 21916 25356 21968 25362
rect 21376 25294 21404 25327
rect 21364 25288 21416 25294
rect 21364 25230 21416 25236
rect 21376 24410 21404 25230
rect 21364 24404 21416 24410
rect 21364 24346 21416 24352
rect 21376 23322 21404 24346
rect 21364 23316 21416 23322
rect 21364 23258 21416 23264
rect 21272 22092 21324 22098
rect 21272 22034 21324 22040
rect 21284 21690 21312 22034
rect 21364 22024 21416 22030
rect 21364 21966 21416 21972
rect 21272 21684 21324 21690
rect 21272 21626 21324 21632
rect 21272 21412 21324 21418
rect 21272 21354 21324 21360
rect 21178 20632 21234 20641
rect 21178 20567 21234 20576
rect 21192 16590 21220 20567
rect 21284 19553 21312 21354
rect 21376 20777 21404 21966
rect 21362 20768 21418 20777
rect 21362 20703 21418 20712
rect 21270 19544 21326 19553
rect 21270 19479 21326 19488
rect 21364 19236 21416 19242
rect 21364 19178 21416 19184
rect 21376 18970 21404 19178
rect 21364 18964 21416 18970
rect 21364 18906 21416 18912
rect 21468 17218 21496 25350
rect 21916 25298 21968 25304
rect 21732 25288 21784 25294
rect 21732 25230 21784 25236
rect 21744 24614 21772 25230
rect 21928 24818 21956 25298
rect 21916 24812 21968 24818
rect 21916 24754 21968 24760
rect 21732 24608 21784 24614
rect 21732 24550 21784 24556
rect 21548 24132 21600 24138
rect 21548 24074 21600 24080
rect 21560 23662 21588 24074
rect 21732 23724 21784 23730
rect 21732 23666 21784 23672
rect 21548 23656 21600 23662
rect 21548 23598 21600 23604
rect 21560 22778 21588 23598
rect 21548 22772 21600 22778
rect 21548 22714 21600 22720
rect 21546 21720 21602 21729
rect 21546 21655 21602 21664
rect 21284 17190 21496 17218
rect 21180 16584 21232 16590
rect 21180 16526 21232 16532
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 21192 9897 21220 16186
rect 21178 9888 21234 9897
rect 21178 9823 21234 9832
rect 21088 8016 21140 8022
rect 21088 7958 21140 7964
rect 21192 7954 21220 9823
rect 21180 7948 21232 7954
rect 21180 7890 21232 7896
rect 21192 7834 21220 7890
rect 21100 7806 21220 7834
rect 21100 7002 21128 7806
rect 21180 7744 21232 7750
rect 21180 7686 21232 7692
rect 21088 6996 21140 7002
rect 21088 6938 21140 6944
rect 20902 6352 20958 6361
rect 20902 6287 20958 6296
rect 20442 5944 20498 5953
rect 20442 5879 20498 5888
rect 19982 4584 20038 4593
rect 19982 4519 20038 4528
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 19996 3398 20024 3674
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19996 2990 20024 3334
rect 19984 2984 20036 2990
rect 20168 2984 20220 2990
rect 19984 2926 20036 2932
rect 20166 2952 20168 2961
rect 20220 2952 20222 2961
rect 19432 2848 19484 2854
rect 19430 2816 19432 2825
rect 19484 2816 19486 2825
rect 19430 2751 19486 2760
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 19996 2650 20024 2926
rect 20166 2887 20222 2896
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 19996 2446 20024 2586
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 19800 2304 19852 2310
rect 19800 2246 19852 2252
rect 19812 800 19840 2246
rect 20548 898 20576 4082
rect 20548 870 20760 898
rect 20732 800 20760 870
rect 21192 800 21220 7686
rect 21284 4146 21312 17190
rect 21364 17128 21416 17134
rect 21560 17082 21588 21655
rect 21640 21480 21692 21486
rect 21640 21422 21692 21428
rect 21652 20942 21680 21422
rect 21640 20936 21692 20942
rect 21638 20904 21640 20913
rect 21692 20904 21694 20913
rect 21638 20839 21694 20848
rect 21744 19938 21772 23666
rect 21364 17070 21416 17076
rect 21376 16998 21404 17070
rect 21468 17054 21588 17082
rect 21652 19910 21772 19938
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21364 16584 21416 16590
rect 21364 16526 21416 16532
rect 21376 16114 21404 16526
rect 21364 16108 21416 16114
rect 21364 16050 21416 16056
rect 21364 14000 21416 14006
rect 21364 13942 21416 13948
rect 21376 5137 21404 13942
rect 21468 13394 21496 17054
rect 21652 16590 21680 19910
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 21744 19514 21772 19790
rect 22020 19786 22048 25894
rect 22284 22092 22336 22098
rect 22284 22034 22336 22040
rect 22296 20806 22324 22034
rect 22388 22030 22416 29951
rect 22558 29744 22614 29753
rect 22558 29679 22560 29688
rect 22612 29679 22614 29688
rect 22744 29708 22796 29714
rect 22560 29650 22612 29656
rect 22744 29650 22796 29656
rect 22756 29306 22784 29650
rect 22836 29640 22888 29646
rect 22836 29582 22888 29588
rect 22744 29300 22796 29306
rect 22744 29242 22796 29248
rect 22848 29186 22876 29582
rect 22940 29510 22968 33816
rect 23018 30832 23074 30841
rect 23018 30767 23020 30776
rect 23072 30767 23074 30776
rect 23020 30738 23072 30744
rect 23216 30598 23244 36230
rect 23294 34912 23350 34921
rect 23294 34847 23350 34856
rect 23308 32910 23336 34847
rect 23296 32904 23348 32910
rect 23296 32846 23348 32852
rect 23296 32768 23348 32774
rect 23296 32710 23348 32716
rect 23204 30592 23256 30598
rect 23204 30534 23256 30540
rect 23216 29714 23244 30534
rect 23308 29850 23336 32710
rect 23480 30048 23532 30054
rect 23480 29990 23532 29996
rect 23296 29844 23348 29850
rect 23296 29786 23348 29792
rect 23492 29753 23520 29990
rect 23478 29744 23534 29753
rect 23204 29708 23256 29714
rect 23478 29679 23534 29688
rect 23204 29650 23256 29656
rect 23480 29640 23532 29646
rect 23480 29582 23532 29588
rect 22928 29504 22980 29510
rect 22928 29446 22980 29452
rect 23296 29504 23348 29510
rect 23296 29446 23348 29452
rect 22756 29158 22876 29186
rect 22756 28966 22784 29158
rect 23112 29028 23164 29034
rect 23112 28970 23164 28976
rect 22744 28960 22796 28966
rect 22744 28902 22796 28908
rect 22756 28558 22784 28902
rect 22926 28656 22982 28665
rect 22926 28591 22928 28600
rect 22980 28591 22982 28600
rect 22928 28562 22980 28568
rect 22744 28552 22796 28558
rect 22744 28494 22796 28500
rect 22940 27674 22968 28562
rect 23020 28552 23072 28558
rect 23020 28494 23072 28500
rect 23032 28082 23060 28494
rect 23020 28076 23072 28082
rect 23020 28018 23072 28024
rect 22928 27668 22980 27674
rect 22928 27610 22980 27616
rect 22836 27532 22888 27538
rect 22836 27474 22888 27480
rect 22848 27130 22876 27474
rect 22836 27124 22888 27130
rect 22836 27066 22888 27072
rect 22468 26920 22520 26926
rect 22468 26862 22520 26868
rect 22480 26042 22508 26862
rect 22834 26480 22890 26489
rect 22834 26415 22890 26424
rect 22848 26246 22876 26415
rect 22836 26240 22888 26246
rect 22836 26182 22888 26188
rect 22468 26036 22520 26042
rect 22468 25978 22520 25984
rect 22848 25838 22876 26182
rect 22836 25832 22888 25838
rect 22836 25774 22888 25780
rect 22560 23180 22612 23186
rect 22560 23122 22612 23128
rect 22572 22778 22600 23122
rect 22560 22772 22612 22778
rect 22560 22714 22612 22720
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 22388 21622 22416 21966
rect 22376 21616 22428 21622
rect 22376 21558 22428 21564
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 22652 21344 22704 21350
rect 22652 21286 22704 21292
rect 22388 21146 22416 21286
rect 22376 21140 22428 21146
rect 22376 21082 22428 21088
rect 22664 21010 22692 21286
rect 22652 21004 22704 21010
rect 22652 20946 22704 20952
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22284 20800 22336 20806
rect 22284 20742 22336 20748
rect 22100 20256 22152 20262
rect 22100 20198 22152 20204
rect 22112 19922 22140 20198
rect 22100 19916 22152 19922
rect 22100 19858 22152 19864
rect 22008 19780 22060 19786
rect 22008 19722 22060 19728
rect 21732 19508 21784 19514
rect 21732 19450 21784 19456
rect 21744 17649 21772 19450
rect 22112 19174 22140 19858
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21730 17640 21786 17649
rect 21730 17575 21786 17584
rect 21640 16584 21692 16590
rect 21640 16526 21692 16532
rect 21548 16448 21600 16454
rect 21548 16390 21600 16396
rect 21560 15722 21588 16390
rect 21652 16250 21680 16526
rect 21640 16244 21692 16250
rect 21640 16186 21692 16192
rect 21560 15694 21680 15722
rect 21548 15632 21600 15638
rect 21548 15574 21600 15580
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 21468 12170 21496 13330
rect 21456 12164 21508 12170
rect 21456 12106 21508 12112
rect 21560 7954 21588 15574
rect 21652 9722 21680 15694
rect 21744 15638 21772 17575
rect 21836 16046 21864 18226
rect 21916 18148 21968 18154
rect 21916 18090 21968 18096
rect 21928 16658 21956 18090
rect 22112 18086 22140 19110
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 22020 17882 22048 18022
rect 22008 17876 22060 17882
rect 22008 17818 22060 17824
rect 22020 17270 22048 17818
rect 22008 17264 22060 17270
rect 22008 17206 22060 17212
rect 22192 17264 22244 17270
rect 22192 17206 22244 17212
rect 21916 16652 21968 16658
rect 21916 16594 21968 16600
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 22112 16114 22140 16594
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 21824 16040 21876 16046
rect 21824 15982 21876 15988
rect 21836 15706 21864 15982
rect 21824 15700 21876 15706
rect 21824 15642 21876 15648
rect 21732 15632 21784 15638
rect 21732 15574 21784 15580
rect 21744 14618 21772 15574
rect 21824 15564 21876 15570
rect 21824 15506 21876 15512
rect 21836 15201 21864 15506
rect 21822 15192 21878 15201
rect 21822 15127 21824 15136
rect 21876 15127 21878 15136
rect 21824 15098 21876 15104
rect 21836 15067 21864 15098
rect 21824 14816 21876 14822
rect 21824 14758 21876 14764
rect 21732 14612 21784 14618
rect 21732 14554 21784 14560
rect 21744 13870 21772 14554
rect 21732 13864 21784 13870
rect 21732 13806 21784 13812
rect 21836 13734 21864 14758
rect 21916 14476 21968 14482
rect 21916 14418 21968 14424
rect 21824 13728 21876 13734
rect 21824 13670 21876 13676
rect 21836 12782 21864 13670
rect 21928 13190 21956 14418
rect 22112 13530 22140 16050
rect 22100 13524 22152 13530
rect 22100 13466 22152 13472
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 22112 12782 22140 13466
rect 21824 12776 21876 12782
rect 21824 12718 21876 12724
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 21836 11694 21864 12718
rect 22112 12442 22140 12718
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22100 12300 22152 12306
rect 22100 12242 22152 12248
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 22020 11694 22048 12174
rect 22112 11694 22140 12242
rect 21824 11688 21876 11694
rect 21824 11630 21876 11636
rect 22008 11688 22060 11694
rect 22008 11630 22060 11636
rect 22100 11688 22152 11694
rect 22100 11630 22152 11636
rect 21836 11393 21864 11630
rect 21822 11384 21878 11393
rect 22020 11354 22048 11630
rect 22112 11354 22140 11630
rect 21822 11319 21878 11328
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 21916 10124 21968 10130
rect 21916 10066 21968 10072
rect 21928 9722 21956 10066
rect 21640 9716 21692 9722
rect 21640 9658 21692 9664
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 21928 9450 21956 9658
rect 21916 9444 21968 9450
rect 21916 9386 21968 9392
rect 21548 7948 21600 7954
rect 21548 7890 21600 7896
rect 21916 7948 21968 7954
rect 21916 7890 21968 7896
rect 21560 7546 21588 7890
rect 21928 7546 21956 7890
rect 22204 7857 22232 17206
rect 22296 15858 22324 20742
rect 22388 20602 22416 20878
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22560 20324 22612 20330
rect 22560 20266 22612 20272
rect 22572 19922 22600 20266
rect 22664 20262 22692 20946
rect 22744 20596 22796 20602
rect 22744 20538 22796 20544
rect 22652 20256 22704 20262
rect 22652 20198 22704 20204
rect 22560 19916 22612 19922
rect 22560 19858 22612 19864
rect 22572 19174 22600 19858
rect 22560 19168 22612 19174
rect 22560 19110 22612 19116
rect 22572 17814 22600 19110
rect 22560 17808 22612 17814
rect 22560 17750 22612 17756
rect 22466 16552 22522 16561
rect 22466 16487 22522 16496
rect 22376 16176 22428 16182
rect 22376 16118 22428 16124
rect 22388 16017 22416 16118
rect 22374 16008 22430 16017
rect 22374 15943 22430 15952
rect 22296 15830 22416 15858
rect 22284 15700 22336 15706
rect 22284 15642 22336 15648
rect 22296 14958 22324 15642
rect 22284 14952 22336 14958
rect 22284 14894 22336 14900
rect 22296 14278 22324 14894
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22388 12764 22416 15830
rect 22480 15094 22508 16487
rect 22756 15706 22784 20538
rect 22744 15700 22796 15706
rect 22744 15642 22796 15648
rect 22560 15428 22612 15434
rect 22560 15370 22612 15376
rect 22744 15428 22796 15434
rect 22744 15370 22796 15376
rect 22572 15337 22600 15370
rect 22558 15328 22614 15337
rect 22558 15263 22614 15272
rect 22468 15088 22520 15094
rect 22468 15030 22520 15036
rect 22572 14958 22600 15263
rect 22560 14952 22612 14958
rect 22560 14894 22612 14900
rect 22572 13870 22600 14894
rect 22756 14618 22784 15370
rect 22744 14612 22796 14618
rect 22744 14554 22796 14560
rect 22560 13864 22612 13870
rect 22560 13806 22612 13812
rect 22572 13394 22600 13806
rect 22560 13388 22612 13394
rect 22560 13330 22612 13336
rect 22558 13016 22614 13025
rect 22558 12951 22614 12960
rect 22468 12912 22520 12918
rect 22466 12880 22468 12889
rect 22520 12880 22522 12889
rect 22466 12815 22522 12824
rect 22572 12782 22600 12951
rect 22560 12776 22612 12782
rect 22388 12736 22508 12764
rect 22376 12300 22428 12306
rect 22376 12242 22428 12248
rect 22388 11830 22416 12242
rect 22376 11824 22428 11830
rect 22376 11766 22428 11772
rect 22376 10124 22428 10130
rect 22296 10084 22376 10112
rect 22296 9382 22324 10084
rect 22376 10066 22428 10072
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 22190 7848 22246 7857
rect 22190 7783 22246 7792
rect 21548 7540 21600 7546
rect 21548 7482 21600 7488
rect 21916 7540 21968 7546
rect 21916 7482 21968 7488
rect 21928 7002 21956 7482
rect 22296 7313 22324 9318
rect 22480 7721 22508 12736
rect 22560 12718 22612 12724
rect 22572 12374 22600 12718
rect 22560 12368 22612 12374
rect 22560 12310 22612 12316
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 22466 7712 22522 7721
rect 22466 7647 22522 7656
rect 22282 7304 22338 7313
rect 22282 7239 22338 7248
rect 21916 6996 21968 7002
rect 21916 6938 21968 6944
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 22468 6792 22520 6798
rect 22468 6734 22520 6740
rect 22204 6458 22232 6734
rect 22192 6452 22244 6458
rect 22192 6394 22244 6400
rect 22480 6186 22508 6734
rect 22572 6633 22600 11698
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22664 9382 22692 9998
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22558 6624 22614 6633
rect 22558 6559 22614 6568
rect 22664 6458 22692 9318
rect 22652 6452 22704 6458
rect 22652 6394 22704 6400
rect 22468 6180 22520 6186
rect 22468 6122 22520 6128
rect 21362 5128 21418 5137
rect 21362 5063 21418 5072
rect 21640 5024 21692 5030
rect 21640 4966 21692 4972
rect 21272 4140 21324 4146
rect 21272 4082 21324 4088
rect 21270 3360 21326 3369
rect 21270 3295 21326 3304
rect 21284 3194 21312 3295
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 21652 2446 21680 4966
rect 22558 2952 22614 2961
rect 22558 2887 22614 2896
rect 21824 2508 21876 2514
rect 21824 2450 21876 2456
rect 21640 2440 21692 2446
rect 21640 2382 21692 2388
rect 21836 2258 21864 2450
rect 22020 2366 22140 2394
rect 22020 2258 22048 2366
rect 21836 2230 22048 2258
rect 22112 800 22140 2366
rect 22572 800 22600 2887
rect 22848 2650 22876 25774
rect 22928 24200 22980 24206
rect 22928 24142 22980 24148
rect 22940 23594 22968 24142
rect 22928 23588 22980 23594
rect 22928 23530 22980 23536
rect 23020 21004 23072 21010
rect 23020 20946 23072 20952
rect 23032 20330 23060 20946
rect 23124 20874 23152 28970
rect 23202 28248 23258 28257
rect 23202 28183 23204 28192
rect 23256 28183 23258 28192
rect 23204 28154 23256 28160
rect 23204 25492 23256 25498
rect 23204 25434 23256 25440
rect 23216 24274 23244 25434
rect 23204 24268 23256 24274
rect 23204 24210 23256 24216
rect 23216 23866 23244 24210
rect 23204 23860 23256 23866
rect 23204 23802 23256 23808
rect 23216 23118 23244 23802
rect 23308 23236 23336 29446
rect 23492 29306 23520 29582
rect 23480 29300 23532 29306
rect 23480 29242 23532 29248
rect 23480 27940 23532 27946
rect 23480 27882 23532 27888
rect 23492 27674 23520 27882
rect 23480 27668 23532 27674
rect 23480 27610 23532 27616
rect 23388 23588 23440 23594
rect 23388 23530 23440 23536
rect 23400 23474 23428 23530
rect 23400 23446 23520 23474
rect 23492 23322 23520 23446
rect 23480 23316 23532 23322
rect 23480 23258 23532 23264
rect 23308 23208 23428 23236
rect 23204 23112 23256 23118
rect 23204 23054 23256 23060
rect 23216 22778 23244 23054
rect 23204 22772 23256 22778
rect 23204 22714 23256 22720
rect 23296 22024 23348 22030
rect 23296 21966 23348 21972
rect 23308 21350 23336 21966
rect 23296 21344 23348 21350
rect 23296 21286 23348 21292
rect 23112 20868 23164 20874
rect 23112 20810 23164 20816
rect 23308 20641 23336 21286
rect 23294 20632 23350 20641
rect 23294 20567 23350 20576
rect 23020 20324 23072 20330
rect 23020 20266 23072 20272
rect 23296 19508 23348 19514
rect 23296 19450 23348 19456
rect 23112 19168 23164 19174
rect 23112 19110 23164 19116
rect 23124 18902 23152 19110
rect 23112 18896 23164 18902
rect 23112 18838 23164 18844
rect 23204 18760 23256 18766
rect 23204 18702 23256 18708
rect 23216 18426 23244 18702
rect 23204 18420 23256 18426
rect 23204 18362 23256 18368
rect 23110 17776 23166 17785
rect 23110 17711 23112 17720
rect 23164 17711 23166 17720
rect 23204 17740 23256 17746
rect 23112 17682 23164 17688
rect 23204 17682 23256 17688
rect 22928 17672 22980 17678
rect 22928 17614 22980 17620
rect 22940 17338 22968 17614
rect 22928 17332 22980 17338
rect 22928 17274 22980 17280
rect 22928 17060 22980 17066
rect 22928 17002 22980 17008
rect 22940 16726 22968 17002
rect 22928 16720 22980 16726
rect 22928 16662 22980 16668
rect 22940 16046 22968 16662
rect 23124 16590 23152 17682
rect 23216 16998 23244 17682
rect 23204 16992 23256 16998
rect 23204 16934 23256 16940
rect 23112 16584 23164 16590
rect 23112 16526 23164 16532
rect 22928 16040 22980 16046
rect 22928 15982 22980 15988
rect 23124 15638 23152 16526
rect 23112 15632 23164 15638
rect 23112 15574 23164 15580
rect 23112 14408 23164 14414
rect 23112 14350 23164 14356
rect 23124 14074 23152 14350
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 22928 13252 22980 13258
rect 22928 13194 22980 13200
rect 22940 12442 22968 13194
rect 23216 12442 23244 16934
rect 23308 15706 23336 19450
rect 23296 15700 23348 15706
rect 23296 15642 23348 15648
rect 23296 15496 23348 15502
rect 23296 15438 23348 15444
rect 23308 15162 23336 15438
rect 23296 15156 23348 15162
rect 23296 15098 23348 15104
rect 23296 12640 23348 12646
rect 23296 12582 23348 12588
rect 22928 12436 22980 12442
rect 22928 12378 22980 12384
rect 23204 12436 23256 12442
rect 23204 12378 23256 12384
rect 23308 12102 23336 12582
rect 23296 12096 23348 12102
rect 23296 12038 23348 12044
rect 23110 10976 23166 10985
rect 23110 10911 23166 10920
rect 23124 7954 23152 10911
rect 23296 9376 23348 9382
rect 23296 9318 23348 9324
rect 23308 9217 23336 9318
rect 23294 9208 23350 9217
rect 23294 9143 23350 9152
rect 23112 7948 23164 7954
rect 23112 7890 23164 7896
rect 23124 7546 23152 7890
rect 23112 7540 23164 7546
rect 23112 7482 23164 7488
rect 23020 6180 23072 6186
rect 23020 6122 23072 6128
rect 22836 2644 22888 2650
rect 22836 2586 22888 2592
rect 23032 800 23060 6122
rect 23202 4448 23258 4457
rect 23202 4383 23258 4392
rect 23216 3602 23244 4383
rect 23204 3596 23256 3602
rect 23204 3538 23256 3544
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 23124 3194 23152 3470
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 23124 2446 23152 3130
rect 23216 3126 23244 3538
rect 23204 3120 23256 3126
rect 23204 3062 23256 3068
rect 23400 2689 23428 23208
rect 23584 21622 23612 37431
rect 24320 37369 24348 38150
rect 24872 37505 24900 40996
rect 25228 38004 25280 38010
rect 25228 37946 25280 37952
rect 24858 37496 24914 37505
rect 24858 37431 24914 37440
rect 24306 37360 24362 37369
rect 24306 37295 24362 37304
rect 25134 36816 25190 36825
rect 25134 36751 25136 36760
rect 25188 36751 25190 36760
rect 25136 36722 25188 36728
rect 25136 36644 25188 36650
rect 25136 36586 25188 36592
rect 24030 36544 24086 36553
rect 24030 36479 24086 36488
rect 23846 35048 23902 35057
rect 23846 34983 23902 34992
rect 23664 34060 23716 34066
rect 23664 34002 23716 34008
rect 23676 33386 23704 34002
rect 23756 33992 23808 33998
rect 23756 33934 23808 33940
rect 23664 33380 23716 33386
rect 23664 33322 23716 33328
rect 23676 33153 23704 33322
rect 23768 33318 23796 33934
rect 23756 33312 23808 33318
rect 23756 33254 23808 33260
rect 23662 33144 23718 33153
rect 23662 33079 23718 33088
rect 23768 32434 23796 33254
rect 23756 32428 23808 32434
rect 23756 32370 23808 32376
rect 23664 31680 23716 31686
rect 23662 31648 23664 31657
rect 23716 31648 23718 31657
rect 23662 31583 23718 31592
rect 23676 31414 23704 31583
rect 23664 31408 23716 31414
rect 23664 31350 23716 31356
rect 23754 31376 23810 31385
rect 23860 31346 23888 34983
rect 23938 33280 23994 33289
rect 23938 33215 23994 33224
rect 23754 31311 23810 31320
rect 23848 31340 23900 31346
rect 23768 31278 23796 31311
rect 23848 31282 23900 31288
rect 23756 31272 23808 31278
rect 23756 31214 23808 31220
rect 23664 31136 23716 31142
rect 23664 31078 23716 31084
rect 23676 29714 23704 31078
rect 23768 30938 23796 31214
rect 23756 30932 23808 30938
rect 23756 30874 23808 30880
rect 23664 29708 23716 29714
rect 23664 29650 23716 29656
rect 23756 27872 23808 27878
rect 23756 27814 23808 27820
rect 23768 27538 23796 27814
rect 23952 27606 23980 33215
rect 24044 29034 24072 36479
rect 25148 36038 25176 36586
rect 25136 36032 25188 36038
rect 25136 35974 25188 35980
rect 24950 35864 25006 35873
rect 24950 35799 24952 35808
rect 25004 35799 25006 35808
rect 24952 35770 25004 35776
rect 25148 35630 25176 35974
rect 25136 35624 25188 35630
rect 25136 35566 25188 35572
rect 25148 34950 25176 35566
rect 24584 34944 24636 34950
rect 25136 34944 25188 34950
rect 24584 34886 24636 34892
rect 25134 34912 25136 34921
rect 25188 34912 25190 34921
rect 24596 34649 24624 34886
rect 25134 34847 25190 34856
rect 25148 34746 25176 34847
rect 25136 34740 25188 34746
rect 25136 34682 25188 34688
rect 24582 34640 24638 34649
rect 24582 34575 24638 34584
rect 24596 34542 24624 34575
rect 24584 34536 24636 34542
rect 24584 34478 24636 34484
rect 24400 34400 24452 34406
rect 24400 34342 24452 34348
rect 24412 34066 24440 34342
rect 24400 34060 24452 34066
rect 24400 34002 24452 34008
rect 24412 33658 24440 34002
rect 24400 33652 24452 33658
rect 24400 33594 24452 33600
rect 24584 33108 24636 33114
rect 24584 33050 24636 33056
rect 24398 32736 24454 32745
rect 24398 32671 24454 32680
rect 24412 31958 24440 32671
rect 24400 31952 24452 31958
rect 24400 31894 24452 31900
rect 24596 31822 24624 33050
rect 24952 32972 25004 32978
rect 24952 32914 25004 32920
rect 24964 32230 24992 32914
rect 25240 32502 25268 37946
rect 25412 33856 25464 33862
rect 25412 33798 25464 33804
rect 25424 33454 25452 33798
rect 25502 33688 25558 33697
rect 25502 33623 25558 33632
rect 25516 33522 25544 33623
rect 25504 33516 25556 33522
rect 25504 33458 25556 33464
rect 25412 33448 25464 33454
rect 25412 33390 25464 33396
rect 25424 33114 25452 33390
rect 25412 33108 25464 33114
rect 25412 33050 25464 33056
rect 25320 32972 25372 32978
rect 25320 32914 25372 32920
rect 25332 32570 25360 32914
rect 25320 32564 25372 32570
rect 25320 32506 25372 32512
rect 25228 32496 25280 32502
rect 25280 32444 25360 32450
rect 25228 32438 25360 32444
rect 25240 32422 25360 32438
rect 25240 32373 25268 32422
rect 24952 32224 25004 32230
rect 24952 32166 25004 32172
rect 24964 31929 24992 32166
rect 24674 31920 24730 31929
rect 24674 31855 24676 31864
rect 24728 31855 24730 31864
rect 24950 31920 25006 31929
rect 24950 31855 25006 31864
rect 24676 31826 24728 31832
rect 24584 31816 24636 31822
rect 24584 31758 24636 31764
rect 24596 30938 24624 31758
rect 25044 31136 25096 31142
rect 25044 31078 25096 31084
rect 24584 30932 24636 30938
rect 24584 30874 24636 30880
rect 25056 30802 25084 31078
rect 25044 30796 25096 30802
rect 25044 30738 25096 30744
rect 24860 30728 24912 30734
rect 24860 30670 24912 30676
rect 24872 30258 24900 30670
rect 24860 30252 24912 30258
rect 24860 30194 24912 30200
rect 24216 30184 24268 30190
rect 24216 30126 24268 30132
rect 24124 30048 24176 30054
rect 24124 29990 24176 29996
rect 24136 29170 24164 29990
rect 24228 29850 24256 30126
rect 24216 29844 24268 29850
rect 24216 29786 24268 29792
rect 24584 29640 24636 29646
rect 24584 29582 24636 29588
rect 24768 29640 24820 29646
rect 24768 29582 24820 29588
rect 24124 29164 24176 29170
rect 24124 29106 24176 29112
rect 24032 29028 24084 29034
rect 24032 28970 24084 28976
rect 24216 28552 24268 28558
rect 24216 28494 24268 28500
rect 24228 28014 24256 28494
rect 24216 28008 24268 28014
rect 24216 27950 24268 27956
rect 23940 27600 23992 27606
rect 23940 27542 23992 27548
rect 24030 27568 24086 27577
rect 23756 27532 23808 27538
rect 24030 27503 24086 27512
rect 23756 27474 23808 27480
rect 23768 26994 23796 27474
rect 23756 26988 23808 26994
rect 23808 26948 23888 26976
rect 23756 26930 23808 26936
rect 23756 26784 23808 26790
rect 23756 26726 23808 26732
rect 23662 26616 23718 26625
rect 23662 26551 23718 26560
rect 23676 25838 23704 26551
rect 23664 25832 23716 25838
rect 23664 25774 23716 25780
rect 23676 25498 23704 25774
rect 23664 25492 23716 25498
rect 23664 25434 23716 25440
rect 23662 24984 23718 24993
rect 23662 24919 23718 24928
rect 23676 21962 23704 24919
rect 23664 21956 23716 21962
rect 23664 21898 23716 21904
rect 23572 21616 23624 21622
rect 23572 21558 23624 21564
rect 23570 19952 23626 19961
rect 23570 19887 23626 19896
rect 23480 18964 23532 18970
rect 23480 18906 23532 18912
rect 23492 17134 23520 18906
rect 23480 17128 23532 17134
rect 23480 17070 23532 17076
rect 23480 15904 23532 15910
rect 23480 15846 23532 15852
rect 23492 15638 23520 15846
rect 23480 15632 23532 15638
rect 23480 15574 23532 15580
rect 23492 14958 23520 15574
rect 23480 14952 23532 14958
rect 23480 14894 23532 14900
rect 23492 14550 23520 14894
rect 23480 14544 23532 14550
rect 23480 14486 23532 14492
rect 23584 12714 23612 19887
rect 23664 18080 23716 18086
rect 23664 18022 23716 18028
rect 23676 17746 23704 18022
rect 23664 17740 23716 17746
rect 23664 17682 23716 17688
rect 23768 17252 23796 26726
rect 23860 26586 23888 26948
rect 23848 26580 23900 26586
rect 23848 26522 23900 26528
rect 23940 25832 23992 25838
rect 23940 25774 23992 25780
rect 23952 25401 23980 25774
rect 23938 25392 23994 25401
rect 23938 25327 23994 25336
rect 24044 24410 24072 27503
rect 24490 27432 24546 27441
rect 24490 27367 24546 27376
rect 24504 26926 24532 27367
rect 24492 26920 24544 26926
rect 24492 26862 24544 26868
rect 24306 24712 24362 24721
rect 24306 24647 24362 24656
rect 24032 24404 24084 24410
rect 24032 24346 24084 24352
rect 24032 21956 24084 21962
rect 24032 21898 24084 21904
rect 23846 21584 23902 21593
rect 23846 21519 23848 21528
rect 23900 21519 23902 21528
rect 23848 21490 23900 21496
rect 24044 21486 24072 21898
rect 24032 21480 24084 21486
rect 24032 21422 24084 21428
rect 24044 20942 24072 21422
rect 24032 20936 24084 20942
rect 24032 20878 24084 20884
rect 24032 19916 24084 19922
rect 24032 19858 24084 19864
rect 23940 19848 23992 19854
rect 23940 19790 23992 19796
rect 23952 19553 23980 19790
rect 23938 19544 23994 19553
rect 23938 19479 23940 19488
rect 23992 19479 23994 19488
rect 23940 19450 23992 19456
rect 24044 19446 24072 19858
rect 24320 19786 24348 24647
rect 24400 24608 24452 24614
rect 24400 24550 24452 24556
rect 24412 23361 24440 24550
rect 24398 23352 24454 23361
rect 24398 23287 24454 23296
rect 24412 20058 24440 23287
rect 24492 22092 24544 22098
rect 24492 22034 24544 22040
rect 24504 21486 24532 22034
rect 24492 21480 24544 21486
rect 24492 21422 24544 21428
rect 24504 21146 24532 21422
rect 24492 21140 24544 21146
rect 24492 21082 24544 21088
rect 24492 20256 24544 20262
rect 24490 20224 24492 20233
rect 24544 20224 24546 20233
rect 24490 20159 24546 20168
rect 24400 20052 24452 20058
rect 24400 19994 24452 20000
rect 24400 19916 24452 19922
rect 24400 19858 24452 19864
rect 24308 19780 24360 19786
rect 24308 19722 24360 19728
rect 24032 19440 24084 19446
rect 24032 19382 24084 19388
rect 24044 18850 24072 19382
rect 24308 19304 24360 19310
rect 24306 19272 24308 19281
rect 24360 19272 24362 19281
rect 24306 19207 24362 19216
rect 24320 18986 24348 19207
rect 23952 18834 24072 18850
rect 23940 18828 24072 18834
rect 23992 18822 24072 18828
rect 23940 18770 23992 18776
rect 23940 18692 23992 18698
rect 23940 18634 23992 18640
rect 23952 18193 23980 18634
rect 24044 18426 24072 18822
rect 24228 18970 24348 18986
rect 24228 18964 24360 18970
rect 24228 18958 24308 18964
rect 24032 18420 24084 18426
rect 24032 18362 24084 18368
rect 24228 18358 24256 18958
rect 24308 18906 24360 18912
rect 24306 18864 24362 18873
rect 24412 18834 24440 19858
rect 24306 18799 24362 18808
rect 24400 18828 24452 18834
rect 24320 18766 24348 18799
rect 24400 18770 24452 18776
rect 24308 18760 24360 18766
rect 24308 18702 24360 18708
rect 24320 18426 24348 18702
rect 24308 18420 24360 18426
rect 24308 18362 24360 18368
rect 24216 18352 24268 18358
rect 24216 18294 24268 18300
rect 23938 18184 23994 18193
rect 23938 18119 23994 18128
rect 24412 17814 24440 18770
rect 24504 18086 24532 20159
rect 24492 18080 24544 18086
rect 24492 18022 24544 18028
rect 24400 17808 24452 17814
rect 24400 17750 24452 17756
rect 23940 17740 23992 17746
rect 23940 17682 23992 17688
rect 23676 17224 23796 17252
rect 23572 12708 23624 12714
rect 23572 12650 23624 12656
rect 23480 12300 23532 12306
rect 23480 12242 23532 12248
rect 23492 11898 23520 12242
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23570 10160 23626 10169
rect 23570 10095 23626 10104
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 23492 7750 23520 9318
rect 23480 7744 23532 7750
rect 23480 7686 23532 7692
rect 23492 5778 23520 7686
rect 23584 6798 23612 10095
rect 23676 7993 23704 17224
rect 23952 16590 23980 17682
rect 24214 17640 24270 17649
rect 24214 17575 24216 17584
rect 24268 17575 24270 17584
rect 24216 17546 24268 17552
rect 24032 17128 24084 17134
rect 24032 17070 24084 17076
rect 23940 16584 23992 16590
rect 23940 16526 23992 16532
rect 23754 16416 23810 16425
rect 23754 16351 23810 16360
rect 23768 16046 23796 16351
rect 23952 16250 23980 16526
rect 23940 16244 23992 16250
rect 23940 16186 23992 16192
rect 23756 16040 23808 16046
rect 23756 15982 23808 15988
rect 23768 15881 23796 15982
rect 23940 15904 23992 15910
rect 23754 15872 23810 15881
rect 23940 15846 23992 15852
rect 23754 15807 23810 15816
rect 23952 15570 23980 15846
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 23848 15360 23900 15366
rect 23848 15302 23900 15308
rect 23860 15026 23888 15302
rect 23848 15020 23900 15026
rect 23848 14962 23900 14968
rect 23860 14278 23888 14962
rect 23940 14476 23992 14482
rect 23940 14418 23992 14424
rect 23848 14272 23900 14278
rect 23846 14240 23848 14249
rect 23900 14240 23902 14249
rect 23846 14175 23902 14184
rect 23756 13728 23808 13734
rect 23756 13670 23808 13676
rect 23768 13190 23796 13670
rect 23848 13524 23900 13530
rect 23952 13512 23980 14418
rect 24044 13938 24072 17070
rect 24124 16992 24176 16998
rect 24124 16934 24176 16940
rect 24308 16992 24360 16998
rect 24308 16934 24360 16940
rect 24136 16658 24164 16934
rect 24124 16652 24176 16658
rect 24124 16594 24176 16600
rect 24320 15910 24348 16934
rect 24400 16584 24452 16590
rect 24400 16526 24452 16532
rect 24308 15904 24360 15910
rect 24308 15846 24360 15852
rect 24320 15706 24348 15846
rect 24308 15700 24360 15706
rect 24308 15642 24360 15648
rect 24216 15360 24268 15366
rect 24216 15302 24268 15308
rect 24124 14952 24176 14958
rect 24124 14894 24176 14900
rect 24136 14482 24164 14894
rect 24228 14822 24256 15302
rect 24320 15162 24348 15642
rect 24412 15502 24440 16526
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24308 15156 24360 15162
rect 24308 15098 24360 15104
rect 24412 15026 24440 15438
rect 24490 15192 24546 15201
rect 24490 15127 24492 15136
rect 24544 15127 24546 15136
rect 24492 15098 24544 15104
rect 24400 15020 24452 15026
rect 24400 14962 24452 14968
rect 24216 14816 24268 14822
rect 24216 14758 24268 14764
rect 24124 14476 24176 14482
rect 24124 14418 24176 14424
rect 24032 13932 24084 13938
rect 24032 13874 24084 13880
rect 23900 13484 23980 13512
rect 23848 13466 23900 13472
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23768 12374 23796 13126
rect 23860 12782 23888 13466
rect 24136 13394 24164 14418
rect 24228 14278 24256 14758
rect 24308 14408 24360 14414
rect 24308 14350 24360 14356
rect 24216 14272 24268 14278
rect 24216 14214 24268 14220
rect 24228 13734 24256 14214
rect 24320 14074 24348 14350
rect 24308 14068 24360 14074
rect 24308 14010 24360 14016
rect 24400 13864 24452 13870
rect 24400 13806 24452 13812
rect 24216 13728 24268 13734
rect 24216 13670 24268 13676
rect 24124 13388 24176 13394
rect 24044 13348 24124 13376
rect 24044 12918 24072 13348
rect 24124 13330 24176 13336
rect 24216 13320 24268 13326
rect 24216 13262 24268 13268
rect 24124 12980 24176 12986
rect 24124 12922 24176 12928
rect 24032 12912 24084 12918
rect 24032 12854 24084 12860
rect 23848 12776 23900 12782
rect 23848 12718 23900 12724
rect 23756 12368 23808 12374
rect 23756 12310 23808 12316
rect 23756 12164 23808 12170
rect 23756 12106 23808 12112
rect 23768 11354 23796 12106
rect 23860 11898 23888 12718
rect 23940 12708 23992 12714
rect 23940 12650 23992 12656
rect 23848 11892 23900 11898
rect 23848 11834 23900 11840
rect 23756 11348 23808 11354
rect 23756 11290 23808 11296
rect 23768 11150 23796 11290
rect 23756 11144 23808 11150
rect 23756 11086 23808 11092
rect 23662 7984 23718 7993
rect 23662 7919 23718 7928
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23480 5772 23532 5778
rect 23480 5714 23532 5720
rect 23848 5772 23900 5778
rect 23848 5714 23900 5720
rect 23480 5568 23532 5574
rect 23480 5510 23532 5516
rect 23492 5166 23520 5510
rect 23860 5370 23888 5714
rect 23848 5364 23900 5370
rect 23848 5306 23900 5312
rect 23480 5160 23532 5166
rect 23480 5102 23532 5108
rect 23386 2680 23442 2689
rect 23386 2615 23442 2624
rect 23112 2440 23164 2446
rect 23112 2382 23164 2388
rect 23952 800 23980 12650
rect 24136 12170 24164 12922
rect 24228 12850 24256 13262
rect 24216 12844 24268 12850
rect 24216 12786 24268 12792
rect 24124 12164 24176 12170
rect 24124 12106 24176 12112
rect 24124 11892 24176 11898
rect 24124 11834 24176 11840
rect 24032 11688 24084 11694
rect 24032 11630 24084 11636
rect 24044 11354 24072 11630
rect 24032 11348 24084 11354
rect 24032 11290 24084 11296
rect 24136 11218 24164 11834
rect 24124 11212 24176 11218
rect 24124 11154 24176 11160
rect 24136 10810 24164 11154
rect 24124 10804 24176 10810
rect 24124 10746 24176 10752
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 24136 10198 24164 10542
rect 24124 10192 24176 10198
rect 24124 10134 24176 10140
rect 24412 10130 24440 13806
rect 24492 12640 24544 12646
rect 24492 12582 24544 12588
rect 24504 12306 24532 12582
rect 24492 12300 24544 12306
rect 24492 12242 24544 12248
rect 24400 10124 24452 10130
rect 24400 10066 24452 10072
rect 24400 9512 24452 9518
rect 24400 9454 24452 9460
rect 24412 9178 24440 9454
rect 24400 9172 24452 9178
rect 24400 9114 24452 9120
rect 24596 5681 24624 29582
rect 24780 29034 24808 29582
rect 24872 29238 24900 30194
rect 24860 29232 24912 29238
rect 24860 29174 24912 29180
rect 24872 29102 24900 29174
rect 25056 29170 25084 30738
rect 25136 29572 25188 29578
rect 25136 29514 25188 29520
rect 25044 29164 25096 29170
rect 25044 29106 25096 29112
rect 24860 29096 24912 29102
rect 24860 29038 24912 29044
rect 24952 29096 25004 29102
rect 24952 29038 25004 29044
rect 24768 29028 24820 29034
rect 24768 28970 24820 28976
rect 24674 27568 24730 27577
rect 24674 27503 24676 27512
rect 24728 27503 24730 27512
rect 24676 27474 24728 27480
rect 24780 27470 24808 28970
rect 24964 28626 24992 29038
rect 25056 29034 25084 29106
rect 25044 29028 25096 29034
rect 25044 28970 25096 28976
rect 25148 28966 25176 29514
rect 25228 29028 25280 29034
rect 25228 28970 25280 28976
rect 25136 28960 25188 28966
rect 25136 28902 25188 28908
rect 24952 28620 25004 28626
rect 24952 28562 25004 28568
rect 24860 28076 24912 28082
rect 24860 28018 24912 28024
rect 24872 27985 24900 28018
rect 24858 27976 24914 27985
rect 24858 27911 24914 27920
rect 24768 27464 24820 27470
rect 24768 27406 24820 27412
rect 24780 27130 24808 27406
rect 24768 27124 24820 27130
rect 24768 27066 24820 27072
rect 24780 27033 24808 27066
rect 24766 27024 24822 27033
rect 24766 26959 24822 26968
rect 24872 26926 24900 27911
rect 25240 26994 25268 28970
rect 25332 28744 25360 32422
rect 25502 32056 25558 32065
rect 25502 31991 25558 32000
rect 25516 31890 25544 31991
rect 25412 31884 25464 31890
rect 25412 31826 25464 31832
rect 25504 31884 25556 31890
rect 25504 31826 25556 31832
rect 25424 31482 25452 31826
rect 25792 31793 25820 40996
rect 26252 39098 26280 40996
rect 26240 39092 26292 39098
rect 26240 39034 26292 39040
rect 26148 38820 26200 38826
rect 26148 38762 26200 38768
rect 26056 38752 26108 38758
rect 26056 38694 26108 38700
rect 26160 38706 26188 38762
rect 26068 38350 26096 38694
rect 26160 38678 26280 38706
rect 26056 38344 26108 38350
rect 26056 38286 26108 38292
rect 26068 37670 26096 38286
rect 26056 37664 26108 37670
rect 26056 37606 26108 37612
rect 26068 37330 26096 37606
rect 26056 37324 26108 37330
rect 26056 37266 26108 37272
rect 26068 36718 26096 37266
rect 26056 36712 26108 36718
rect 26056 36654 26108 36660
rect 26252 33658 26280 38678
rect 26712 37874 26740 40996
rect 26884 40112 26936 40118
rect 26884 40054 26936 40060
rect 26790 38584 26846 38593
rect 26790 38519 26846 38528
rect 26804 38418 26832 38519
rect 26792 38412 26844 38418
rect 26792 38354 26844 38360
rect 26700 37868 26752 37874
rect 26700 37810 26752 37816
rect 26804 37466 26832 38354
rect 26792 37460 26844 37466
rect 26792 37402 26844 37408
rect 26792 35556 26844 35562
rect 26792 35498 26844 35504
rect 26424 34400 26476 34406
rect 26424 34342 26476 34348
rect 26240 33652 26292 33658
rect 26240 33594 26292 33600
rect 26436 33522 26464 34342
rect 26424 33516 26476 33522
rect 26424 33458 26476 33464
rect 26436 32026 26464 33458
rect 26424 32020 26476 32026
rect 26424 31962 26476 31968
rect 26700 31884 26752 31890
rect 26700 31826 26752 31832
rect 26516 31816 26568 31822
rect 25778 31784 25834 31793
rect 26516 31758 26568 31764
rect 25778 31719 25834 31728
rect 25964 31680 26016 31686
rect 25964 31622 26016 31628
rect 25412 31476 25464 31482
rect 25412 31418 25464 31424
rect 25424 28937 25452 31418
rect 25976 31210 26004 31622
rect 26528 31346 26556 31758
rect 26516 31340 26568 31346
rect 26516 31282 26568 31288
rect 25964 31204 26016 31210
rect 25964 31146 26016 31152
rect 26528 31142 26556 31282
rect 26056 31136 26108 31142
rect 26056 31078 26108 31084
rect 26516 31136 26568 31142
rect 26516 31078 26568 31084
rect 25596 30728 25648 30734
rect 25596 30670 25648 30676
rect 25608 30190 25636 30670
rect 26068 30598 26096 31078
rect 26056 30592 26108 30598
rect 26056 30534 26108 30540
rect 25596 30184 25648 30190
rect 25596 30126 25648 30132
rect 26068 29578 26096 30534
rect 26148 30184 26200 30190
rect 26148 30126 26200 30132
rect 26056 29572 26108 29578
rect 26056 29514 26108 29520
rect 26068 29102 26096 29514
rect 26160 29510 26188 30126
rect 26424 30048 26476 30054
rect 26424 29990 26476 29996
rect 26238 29744 26294 29753
rect 26238 29679 26294 29688
rect 26148 29504 26200 29510
rect 26146 29472 26148 29481
rect 26200 29472 26202 29481
rect 26146 29407 26202 29416
rect 26056 29096 26108 29102
rect 26056 29038 26108 29044
rect 25410 28928 25466 28937
rect 25410 28863 25466 28872
rect 25332 28716 25636 28744
rect 25320 28620 25372 28626
rect 25320 28562 25372 28568
rect 25412 28620 25464 28626
rect 25412 28562 25464 28568
rect 25332 28257 25360 28562
rect 25318 28248 25374 28257
rect 25424 28218 25452 28562
rect 25318 28183 25374 28192
rect 25412 28212 25464 28218
rect 25412 28154 25464 28160
rect 25412 28008 25464 28014
rect 25412 27950 25464 27956
rect 25320 27872 25372 27878
rect 25320 27814 25372 27820
rect 25332 27305 25360 27814
rect 25424 27334 25452 27950
rect 25504 27940 25556 27946
rect 25504 27882 25556 27888
rect 25516 27441 25544 27882
rect 25502 27432 25558 27441
rect 25502 27367 25558 27376
rect 25412 27328 25464 27334
rect 25318 27296 25374 27305
rect 25412 27270 25464 27276
rect 25318 27231 25374 27240
rect 25228 26988 25280 26994
rect 25228 26930 25280 26936
rect 24860 26920 24912 26926
rect 24860 26862 24912 26868
rect 24872 26518 24900 26862
rect 24860 26512 24912 26518
rect 24860 26454 24912 26460
rect 25332 26042 25360 27231
rect 25424 26994 25452 27270
rect 25412 26988 25464 26994
rect 25412 26930 25464 26936
rect 25320 26036 25372 26042
rect 25320 25978 25372 25984
rect 25044 25696 25096 25702
rect 25044 25638 25096 25644
rect 25056 25265 25084 25638
rect 25608 25362 25636 28716
rect 25964 26920 26016 26926
rect 25964 26862 26016 26868
rect 25976 26586 26004 26862
rect 25964 26580 26016 26586
rect 25964 26522 26016 26528
rect 25778 25800 25834 25809
rect 25778 25735 25834 25744
rect 25596 25356 25648 25362
rect 25596 25298 25648 25304
rect 25042 25256 25098 25265
rect 25042 25191 25098 25200
rect 25688 25220 25740 25226
rect 25688 25162 25740 25168
rect 25700 24750 25728 25162
rect 25596 24744 25648 24750
rect 25596 24686 25648 24692
rect 25688 24744 25740 24750
rect 25688 24686 25740 24692
rect 25502 24304 25558 24313
rect 25502 24239 25504 24248
rect 25556 24239 25558 24248
rect 25504 24210 25556 24216
rect 24860 23792 24912 23798
rect 24858 23760 24860 23769
rect 24912 23760 24914 23769
rect 24858 23695 24914 23704
rect 25318 23624 25374 23633
rect 25318 23559 25374 23568
rect 25332 23526 25360 23559
rect 25516 23526 25544 24210
rect 25320 23520 25372 23526
rect 25320 23462 25372 23468
rect 25504 23520 25556 23526
rect 25504 23462 25556 23468
rect 25516 22642 25544 23462
rect 25608 23322 25636 24686
rect 25596 23316 25648 23322
rect 25596 23258 25648 23264
rect 25608 22710 25636 23258
rect 25596 22704 25648 22710
rect 25596 22646 25648 22652
rect 25504 22636 25556 22642
rect 25504 22578 25556 22584
rect 25504 21480 25556 21486
rect 25504 21422 25556 21428
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24688 20602 24716 20946
rect 24768 20936 24820 20942
rect 24768 20878 24820 20884
rect 25228 20936 25280 20942
rect 25228 20878 25280 20884
rect 24676 20596 24728 20602
rect 24676 20538 24728 20544
rect 24780 20330 24808 20878
rect 24768 20324 24820 20330
rect 24768 20266 24820 20272
rect 24676 20052 24728 20058
rect 24676 19994 24728 20000
rect 24688 17898 24716 19994
rect 24780 19961 24808 20266
rect 25240 20233 25268 20878
rect 25226 20224 25282 20233
rect 25226 20159 25282 20168
rect 24766 19952 24822 19961
rect 24766 19887 24822 19896
rect 25228 19916 25280 19922
rect 25228 19858 25280 19864
rect 25240 19242 25268 19858
rect 25410 19680 25466 19689
rect 25410 19615 25466 19624
rect 25320 19304 25372 19310
rect 25320 19246 25372 19252
rect 25228 19236 25280 19242
rect 25228 19178 25280 19184
rect 25136 18216 25188 18222
rect 25136 18158 25188 18164
rect 24768 18080 24820 18086
rect 24820 18040 24900 18068
rect 24768 18022 24820 18028
rect 24688 17870 24808 17898
rect 24676 16652 24728 16658
rect 24676 16594 24728 16600
rect 24688 15978 24716 16594
rect 24676 15972 24728 15978
rect 24676 15914 24728 15920
rect 24688 15638 24716 15914
rect 24676 15632 24728 15638
rect 24676 15574 24728 15580
rect 24676 12912 24728 12918
rect 24676 12854 24728 12860
rect 24688 12442 24716 12854
rect 24676 12436 24728 12442
rect 24676 12378 24728 12384
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 24688 9353 24716 9454
rect 24674 9344 24730 9353
rect 24674 9279 24730 9288
rect 24780 7936 24808 17870
rect 24872 16794 24900 18040
rect 24952 16992 25004 16998
rect 24952 16934 25004 16940
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 24964 16658 24992 16934
rect 24952 16652 25004 16658
rect 24952 16594 25004 16600
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 25044 16448 25096 16454
rect 25044 16390 25096 16396
rect 24872 16046 24900 16390
rect 25056 16182 25084 16390
rect 25044 16176 25096 16182
rect 25044 16118 25096 16124
rect 24860 16040 24912 16046
rect 24860 15982 24912 15988
rect 25056 15706 25084 16118
rect 25044 15700 25096 15706
rect 25044 15642 25096 15648
rect 25148 15201 25176 18158
rect 25240 16250 25268 19178
rect 25332 16946 25360 19246
rect 25424 17882 25452 19615
rect 25412 17876 25464 17882
rect 25412 17818 25464 17824
rect 25424 17678 25452 17818
rect 25412 17672 25464 17678
rect 25412 17614 25464 17620
rect 25516 17513 25544 21422
rect 25688 20800 25740 20806
rect 25688 20742 25740 20748
rect 25594 20632 25650 20641
rect 25594 20567 25650 20576
rect 25608 20466 25636 20567
rect 25596 20460 25648 20466
rect 25596 20402 25648 20408
rect 25608 18698 25636 20402
rect 25700 20398 25728 20742
rect 25688 20392 25740 20398
rect 25688 20334 25740 20340
rect 25700 19990 25728 20334
rect 25688 19984 25740 19990
rect 25688 19926 25740 19932
rect 25700 19446 25728 19926
rect 25792 19446 25820 25735
rect 25964 25356 26016 25362
rect 25964 25298 26016 25304
rect 25872 25152 25924 25158
rect 25872 25094 25924 25100
rect 25884 24818 25912 25094
rect 25872 24812 25924 24818
rect 25872 24754 25924 24760
rect 25884 23866 25912 24754
rect 25976 24614 26004 25298
rect 25964 24608 26016 24614
rect 25964 24550 26016 24556
rect 25976 24342 26004 24550
rect 25964 24336 26016 24342
rect 25964 24278 26016 24284
rect 26068 24138 26096 29038
rect 26252 28762 26280 29679
rect 26332 29504 26384 29510
rect 26332 29446 26384 29452
rect 26240 28756 26292 28762
rect 26240 28698 26292 28704
rect 26344 28558 26372 29446
rect 26436 28966 26464 29990
rect 26528 29714 26556 31078
rect 26712 30598 26740 31826
rect 26804 30666 26832 35498
rect 26896 34610 26924 40054
rect 27344 39092 27396 39098
rect 27344 39034 27396 39040
rect 27356 38894 27384 39034
rect 27344 38888 27396 38894
rect 27344 38830 27396 38836
rect 27632 37346 27660 40996
rect 27896 38208 27948 38214
rect 27896 38150 27948 38156
rect 27540 37318 27660 37346
rect 27540 36922 27568 37318
rect 27528 36916 27580 36922
rect 27528 36858 27580 36864
rect 27618 35184 27674 35193
rect 27618 35119 27674 35128
rect 27342 34640 27398 34649
rect 26884 34604 26936 34610
rect 27342 34575 27398 34584
rect 26884 34546 26936 34552
rect 27160 34536 27212 34542
rect 27160 34478 27212 34484
rect 27172 34202 27200 34478
rect 27160 34196 27212 34202
rect 27160 34138 27212 34144
rect 27068 33516 27120 33522
rect 27068 33458 27120 33464
rect 26976 32972 27028 32978
rect 26976 32914 27028 32920
rect 26988 32366 27016 32914
rect 26976 32360 27028 32366
rect 26976 32302 27028 32308
rect 26988 31958 27016 32302
rect 26976 31952 27028 31958
rect 26976 31894 27028 31900
rect 26976 31136 27028 31142
rect 26976 31078 27028 31084
rect 26988 30734 27016 31078
rect 26976 30728 27028 30734
rect 26976 30670 27028 30676
rect 26792 30660 26844 30666
rect 26792 30602 26844 30608
rect 26700 30592 26752 30598
rect 26700 30534 26752 30540
rect 26608 30252 26660 30258
rect 26608 30194 26660 30200
rect 26516 29708 26568 29714
rect 26516 29650 26568 29656
rect 26528 29170 26556 29650
rect 26516 29164 26568 29170
rect 26516 29106 26568 29112
rect 26424 28960 26476 28966
rect 26424 28902 26476 28908
rect 26436 28626 26464 28902
rect 26620 28694 26648 30194
rect 26712 29034 26740 30534
rect 26988 29510 27016 30670
rect 26976 29504 27028 29510
rect 26976 29446 27028 29452
rect 26700 29028 26752 29034
rect 26700 28970 26752 28976
rect 26608 28688 26660 28694
rect 26884 28688 26936 28694
rect 26608 28630 26660 28636
rect 26804 28648 26884 28676
rect 26424 28620 26476 28626
rect 26424 28562 26476 28568
rect 26332 28552 26384 28558
rect 26332 28494 26384 28500
rect 26344 27878 26372 28494
rect 26436 28014 26464 28562
rect 26424 28008 26476 28014
rect 26424 27950 26476 27956
rect 26332 27872 26384 27878
rect 26332 27814 26384 27820
rect 26148 26784 26200 26790
rect 26148 26726 26200 26732
rect 26240 26784 26292 26790
rect 26240 26726 26292 26732
rect 26160 26625 26188 26726
rect 26146 26616 26202 26625
rect 26146 26551 26202 26560
rect 26252 26518 26280 26726
rect 26240 26512 26292 26518
rect 26238 26480 26240 26489
rect 26292 26480 26294 26489
rect 26238 26415 26294 26424
rect 26240 26376 26292 26382
rect 26160 26324 26240 26330
rect 26160 26318 26292 26324
rect 26160 26302 26280 26318
rect 26160 26042 26188 26302
rect 26344 26194 26372 27814
rect 26436 27334 26464 27950
rect 26620 27538 26648 28630
rect 26608 27532 26660 27538
rect 26608 27474 26660 27480
rect 26804 27402 26832 28648
rect 26884 28630 26936 28636
rect 26884 28552 26936 28558
rect 26884 28494 26936 28500
rect 26792 27396 26844 27402
rect 26792 27338 26844 27344
rect 26424 27328 26476 27334
rect 26424 27270 26476 27276
rect 26252 26166 26372 26194
rect 26148 26036 26200 26042
rect 26148 25978 26200 25984
rect 26252 24750 26280 26166
rect 26436 25226 26464 27270
rect 26608 26512 26660 26518
rect 26608 26454 26660 26460
rect 26514 25936 26570 25945
rect 26514 25871 26570 25880
rect 26424 25220 26476 25226
rect 26424 25162 26476 25168
rect 26240 24744 26292 24750
rect 26240 24686 26292 24692
rect 26252 24410 26280 24686
rect 26424 24676 26476 24682
rect 26424 24618 26476 24624
rect 26240 24404 26292 24410
rect 26240 24346 26292 24352
rect 26056 24132 26108 24138
rect 26056 24074 26108 24080
rect 25872 23860 25924 23866
rect 25872 23802 25924 23808
rect 25884 23662 25912 23802
rect 25872 23656 25924 23662
rect 25872 23598 25924 23604
rect 25964 23180 26016 23186
rect 25964 23122 26016 23128
rect 25976 22982 26004 23122
rect 26068 22982 26096 24074
rect 26238 23352 26294 23361
rect 26238 23287 26240 23296
rect 26292 23287 26294 23296
rect 26240 23258 26292 23264
rect 25964 22976 26016 22982
rect 25964 22918 26016 22924
rect 26056 22976 26108 22982
rect 26056 22918 26108 22924
rect 26332 22976 26384 22982
rect 26332 22918 26384 22924
rect 25976 22574 26004 22918
rect 25964 22568 26016 22574
rect 25962 22536 25964 22545
rect 26016 22536 26018 22545
rect 25962 22471 26018 22480
rect 25976 22445 26004 22471
rect 26344 22234 26372 22918
rect 26332 22228 26384 22234
rect 26332 22170 26384 22176
rect 25872 21888 25924 21894
rect 25872 21830 25924 21836
rect 25884 21554 25912 21830
rect 26056 21684 26108 21690
rect 26056 21626 26108 21632
rect 26068 21593 26096 21626
rect 26054 21584 26110 21593
rect 25872 21548 25924 21554
rect 26054 21519 26110 21528
rect 25872 21490 25924 21496
rect 25884 20346 25912 21490
rect 25964 21480 26016 21486
rect 25964 21422 26016 21428
rect 25976 21146 26004 21422
rect 25964 21140 26016 21146
rect 25964 21082 26016 21088
rect 25964 20528 26016 20534
rect 25962 20496 25964 20505
rect 26016 20496 26018 20505
rect 25962 20431 26018 20440
rect 25964 20392 26016 20398
rect 25884 20340 25964 20346
rect 25884 20334 26016 20340
rect 25884 20318 26004 20334
rect 25976 20058 26004 20318
rect 25964 20052 26016 20058
rect 25964 19994 26016 20000
rect 25962 19952 26018 19961
rect 25962 19887 26018 19896
rect 25688 19440 25740 19446
rect 25688 19382 25740 19388
rect 25780 19440 25832 19446
rect 25780 19382 25832 19388
rect 25700 19310 25728 19382
rect 25688 19304 25740 19310
rect 25688 19246 25740 19252
rect 25700 18902 25728 19246
rect 25976 19174 26004 19887
rect 26068 19786 26096 21519
rect 26436 21010 26464 24618
rect 26528 21622 26556 25871
rect 26516 21616 26568 21622
rect 26516 21558 26568 21564
rect 26424 21004 26476 21010
rect 26424 20946 26476 20952
rect 26436 20602 26464 20946
rect 26424 20596 26476 20602
rect 26252 20556 26424 20584
rect 26148 20324 26200 20330
rect 26148 20266 26200 20272
rect 26056 19780 26108 19786
rect 26056 19722 26108 19728
rect 26056 19304 26108 19310
rect 26056 19246 26108 19252
rect 25964 19168 26016 19174
rect 25964 19110 26016 19116
rect 25688 18896 25740 18902
rect 25688 18838 25740 18844
rect 25596 18692 25648 18698
rect 25596 18634 25648 18640
rect 25700 18222 25728 18838
rect 25780 18284 25832 18290
rect 25780 18226 25832 18232
rect 25688 18216 25740 18222
rect 25688 18158 25740 18164
rect 25502 17504 25558 17513
rect 25502 17439 25558 17448
rect 25332 16918 25452 16946
rect 25228 16244 25280 16250
rect 25228 16186 25280 16192
rect 25320 16040 25372 16046
rect 25320 15982 25372 15988
rect 25332 15502 25360 15982
rect 25424 15609 25452 16918
rect 25410 15600 25466 15609
rect 25410 15535 25466 15544
rect 25504 15564 25556 15570
rect 25504 15506 25556 15512
rect 25320 15496 25372 15502
rect 25320 15438 25372 15444
rect 25134 15192 25190 15201
rect 25134 15127 25190 15136
rect 25516 14822 25544 15506
rect 25504 14816 25556 14822
rect 25504 14758 25556 14764
rect 25228 14408 25280 14414
rect 25516 14362 25544 14758
rect 25280 14356 25544 14362
rect 25228 14350 25544 14356
rect 25240 14334 25544 14350
rect 25318 14240 25374 14249
rect 25318 14175 25374 14184
rect 25044 13796 25096 13802
rect 25044 13738 25096 13744
rect 25056 13530 25084 13738
rect 25044 13524 25096 13530
rect 25044 13466 25096 13472
rect 24860 12300 24912 12306
rect 24860 12242 24912 12248
rect 24872 11694 24900 12242
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 25056 12186 25084 13466
rect 25228 13388 25280 13394
rect 25228 13330 25280 13336
rect 25240 12986 25268 13330
rect 25228 12980 25280 12986
rect 25228 12922 25280 12928
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 24964 11558 24992 12174
rect 25056 12170 25176 12186
rect 25056 12164 25188 12170
rect 25056 12158 25136 12164
rect 25136 12106 25188 12112
rect 25044 12096 25096 12102
rect 25044 12038 25096 12044
rect 25056 11694 25084 12038
rect 25148 11898 25176 12106
rect 25136 11892 25188 11898
rect 25136 11834 25188 11840
rect 25240 11830 25268 12922
rect 25228 11824 25280 11830
rect 25228 11766 25280 11772
rect 25044 11688 25096 11694
rect 25044 11630 25096 11636
rect 24952 11552 25004 11558
rect 24872 11500 24952 11506
rect 24872 11494 25004 11500
rect 24872 11478 24992 11494
rect 24872 11218 24900 11478
rect 25240 11286 25268 11766
rect 25228 11280 25280 11286
rect 25228 11222 25280 11228
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 24872 10606 24900 11154
rect 25332 10810 25360 14175
rect 25412 13932 25464 13938
rect 25412 13874 25464 13880
rect 25424 13530 25452 13874
rect 25412 13524 25464 13530
rect 25412 13466 25464 13472
rect 25516 12850 25544 14334
rect 25504 12844 25556 12850
rect 25504 12786 25556 12792
rect 25594 12336 25650 12345
rect 25594 12271 25596 12280
rect 25648 12271 25650 12280
rect 25596 12242 25648 12248
rect 25596 12096 25648 12102
rect 25596 12038 25648 12044
rect 25320 10804 25372 10810
rect 25320 10746 25372 10752
rect 24860 10600 24912 10606
rect 24860 10542 24912 10548
rect 25608 10266 25636 12038
rect 25596 10260 25648 10266
rect 25596 10202 25648 10208
rect 25504 10124 25556 10130
rect 25504 10066 25556 10072
rect 25516 9110 25544 10066
rect 25792 9761 25820 18226
rect 25976 17746 26004 19110
rect 26068 18970 26096 19246
rect 26160 18986 26188 20266
rect 26252 19281 26280 20556
rect 26424 20538 26476 20544
rect 26332 20324 26384 20330
rect 26332 20266 26384 20272
rect 26344 20058 26372 20266
rect 26332 20052 26384 20058
rect 26332 19994 26384 20000
rect 26344 19378 26372 19994
rect 26332 19372 26384 19378
rect 26332 19314 26384 19320
rect 26238 19272 26294 19281
rect 26238 19207 26294 19216
rect 26160 18970 26280 18986
rect 26056 18964 26108 18970
rect 26160 18964 26292 18970
rect 26160 18958 26240 18964
rect 26056 18906 26108 18912
rect 26240 18906 26292 18912
rect 26068 18222 26096 18906
rect 26148 18692 26200 18698
rect 26148 18634 26200 18640
rect 26056 18216 26108 18222
rect 26056 18158 26108 18164
rect 25964 17740 26016 17746
rect 25964 17682 26016 17688
rect 25964 17536 26016 17542
rect 25964 17478 26016 17484
rect 25872 17332 25924 17338
rect 25872 17274 25924 17280
rect 25884 16454 25912 17274
rect 25976 17134 26004 17478
rect 26056 17264 26108 17270
rect 26056 17206 26108 17212
rect 25964 17128 26016 17134
rect 25964 17070 26016 17076
rect 25976 16726 26004 17070
rect 25964 16720 26016 16726
rect 25964 16662 26016 16668
rect 25872 16448 25924 16454
rect 25872 16390 25924 16396
rect 25976 15638 26004 16662
rect 26068 16658 26096 17206
rect 26056 16652 26108 16658
rect 26056 16594 26108 16600
rect 26056 16176 26108 16182
rect 26056 16118 26108 16124
rect 25964 15632 26016 15638
rect 25964 15574 26016 15580
rect 25872 15088 25924 15094
rect 25872 15030 25924 15036
rect 25884 14822 25912 15030
rect 25976 14958 26004 15574
rect 26068 15502 26096 16118
rect 26160 16114 26188 18634
rect 26516 17740 26568 17746
rect 26516 17682 26568 17688
rect 26528 17377 26556 17682
rect 26238 17368 26294 17377
rect 26238 17303 26294 17312
rect 26514 17368 26570 17377
rect 26514 17303 26570 17312
rect 26252 16425 26280 17303
rect 26620 17252 26648 26454
rect 26804 26450 26832 27338
rect 26896 26926 26924 28494
rect 26976 27396 27028 27402
rect 26976 27338 27028 27344
rect 26988 27130 27016 27338
rect 26976 27124 27028 27130
rect 26976 27066 27028 27072
rect 26988 26926 27016 27066
rect 26884 26920 26936 26926
rect 26884 26862 26936 26868
rect 26976 26920 27028 26926
rect 26976 26862 27028 26868
rect 26792 26444 26844 26450
rect 26792 26386 26844 26392
rect 26804 25158 26832 26386
rect 26884 26376 26936 26382
rect 26884 26318 26936 26324
rect 26896 26042 26924 26318
rect 27080 26217 27108 33458
rect 27252 33448 27304 33454
rect 27252 33390 27304 33396
rect 27160 33312 27212 33318
rect 27160 33254 27212 33260
rect 27172 30326 27200 33254
rect 27264 32842 27292 33390
rect 27356 32978 27384 34575
rect 27632 34513 27660 35119
rect 27618 34504 27674 34513
rect 27618 34439 27674 34448
rect 27908 34202 27936 38150
rect 27896 34196 27948 34202
rect 27896 34138 27948 34144
rect 27908 33454 27936 34138
rect 27988 34060 28040 34066
rect 27988 34002 28040 34008
rect 28000 33862 28028 34002
rect 27988 33856 28040 33862
rect 27988 33798 28040 33804
rect 27528 33448 27580 33454
rect 27528 33390 27580 33396
rect 27896 33448 27948 33454
rect 27896 33390 27948 33396
rect 27344 32972 27396 32978
rect 27344 32914 27396 32920
rect 27252 32836 27304 32842
rect 27252 32778 27304 32784
rect 27356 32570 27384 32914
rect 27436 32904 27488 32910
rect 27436 32846 27488 32852
rect 27344 32564 27396 32570
rect 27344 32506 27396 32512
rect 27448 32298 27476 32846
rect 27436 32292 27488 32298
rect 27436 32234 27488 32240
rect 27436 31884 27488 31890
rect 27436 31826 27488 31832
rect 27252 31680 27304 31686
rect 27252 31622 27304 31628
rect 27264 31142 27292 31622
rect 27448 31142 27476 31826
rect 27540 31210 27568 33390
rect 27804 32768 27856 32774
rect 27804 32710 27856 32716
rect 27816 32366 27844 32710
rect 27804 32360 27856 32366
rect 27804 32302 27856 32308
rect 27816 31346 27844 32302
rect 28000 32026 28028 33798
rect 28092 33674 28120 40996
rect 28092 33646 28488 33674
rect 28264 33312 28316 33318
rect 28264 33254 28316 33260
rect 28172 33108 28224 33114
rect 28172 33050 28224 33056
rect 28184 32366 28212 33050
rect 28172 32360 28224 32366
rect 28172 32302 28224 32308
rect 27988 32020 28040 32026
rect 27988 31962 28040 31968
rect 27986 31920 28042 31929
rect 28276 31890 28304 33254
rect 28356 32972 28408 32978
rect 28356 32914 28408 32920
rect 28368 32570 28396 32914
rect 28460 32586 28488 33646
rect 28552 32722 28580 40996
rect 28724 38820 28776 38826
rect 28724 38762 28776 38768
rect 28736 32881 28764 38762
rect 29472 38418 29500 40996
rect 29460 38412 29512 38418
rect 29460 38354 29512 38360
rect 29472 38010 29500 38354
rect 29460 38004 29512 38010
rect 29460 37946 29512 37952
rect 29276 35284 29328 35290
rect 29276 35226 29328 35232
rect 29288 34542 29316 35226
rect 29932 34610 29960 40996
rect 30012 38344 30064 38350
rect 30012 38286 30064 38292
rect 30024 38010 30052 38286
rect 30852 38185 30880 40996
rect 31024 38208 31076 38214
rect 30838 38176 30894 38185
rect 31024 38150 31076 38156
rect 30838 38111 30894 38120
rect 30012 38004 30064 38010
rect 30012 37946 30064 37952
rect 30024 35290 30052 37946
rect 30562 37088 30618 37097
rect 30562 37023 30618 37032
rect 30012 35284 30064 35290
rect 30012 35226 30064 35232
rect 29920 34604 29972 34610
rect 29920 34546 29972 34552
rect 29276 34536 29328 34542
rect 29276 34478 29328 34484
rect 30378 34504 30434 34513
rect 29000 33856 29052 33862
rect 29000 33798 29052 33804
rect 29012 33130 29040 33798
rect 28920 33114 29040 33130
rect 29288 33114 29316 34478
rect 30576 34490 30604 37023
rect 30656 34672 30708 34678
rect 30654 34640 30656 34649
rect 30708 34640 30710 34649
rect 30654 34575 30710 34584
rect 30576 34462 30696 34490
rect 30378 34439 30434 34448
rect 30286 34232 30342 34241
rect 30286 34167 30342 34176
rect 30300 34066 30328 34167
rect 30288 34060 30340 34066
rect 30288 34002 30340 34008
rect 29644 33992 29696 33998
rect 29644 33934 29696 33940
rect 30196 33992 30248 33998
rect 30196 33934 30248 33940
rect 29656 33386 29684 33934
rect 30104 33856 30156 33862
rect 30104 33798 30156 33804
rect 30116 33454 30144 33798
rect 30208 33454 30236 33934
rect 30104 33448 30156 33454
rect 30196 33448 30248 33454
rect 30104 33390 30156 33396
rect 30194 33416 30196 33425
rect 30248 33416 30250 33425
rect 29644 33380 29696 33386
rect 29644 33322 29696 33328
rect 30012 33380 30064 33386
rect 30012 33322 30064 33328
rect 28908 33108 29040 33114
rect 28960 33102 29040 33108
rect 29276 33108 29328 33114
rect 28908 33050 28960 33056
rect 29276 33050 29328 33056
rect 29826 33008 29882 33017
rect 29000 32972 29052 32978
rect 29826 32943 29882 32952
rect 29000 32914 29052 32920
rect 28722 32872 28778 32881
rect 28722 32807 28778 32816
rect 28552 32694 28948 32722
rect 28356 32564 28408 32570
rect 28460 32558 28672 32586
rect 28356 32506 28408 32512
rect 27986 31855 28042 31864
rect 28264 31884 28316 31890
rect 27804 31340 27856 31346
rect 27804 31282 27856 31288
rect 27528 31204 27580 31210
rect 27528 31146 27580 31152
rect 27252 31136 27304 31142
rect 27252 31078 27304 31084
rect 27436 31136 27488 31142
rect 27436 31078 27488 31084
rect 27264 30802 27292 31078
rect 27448 30954 27476 31078
rect 27356 30926 27476 30954
rect 27540 30938 27568 31146
rect 27528 30932 27580 30938
rect 27356 30870 27384 30926
rect 27528 30874 27580 30880
rect 27344 30864 27396 30870
rect 27344 30806 27396 30812
rect 27252 30796 27304 30802
rect 27252 30738 27304 30744
rect 27528 30796 27580 30802
rect 27528 30738 27580 30744
rect 27160 30320 27212 30326
rect 27160 30262 27212 30268
rect 27264 30054 27292 30738
rect 27540 30274 27568 30738
rect 27804 30728 27856 30734
rect 27804 30670 27856 30676
rect 27540 30246 27660 30274
rect 27632 30172 27660 30246
rect 27712 30184 27764 30190
rect 27632 30144 27712 30172
rect 27712 30126 27764 30132
rect 27528 30116 27580 30122
rect 27528 30058 27580 30064
rect 27252 30048 27304 30054
rect 27252 29990 27304 29996
rect 27436 29572 27488 29578
rect 27436 29514 27488 29520
rect 27448 29102 27476 29514
rect 27436 29096 27488 29102
rect 27436 29038 27488 29044
rect 27160 29028 27212 29034
rect 27160 28970 27212 28976
rect 27066 26208 27122 26217
rect 27066 26143 27122 26152
rect 26884 26036 26936 26042
rect 26884 25978 26936 25984
rect 27172 25974 27200 28970
rect 27344 28416 27396 28422
rect 27344 28358 27396 28364
rect 27356 28014 27384 28358
rect 27344 28008 27396 28014
rect 27344 27950 27396 27956
rect 27252 27940 27304 27946
rect 27252 27882 27304 27888
rect 27264 27674 27292 27882
rect 27252 27668 27304 27674
rect 27252 27610 27304 27616
rect 27264 26518 27292 27610
rect 27436 26784 27488 26790
rect 27436 26726 27488 26732
rect 27252 26512 27304 26518
rect 27252 26454 27304 26460
rect 27160 25968 27212 25974
rect 27160 25910 27212 25916
rect 26884 25832 26936 25838
rect 26884 25774 26936 25780
rect 26792 25152 26844 25158
rect 26792 25094 26844 25100
rect 26804 22658 26832 25094
rect 26896 24342 26924 25774
rect 27448 25430 27476 26726
rect 27436 25424 27488 25430
rect 27436 25366 27488 25372
rect 27068 25152 27120 25158
rect 27068 25094 27120 25100
rect 27080 24886 27108 25094
rect 27252 24948 27304 24954
rect 27252 24890 27304 24896
rect 27068 24880 27120 24886
rect 27068 24822 27120 24828
rect 26884 24336 26936 24342
rect 26884 24278 26936 24284
rect 26896 23798 26924 24278
rect 26884 23792 26936 23798
rect 27080 23769 27108 24822
rect 27264 24274 27292 24890
rect 27252 24268 27304 24274
rect 27252 24210 27304 24216
rect 27264 23866 27292 24210
rect 27252 23860 27304 23866
rect 27252 23802 27304 23808
rect 26884 23734 26936 23740
rect 27066 23760 27122 23769
rect 27066 23695 27122 23704
rect 26884 23588 26936 23594
rect 26884 23530 26936 23536
rect 26896 23118 26924 23530
rect 27068 23316 27120 23322
rect 27068 23258 27120 23264
rect 26884 23112 26936 23118
rect 26884 23054 26936 23060
rect 26896 22778 26924 23054
rect 26884 22772 26936 22778
rect 26884 22714 26936 22720
rect 26804 22630 26924 22658
rect 26700 21140 26752 21146
rect 26700 21082 26752 21088
rect 26712 20777 26740 21082
rect 26698 20768 26754 20777
rect 26698 20703 26754 20712
rect 26792 19712 26844 19718
rect 26792 19654 26844 19660
rect 26804 19378 26832 19654
rect 26792 19372 26844 19378
rect 26792 19314 26844 19320
rect 26436 17224 26648 17252
rect 26332 16584 26384 16590
rect 26332 16526 26384 16532
rect 26238 16416 26294 16425
rect 26238 16351 26294 16360
rect 26240 16244 26292 16250
rect 26240 16186 26292 16192
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 26252 15910 26280 16186
rect 26240 15904 26292 15910
rect 26240 15846 26292 15852
rect 26056 15496 26108 15502
rect 26056 15438 26108 15444
rect 26068 15162 26096 15438
rect 26056 15156 26108 15162
rect 26056 15098 26108 15104
rect 25964 14952 26016 14958
rect 25964 14894 26016 14900
rect 25872 14816 25924 14822
rect 25872 14758 25924 14764
rect 25884 14006 25912 14758
rect 25976 14618 26004 14894
rect 25964 14612 26016 14618
rect 25964 14554 26016 14560
rect 25976 14074 26004 14554
rect 26068 14414 26096 15098
rect 26056 14408 26108 14414
rect 26056 14350 26108 14356
rect 26148 14272 26200 14278
rect 26148 14214 26200 14220
rect 26160 14074 26188 14214
rect 25964 14068 26016 14074
rect 25964 14010 26016 14016
rect 26148 14068 26200 14074
rect 26148 14010 26200 14016
rect 25872 14000 25924 14006
rect 25872 13942 25924 13948
rect 25976 13870 26004 14010
rect 25964 13864 26016 13870
rect 25964 13806 26016 13812
rect 26056 13388 26108 13394
rect 26056 13330 26108 13336
rect 25872 12844 25924 12850
rect 25872 12786 25924 12792
rect 25884 10810 25912 12786
rect 26068 12782 26096 13330
rect 26252 12866 26280 15846
rect 26344 15570 26372 16526
rect 26332 15564 26384 15570
rect 26332 15506 26384 15512
rect 26344 15162 26372 15506
rect 26332 15156 26384 15162
rect 26332 15098 26384 15104
rect 26332 15020 26384 15026
rect 26332 14962 26384 14968
rect 26344 14550 26372 14962
rect 26332 14544 26384 14550
rect 26332 14486 26384 14492
rect 26344 13938 26372 14486
rect 26332 13932 26384 13938
rect 26332 13874 26384 13880
rect 26332 12912 26384 12918
rect 26252 12860 26332 12866
rect 26252 12854 26384 12860
rect 26252 12838 26372 12854
rect 26056 12776 26108 12782
rect 26252 12764 26280 12838
rect 26056 12718 26108 12724
rect 26160 12736 26280 12764
rect 26332 12776 26384 12782
rect 26160 12102 26188 12736
rect 26332 12718 26384 12724
rect 26240 12640 26292 12646
rect 26240 12582 26292 12588
rect 26148 12096 26200 12102
rect 26148 12038 26200 12044
rect 26252 11354 26280 12582
rect 26344 12442 26372 12718
rect 26332 12436 26384 12442
rect 26332 12378 26384 12384
rect 26344 12306 26372 12378
rect 26332 12300 26384 12306
rect 26332 12242 26384 12248
rect 26240 11348 26292 11354
rect 26240 11290 26292 11296
rect 26240 11212 26292 11218
rect 26240 11154 26292 11160
rect 26252 10962 26280 11154
rect 26160 10934 26280 10962
rect 25872 10804 25924 10810
rect 25872 10746 25924 10752
rect 26160 10470 26188 10934
rect 26148 10464 26200 10470
rect 26148 10406 26200 10412
rect 26160 10130 26188 10406
rect 26148 10124 26200 10130
rect 26148 10066 26200 10072
rect 25778 9752 25834 9761
rect 25778 9687 25834 9696
rect 25780 9648 25832 9654
rect 25778 9616 25780 9625
rect 25832 9616 25834 9625
rect 25778 9551 25834 9560
rect 25962 9616 26018 9625
rect 25962 9551 26018 9560
rect 25976 9178 26004 9551
rect 26146 9208 26202 9217
rect 25964 9172 26016 9178
rect 26146 9143 26202 9152
rect 25964 9114 26016 9120
rect 25504 9104 25556 9110
rect 25504 9046 25556 9052
rect 26160 9042 26188 9143
rect 26148 9036 26200 9042
rect 26148 8978 26200 8984
rect 26160 8634 26188 8978
rect 26148 8628 26200 8634
rect 26148 8570 26200 8576
rect 24688 7908 24808 7936
rect 24582 5672 24638 5681
rect 24582 5607 24638 5616
rect 24688 3738 24716 7908
rect 24950 6216 25006 6225
rect 24950 6151 25006 6160
rect 24676 3732 24728 3738
rect 24676 3674 24728 3680
rect 24582 3632 24638 3641
rect 24582 3567 24638 3576
rect 24596 3194 24624 3567
rect 24584 3188 24636 3194
rect 24584 3130 24636 3136
rect 24860 2984 24912 2990
rect 24860 2926 24912 2932
rect 24398 2816 24454 2825
rect 24398 2751 24454 2760
rect 24412 800 24440 2751
rect 24872 2446 24900 2926
rect 24860 2440 24912 2446
rect 24860 2382 24912 2388
rect 24964 1442 24992 6151
rect 26238 5808 26294 5817
rect 26238 5743 26294 5752
rect 25412 5024 25464 5030
rect 25412 4966 25464 4972
rect 25424 4078 25452 4966
rect 25412 4072 25464 4078
rect 25412 4014 25464 4020
rect 25780 4072 25832 4078
rect 25780 4014 25832 4020
rect 25424 3398 25452 4014
rect 25412 3392 25464 3398
rect 25412 3334 25464 3340
rect 24872 1414 24992 1442
rect 24872 800 24900 1414
rect 25792 800 25820 4014
rect 26252 800 26280 5743
rect 26436 3194 26464 17224
rect 26792 17196 26844 17202
rect 26792 17138 26844 17144
rect 26516 16992 26568 16998
rect 26516 16934 26568 16940
rect 26528 16182 26556 16934
rect 26608 16788 26660 16794
rect 26608 16730 26660 16736
rect 26620 16454 26648 16730
rect 26700 16584 26752 16590
rect 26700 16526 26752 16532
rect 26608 16448 26660 16454
rect 26608 16390 26660 16396
rect 26516 16176 26568 16182
rect 26516 16118 26568 16124
rect 26712 16114 26740 16526
rect 26700 16108 26752 16114
rect 26700 16050 26752 16056
rect 26712 15026 26740 16050
rect 26804 15502 26832 17138
rect 26792 15496 26844 15502
rect 26792 15438 26844 15444
rect 26792 15360 26844 15366
rect 26792 15302 26844 15308
rect 26804 15094 26832 15302
rect 26792 15088 26844 15094
rect 26792 15030 26844 15036
rect 26700 15020 26752 15026
rect 26700 14962 26752 14968
rect 26608 14952 26660 14958
rect 26608 14894 26660 14900
rect 26516 14340 26568 14346
rect 26516 14282 26568 14288
rect 26528 14006 26556 14282
rect 26620 14074 26648 14894
rect 26700 14884 26752 14890
rect 26700 14826 26752 14832
rect 26712 14521 26740 14826
rect 26698 14512 26754 14521
rect 26698 14447 26754 14456
rect 26792 14476 26844 14482
rect 26792 14418 26844 14424
rect 26804 14074 26832 14418
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 26792 14068 26844 14074
rect 26792 14010 26844 14016
rect 26516 14000 26568 14006
rect 26516 13942 26568 13948
rect 26528 12646 26556 13942
rect 26700 13864 26752 13870
rect 26700 13806 26752 13812
rect 26712 13530 26740 13806
rect 26804 13530 26832 14010
rect 26700 13524 26752 13530
rect 26700 13466 26752 13472
rect 26792 13524 26844 13530
rect 26792 13466 26844 13472
rect 26700 12980 26752 12986
rect 26700 12922 26752 12928
rect 26608 12708 26660 12714
rect 26608 12650 26660 12656
rect 26516 12640 26568 12646
rect 26516 12582 26568 12588
rect 26620 12238 26648 12650
rect 26712 12442 26740 12922
rect 26792 12708 26844 12714
rect 26792 12650 26844 12656
rect 26700 12436 26752 12442
rect 26700 12378 26752 12384
rect 26608 12232 26660 12238
rect 26608 12174 26660 12180
rect 26712 11694 26740 12378
rect 26804 12073 26832 12650
rect 26790 12064 26846 12073
rect 26790 11999 26846 12008
rect 26792 11756 26844 11762
rect 26792 11698 26844 11704
rect 26700 11688 26752 11694
rect 26700 11630 26752 11636
rect 26804 10130 26832 11698
rect 26792 10124 26844 10130
rect 26792 10066 26844 10072
rect 26804 9722 26832 10066
rect 26792 9716 26844 9722
rect 26792 9658 26844 9664
rect 26516 4616 26568 4622
rect 26516 4558 26568 4564
rect 26792 4616 26844 4622
rect 26792 4558 26844 4564
rect 26528 3398 26556 4558
rect 26804 4321 26832 4558
rect 26790 4312 26846 4321
rect 26790 4247 26792 4256
rect 26844 4247 26846 4256
rect 26792 4218 26844 4224
rect 26804 4187 26832 4218
rect 26896 4146 26924 22630
rect 27080 22574 27108 23258
rect 27264 23050 27292 23802
rect 27252 23044 27304 23050
rect 27252 22986 27304 22992
rect 27160 22976 27212 22982
rect 27160 22918 27212 22924
rect 27068 22568 27120 22574
rect 27068 22510 27120 22516
rect 27172 22409 27200 22918
rect 27264 22778 27292 22986
rect 27252 22772 27304 22778
rect 27252 22714 27304 22720
rect 27264 22506 27292 22714
rect 27252 22500 27304 22506
rect 27252 22442 27304 22448
rect 27158 22400 27214 22409
rect 27158 22335 27214 22344
rect 27344 22092 27396 22098
rect 27344 22034 27396 22040
rect 27160 22024 27212 22030
rect 27160 21966 27212 21972
rect 27172 21350 27200 21966
rect 27356 21865 27384 22034
rect 27342 21856 27398 21865
rect 27342 21791 27398 21800
rect 27356 21690 27384 21791
rect 27344 21684 27396 21690
rect 27344 21626 27396 21632
rect 27160 21344 27212 21350
rect 27160 21286 27212 21292
rect 27172 20330 27200 21286
rect 27160 20324 27212 20330
rect 27160 20266 27212 20272
rect 27172 20210 27200 20266
rect 27080 20182 27200 20210
rect 27080 19718 27108 20182
rect 27436 19916 27488 19922
rect 27436 19858 27488 19864
rect 27068 19712 27120 19718
rect 27066 19680 27068 19689
rect 27120 19680 27122 19689
rect 27066 19615 27122 19624
rect 27448 19310 27476 19858
rect 27436 19304 27488 19310
rect 27436 19246 27488 19252
rect 26974 19000 27030 19009
rect 26974 18935 26976 18944
rect 27028 18935 27030 18944
rect 26976 18906 27028 18912
rect 27436 18896 27488 18902
rect 27436 18838 27488 18844
rect 26976 18828 27028 18834
rect 26976 18770 27028 18776
rect 26988 18086 27016 18770
rect 27448 18086 27476 18838
rect 26976 18080 27028 18086
rect 26976 18022 27028 18028
rect 27436 18080 27488 18086
rect 27436 18022 27488 18028
rect 26988 15706 27016 18022
rect 27434 17640 27490 17649
rect 27434 17575 27490 17584
rect 27068 17536 27120 17542
rect 27068 17478 27120 17484
rect 27080 17066 27108 17478
rect 27448 17338 27476 17575
rect 27436 17332 27488 17338
rect 27436 17274 27488 17280
rect 27068 17060 27120 17066
rect 27068 17002 27120 17008
rect 27252 16720 27304 16726
rect 27250 16688 27252 16697
rect 27304 16688 27306 16697
rect 27250 16623 27306 16632
rect 27066 16416 27122 16425
rect 27066 16351 27122 16360
rect 26976 15700 27028 15706
rect 26976 15642 27028 15648
rect 27080 15314 27108 16351
rect 27344 15496 27396 15502
rect 27344 15438 27396 15444
rect 26988 15286 27108 15314
rect 26988 12986 27016 15286
rect 27068 15156 27120 15162
rect 27068 15098 27120 15104
rect 26976 12980 27028 12986
rect 26976 12922 27028 12928
rect 26976 12300 27028 12306
rect 26976 12242 27028 12248
rect 26988 11082 27016 12242
rect 26976 11076 27028 11082
rect 26976 11018 27028 11024
rect 26976 10600 27028 10606
rect 26976 10542 27028 10548
rect 26988 5545 27016 10542
rect 27080 10266 27108 15098
rect 27356 14618 27384 15438
rect 27436 15360 27488 15366
rect 27436 15302 27488 15308
rect 27448 14958 27476 15302
rect 27436 14952 27488 14958
rect 27436 14894 27488 14900
rect 27344 14612 27396 14618
rect 27344 14554 27396 14560
rect 27436 13864 27488 13870
rect 27436 13806 27488 13812
rect 27252 13320 27304 13326
rect 27252 13262 27304 13268
rect 27264 12238 27292 13262
rect 27344 12708 27396 12714
rect 27344 12650 27396 12656
rect 27252 12232 27304 12238
rect 27252 12174 27304 12180
rect 27264 11898 27292 12174
rect 27356 12102 27384 12650
rect 27448 12442 27476 13806
rect 27436 12436 27488 12442
rect 27436 12378 27488 12384
rect 27344 12096 27396 12102
rect 27344 12038 27396 12044
rect 27252 11892 27304 11898
rect 27252 11834 27304 11840
rect 27356 11150 27384 12038
rect 27344 11144 27396 11150
rect 27344 11086 27396 11092
rect 27344 10464 27396 10470
rect 27344 10406 27396 10412
rect 27068 10260 27120 10266
rect 27068 10202 27120 10208
rect 27356 9926 27384 10406
rect 27344 9920 27396 9926
rect 27344 9862 27396 9868
rect 27356 9625 27384 9862
rect 27342 9616 27398 9625
rect 27264 9574 27342 9602
rect 27160 6860 27212 6866
rect 27160 6802 27212 6808
rect 27172 6746 27200 6802
rect 27264 6798 27292 9574
rect 27342 9551 27398 9560
rect 27080 6718 27200 6746
rect 27252 6792 27304 6798
rect 27252 6734 27304 6740
rect 27080 6118 27108 6718
rect 27264 6458 27292 6734
rect 27252 6452 27304 6458
rect 27252 6394 27304 6400
rect 27068 6112 27120 6118
rect 27066 6080 27068 6089
rect 27120 6080 27122 6089
rect 27066 6015 27122 6024
rect 26974 5536 27030 5545
rect 26974 5471 27030 5480
rect 27540 5012 27568 30058
rect 27724 29753 27752 30126
rect 27816 29850 27844 30670
rect 27896 30320 27948 30326
rect 27896 30262 27948 30268
rect 27908 30190 27936 30262
rect 27896 30184 27948 30190
rect 27896 30126 27948 30132
rect 27804 29844 27856 29850
rect 27804 29786 27856 29792
rect 27710 29744 27766 29753
rect 27710 29679 27766 29688
rect 27804 29164 27856 29170
rect 27804 29106 27856 29112
rect 27620 28144 27672 28150
rect 27620 28086 27672 28092
rect 27632 26994 27660 28086
rect 27712 28008 27764 28014
rect 27712 27950 27764 27956
rect 27724 27674 27752 27950
rect 27712 27668 27764 27674
rect 27712 27610 27764 27616
rect 27620 26988 27672 26994
rect 27620 26930 27672 26936
rect 27632 26489 27660 26930
rect 27618 26480 27674 26489
rect 27618 26415 27674 26424
rect 27816 26042 27844 29106
rect 27908 27402 27936 30126
rect 28000 29646 28028 31855
rect 28264 31826 28316 31832
rect 28172 31136 28224 31142
rect 28172 31078 28224 31084
rect 28184 30394 28212 31078
rect 28276 30410 28304 31826
rect 28538 31784 28594 31793
rect 28538 31719 28594 31728
rect 28552 30938 28580 31719
rect 28540 30932 28592 30938
rect 28540 30874 28592 30880
rect 28172 30388 28224 30394
rect 28276 30382 28396 30410
rect 28172 30330 28224 30336
rect 27988 29640 28040 29646
rect 27988 29582 28040 29588
rect 28000 29306 28028 29582
rect 27988 29300 28040 29306
rect 27988 29242 28040 29248
rect 28184 29238 28212 30330
rect 28368 30326 28396 30382
rect 28356 30320 28408 30326
rect 28356 30262 28408 30268
rect 28264 30252 28316 30258
rect 28264 30194 28316 30200
rect 28276 29850 28304 30194
rect 28264 29844 28316 29850
rect 28264 29786 28316 29792
rect 28262 29744 28318 29753
rect 28262 29679 28264 29688
rect 28316 29679 28318 29688
rect 28264 29650 28316 29656
rect 28172 29232 28224 29238
rect 28172 29174 28224 29180
rect 28184 28626 28212 29174
rect 28276 28762 28304 29650
rect 28264 28756 28316 28762
rect 28644 28744 28672 32558
rect 28724 32360 28776 32366
rect 28724 32302 28776 32308
rect 28736 31958 28764 32302
rect 28724 31952 28776 31958
rect 28724 31894 28776 31900
rect 28736 31482 28764 31894
rect 28816 31884 28868 31890
rect 28816 31826 28868 31832
rect 28724 31476 28776 31482
rect 28724 31418 28776 31424
rect 28264 28698 28316 28704
rect 28552 28716 28672 28744
rect 28172 28620 28224 28626
rect 28172 28562 28224 28568
rect 28184 28218 28212 28562
rect 28172 28212 28224 28218
rect 28172 28154 28224 28160
rect 28264 28212 28316 28218
rect 28264 28154 28316 28160
rect 27986 28112 28042 28121
rect 27986 28047 28042 28056
rect 28000 27538 28028 28047
rect 28184 28014 28212 28154
rect 28172 28008 28224 28014
rect 28172 27950 28224 27956
rect 28276 27674 28304 28154
rect 28264 27668 28316 27674
rect 28264 27610 28316 27616
rect 27988 27532 28040 27538
rect 27988 27474 28040 27480
rect 27896 27396 27948 27402
rect 27896 27338 27948 27344
rect 27908 27130 27936 27338
rect 27896 27124 27948 27130
rect 27896 27066 27948 27072
rect 27908 26450 27936 27066
rect 28000 26586 28028 27474
rect 28080 27464 28132 27470
rect 28080 27406 28132 27412
rect 27988 26580 28040 26586
rect 27988 26522 28040 26528
rect 27896 26444 27948 26450
rect 27896 26386 27948 26392
rect 27988 26240 28040 26246
rect 27988 26182 28040 26188
rect 27804 26036 27856 26042
rect 27804 25978 27856 25984
rect 27620 25288 27672 25294
rect 27620 25230 27672 25236
rect 27632 24750 27660 25230
rect 27712 24880 27764 24886
rect 27712 24822 27764 24828
rect 27620 24744 27672 24750
rect 27620 24686 27672 24692
rect 27632 24614 27660 24686
rect 27620 24608 27672 24614
rect 27620 24550 27672 24556
rect 27632 24070 27660 24550
rect 27724 24206 27752 24822
rect 27712 24200 27764 24206
rect 27712 24142 27764 24148
rect 27620 24064 27672 24070
rect 27620 24006 27672 24012
rect 27632 23662 27660 24006
rect 27896 23792 27948 23798
rect 27896 23734 27948 23740
rect 27620 23656 27672 23662
rect 27620 23598 27672 23604
rect 27632 23322 27660 23598
rect 27908 23322 27936 23734
rect 27620 23316 27672 23322
rect 27620 23258 27672 23264
rect 27896 23316 27948 23322
rect 27896 23258 27948 23264
rect 27620 21956 27672 21962
rect 27620 21898 27672 21904
rect 27632 21350 27660 21898
rect 27620 21344 27672 21350
rect 27620 21286 27672 21292
rect 27632 20874 27660 21286
rect 27620 20868 27672 20874
rect 27620 20810 27672 20816
rect 27632 20398 27660 20810
rect 27804 20800 27856 20806
rect 27804 20742 27856 20748
rect 27620 20392 27672 20398
rect 27620 20334 27672 20340
rect 27632 20058 27660 20334
rect 27620 20052 27672 20058
rect 27620 19994 27672 20000
rect 27712 18964 27764 18970
rect 27712 18906 27764 18912
rect 27620 18624 27672 18630
rect 27620 18566 27672 18572
rect 27632 18222 27660 18566
rect 27620 18216 27672 18222
rect 27620 18158 27672 18164
rect 27632 17746 27660 18158
rect 27724 17785 27752 18906
rect 27816 18902 27844 20742
rect 27894 20496 27950 20505
rect 27894 20431 27950 20440
rect 27908 20398 27936 20431
rect 27896 20392 27948 20398
rect 27896 20334 27948 20340
rect 27804 18896 27856 18902
rect 27804 18838 27856 18844
rect 27802 18456 27858 18465
rect 27802 18391 27858 18400
rect 27816 18154 27844 18391
rect 27804 18148 27856 18154
rect 27804 18090 27856 18096
rect 27710 17776 27766 17785
rect 27620 17740 27672 17746
rect 27710 17711 27766 17720
rect 27620 17682 27672 17688
rect 27632 17066 27660 17682
rect 27712 17536 27764 17542
rect 27712 17478 27764 17484
rect 27724 17066 27752 17478
rect 27620 17060 27672 17066
rect 27620 17002 27672 17008
rect 27712 17060 27764 17066
rect 27712 17002 27764 17008
rect 27632 15502 27660 17002
rect 27816 16250 27844 18090
rect 27896 18080 27948 18086
rect 27896 18022 27948 18028
rect 27908 17678 27936 18022
rect 27896 17672 27948 17678
rect 27896 17614 27948 17620
rect 27908 17134 27936 17614
rect 27896 17128 27948 17134
rect 27896 17070 27948 17076
rect 27908 16794 27936 17070
rect 27896 16788 27948 16794
rect 27896 16730 27948 16736
rect 27804 16244 27856 16250
rect 27804 16186 27856 16192
rect 27896 15972 27948 15978
rect 27896 15914 27948 15920
rect 27908 15706 27936 15914
rect 27896 15700 27948 15706
rect 27896 15642 27948 15648
rect 27802 15600 27858 15609
rect 27802 15535 27858 15544
rect 27620 15496 27672 15502
rect 27620 15438 27672 15444
rect 27710 15192 27766 15201
rect 27710 15127 27766 15136
rect 27724 15094 27752 15127
rect 27712 15088 27764 15094
rect 27712 15030 27764 15036
rect 27816 14074 27844 15535
rect 27896 15428 27948 15434
rect 27896 15370 27948 15376
rect 27908 14618 27936 15370
rect 27896 14612 27948 14618
rect 27896 14554 27948 14560
rect 27804 14068 27856 14074
rect 27804 14010 27856 14016
rect 27896 13796 27948 13802
rect 27896 13738 27948 13744
rect 27712 13524 27764 13530
rect 27712 13466 27764 13472
rect 27620 13252 27672 13258
rect 27620 13194 27672 13200
rect 27632 12850 27660 13194
rect 27620 12844 27672 12850
rect 27620 12786 27672 12792
rect 27724 12782 27752 13466
rect 27804 13388 27856 13394
rect 27804 13330 27856 13336
rect 27712 12776 27764 12782
rect 27712 12718 27764 12724
rect 27724 12170 27752 12718
rect 27816 12714 27844 13330
rect 27908 12986 27936 13738
rect 27896 12980 27948 12986
rect 27896 12922 27948 12928
rect 27804 12708 27856 12714
rect 27804 12650 27856 12656
rect 28000 12209 28028 26182
rect 28092 22273 28120 27406
rect 28354 26208 28410 26217
rect 28354 26143 28410 26152
rect 28264 25696 28316 25702
rect 28264 25638 28316 25644
rect 28276 25294 28304 25638
rect 28264 25288 28316 25294
rect 28264 25230 28316 25236
rect 28276 24818 28304 25230
rect 28264 24812 28316 24818
rect 28264 24754 28316 24760
rect 28264 24676 28316 24682
rect 28264 24618 28316 24624
rect 28276 24410 28304 24618
rect 28264 24404 28316 24410
rect 28264 24346 28316 24352
rect 28276 23322 28304 24346
rect 28264 23316 28316 23322
rect 28264 23258 28316 23264
rect 28078 22264 28134 22273
rect 28078 22199 28134 22208
rect 28264 21548 28316 21554
rect 28264 21490 28316 21496
rect 28078 20632 28134 20641
rect 28078 20567 28134 20576
rect 28092 20398 28120 20567
rect 28080 20392 28132 20398
rect 28080 20334 28132 20340
rect 28172 19304 28224 19310
rect 28172 19246 28224 19252
rect 28080 19168 28132 19174
rect 28080 19110 28132 19116
rect 28092 18329 28120 19110
rect 28184 18834 28212 19246
rect 28172 18828 28224 18834
rect 28172 18770 28224 18776
rect 28078 18320 28134 18329
rect 28184 18290 28212 18770
rect 28078 18255 28080 18264
rect 28132 18255 28134 18264
rect 28172 18284 28224 18290
rect 28080 18226 28132 18232
rect 28172 18226 28224 18232
rect 28080 17740 28132 17746
rect 28080 17682 28132 17688
rect 28092 16998 28120 17682
rect 28184 17610 28212 18226
rect 28276 17746 28304 21490
rect 28264 17740 28316 17746
rect 28264 17682 28316 17688
rect 28172 17604 28224 17610
rect 28172 17546 28224 17552
rect 28276 17338 28304 17682
rect 28264 17332 28316 17338
rect 28264 17274 28316 17280
rect 28080 16992 28132 16998
rect 28080 16934 28132 16940
rect 28092 16454 28120 16934
rect 28080 16448 28132 16454
rect 28080 16390 28132 16396
rect 28092 15910 28120 16390
rect 28080 15904 28132 15910
rect 28080 15846 28132 15852
rect 28092 14822 28120 15846
rect 28080 14816 28132 14822
rect 28080 14758 28132 14764
rect 27986 12200 28042 12209
rect 27712 12164 27764 12170
rect 27986 12135 28042 12144
rect 27712 12106 27764 12112
rect 27724 11898 27752 12106
rect 27712 11892 27764 11898
rect 27712 11834 27764 11840
rect 27804 11688 27856 11694
rect 27804 11630 27856 11636
rect 27816 11218 27844 11630
rect 27804 11212 27856 11218
rect 27804 11154 27856 11160
rect 27620 11144 27672 11150
rect 27620 11086 27672 11092
rect 27632 10130 27660 11086
rect 27712 11008 27764 11014
rect 27712 10950 27764 10956
rect 27724 10810 27752 10950
rect 27712 10804 27764 10810
rect 27712 10746 27764 10752
rect 28092 10266 28120 14758
rect 28276 14550 28304 17274
rect 28368 17252 28396 26143
rect 28552 25809 28580 28716
rect 28736 28626 28764 31418
rect 28828 31278 28856 31826
rect 28816 31272 28868 31278
rect 28816 31214 28868 31220
rect 28828 30870 28856 31214
rect 28816 30864 28868 30870
rect 28816 30806 28868 30812
rect 28816 30320 28868 30326
rect 28816 30262 28868 30268
rect 28632 28620 28684 28626
rect 28632 28562 28684 28568
rect 28724 28620 28776 28626
rect 28724 28562 28776 28568
rect 28644 27946 28672 28562
rect 28736 28218 28764 28562
rect 28724 28212 28776 28218
rect 28724 28154 28776 28160
rect 28828 28014 28856 30262
rect 28920 29306 28948 32694
rect 29012 32502 29040 32914
rect 29840 32910 29868 32943
rect 29828 32904 29880 32910
rect 29182 32872 29238 32881
rect 29828 32846 29880 32852
rect 29182 32807 29238 32816
rect 29000 32496 29052 32502
rect 29000 32438 29052 32444
rect 29196 31890 29224 32807
rect 29840 32570 29868 32846
rect 29552 32564 29604 32570
rect 29552 32506 29604 32512
rect 29828 32564 29880 32570
rect 29828 32506 29880 32512
rect 29564 32366 29592 32506
rect 29552 32360 29604 32366
rect 29552 32302 29604 32308
rect 29184 31884 29236 31890
rect 29184 31826 29236 31832
rect 29196 31793 29224 31826
rect 29182 31784 29238 31793
rect 29182 31719 29238 31728
rect 29276 30592 29328 30598
rect 29276 30534 29328 30540
rect 28998 30288 29054 30297
rect 29288 30258 29316 30534
rect 28998 30223 29054 30232
rect 29276 30252 29328 30258
rect 29012 30190 29040 30223
rect 29276 30194 29328 30200
rect 29000 30184 29052 30190
rect 29564 30161 29592 32302
rect 30024 32026 30052 33322
rect 30116 33300 30144 33390
rect 30194 33351 30250 33360
rect 30116 33272 30236 33300
rect 30104 32972 30156 32978
rect 30104 32914 30156 32920
rect 30116 32570 30144 32914
rect 30104 32564 30156 32570
rect 30104 32506 30156 32512
rect 30012 32020 30064 32026
rect 30012 31962 30064 31968
rect 30116 31958 30144 32506
rect 30104 31952 30156 31958
rect 30104 31894 30156 31900
rect 30208 31770 30236 33272
rect 30300 33046 30328 34002
rect 30392 33998 30420 34439
rect 30380 33992 30432 33998
rect 30380 33934 30432 33940
rect 30288 33040 30340 33046
rect 30288 32982 30340 32988
rect 30564 32904 30616 32910
rect 30564 32846 30616 32852
rect 29736 31748 29788 31754
rect 29736 31690 29788 31696
rect 30116 31742 30236 31770
rect 29748 31278 29776 31690
rect 30116 31668 30144 31742
rect 30116 31640 30236 31668
rect 30010 31376 30066 31385
rect 30010 31311 30012 31320
rect 30064 31311 30066 31320
rect 30012 31282 30064 31288
rect 29736 31272 29788 31278
rect 29736 31214 29788 31220
rect 29748 30938 29776 31214
rect 29736 30932 29788 30938
rect 29736 30874 29788 30880
rect 30010 30832 30066 30841
rect 30010 30767 30012 30776
rect 30064 30767 30066 30776
rect 30012 30738 30064 30744
rect 29736 30252 29788 30258
rect 29736 30194 29788 30200
rect 29000 30126 29052 30132
rect 29550 30152 29606 30161
rect 29368 30116 29420 30122
rect 29550 30087 29606 30096
rect 29368 30058 29420 30064
rect 29276 29640 29328 29646
rect 29276 29582 29328 29588
rect 28908 29300 28960 29306
rect 28908 29242 28960 29248
rect 29288 29170 29316 29582
rect 29276 29164 29328 29170
rect 29276 29106 29328 29112
rect 29184 29096 29236 29102
rect 29184 29038 29236 29044
rect 28908 28960 28960 28966
rect 28908 28902 28960 28908
rect 28816 28008 28868 28014
rect 28816 27950 28868 27956
rect 28632 27940 28684 27946
rect 28632 27882 28684 27888
rect 28644 27674 28672 27882
rect 28632 27668 28684 27674
rect 28632 27610 28684 27616
rect 28816 27532 28868 27538
rect 28816 27474 28868 27480
rect 28724 27056 28776 27062
rect 28722 27024 28724 27033
rect 28776 27024 28778 27033
rect 28722 26959 28778 26968
rect 28828 26518 28856 27474
rect 28816 26512 28868 26518
rect 28816 26454 28868 26460
rect 28538 25800 28594 25809
rect 28538 25735 28594 25744
rect 28724 25696 28776 25702
rect 28722 25664 28724 25673
rect 28776 25664 28778 25673
rect 28722 25599 28778 25608
rect 28446 24304 28502 24313
rect 28446 24239 28448 24248
rect 28500 24239 28502 24248
rect 28448 24210 28500 24216
rect 28460 23866 28488 24210
rect 28448 23860 28500 23866
rect 28448 23802 28500 23808
rect 28816 23588 28868 23594
rect 28816 23530 28868 23536
rect 28724 23248 28776 23254
rect 28724 23190 28776 23196
rect 28540 23112 28592 23118
rect 28540 23054 28592 23060
rect 28448 22568 28500 22574
rect 28448 22510 28500 22516
rect 28460 21010 28488 22510
rect 28552 21010 28580 23054
rect 28736 22710 28764 23190
rect 28724 22704 28776 22710
rect 28724 22646 28776 22652
rect 28828 22098 28856 23530
rect 28816 22092 28868 22098
rect 28816 22034 28868 22040
rect 28632 21888 28684 21894
rect 28632 21830 28684 21836
rect 28644 21554 28672 21830
rect 28828 21690 28856 22034
rect 28816 21684 28868 21690
rect 28816 21626 28868 21632
rect 28632 21548 28684 21554
rect 28632 21490 28684 21496
rect 28816 21072 28868 21078
rect 28816 21014 28868 21020
rect 28448 21004 28500 21010
rect 28448 20946 28500 20952
rect 28540 21004 28592 21010
rect 28540 20946 28592 20952
rect 28460 20602 28488 20946
rect 28724 20868 28776 20874
rect 28724 20810 28776 20816
rect 28448 20596 28500 20602
rect 28448 20538 28500 20544
rect 28736 19854 28764 20810
rect 28828 19922 28856 21014
rect 28816 19916 28868 19922
rect 28816 19858 28868 19864
rect 28724 19848 28776 19854
rect 28724 19790 28776 19796
rect 28736 19378 28764 19790
rect 28724 19372 28776 19378
rect 28724 19314 28776 19320
rect 28632 19168 28684 19174
rect 28632 19110 28684 19116
rect 28644 18222 28672 19110
rect 28736 18834 28764 19314
rect 28724 18828 28776 18834
rect 28724 18770 28776 18776
rect 28736 18426 28764 18770
rect 28724 18420 28776 18426
rect 28724 18362 28776 18368
rect 28632 18216 28684 18222
rect 28632 18158 28684 18164
rect 28368 17224 28764 17252
rect 28540 17060 28592 17066
rect 28540 17002 28592 17008
rect 28552 16794 28580 17002
rect 28540 16788 28592 16794
rect 28540 16730 28592 16736
rect 28552 16454 28580 16730
rect 28540 16448 28592 16454
rect 28540 16390 28592 16396
rect 28552 15910 28580 16390
rect 28540 15904 28592 15910
rect 28540 15846 28592 15852
rect 28448 15700 28500 15706
rect 28448 15642 28500 15648
rect 28356 15564 28408 15570
rect 28356 15506 28408 15512
rect 28264 14544 28316 14550
rect 28264 14486 28316 14492
rect 28276 14074 28304 14486
rect 28264 14068 28316 14074
rect 28264 14010 28316 14016
rect 28276 13462 28304 14010
rect 28368 13716 28396 15506
rect 28460 15434 28488 15642
rect 28552 15620 28580 15846
rect 28632 15632 28684 15638
rect 28552 15592 28632 15620
rect 28632 15574 28684 15580
rect 28448 15428 28500 15434
rect 28448 15370 28500 15376
rect 28460 15162 28488 15370
rect 28644 15162 28672 15574
rect 28448 15156 28500 15162
rect 28448 15098 28500 15104
rect 28632 15156 28684 15162
rect 28632 15098 28684 15104
rect 28448 14272 28500 14278
rect 28448 14214 28500 14220
rect 28460 13870 28488 14214
rect 28448 13864 28500 13870
rect 28448 13806 28500 13812
rect 28368 13688 28488 13716
rect 28264 13456 28316 13462
rect 28264 13398 28316 13404
rect 28276 12850 28304 13398
rect 28356 13388 28408 13394
rect 28356 13330 28408 13336
rect 28264 12844 28316 12850
rect 28264 12786 28316 12792
rect 28264 12640 28316 12646
rect 28264 12582 28316 12588
rect 28276 11898 28304 12582
rect 28368 12442 28396 13330
rect 28460 12646 28488 13688
rect 28632 12980 28684 12986
rect 28632 12922 28684 12928
rect 28448 12640 28500 12646
rect 28448 12582 28500 12588
rect 28356 12436 28408 12442
rect 28356 12378 28408 12384
rect 28644 12306 28672 12922
rect 28632 12300 28684 12306
rect 28632 12242 28684 12248
rect 28644 11898 28672 12242
rect 28264 11892 28316 11898
rect 28264 11834 28316 11840
rect 28632 11892 28684 11898
rect 28632 11834 28684 11840
rect 28736 11665 28764 17224
rect 28828 16454 28856 19858
rect 28816 16448 28868 16454
rect 28816 16390 28868 16396
rect 28816 16244 28868 16250
rect 28816 16186 28868 16192
rect 28828 13802 28856 16186
rect 28816 13796 28868 13802
rect 28816 13738 28868 13744
rect 28816 13184 28868 13190
rect 28816 13126 28868 13132
rect 28828 12442 28856 13126
rect 28816 12436 28868 12442
rect 28816 12378 28868 12384
rect 28722 11656 28778 11665
rect 28722 11591 28778 11600
rect 28538 11384 28594 11393
rect 28538 11319 28594 11328
rect 28552 11218 28580 11319
rect 28540 11212 28592 11218
rect 28540 11154 28592 11160
rect 28552 10810 28580 11154
rect 28540 10804 28592 10810
rect 28540 10746 28592 10752
rect 28080 10260 28132 10266
rect 28080 10202 28132 10208
rect 27620 10124 27672 10130
rect 27620 10066 27672 10072
rect 27632 9722 27660 10066
rect 27620 9716 27672 9722
rect 27620 9658 27672 9664
rect 28722 6896 28778 6905
rect 28722 6831 28724 6840
rect 28776 6831 28778 6840
rect 28724 6802 28776 6808
rect 28078 5944 28134 5953
rect 28078 5879 28134 5888
rect 27172 4984 27568 5012
rect 26884 4140 26936 4146
rect 26884 4082 26936 4088
rect 26516 3392 26568 3398
rect 26516 3334 26568 3340
rect 26424 3188 26476 3194
rect 26424 3130 26476 3136
rect 27172 800 27200 4984
rect 27344 3392 27396 3398
rect 27344 3334 27396 3340
rect 27356 2825 27384 3334
rect 27526 3224 27582 3233
rect 27526 3159 27582 3168
rect 27540 2854 27568 3159
rect 27528 2848 27580 2854
rect 27342 2816 27398 2825
rect 27528 2790 27580 2796
rect 27342 2751 27398 2760
rect 27356 2446 27384 2751
rect 27344 2440 27396 2446
rect 27344 2382 27396 2388
rect 27528 2440 27580 2446
rect 27580 2400 27660 2428
rect 27528 2382 27580 2388
rect 27632 800 27660 2400
rect 28092 800 28120 5879
rect 28920 4758 28948 28902
rect 29000 27668 29052 27674
rect 29000 27610 29052 27616
rect 29012 27538 29040 27610
rect 29000 27532 29052 27538
rect 29000 27474 29052 27480
rect 29090 27432 29146 27441
rect 29090 27367 29146 27376
rect 29104 26518 29132 27367
rect 29092 26512 29144 26518
rect 29092 26454 29144 26460
rect 29090 26344 29146 26353
rect 29090 26279 29092 26288
rect 29144 26279 29146 26288
rect 29092 26250 29144 26256
rect 29104 25838 29132 26250
rect 29196 25974 29224 29038
rect 29274 28928 29330 28937
rect 29274 28863 29330 28872
rect 29184 25968 29236 25974
rect 29184 25910 29236 25916
rect 29092 25832 29144 25838
rect 29288 25786 29316 28863
rect 29380 27674 29408 30058
rect 29460 29504 29512 29510
rect 29460 29446 29512 29452
rect 29472 29170 29500 29446
rect 29460 29164 29512 29170
rect 29460 29106 29512 29112
rect 29368 27668 29420 27674
rect 29368 27610 29420 27616
rect 29368 27532 29420 27538
rect 29368 27474 29420 27480
rect 29380 25945 29408 27474
rect 29564 27130 29592 30087
rect 29748 30025 29776 30194
rect 30024 30190 30052 30738
rect 30012 30184 30064 30190
rect 30012 30126 30064 30132
rect 29734 30016 29790 30025
rect 29734 29951 29790 29960
rect 29748 29850 29776 29951
rect 29736 29844 29788 29850
rect 29788 29804 29868 29832
rect 29736 29786 29788 29792
rect 29736 29708 29788 29714
rect 29736 29650 29788 29656
rect 29644 28008 29696 28014
rect 29644 27950 29696 27956
rect 29656 27674 29684 27950
rect 29644 27668 29696 27674
rect 29644 27610 29696 27616
rect 29748 27334 29776 29650
rect 29840 29617 29868 29804
rect 29920 29640 29972 29646
rect 29826 29608 29882 29617
rect 29920 29582 29972 29588
rect 29826 29543 29882 29552
rect 29932 29238 29960 29582
rect 29920 29232 29972 29238
rect 29920 29174 29972 29180
rect 30104 29096 30156 29102
rect 30104 29038 30156 29044
rect 30116 27946 30144 29038
rect 30104 27940 30156 27946
rect 30104 27882 30156 27888
rect 29736 27328 29788 27334
rect 29736 27270 29788 27276
rect 29828 27328 29880 27334
rect 29828 27270 29880 27276
rect 29552 27124 29604 27130
rect 29552 27066 29604 27072
rect 29552 26444 29604 26450
rect 29552 26386 29604 26392
rect 29564 26042 29592 26386
rect 29552 26036 29604 26042
rect 29552 25978 29604 25984
rect 29366 25936 29422 25945
rect 29366 25871 29422 25880
rect 29092 25774 29144 25780
rect 29196 25758 29316 25786
rect 29368 25832 29420 25838
rect 29368 25774 29420 25780
rect 29196 24342 29224 25758
rect 29276 25356 29328 25362
rect 29276 25298 29328 25304
rect 29288 24954 29316 25298
rect 29276 24948 29328 24954
rect 29276 24890 29328 24896
rect 29380 24750 29408 25774
rect 29564 25498 29592 25978
rect 29748 25922 29776 27270
rect 29840 26450 29868 27270
rect 29828 26444 29880 26450
rect 29828 26386 29880 26392
rect 30012 26444 30064 26450
rect 30012 26386 30064 26392
rect 29840 26042 29868 26386
rect 29828 26036 29880 26042
rect 29828 25978 29880 25984
rect 30024 25974 30052 26386
rect 30012 25968 30064 25974
rect 29644 25900 29696 25906
rect 29748 25894 29868 25922
rect 30012 25910 30064 25916
rect 30208 25906 30236 31640
rect 30576 31346 30604 32846
rect 30564 31340 30616 31346
rect 30564 31282 30616 31288
rect 30470 29744 30526 29753
rect 30470 29679 30472 29688
rect 30524 29679 30526 29688
rect 30472 29650 30524 29656
rect 30380 29164 30432 29170
rect 30380 29106 30432 29112
rect 30392 28762 30420 29106
rect 30380 28756 30432 28762
rect 30380 28698 30432 28704
rect 30564 28688 30616 28694
rect 30564 28630 30616 28636
rect 30288 28620 30340 28626
rect 30288 28562 30340 28568
rect 30300 28150 30328 28562
rect 30288 28144 30340 28150
rect 30576 28121 30604 28630
rect 30288 28086 30340 28092
rect 30562 28112 30618 28121
rect 30562 28047 30618 28056
rect 30472 28008 30524 28014
rect 30472 27950 30524 27956
rect 30564 28008 30616 28014
rect 30564 27950 30616 27956
rect 30484 27334 30512 27950
rect 30472 27328 30524 27334
rect 30472 27270 30524 27276
rect 30472 27056 30524 27062
rect 30472 26998 30524 27004
rect 30484 26450 30512 26998
rect 30472 26444 30524 26450
rect 30472 26386 30524 26392
rect 29644 25842 29696 25848
rect 29656 25786 29684 25842
rect 29656 25758 29776 25786
rect 29552 25492 29604 25498
rect 29552 25434 29604 25440
rect 29460 25356 29512 25362
rect 29460 25298 29512 25304
rect 29472 24750 29500 25298
rect 29368 24744 29420 24750
rect 29368 24686 29420 24692
rect 29460 24744 29512 24750
rect 29460 24686 29512 24692
rect 29184 24336 29236 24342
rect 29184 24278 29236 24284
rect 29184 24200 29236 24206
rect 29184 24142 29236 24148
rect 29092 23724 29144 23730
rect 29092 23666 29144 23672
rect 29104 22574 29132 23666
rect 29196 22574 29224 24142
rect 29276 24132 29328 24138
rect 29276 24074 29328 24080
rect 29288 23186 29316 24074
rect 29368 24064 29420 24070
rect 29368 24006 29420 24012
rect 29380 23322 29408 24006
rect 29472 23866 29500 24686
rect 29644 24336 29696 24342
rect 29644 24278 29696 24284
rect 29552 24064 29604 24070
rect 29552 24006 29604 24012
rect 29460 23860 29512 23866
rect 29460 23802 29512 23808
rect 29368 23316 29420 23322
rect 29368 23258 29420 23264
rect 29472 23186 29500 23802
rect 29564 23662 29592 24006
rect 29552 23656 29604 23662
rect 29552 23598 29604 23604
rect 29276 23180 29328 23186
rect 29276 23122 29328 23128
rect 29460 23180 29512 23186
rect 29460 23122 29512 23128
rect 29288 22778 29316 23122
rect 29276 22772 29328 22778
rect 29276 22714 29328 22720
rect 29092 22568 29144 22574
rect 29092 22510 29144 22516
rect 29184 22568 29236 22574
rect 29184 22510 29236 22516
rect 29472 22506 29500 23122
rect 29552 22704 29604 22710
rect 29552 22646 29604 22652
rect 29460 22500 29512 22506
rect 29460 22442 29512 22448
rect 29460 22228 29512 22234
rect 29460 22170 29512 22176
rect 29472 21622 29500 22170
rect 29184 21616 29236 21622
rect 29184 21558 29236 21564
rect 29460 21616 29512 21622
rect 29460 21558 29512 21564
rect 29092 21004 29144 21010
rect 29092 20946 29144 20952
rect 29104 20330 29132 20946
rect 29092 20324 29144 20330
rect 29092 20266 29144 20272
rect 29104 20058 29132 20266
rect 29092 20052 29144 20058
rect 29092 19994 29144 20000
rect 29196 19242 29224 21558
rect 29564 21486 29592 22646
rect 29656 22001 29684 24278
rect 29642 21992 29698 22001
rect 29642 21927 29698 21936
rect 29644 21616 29696 21622
rect 29644 21558 29696 21564
rect 29552 21480 29604 21486
rect 29552 21422 29604 21428
rect 29552 21344 29604 21350
rect 29552 21286 29604 21292
rect 29368 20392 29420 20398
rect 29368 20334 29420 20340
rect 29380 19718 29408 20334
rect 29564 20233 29592 21286
rect 29550 20224 29606 20233
rect 29550 20159 29606 20168
rect 29368 19712 29420 19718
rect 29368 19654 29420 19660
rect 29276 19304 29328 19310
rect 29276 19246 29328 19252
rect 29184 19236 29236 19242
rect 29184 19178 29236 19184
rect 29288 19174 29316 19246
rect 29276 19168 29328 19174
rect 29276 19110 29328 19116
rect 29092 18760 29144 18766
rect 29092 18702 29144 18708
rect 28998 18048 29054 18057
rect 28998 17983 29054 17992
rect 29012 12356 29040 17983
rect 29104 17785 29132 18702
rect 29184 17876 29236 17882
rect 29184 17818 29236 17824
rect 29090 17776 29146 17785
rect 29090 17711 29146 17720
rect 29104 17202 29132 17711
rect 29092 17196 29144 17202
rect 29092 17138 29144 17144
rect 29092 15972 29144 15978
rect 29092 15914 29144 15920
rect 29104 15638 29132 15914
rect 29092 15632 29144 15638
rect 29092 15574 29144 15580
rect 29012 12328 29132 12356
rect 29000 11076 29052 11082
rect 29000 11018 29052 11024
rect 29012 10810 29040 11018
rect 29000 10804 29052 10810
rect 29000 10746 29052 10752
rect 28908 4752 28960 4758
rect 28908 4694 28960 4700
rect 29104 2106 29132 12328
rect 29196 2582 29224 17818
rect 29380 17814 29408 19654
rect 29564 18714 29592 20159
rect 29472 18686 29592 18714
rect 29368 17808 29420 17814
rect 29368 17750 29420 17756
rect 29368 17536 29420 17542
rect 29368 17478 29420 17484
rect 29380 17134 29408 17478
rect 29472 17218 29500 18686
rect 29656 18465 29684 21558
rect 29642 18456 29698 18465
rect 29642 18391 29698 18400
rect 29644 18080 29696 18086
rect 29644 18022 29696 18028
rect 29552 17740 29604 17746
rect 29552 17682 29604 17688
rect 29564 17649 29592 17682
rect 29550 17640 29606 17649
rect 29550 17575 29606 17584
rect 29564 17338 29592 17575
rect 29552 17332 29604 17338
rect 29552 17274 29604 17280
rect 29472 17190 29592 17218
rect 29368 17128 29420 17134
rect 29368 17070 29420 17076
rect 29276 17060 29328 17066
rect 29276 17002 29328 17008
rect 29288 16590 29316 17002
rect 29380 16658 29408 17070
rect 29460 16992 29512 16998
rect 29460 16934 29512 16940
rect 29472 16726 29500 16934
rect 29460 16720 29512 16726
rect 29460 16662 29512 16668
rect 29368 16652 29420 16658
rect 29368 16594 29420 16600
rect 29276 16584 29328 16590
rect 29276 16526 29328 16532
rect 29288 16250 29316 16526
rect 29276 16244 29328 16250
rect 29276 16186 29328 16192
rect 29288 15502 29316 16186
rect 29380 15638 29408 16594
rect 29368 15632 29420 15638
rect 29368 15574 29420 15580
rect 29472 15570 29500 16662
rect 29564 16561 29592 17190
rect 29550 16552 29606 16561
rect 29550 16487 29606 16496
rect 29460 15564 29512 15570
rect 29460 15506 29512 15512
rect 29276 15496 29328 15502
rect 29276 15438 29328 15444
rect 29288 15162 29316 15438
rect 29276 15156 29328 15162
rect 29276 15098 29328 15104
rect 29288 13870 29316 15098
rect 29460 14340 29512 14346
rect 29460 14282 29512 14288
rect 29472 13870 29500 14282
rect 29276 13864 29328 13870
rect 29276 13806 29328 13812
rect 29460 13864 29512 13870
rect 29460 13806 29512 13812
rect 29288 13530 29316 13806
rect 29656 13682 29684 18022
rect 29748 17882 29776 25758
rect 29840 22234 29868 25894
rect 30196 25900 30248 25906
rect 30196 25842 30248 25848
rect 30196 25764 30248 25770
rect 30196 25706 30248 25712
rect 30208 25498 30236 25706
rect 30484 25673 30512 26386
rect 30470 25664 30526 25673
rect 30470 25599 30526 25608
rect 30196 25492 30248 25498
rect 30196 25434 30248 25440
rect 30484 25344 30512 25599
rect 30576 25498 30604 27950
rect 30564 25492 30616 25498
rect 30564 25434 30616 25440
rect 30564 25356 30616 25362
rect 30484 25316 30564 25344
rect 30564 25298 30616 25304
rect 30472 25220 30524 25226
rect 30472 25162 30524 25168
rect 30012 24676 30064 24682
rect 30012 24618 30064 24624
rect 29920 24608 29972 24614
rect 29920 24550 29972 24556
rect 29828 22228 29880 22234
rect 29828 22170 29880 22176
rect 29932 21622 29960 24550
rect 30024 24274 30052 24618
rect 30484 24614 30512 25162
rect 30472 24608 30524 24614
rect 30472 24550 30524 24556
rect 30012 24268 30064 24274
rect 30012 24210 30064 24216
rect 30024 23866 30052 24210
rect 30576 24070 30604 25298
rect 30564 24064 30616 24070
rect 30564 24006 30616 24012
rect 30012 23860 30064 23866
rect 30012 23802 30064 23808
rect 30194 23216 30250 23225
rect 30194 23151 30250 23160
rect 29920 21616 29972 21622
rect 29920 21558 29972 21564
rect 29920 21480 29972 21486
rect 29920 21422 29972 21428
rect 29828 21344 29880 21350
rect 29828 21286 29880 21292
rect 29840 21010 29868 21286
rect 29828 21004 29880 21010
rect 29828 20946 29880 20952
rect 29828 20528 29880 20534
rect 29828 20470 29880 20476
rect 29736 17876 29788 17882
rect 29736 17818 29788 17824
rect 29736 17672 29788 17678
rect 29736 17614 29788 17620
rect 29748 17066 29776 17614
rect 29736 17060 29788 17066
rect 29736 17002 29788 17008
rect 29748 16794 29776 17002
rect 29840 16794 29868 20470
rect 29932 18426 29960 21422
rect 30208 20913 30236 23151
rect 30288 22976 30340 22982
rect 30288 22918 30340 22924
rect 30300 22642 30328 22918
rect 30288 22636 30340 22642
rect 30288 22578 30340 22584
rect 30378 22400 30434 22409
rect 30378 22335 30434 22344
rect 30288 22024 30340 22030
rect 30288 21966 30340 21972
rect 30300 21622 30328 21966
rect 30288 21616 30340 21622
rect 30288 21558 30340 21564
rect 30392 21486 30420 22335
rect 30472 22092 30524 22098
rect 30472 22034 30524 22040
rect 30484 21865 30512 22034
rect 30668 22030 30696 34462
rect 30748 32904 30800 32910
rect 30748 32846 30800 32852
rect 30760 32298 30788 32846
rect 30748 32292 30800 32298
rect 30748 32234 30800 32240
rect 30932 31680 30984 31686
rect 30932 31622 30984 31628
rect 30944 31482 30972 31622
rect 30932 31476 30984 31482
rect 30932 31418 30984 31424
rect 30932 31340 30984 31346
rect 30932 31282 30984 31288
rect 30748 31204 30800 31210
rect 30748 31146 30800 31152
rect 30760 30802 30788 31146
rect 30748 30796 30800 30802
rect 30748 30738 30800 30744
rect 30760 30054 30788 30738
rect 30748 30048 30800 30054
rect 30748 29990 30800 29996
rect 30760 28150 30788 29990
rect 30840 28416 30892 28422
rect 30840 28358 30892 28364
rect 30748 28144 30800 28150
rect 30748 28086 30800 28092
rect 30852 28014 30880 28358
rect 30840 28008 30892 28014
rect 30840 27950 30892 27956
rect 30852 27334 30880 27365
rect 30840 27328 30892 27334
rect 30838 27296 30840 27305
rect 30892 27296 30894 27305
rect 30838 27231 30894 27240
rect 30852 26994 30880 27231
rect 30840 26988 30892 26994
rect 30840 26930 30892 26936
rect 30748 26920 30800 26926
rect 30748 26862 30800 26868
rect 30760 26042 30788 26862
rect 30840 26852 30892 26858
rect 30840 26794 30892 26800
rect 30852 26246 30880 26794
rect 30840 26240 30892 26246
rect 30840 26182 30892 26188
rect 30748 26036 30800 26042
rect 30748 25978 30800 25984
rect 30852 25922 30880 26182
rect 30760 25894 30880 25922
rect 30656 22024 30708 22030
rect 30656 21966 30708 21972
rect 30470 21856 30526 21865
rect 30470 21791 30526 21800
rect 30380 21480 30432 21486
rect 30380 21422 30432 21428
rect 30484 21146 30512 21791
rect 30472 21140 30524 21146
rect 30472 21082 30524 21088
rect 30656 21004 30708 21010
rect 30656 20946 30708 20952
rect 30194 20904 30250 20913
rect 30194 20839 30250 20848
rect 30472 20800 30524 20806
rect 30472 20742 30524 20748
rect 30484 20641 30512 20742
rect 30470 20632 30526 20641
rect 30668 20602 30696 20946
rect 30470 20567 30526 20576
rect 30656 20596 30708 20602
rect 30656 20538 30708 20544
rect 30012 19916 30064 19922
rect 30012 19858 30064 19864
rect 30104 19916 30156 19922
rect 30104 19858 30156 19864
rect 30024 19378 30052 19858
rect 30012 19372 30064 19378
rect 30012 19314 30064 19320
rect 29920 18420 29972 18426
rect 29920 18362 29972 18368
rect 29932 18222 29960 18362
rect 29920 18216 29972 18222
rect 29920 18158 29972 18164
rect 29920 17536 29972 17542
rect 29918 17504 29920 17513
rect 29972 17504 29974 17513
rect 29918 17439 29974 17448
rect 30024 17202 30052 19314
rect 30116 19242 30144 19858
rect 30196 19848 30248 19854
rect 30196 19790 30248 19796
rect 30104 19236 30156 19242
rect 30104 19178 30156 19184
rect 30116 18970 30144 19178
rect 30208 18970 30236 19790
rect 30288 19780 30340 19786
rect 30288 19722 30340 19728
rect 30300 19281 30328 19722
rect 30286 19272 30342 19281
rect 30286 19207 30342 19216
rect 30288 19168 30340 19174
rect 30288 19110 30340 19116
rect 30104 18964 30156 18970
rect 30104 18906 30156 18912
rect 30196 18964 30248 18970
rect 30196 18906 30248 18912
rect 30300 18630 30328 19110
rect 30288 18624 30340 18630
rect 30288 18566 30340 18572
rect 30656 18624 30708 18630
rect 30656 18566 30708 18572
rect 30012 17196 30064 17202
rect 30012 17138 30064 17144
rect 29736 16788 29788 16794
rect 29736 16730 29788 16736
rect 29828 16788 29880 16794
rect 29828 16730 29880 16736
rect 29840 16046 29868 16730
rect 30300 16726 30328 18566
rect 30472 18420 30524 18426
rect 30472 18362 30524 18368
rect 30380 17808 30432 17814
rect 30378 17776 30380 17785
rect 30432 17776 30434 17785
rect 30484 17746 30512 18362
rect 30668 18329 30696 18566
rect 30654 18320 30710 18329
rect 30654 18255 30710 18264
rect 30378 17711 30434 17720
rect 30472 17740 30524 17746
rect 30472 17682 30524 17688
rect 30484 17338 30512 17682
rect 30472 17332 30524 17338
rect 30472 17274 30524 17280
rect 30760 16776 30788 25894
rect 30944 24410 30972 31282
rect 31036 26586 31064 38150
rect 31206 36952 31262 36961
rect 31206 36887 31262 36896
rect 31220 36258 31248 36887
rect 31312 36360 31340 40996
rect 31484 38548 31536 38554
rect 31484 38490 31536 38496
rect 31496 38457 31524 38490
rect 31482 38448 31538 38457
rect 31772 38418 31800 40996
rect 31482 38383 31538 38392
rect 31760 38412 31812 38418
rect 31760 38354 31812 38360
rect 31390 38040 31446 38049
rect 31772 38010 31800 38354
rect 32128 38344 32180 38350
rect 32128 38286 32180 38292
rect 32402 38312 32458 38321
rect 31390 37975 31392 37984
rect 31444 37975 31446 37984
rect 31760 38004 31812 38010
rect 31392 37946 31444 37952
rect 31760 37946 31812 37952
rect 31852 37664 31904 37670
rect 31852 37606 31904 37612
rect 31312 36332 31616 36360
rect 31220 36230 31340 36258
rect 31208 32904 31260 32910
rect 31208 32846 31260 32852
rect 31220 32026 31248 32846
rect 31208 32020 31260 32026
rect 31208 31962 31260 31968
rect 31208 29504 31260 29510
rect 31208 29446 31260 29452
rect 31220 29102 31248 29446
rect 31312 29170 31340 36230
rect 31392 32224 31444 32230
rect 31392 32166 31444 32172
rect 31300 29164 31352 29170
rect 31300 29106 31352 29112
rect 31208 29096 31260 29102
rect 31208 29038 31260 29044
rect 31208 28756 31260 28762
rect 31208 28698 31260 28704
rect 31220 28422 31248 28698
rect 31208 28416 31260 28422
rect 31208 28358 31260 28364
rect 31116 28008 31168 28014
rect 31116 27950 31168 27956
rect 31128 27538 31156 27950
rect 31116 27532 31168 27538
rect 31116 27474 31168 27480
rect 31128 26926 31156 27474
rect 31208 27328 31260 27334
rect 31208 27270 31260 27276
rect 31116 26920 31168 26926
rect 31116 26862 31168 26868
rect 31024 26580 31076 26586
rect 31024 26522 31076 26528
rect 31220 26489 31248 27270
rect 31206 26480 31262 26489
rect 31206 26415 31208 26424
rect 31260 26415 31262 26424
rect 31208 26386 31260 26392
rect 31116 25152 31168 25158
rect 31116 25094 31168 25100
rect 30932 24404 30984 24410
rect 30932 24346 30984 24352
rect 31024 24268 31076 24274
rect 31024 24210 31076 24216
rect 30840 24064 30892 24070
rect 30840 24006 30892 24012
rect 30852 22506 30880 24006
rect 30932 23724 30984 23730
rect 31036 23712 31064 24210
rect 31128 23730 31156 25094
rect 31404 24818 31432 32166
rect 31484 31272 31536 31278
rect 31484 31214 31536 31220
rect 31496 30802 31524 31214
rect 31484 30796 31536 30802
rect 31484 30738 31536 30744
rect 31588 25242 31616 36332
rect 31668 31136 31720 31142
rect 31668 31078 31720 31084
rect 31680 29866 31708 31078
rect 31680 29850 31800 29866
rect 31680 29844 31812 29850
rect 31680 29838 31760 29844
rect 31760 29786 31812 29792
rect 31760 29096 31812 29102
rect 31760 29038 31812 29044
rect 31668 28484 31720 28490
rect 31668 28426 31720 28432
rect 31680 28218 31708 28426
rect 31772 28218 31800 29038
rect 31864 28694 31892 37606
rect 32140 37398 32168 38286
rect 32402 38247 32458 38256
rect 32416 37874 32444 38247
rect 32404 37868 32456 37874
rect 32404 37810 32456 37816
rect 32128 37392 32180 37398
rect 32128 37334 32180 37340
rect 32692 36689 32720 40996
rect 33152 37346 33180 40996
rect 33612 39438 33640 40996
rect 34426 39536 34482 39545
rect 34426 39471 34482 39480
rect 33600 39432 33652 39438
rect 33600 39374 33652 39380
rect 33232 38208 33284 38214
rect 33232 38150 33284 38156
rect 33244 38049 33272 38150
rect 33230 38040 33286 38049
rect 33230 37975 33286 37984
rect 33244 37942 33272 37975
rect 33232 37936 33284 37942
rect 33232 37878 33284 37884
rect 33232 37800 33284 37806
rect 33232 37742 33284 37748
rect 33060 37318 33180 37346
rect 33244 37330 33272 37742
rect 34440 37330 34468 39471
rect 34532 39302 34560 40996
rect 34992 39386 35020 40996
rect 35254 40216 35310 40225
rect 35254 40151 35310 40160
rect 35268 40118 35296 40151
rect 35256 40112 35308 40118
rect 35256 40054 35308 40060
rect 34808 39358 35020 39386
rect 34520 39296 34572 39302
rect 34520 39238 34572 39244
rect 34808 37777 34836 39358
rect 34940 39196 35236 39216
rect 34996 39194 35020 39196
rect 35076 39194 35100 39196
rect 35156 39194 35180 39196
rect 35018 39142 35020 39194
rect 35082 39142 35094 39194
rect 35156 39142 35158 39194
rect 34996 39140 35020 39142
rect 35076 39140 35100 39142
rect 35156 39140 35180 39142
rect 34940 39120 35236 39140
rect 35256 38956 35308 38962
rect 35256 38898 35308 38904
rect 35268 38865 35296 38898
rect 35254 38856 35310 38865
rect 35254 38791 35310 38800
rect 34940 38108 35236 38128
rect 34996 38106 35020 38108
rect 35076 38106 35100 38108
rect 35156 38106 35180 38108
rect 35018 38054 35020 38106
rect 35082 38054 35094 38106
rect 35156 38054 35158 38106
rect 34996 38052 35020 38054
rect 35076 38052 35100 38054
rect 35156 38052 35180 38054
rect 34940 38032 35236 38052
rect 34794 37768 34850 37777
rect 34794 37703 34850 37712
rect 34796 37460 34848 37466
rect 34796 37402 34848 37408
rect 33232 37324 33284 37330
rect 32678 36680 32734 36689
rect 32678 36615 32734 36624
rect 31942 35320 31998 35329
rect 31942 35255 31998 35264
rect 31852 28688 31904 28694
rect 31852 28630 31904 28636
rect 31668 28212 31720 28218
rect 31668 28154 31720 28160
rect 31760 28212 31812 28218
rect 31760 28154 31812 28160
rect 31852 27464 31904 27470
rect 31852 27406 31904 27412
rect 31864 27130 31892 27406
rect 31852 27124 31904 27130
rect 31852 27066 31904 27072
rect 31852 25900 31904 25906
rect 31852 25842 31904 25848
rect 31864 25498 31892 25842
rect 31852 25492 31904 25498
rect 31852 25434 31904 25440
rect 31588 25214 31892 25242
rect 31576 25152 31628 25158
rect 31576 25094 31628 25100
rect 31588 24886 31616 25094
rect 31576 24880 31628 24886
rect 31576 24822 31628 24828
rect 31392 24812 31444 24818
rect 31392 24754 31444 24760
rect 31404 24410 31432 24754
rect 31484 24744 31536 24750
rect 31484 24686 31536 24692
rect 31392 24404 31444 24410
rect 31392 24346 31444 24352
rect 31496 24274 31524 24686
rect 31760 24676 31812 24682
rect 31760 24618 31812 24624
rect 31574 24576 31630 24585
rect 31574 24511 31630 24520
rect 31484 24268 31536 24274
rect 31484 24210 31536 24216
rect 31588 24138 31616 24511
rect 31576 24132 31628 24138
rect 31576 24074 31628 24080
rect 30984 23684 31064 23712
rect 30932 23666 30984 23672
rect 31036 23322 31064 23684
rect 31116 23724 31168 23730
rect 31116 23666 31168 23672
rect 31128 23322 31156 23666
rect 31588 23662 31616 24074
rect 31772 23662 31800 24618
rect 31576 23656 31628 23662
rect 31576 23598 31628 23604
rect 31760 23656 31812 23662
rect 31760 23598 31812 23604
rect 31772 23322 31800 23598
rect 31024 23316 31076 23322
rect 31024 23258 31076 23264
rect 31116 23316 31168 23322
rect 31116 23258 31168 23264
rect 31760 23316 31812 23322
rect 31760 23258 31812 23264
rect 31760 23112 31812 23118
rect 31760 23054 31812 23060
rect 30840 22500 30892 22506
rect 30840 22442 30892 22448
rect 31576 22500 31628 22506
rect 31576 22442 31628 22448
rect 31300 22092 31352 22098
rect 31300 22034 31352 22040
rect 31312 21554 31340 22034
rect 31300 21548 31352 21554
rect 31300 21490 31352 21496
rect 31312 20806 31340 21490
rect 31392 21480 31444 21486
rect 31392 21422 31444 21428
rect 31300 20800 31352 20806
rect 31300 20742 31352 20748
rect 31116 20256 31168 20262
rect 31116 20198 31168 20204
rect 30932 19168 30984 19174
rect 30852 19128 30932 19156
rect 30852 18290 30880 19128
rect 30932 19110 30984 19116
rect 30932 18624 30984 18630
rect 30932 18566 30984 18572
rect 30840 18284 30892 18290
rect 30840 18226 30892 18232
rect 30852 17882 30880 18226
rect 30840 17876 30892 17882
rect 30840 17818 30892 17824
rect 30760 16748 30880 16776
rect 30288 16720 30340 16726
rect 30288 16662 30340 16668
rect 30746 16688 30802 16697
rect 30196 16652 30248 16658
rect 30196 16594 30248 16600
rect 30208 16114 30236 16594
rect 30196 16108 30248 16114
rect 30196 16050 30248 16056
rect 29828 16040 29880 16046
rect 29828 15982 29880 15988
rect 29840 15026 29868 15982
rect 30012 15564 30064 15570
rect 30012 15506 30064 15512
rect 29920 15428 29972 15434
rect 29920 15370 29972 15376
rect 29828 15020 29880 15026
rect 29828 14962 29880 14968
rect 29840 14482 29868 14962
rect 29932 14618 29960 15370
rect 30024 14890 30052 15506
rect 30208 15450 30236 16050
rect 30300 15722 30328 16662
rect 30746 16623 30748 16632
rect 30800 16623 30802 16632
rect 30748 16594 30800 16600
rect 30760 16250 30788 16594
rect 30748 16244 30800 16250
rect 30748 16186 30800 16192
rect 30300 15706 30512 15722
rect 30300 15700 30524 15706
rect 30300 15694 30472 15700
rect 30472 15642 30524 15648
rect 30288 15632 30340 15638
rect 30340 15592 30420 15620
rect 30288 15574 30340 15580
rect 30116 15422 30236 15450
rect 30012 14884 30064 14890
rect 30012 14826 30064 14832
rect 29920 14612 29972 14618
rect 29920 14554 29972 14560
rect 29828 14476 29880 14482
rect 29828 14418 29880 14424
rect 29840 14074 29868 14418
rect 29828 14068 29880 14074
rect 29828 14010 29880 14016
rect 29472 13654 29684 13682
rect 29276 13524 29328 13530
rect 29276 13466 29328 13472
rect 29288 13190 29316 13466
rect 29276 13184 29328 13190
rect 29276 13126 29328 13132
rect 29472 11393 29500 13654
rect 29552 13456 29604 13462
rect 29552 13398 29604 13404
rect 29564 12782 29592 13398
rect 29840 13394 29868 14010
rect 29932 14006 29960 14554
rect 29920 14000 29972 14006
rect 29920 13942 29972 13948
rect 30012 13796 30064 13802
rect 30012 13738 30064 13744
rect 29828 13388 29880 13394
rect 29828 13330 29880 13336
rect 30024 13258 30052 13738
rect 30116 13462 30144 15422
rect 30196 15360 30248 15366
rect 30196 15302 30248 15308
rect 30208 14958 30236 15302
rect 30196 14952 30248 14958
rect 30196 14894 30248 14900
rect 30208 14414 30236 14894
rect 30392 14890 30420 15592
rect 30564 15496 30616 15502
rect 30564 15438 30616 15444
rect 30470 15328 30526 15337
rect 30470 15263 30526 15272
rect 30380 14884 30432 14890
rect 30380 14826 30432 14832
rect 30484 14618 30512 15263
rect 30576 15026 30604 15438
rect 30564 15020 30616 15026
rect 30564 14962 30616 14968
rect 30472 14612 30524 14618
rect 30472 14554 30524 14560
rect 30380 14476 30432 14482
rect 30380 14418 30432 14424
rect 30196 14408 30248 14414
rect 30196 14350 30248 14356
rect 30104 13456 30156 13462
rect 30104 13398 30156 13404
rect 30208 13394 30236 14350
rect 30196 13388 30248 13394
rect 30196 13330 30248 13336
rect 30012 13252 30064 13258
rect 30012 13194 30064 13200
rect 30208 12986 30236 13330
rect 30392 13161 30420 14418
rect 30472 14068 30524 14074
rect 30472 14010 30524 14016
rect 30378 13152 30434 13161
rect 30378 13087 30434 13096
rect 30196 12980 30248 12986
rect 30196 12922 30248 12928
rect 30392 12850 30420 13087
rect 30380 12844 30432 12850
rect 30380 12786 30432 12792
rect 29552 12776 29604 12782
rect 29552 12718 29604 12724
rect 29564 12442 29592 12718
rect 30484 12442 30512 14010
rect 30564 13252 30616 13258
rect 30564 13194 30616 13200
rect 30576 12986 30604 13194
rect 30564 12980 30616 12986
rect 30564 12922 30616 12928
rect 30656 12776 30708 12782
rect 30656 12718 30708 12724
rect 30564 12708 30616 12714
rect 30564 12650 30616 12656
rect 30576 12442 30604 12650
rect 29552 12436 29604 12442
rect 29552 12378 29604 12384
rect 30472 12436 30524 12442
rect 30472 12378 30524 12384
rect 30564 12436 30616 12442
rect 30564 12378 30616 12384
rect 29642 12336 29698 12345
rect 29642 12271 29644 12280
rect 29696 12271 29698 12280
rect 29644 12242 29696 12248
rect 29656 11898 29684 12242
rect 29644 11892 29696 11898
rect 29644 11834 29696 11840
rect 30380 11552 30432 11558
rect 30380 11494 30432 11500
rect 29458 11384 29514 11393
rect 29458 11319 29514 11328
rect 29920 11144 29972 11150
rect 29920 11086 29972 11092
rect 29550 10840 29606 10849
rect 29550 10775 29606 10784
rect 29458 5536 29514 5545
rect 29458 5471 29514 5480
rect 29274 4448 29330 4457
rect 29274 4383 29330 4392
rect 29184 2576 29236 2582
rect 29184 2518 29236 2524
rect 29092 2100 29144 2106
rect 29092 2042 29144 2048
rect 29288 1442 29316 4383
rect 29368 2984 29420 2990
rect 29368 2926 29420 2932
rect 29380 2825 29408 2926
rect 29366 2816 29422 2825
rect 29366 2751 29422 2760
rect 29380 2650 29408 2751
rect 29368 2644 29420 2650
rect 29368 2586 29420 2592
rect 29012 1414 29316 1442
rect 29012 800 29040 1414
rect 29472 800 29500 5471
rect 29564 3194 29592 10775
rect 29552 3188 29604 3194
rect 29552 3130 29604 3136
rect 29564 2990 29592 3130
rect 29552 2984 29604 2990
rect 29552 2926 29604 2932
rect 29932 800 29960 11086
rect 30196 10804 30248 10810
rect 30196 10746 30248 10752
rect 30208 10266 30236 10746
rect 30392 10742 30420 11494
rect 30668 11218 30696 12718
rect 30748 11892 30800 11898
rect 30748 11834 30800 11840
rect 30760 11218 30788 11834
rect 30656 11212 30708 11218
rect 30656 11154 30708 11160
rect 30748 11212 30800 11218
rect 30748 11154 30800 11160
rect 30380 10736 30432 10742
rect 30380 10678 30432 10684
rect 30668 10606 30696 11154
rect 30760 10674 30788 11154
rect 30748 10668 30800 10674
rect 30748 10610 30800 10616
rect 30656 10600 30708 10606
rect 30656 10542 30708 10548
rect 30668 10470 30696 10542
rect 30656 10464 30708 10470
rect 30656 10406 30708 10412
rect 30196 10260 30248 10266
rect 30196 10202 30248 10208
rect 30668 10130 30696 10406
rect 30760 10266 30788 10610
rect 30748 10260 30800 10266
rect 30748 10202 30800 10208
rect 30656 10124 30708 10130
rect 30656 10066 30708 10072
rect 30852 6905 30880 16748
rect 30944 16454 30972 18566
rect 31024 16720 31076 16726
rect 31024 16662 31076 16668
rect 30932 16448 30984 16454
rect 30932 16390 30984 16396
rect 30944 16114 30972 16390
rect 31036 16182 31064 16662
rect 31024 16176 31076 16182
rect 31024 16118 31076 16124
rect 30932 16108 30984 16114
rect 30932 16050 30984 16056
rect 31024 14476 31076 14482
rect 31024 14418 31076 14424
rect 30932 13864 30984 13870
rect 30932 13806 30984 13812
rect 30944 13025 30972 13806
rect 31036 13530 31064 14418
rect 31024 13524 31076 13530
rect 31024 13466 31076 13472
rect 31128 13410 31156 20198
rect 31206 19000 31262 19009
rect 31206 18935 31208 18944
rect 31260 18935 31262 18944
rect 31208 18906 31260 18912
rect 31220 18222 31248 18906
rect 31208 18216 31260 18222
rect 31208 18158 31260 18164
rect 31208 17536 31260 17542
rect 31208 17478 31260 17484
rect 31220 17202 31248 17478
rect 31312 17270 31340 20742
rect 31404 17921 31432 21422
rect 31482 20768 31538 20777
rect 31482 20703 31538 20712
rect 31496 20398 31524 20703
rect 31484 20392 31536 20398
rect 31484 20334 31536 20340
rect 31496 20058 31524 20334
rect 31484 20052 31536 20058
rect 31484 19994 31536 20000
rect 31484 19712 31536 19718
rect 31484 19654 31536 19660
rect 31496 19446 31524 19654
rect 31484 19440 31536 19446
rect 31484 19382 31536 19388
rect 31496 18086 31524 19382
rect 31484 18080 31536 18086
rect 31484 18022 31536 18028
rect 31390 17912 31446 17921
rect 31390 17847 31446 17856
rect 31390 17368 31446 17377
rect 31390 17303 31446 17312
rect 31300 17264 31352 17270
rect 31300 17206 31352 17212
rect 31208 17196 31260 17202
rect 31208 17138 31260 17144
rect 31300 17060 31352 17066
rect 31300 17002 31352 17008
rect 31312 16794 31340 17002
rect 31404 16794 31432 17303
rect 31300 16788 31352 16794
rect 31300 16730 31352 16736
rect 31392 16788 31444 16794
rect 31392 16730 31444 16736
rect 31390 15192 31446 15201
rect 31390 15127 31446 15136
rect 31404 14550 31432 15127
rect 31392 14544 31444 14550
rect 31392 14486 31444 14492
rect 31404 14414 31432 14486
rect 31392 14408 31444 14414
rect 31392 14350 31444 14356
rect 31588 14362 31616 22442
rect 31668 21888 31720 21894
rect 31668 21830 31720 21836
rect 31680 21486 31708 21830
rect 31668 21480 31720 21486
rect 31668 21422 31720 21428
rect 31680 20505 31708 21422
rect 31666 20496 31722 20505
rect 31666 20431 31722 20440
rect 31668 19236 31720 19242
rect 31668 19178 31720 19184
rect 31680 18630 31708 19178
rect 31668 18624 31720 18630
rect 31668 18566 31720 18572
rect 31772 18306 31800 23054
rect 31864 20534 31892 25214
rect 31852 20528 31904 20534
rect 31852 20470 31904 20476
rect 31956 18358 31984 35255
rect 32036 33312 32088 33318
rect 32036 33254 32088 33260
rect 32048 30190 32076 33254
rect 32770 32056 32826 32065
rect 32770 31991 32826 32000
rect 32128 31340 32180 31346
rect 32128 31282 32180 31288
rect 32140 30394 32168 31282
rect 32128 30388 32180 30394
rect 32128 30330 32180 30336
rect 32036 30184 32088 30190
rect 32036 30126 32088 30132
rect 32126 29472 32182 29481
rect 32126 29407 32182 29416
rect 32034 26072 32090 26081
rect 32034 26007 32090 26016
rect 32048 19378 32076 26007
rect 32140 24818 32168 29407
rect 32220 29096 32272 29102
rect 32220 29038 32272 29044
rect 32232 28422 32260 29038
rect 32220 28416 32272 28422
rect 32220 28358 32272 28364
rect 32232 27538 32260 28358
rect 32680 28008 32732 28014
rect 32680 27950 32732 27956
rect 32692 27606 32720 27950
rect 32680 27600 32732 27606
rect 32680 27542 32732 27548
rect 32220 27532 32272 27538
rect 32220 27474 32272 27480
rect 32232 26790 32260 27474
rect 32678 27432 32734 27441
rect 32678 27367 32734 27376
rect 32496 27124 32548 27130
rect 32496 27066 32548 27072
rect 32404 26920 32456 26926
rect 32404 26862 32456 26868
rect 32220 26784 32272 26790
rect 32220 26726 32272 26732
rect 32232 25362 32260 26726
rect 32416 26586 32444 26862
rect 32404 26580 32456 26586
rect 32404 26522 32456 26528
rect 32312 25968 32364 25974
rect 32312 25910 32364 25916
rect 32324 25702 32352 25910
rect 32404 25764 32456 25770
rect 32404 25706 32456 25712
rect 32312 25696 32364 25702
rect 32312 25638 32364 25644
rect 32220 25356 32272 25362
rect 32220 25298 32272 25304
rect 32220 25220 32272 25226
rect 32220 25162 32272 25168
rect 32128 24812 32180 24818
rect 32128 24754 32180 24760
rect 32232 24614 32260 25162
rect 32220 24608 32272 24614
rect 32220 24550 32272 24556
rect 32232 24274 32260 24550
rect 32324 24410 32352 25638
rect 32312 24404 32364 24410
rect 32312 24346 32364 24352
rect 32220 24268 32272 24274
rect 32220 24210 32272 24216
rect 32128 23112 32180 23118
rect 32128 23054 32180 23060
rect 32140 22778 32168 23054
rect 32128 22772 32180 22778
rect 32128 22714 32180 22720
rect 32312 20936 32364 20942
rect 32312 20878 32364 20884
rect 32128 20800 32180 20806
rect 32128 20742 32180 20748
rect 32140 20398 32168 20742
rect 32128 20392 32180 20398
rect 32128 20334 32180 20340
rect 32140 19854 32168 20334
rect 32324 20262 32352 20878
rect 32312 20256 32364 20262
rect 32312 20198 32364 20204
rect 32128 19848 32180 19854
rect 32128 19790 32180 19796
rect 32036 19372 32088 19378
rect 32036 19314 32088 19320
rect 31944 18352 31996 18358
rect 31772 18278 31892 18306
rect 31944 18294 31996 18300
rect 31760 18216 31812 18222
rect 31760 18158 31812 18164
rect 31668 17536 31720 17542
rect 31668 17478 31720 17484
rect 31680 17134 31708 17478
rect 31668 17128 31720 17134
rect 31668 17070 31720 17076
rect 31680 16726 31708 17070
rect 31772 17066 31800 18158
rect 31864 17762 31892 18278
rect 32220 18148 32272 18154
rect 32220 18090 32272 18096
rect 31864 17734 32076 17762
rect 31760 17060 31812 17066
rect 31760 17002 31812 17008
rect 31668 16720 31720 16726
rect 31668 16662 31720 16668
rect 31942 16552 31998 16561
rect 31942 16487 31998 16496
rect 31852 16040 31904 16046
rect 31956 16017 31984 16487
rect 31852 15982 31904 15988
rect 31942 16008 31998 16017
rect 31760 15700 31812 15706
rect 31760 15642 31812 15648
rect 31772 14498 31800 15642
rect 31864 15162 31892 15982
rect 31942 15943 31998 15952
rect 31956 15570 31984 15943
rect 31944 15564 31996 15570
rect 31944 15506 31996 15512
rect 31956 15162 31984 15506
rect 31852 15156 31904 15162
rect 31852 15098 31904 15104
rect 31944 15156 31996 15162
rect 31944 15098 31996 15104
rect 31680 14482 31800 14498
rect 31668 14476 31800 14482
rect 31720 14470 31800 14476
rect 31668 14418 31720 14424
rect 31404 13870 31432 14350
rect 31588 14334 31708 14362
rect 31392 13864 31444 13870
rect 31392 13806 31444 13812
rect 31576 13796 31628 13802
rect 31576 13738 31628 13744
rect 31588 13530 31616 13738
rect 31576 13524 31628 13530
rect 31576 13466 31628 13472
rect 31036 13382 31156 13410
rect 30930 13016 30986 13025
rect 30930 12951 30986 12960
rect 30932 12300 30984 12306
rect 30932 12242 30984 12248
rect 30944 12073 30972 12242
rect 31036 12170 31064 13382
rect 31116 13320 31168 13326
rect 31116 13262 31168 13268
rect 31128 12782 31156 13262
rect 31680 12782 31708 14334
rect 31944 14272 31996 14278
rect 31944 14214 31996 14220
rect 31760 14068 31812 14074
rect 31760 14010 31812 14016
rect 31772 13394 31800 14010
rect 31956 14006 31984 14214
rect 31944 14000 31996 14006
rect 31944 13942 31996 13948
rect 31956 13530 31984 13942
rect 31944 13524 31996 13530
rect 31944 13466 31996 13472
rect 31760 13388 31812 13394
rect 31760 13330 31812 13336
rect 31852 13184 31904 13190
rect 31850 13152 31852 13161
rect 31904 13152 31906 13161
rect 31850 13087 31906 13096
rect 31116 12776 31168 12782
rect 31116 12718 31168 12724
rect 31668 12776 31720 12782
rect 31668 12718 31720 12724
rect 31944 12776 31996 12782
rect 31944 12718 31996 12724
rect 31024 12164 31076 12170
rect 31024 12106 31076 12112
rect 30930 12064 30986 12073
rect 30930 11999 30986 12008
rect 30944 11830 30972 11999
rect 30932 11824 30984 11830
rect 30932 11766 30984 11772
rect 31036 11694 31064 12106
rect 31484 12096 31536 12102
rect 31484 12038 31536 12044
rect 31024 11688 31076 11694
rect 31024 11630 31076 11636
rect 31496 11286 31524 12038
rect 31680 11762 31708 12718
rect 31956 12102 31984 12718
rect 31944 12096 31996 12102
rect 31944 12038 31996 12044
rect 31668 11756 31720 11762
rect 31668 11698 31720 11704
rect 31484 11280 31536 11286
rect 31484 11222 31536 11228
rect 31024 11212 31076 11218
rect 31024 11154 31076 11160
rect 31036 10810 31064 11154
rect 31024 10804 31076 10810
rect 31024 10746 31076 10752
rect 32048 10713 32076 17734
rect 32232 16522 32260 18090
rect 32220 16516 32272 16522
rect 32220 16458 32272 16464
rect 32232 15978 32260 16458
rect 32220 15972 32272 15978
rect 32220 15914 32272 15920
rect 32220 15564 32272 15570
rect 32220 15506 32272 15512
rect 32126 14512 32182 14521
rect 32126 14447 32128 14456
rect 32180 14447 32182 14456
rect 32128 14418 32180 14424
rect 32140 14074 32168 14418
rect 32128 14068 32180 14074
rect 32128 14010 32180 14016
rect 32034 10704 32090 10713
rect 32034 10639 32090 10648
rect 31392 10532 31444 10538
rect 31392 10474 31444 10480
rect 30838 6896 30894 6905
rect 30838 6831 30894 6840
rect 31404 5001 31432 10474
rect 32232 7857 32260 15506
rect 32324 12764 32352 20198
rect 32416 15570 32444 25706
rect 32508 23118 32536 27066
rect 32692 25430 32720 27367
rect 32680 25424 32732 25430
rect 32680 25366 32732 25372
rect 32588 25356 32640 25362
rect 32588 25298 32640 25304
rect 32600 24410 32628 25298
rect 32588 24404 32640 24410
rect 32588 24346 32640 24352
rect 32680 24268 32732 24274
rect 32680 24210 32732 24216
rect 32692 23526 32720 24210
rect 32680 23520 32732 23526
rect 32680 23462 32732 23468
rect 32496 23112 32548 23118
rect 32496 23054 32548 23060
rect 32508 22778 32536 23054
rect 32496 22772 32548 22778
rect 32496 22714 32548 22720
rect 32496 21004 32548 21010
rect 32496 20946 32548 20952
rect 32508 20466 32536 20946
rect 32496 20460 32548 20466
rect 32496 20402 32548 20408
rect 32508 20330 32536 20402
rect 32496 20324 32548 20330
rect 32496 20266 32548 20272
rect 32508 19990 32536 20266
rect 32496 19984 32548 19990
rect 32496 19926 32548 19932
rect 32508 19174 32536 19926
rect 32496 19168 32548 19174
rect 32496 19110 32548 19116
rect 32588 19168 32640 19174
rect 32588 19110 32640 19116
rect 32508 17746 32536 19110
rect 32600 18630 32628 19110
rect 32588 18624 32640 18630
rect 32588 18566 32640 18572
rect 32496 17740 32548 17746
rect 32496 17682 32548 17688
rect 32588 17672 32640 17678
rect 32588 17614 32640 17620
rect 32600 17338 32628 17614
rect 32588 17332 32640 17338
rect 32588 17274 32640 17280
rect 32496 17128 32548 17134
rect 32496 17070 32548 17076
rect 32508 16658 32536 17070
rect 32496 16652 32548 16658
rect 32496 16594 32548 16600
rect 32494 15600 32550 15609
rect 32404 15564 32456 15570
rect 32494 15535 32496 15544
rect 32404 15506 32456 15512
rect 32548 15535 32550 15544
rect 32496 15506 32548 15512
rect 32600 15162 32628 17274
rect 32588 15156 32640 15162
rect 32588 15098 32640 15104
rect 32600 14958 32628 15098
rect 32588 14952 32640 14958
rect 32588 14894 32640 14900
rect 32600 14618 32628 14894
rect 32588 14612 32640 14618
rect 32588 14554 32640 14560
rect 32588 14272 32640 14278
rect 32588 14214 32640 14220
rect 32600 13870 32628 14214
rect 32588 13864 32640 13870
rect 32588 13806 32640 13812
rect 32496 13388 32548 13394
rect 32496 13330 32548 13336
rect 32508 12986 32536 13330
rect 32496 12980 32548 12986
rect 32496 12922 32548 12928
rect 32324 12736 32536 12764
rect 32508 12442 32536 12736
rect 32496 12436 32548 12442
rect 32496 12378 32548 12384
rect 32508 12306 32536 12378
rect 32496 12300 32548 12306
rect 32496 12242 32548 12248
rect 32218 7848 32274 7857
rect 32218 7783 32274 7792
rect 31390 4992 31446 5001
rect 31390 4927 31446 4936
rect 32692 4808 32720 23462
rect 32784 21554 32812 31991
rect 32864 30184 32916 30190
rect 32864 30126 32916 30132
rect 32956 30184 33008 30190
rect 32956 30126 33008 30132
rect 32876 25498 32904 30126
rect 32968 29850 32996 30126
rect 32956 29844 33008 29850
rect 32956 29786 33008 29792
rect 32968 29646 32996 29786
rect 32956 29640 33008 29646
rect 32956 29582 33008 29588
rect 32956 26852 33008 26858
rect 32956 26794 33008 26800
rect 32968 25838 32996 26794
rect 32956 25832 33008 25838
rect 32956 25774 33008 25780
rect 32864 25492 32916 25498
rect 32864 25434 32916 25440
rect 32956 24744 33008 24750
rect 32956 24686 33008 24692
rect 32968 24410 32996 24686
rect 32956 24404 33008 24410
rect 32956 24346 33008 24352
rect 32864 23588 32916 23594
rect 32864 23530 32916 23536
rect 32772 21548 32824 21554
rect 32772 21490 32824 21496
rect 32772 18080 32824 18086
rect 32772 18022 32824 18028
rect 32784 12918 32812 18022
rect 32876 17218 32904 23530
rect 32956 23180 33008 23186
rect 32956 23122 33008 23128
rect 32968 22710 32996 23122
rect 32956 22704 33008 22710
rect 32954 22672 32956 22681
rect 33008 22672 33010 22681
rect 32954 22607 33010 22616
rect 33060 22522 33088 37318
rect 33232 37266 33284 37272
rect 33600 37324 33652 37330
rect 33600 37266 33652 37272
rect 33876 37324 33928 37330
rect 33876 37266 33928 37272
rect 34428 37324 34480 37330
rect 34428 37266 34480 37272
rect 34520 37324 34572 37330
rect 34520 37266 34572 37272
rect 33612 31929 33640 37266
rect 33888 36922 33916 37266
rect 34532 36938 34560 37266
rect 34440 36922 34560 36938
rect 33876 36916 33928 36922
rect 33876 36858 33928 36864
rect 34428 36916 34560 36922
rect 34480 36910 34560 36916
rect 34428 36858 34480 36864
rect 34610 33960 34666 33969
rect 34610 33895 34666 33904
rect 33598 31920 33654 31929
rect 33598 31855 33654 31864
rect 33416 30116 33468 30122
rect 33416 30058 33468 30064
rect 33140 28484 33192 28490
rect 33140 28426 33192 28432
rect 33152 28014 33180 28426
rect 33232 28416 33284 28422
rect 33232 28358 33284 28364
rect 33140 28008 33192 28014
rect 33140 27950 33192 27956
rect 33152 27334 33180 27950
rect 33140 27328 33192 27334
rect 33140 27270 33192 27276
rect 33152 27033 33180 27270
rect 33138 27024 33194 27033
rect 33138 26959 33194 26968
rect 32968 22494 33088 22522
rect 32968 22030 32996 22494
rect 33048 22092 33100 22098
rect 33048 22034 33100 22040
rect 32956 22024 33008 22030
rect 32956 21966 33008 21972
rect 32968 21690 32996 21966
rect 33060 21690 33088 22034
rect 32956 21684 33008 21690
rect 32956 21626 33008 21632
rect 33048 21684 33100 21690
rect 33048 21626 33100 21632
rect 33048 21004 33100 21010
rect 33048 20946 33100 20952
rect 33060 19854 33088 20946
rect 33140 19916 33192 19922
rect 33140 19858 33192 19864
rect 33048 19848 33100 19854
rect 33048 19790 33100 19796
rect 33048 19712 33100 19718
rect 33048 19654 33100 19660
rect 33060 19553 33088 19654
rect 33046 19544 33102 19553
rect 33046 19479 33102 19488
rect 32956 19372 33008 19378
rect 32956 19314 33008 19320
rect 32968 18970 32996 19314
rect 33060 19258 33088 19479
rect 33152 19378 33180 19858
rect 33140 19372 33192 19378
rect 33140 19314 33192 19320
rect 33060 19230 33180 19258
rect 33152 19174 33180 19230
rect 33140 19168 33192 19174
rect 33140 19110 33192 19116
rect 32956 18964 33008 18970
rect 32956 18906 33008 18912
rect 32968 18358 32996 18906
rect 33048 18760 33100 18766
rect 33048 18702 33100 18708
rect 33060 18426 33088 18702
rect 33048 18420 33100 18426
rect 33048 18362 33100 18368
rect 32956 18352 33008 18358
rect 33008 18300 33180 18306
rect 32956 18294 33180 18300
rect 32968 18278 33180 18294
rect 33048 18148 33100 18154
rect 33048 18090 33100 18096
rect 32876 17190 32996 17218
rect 32864 17128 32916 17134
rect 32864 17070 32916 17076
rect 32876 16794 32904 17070
rect 32864 16788 32916 16794
rect 32864 16730 32916 16736
rect 32864 16584 32916 16590
rect 32864 16526 32916 16532
rect 32876 15910 32904 16526
rect 32864 15904 32916 15910
rect 32864 15846 32916 15852
rect 32876 13870 32904 15846
rect 32968 14498 32996 17190
rect 33060 16590 33088 18090
rect 33152 17746 33180 18278
rect 33140 17740 33192 17746
rect 33140 17682 33192 17688
rect 33048 16584 33100 16590
rect 33048 16526 33100 16532
rect 33140 15564 33192 15570
rect 33140 15506 33192 15512
rect 33152 15162 33180 15506
rect 33140 15156 33192 15162
rect 33140 15098 33192 15104
rect 33048 15020 33100 15026
rect 33048 14962 33100 14968
rect 33060 14618 33088 14962
rect 33048 14612 33100 14618
rect 33048 14554 33100 14560
rect 32968 14470 33088 14498
rect 32864 13864 32916 13870
rect 32864 13806 32916 13812
rect 32864 13320 32916 13326
rect 32864 13262 32916 13268
rect 32876 12986 32904 13262
rect 32864 12980 32916 12986
rect 32864 12922 32916 12928
rect 32772 12912 32824 12918
rect 32772 12854 32824 12860
rect 32864 12300 32916 12306
rect 32864 12242 32916 12248
rect 32876 11898 32904 12242
rect 32864 11892 32916 11898
rect 32864 11834 32916 11840
rect 32692 4780 32812 4808
rect 32680 4684 32732 4690
rect 32680 4626 32732 4632
rect 32128 4616 32180 4622
rect 32128 4558 32180 4564
rect 32140 3942 32168 4558
rect 32692 4010 32720 4626
rect 32680 4004 32732 4010
rect 32680 3946 32732 3952
rect 32128 3936 32180 3942
rect 32128 3878 32180 3884
rect 32140 3534 32168 3878
rect 32128 3528 32180 3534
rect 32128 3470 32180 3476
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 32140 2990 32168 3470
rect 32220 3052 32272 3058
rect 32220 2994 32272 3000
rect 32128 2984 32180 2990
rect 32128 2926 32180 2932
rect 31300 2916 31352 2922
rect 31300 2858 31352 2864
rect 30838 2816 30894 2825
rect 30838 2751 30894 2760
rect 30852 800 30880 2751
rect 31312 800 31340 2858
rect 32140 2650 32168 2926
rect 32128 2644 32180 2650
rect 32128 2586 32180 2592
rect 32232 800 32260 2994
rect 32416 2310 32444 3470
rect 32404 2304 32456 2310
rect 32404 2246 32456 2252
rect 32416 1766 32444 2246
rect 32404 1760 32456 1766
rect 32404 1702 32456 1708
rect 32692 800 32720 3946
rect 32784 3233 32812 4780
rect 33060 4457 33088 14470
rect 33152 13870 33180 15098
rect 33140 13864 33192 13870
rect 33140 13806 33192 13812
rect 33152 13530 33180 13806
rect 33140 13524 33192 13530
rect 33140 13466 33192 13472
rect 33138 5264 33194 5273
rect 33138 5199 33194 5208
rect 33046 4448 33102 4457
rect 33046 4383 33102 4392
rect 33152 3738 33180 5199
rect 33140 3732 33192 3738
rect 33140 3674 33192 3680
rect 32770 3224 32826 3233
rect 32770 3159 32772 3168
rect 32824 3159 32826 3168
rect 32772 3130 32824 3136
rect 32784 3099 32812 3130
rect 33048 1760 33100 1766
rect 33100 1708 33180 1714
rect 33048 1702 33180 1708
rect 33060 1686 33180 1702
rect 33152 800 33180 1686
rect 1398 776 1454 785
rect 1398 711 1454 720
rect 1858 0 1914 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3698 0 3754 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6918 0 6974 800
rect 7378 0 7434 800
rect 7838 0 7894 800
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 9678 0 9734 800
rect 10598 0 10654 800
rect 11058 0 11114 800
rect 11978 0 12034 800
rect 12438 0 12494 800
rect 12898 0 12954 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 14738 0 14794 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 17958 0 18014 800
rect 18878 0 18934 800
rect 19338 0 19394 800
rect 19798 0 19854 800
rect 20718 0 20774 800
rect 21178 0 21234 800
rect 22098 0 22154 800
rect 22558 0 22614 800
rect 23018 0 23074 800
rect 23938 0 23994 800
rect 24398 0 24454 800
rect 24858 0 24914 800
rect 25778 0 25834 800
rect 26238 0 26294 800
rect 27158 0 27214 800
rect 27618 0 27674 800
rect 28078 0 28134 800
rect 28998 0 29054 800
rect 29458 0 29514 800
rect 29918 0 29974 800
rect 30838 0 30894 800
rect 31298 0 31354 800
rect 32218 0 32274 800
rect 32678 0 32734 800
rect 33138 0 33194 800
rect 33244 105 33272 28358
rect 33322 21312 33378 21321
rect 33322 21247 33378 21256
rect 33336 21078 33364 21247
rect 33324 21072 33376 21078
rect 33324 21014 33376 21020
rect 33324 17196 33376 17202
rect 33324 17138 33376 17144
rect 33336 16726 33364 17138
rect 33324 16720 33376 16726
rect 33324 16662 33376 16668
rect 33336 16046 33364 16662
rect 33324 16040 33376 16046
rect 33324 15982 33376 15988
rect 33428 10305 33456 30058
rect 33612 27606 33640 31855
rect 33692 29708 33744 29714
rect 33692 29650 33744 29656
rect 33704 29306 33732 29650
rect 34348 29646 34376 29677
rect 33968 29640 34020 29646
rect 33968 29582 34020 29588
rect 34152 29640 34204 29646
rect 34336 29640 34388 29646
rect 34152 29582 34204 29588
rect 34334 29608 34336 29617
rect 34388 29608 34390 29617
rect 33980 29306 34008 29582
rect 33692 29300 33744 29306
rect 33692 29242 33744 29248
rect 33968 29300 34020 29306
rect 33968 29242 34020 29248
rect 33784 28620 33836 28626
rect 33784 28562 33836 28568
rect 33692 28552 33744 28558
rect 33692 28494 33744 28500
rect 33704 27878 33732 28494
rect 33796 28082 33824 28562
rect 33784 28076 33836 28082
rect 33784 28018 33836 28024
rect 33692 27872 33744 27878
rect 33692 27814 33744 27820
rect 33600 27600 33652 27606
rect 33600 27542 33652 27548
rect 33612 27334 33640 27542
rect 33704 27441 33732 27814
rect 34164 27441 34192 29582
rect 34334 29543 34390 29552
rect 34348 29306 34376 29543
rect 34336 29300 34388 29306
rect 34336 29242 34388 29248
rect 33690 27432 33746 27441
rect 33690 27367 33746 27376
rect 34150 27432 34206 27441
rect 34150 27367 34206 27376
rect 33600 27328 33652 27334
rect 33600 27270 33652 27276
rect 34348 27130 34376 29242
rect 34520 27532 34572 27538
rect 34520 27474 34572 27480
rect 34336 27124 34388 27130
rect 34336 27066 34388 27072
rect 34532 26790 34560 27474
rect 34520 26784 34572 26790
rect 34520 26726 34572 26732
rect 34532 26450 34560 26726
rect 34520 26444 34572 26450
rect 34520 26386 34572 26392
rect 33508 26308 33560 26314
rect 33508 26250 33560 26256
rect 33520 25838 33548 26250
rect 34532 26042 34560 26386
rect 34520 26036 34572 26042
rect 34520 25978 34572 25984
rect 33508 25832 33560 25838
rect 33508 25774 33560 25780
rect 33520 25362 33548 25774
rect 33508 25356 33560 25362
rect 33508 25298 33560 25304
rect 33520 24614 33548 25298
rect 33508 24608 33560 24614
rect 33506 24576 33508 24585
rect 33560 24576 33562 24585
rect 33506 24511 33562 24520
rect 33874 24576 33930 24585
rect 33874 24511 33930 24520
rect 33888 23633 33916 24511
rect 34518 23760 34574 23769
rect 34518 23695 34574 23704
rect 33874 23624 33930 23633
rect 33874 23559 33930 23568
rect 34532 22794 34560 23695
rect 34440 22766 34560 22794
rect 34060 21888 34112 21894
rect 34060 21830 34112 21836
rect 33874 20632 33930 20641
rect 33874 20567 33930 20576
rect 33888 19310 33916 20567
rect 34072 20369 34100 21830
rect 34058 20360 34114 20369
rect 34058 20295 34114 20304
rect 34440 19990 34468 22766
rect 34428 19984 34480 19990
rect 34428 19926 34480 19932
rect 33968 19916 34020 19922
rect 33968 19858 34020 19864
rect 33980 19446 34008 19858
rect 33968 19440 34020 19446
rect 33968 19382 34020 19388
rect 33508 19304 33560 19310
rect 33506 19272 33508 19281
rect 33784 19304 33836 19310
rect 33560 19272 33562 19281
rect 33784 19246 33836 19252
rect 33876 19304 33928 19310
rect 33876 19246 33928 19252
rect 33506 19207 33562 19216
rect 33796 19174 33824 19246
rect 33784 19168 33836 19174
rect 34428 19168 34480 19174
rect 33784 19110 33836 19116
rect 34058 19136 34114 19145
rect 34428 19110 34480 19116
rect 34058 19071 34114 19080
rect 34072 18902 34100 19071
rect 34060 18896 34112 18902
rect 34060 18838 34112 18844
rect 33508 18828 33560 18834
rect 33508 18770 33560 18776
rect 33784 18828 33836 18834
rect 33784 18770 33836 18776
rect 33520 18358 33548 18770
rect 33508 18352 33560 18358
rect 33508 18294 33560 18300
rect 33520 17678 33548 18294
rect 33796 18086 33824 18770
rect 33784 18080 33836 18086
rect 33784 18022 33836 18028
rect 33508 17672 33560 17678
rect 33508 17614 33560 17620
rect 33968 17672 34020 17678
rect 33968 17614 34020 17620
rect 33782 17504 33838 17513
rect 33782 17439 33838 17448
rect 33796 17134 33824 17439
rect 33784 17128 33836 17134
rect 33704 17088 33784 17116
rect 33600 17060 33652 17066
rect 33600 17002 33652 17008
rect 33612 16794 33640 17002
rect 33600 16788 33652 16794
rect 33600 16730 33652 16736
rect 33704 16658 33732 17088
rect 33784 17070 33836 17076
rect 33692 16652 33744 16658
rect 33692 16594 33744 16600
rect 33508 16040 33560 16046
rect 33508 15982 33560 15988
rect 33520 15910 33548 15982
rect 33508 15904 33560 15910
rect 33508 15846 33560 15852
rect 33520 14958 33548 15846
rect 33704 15706 33732 16594
rect 33876 16584 33928 16590
rect 33876 16526 33928 16532
rect 33888 16250 33916 16526
rect 33876 16244 33928 16250
rect 33876 16186 33928 16192
rect 33692 15700 33744 15706
rect 33692 15642 33744 15648
rect 33508 14952 33560 14958
rect 33508 14894 33560 14900
rect 33520 14278 33548 14894
rect 33600 14884 33652 14890
rect 33600 14826 33652 14832
rect 33612 14550 33640 14826
rect 33600 14544 33652 14550
rect 33600 14486 33652 14492
rect 33508 14272 33560 14278
rect 33508 14214 33560 14220
rect 33612 13870 33640 14486
rect 33876 14408 33928 14414
rect 33876 14350 33928 14356
rect 33600 13864 33652 13870
rect 33600 13806 33652 13812
rect 33612 13530 33640 13806
rect 33888 13530 33916 14350
rect 33600 13524 33652 13530
rect 33600 13466 33652 13472
rect 33876 13524 33928 13530
rect 33876 13466 33928 13472
rect 33414 10296 33470 10305
rect 33414 10231 33470 10240
rect 33980 9081 34008 17614
rect 34336 17332 34388 17338
rect 34336 17274 34388 17280
rect 34060 16584 34112 16590
rect 34058 16552 34060 16561
rect 34112 16552 34114 16561
rect 34058 16487 34114 16496
rect 34348 15502 34376 17274
rect 34440 15570 34468 19110
rect 34518 17912 34574 17921
rect 34518 17847 34574 17856
rect 34532 17746 34560 17847
rect 34520 17740 34572 17746
rect 34520 17682 34572 17688
rect 34532 17338 34560 17682
rect 34520 17332 34572 17338
rect 34520 17274 34572 17280
rect 34428 15564 34480 15570
rect 34428 15506 34480 15512
rect 34336 15496 34388 15502
rect 34336 15438 34388 15444
rect 34348 15162 34376 15438
rect 34336 15156 34388 15162
rect 34336 15098 34388 15104
rect 34152 14476 34204 14482
rect 34152 14418 34204 14424
rect 34164 14074 34192 14418
rect 34348 14414 34376 15098
rect 34440 15094 34468 15506
rect 34428 15088 34480 15094
rect 34428 15030 34480 15036
rect 34336 14408 34388 14414
rect 34336 14350 34388 14356
rect 34244 14340 34296 14346
rect 34244 14282 34296 14288
rect 34152 14068 34204 14074
rect 34152 14010 34204 14016
rect 33966 9072 34022 9081
rect 33966 9007 34022 9016
rect 33506 7712 33562 7721
rect 33506 7647 33562 7656
rect 33520 4826 33548 7647
rect 33508 4820 33560 4826
rect 33508 4762 33560 4768
rect 34256 1465 34284 14282
rect 34428 13864 34480 13870
rect 34428 13806 34480 13812
rect 34440 9602 34468 13806
rect 34440 9574 34560 9602
rect 34532 6905 34560 9574
rect 34624 9489 34652 33895
rect 34808 28626 34836 37402
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 35532 36644 35584 36650
rect 35532 36586 35584 36592
rect 35440 36576 35492 36582
rect 35440 36518 35492 36524
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 35346 34776 35402 34785
rect 35346 34711 35402 34720
rect 35360 34105 35388 34711
rect 35452 34241 35480 36518
rect 35544 36038 35572 36586
rect 35532 36032 35584 36038
rect 35532 35974 35584 35980
rect 35438 34232 35494 34241
rect 35438 34167 35494 34176
rect 35346 34096 35402 34105
rect 35346 34031 35402 34040
rect 35544 33946 35572 35974
rect 35360 33918 35572 33946
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 35254 30696 35310 30705
rect 35254 30631 35310 30640
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 35268 30025 35296 30631
rect 35254 30016 35310 30025
rect 35254 29951 35310 29960
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 34796 28620 34848 28626
rect 34796 28562 34848 28568
rect 34808 28218 34836 28562
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 34796 28212 34848 28218
rect 34796 28154 34848 28160
rect 35360 27985 35388 33918
rect 35636 31482 35664 41511
rect 35898 40996 35954 41796
rect 36358 40996 36414 41796
rect 36818 40996 36874 41796
rect 37738 40996 37794 41796
rect 38198 40996 38254 41796
rect 38658 40996 38714 41796
rect 39578 40996 39634 41796
rect 35912 37913 35940 40996
rect 36372 38321 36400 40996
rect 36358 38312 36414 38321
rect 36358 38247 36414 38256
rect 35898 37904 35954 37913
rect 35898 37839 35954 37848
rect 36082 37904 36138 37913
rect 36082 37839 36084 37848
rect 36136 37839 36138 37848
rect 36084 37810 36136 37816
rect 35716 37732 35768 37738
rect 35716 37674 35768 37680
rect 35728 37330 35756 37674
rect 36544 37664 36596 37670
rect 36544 37606 36596 37612
rect 35806 37496 35862 37505
rect 35806 37431 35862 37440
rect 35716 37324 35768 37330
rect 35716 37266 35768 37272
rect 35728 35850 35756 37266
rect 35820 36786 35848 37431
rect 36556 36922 36584 37606
rect 36544 36916 36596 36922
rect 36544 36858 36596 36864
rect 35808 36780 35860 36786
rect 35808 36722 35860 36728
rect 36556 36718 36584 36858
rect 36544 36712 36596 36718
rect 36544 36654 36596 36660
rect 36832 36553 36860 40996
rect 37752 38554 37780 40996
rect 37740 38548 37792 38554
rect 37740 38490 37792 38496
rect 38212 37913 38240 40996
rect 38198 37904 38254 37913
rect 38198 37839 38254 37848
rect 36818 36544 36874 36553
rect 36818 36479 36874 36488
rect 38672 36378 38700 40996
rect 39592 37233 39620 40996
rect 39578 37224 39634 37233
rect 39578 37159 39634 37168
rect 37464 36372 37516 36378
rect 37464 36314 37516 36320
rect 38660 36372 38712 36378
rect 38660 36314 38712 36320
rect 36082 35864 36138 35873
rect 35728 35822 35940 35850
rect 35912 35630 35940 35822
rect 36082 35799 36138 35808
rect 36096 35698 36124 35799
rect 36084 35692 36136 35698
rect 36084 35634 36136 35640
rect 35900 35624 35952 35630
rect 35900 35566 35952 35572
rect 35912 34950 35940 35566
rect 36084 35488 36136 35494
rect 36084 35430 36136 35436
rect 37370 35456 37426 35465
rect 35900 34944 35952 34950
rect 35900 34886 35952 34892
rect 35912 34542 35940 34886
rect 36096 34610 36124 35430
rect 37370 35391 37426 35400
rect 37384 34746 37412 35391
rect 37372 34740 37424 34746
rect 37372 34682 37424 34688
rect 36084 34604 36136 34610
rect 36084 34546 36136 34552
rect 35900 34536 35952 34542
rect 35900 34478 35952 34484
rect 35912 33862 35940 34478
rect 35900 33856 35952 33862
rect 35900 33798 35952 33804
rect 35624 31476 35676 31482
rect 35624 31418 35676 31424
rect 35622 31376 35678 31385
rect 35622 31311 35678 31320
rect 35806 31376 35862 31385
rect 35806 31311 35862 31320
rect 35438 29336 35494 29345
rect 35438 29271 35494 29280
rect 35452 29170 35480 29271
rect 35440 29164 35492 29170
rect 35440 29106 35492 29112
rect 35452 28762 35480 29106
rect 35440 28756 35492 28762
rect 35440 28698 35492 28704
rect 34702 27976 34758 27985
rect 34702 27911 34758 27920
rect 35346 27976 35402 27985
rect 35346 27911 35402 27920
rect 34716 26586 34744 27911
rect 35636 27538 35664 31311
rect 35820 30326 35848 31311
rect 35912 31278 35940 33798
rect 35900 31272 35952 31278
rect 35900 31214 35952 31220
rect 35912 30938 35940 31214
rect 37280 31136 37332 31142
rect 37280 31078 37332 31084
rect 35900 30932 35952 30938
rect 35900 30874 35952 30880
rect 35808 30320 35860 30326
rect 35808 30262 35860 30268
rect 35900 30184 35952 30190
rect 35900 30126 35952 30132
rect 35912 29510 35940 30126
rect 36544 29708 36596 29714
rect 36544 29650 36596 29656
rect 35900 29504 35952 29510
rect 35900 29446 35952 29452
rect 35912 29102 35940 29446
rect 36556 29306 36584 29650
rect 37292 29617 37320 31078
rect 37372 30048 37424 30054
rect 37372 29990 37424 29996
rect 37278 29608 37334 29617
rect 37278 29543 37334 29552
rect 36544 29300 36596 29306
rect 36544 29242 36596 29248
rect 35900 29096 35952 29102
rect 35900 29038 35952 29044
rect 35808 28416 35860 28422
rect 35912 28404 35940 29038
rect 37384 28801 37412 29990
rect 37370 28792 37426 28801
rect 37370 28727 37426 28736
rect 36082 28656 36138 28665
rect 36082 28591 36138 28600
rect 35860 28376 35940 28404
rect 35808 28358 35860 28364
rect 35820 28014 35848 28358
rect 36096 28082 36124 28591
rect 36084 28076 36136 28082
rect 36084 28018 36136 28024
rect 35808 28008 35860 28014
rect 35808 27950 35860 27956
rect 35624 27532 35676 27538
rect 35624 27474 35676 27480
rect 34796 27328 34848 27334
rect 34796 27270 34848 27276
rect 34808 27010 34836 27270
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 34808 26982 34928 27010
rect 34900 26926 34928 26982
rect 34888 26920 34940 26926
rect 34888 26862 34940 26868
rect 34900 26625 34928 26862
rect 34886 26616 34942 26625
rect 34704 26580 34756 26586
rect 34886 26551 34942 26560
rect 35254 26616 35310 26625
rect 35636 26586 35664 27474
rect 35254 26551 35310 26560
rect 35624 26580 35676 26586
rect 34704 26522 34756 26528
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 35268 25401 35296 26551
rect 35624 26522 35676 26528
rect 35820 26246 35848 27950
rect 37372 27872 37424 27878
rect 37372 27814 37424 27820
rect 36084 27600 36136 27606
rect 36084 27542 36136 27548
rect 36266 27568 36322 27577
rect 35992 27464 36044 27470
rect 35992 27406 36044 27412
rect 35808 26240 35860 26246
rect 35808 26182 35860 26188
rect 35820 25838 35848 26182
rect 35808 25832 35860 25838
rect 35808 25774 35860 25780
rect 35820 25498 35848 25774
rect 35808 25492 35860 25498
rect 35808 25434 35860 25440
rect 35254 25392 35310 25401
rect 35254 25327 35310 25336
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 35820 24750 35848 25434
rect 35808 24744 35860 24750
rect 35808 24686 35860 24692
rect 35820 24410 35848 24686
rect 35808 24404 35860 24410
rect 35808 24346 35860 24352
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 35820 23662 35848 24346
rect 35808 23656 35860 23662
rect 35808 23598 35860 23604
rect 35820 23322 35848 23598
rect 35808 23316 35860 23322
rect 35808 23258 35860 23264
rect 34702 23080 34758 23089
rect 34702 23015 34758 23024
rect 34716 21185 34744 23015
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 35820 22574 35848 23258
rect 35808 22568 35860 22574
rect 35346 22536 35402 22545
rect 35808 22510 35860 22516
rect 35346 22471 35402 22480
rect 35256 22092 35308 22098
rect 35256 22034 35308 22040
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 35268 21690 35296 22034
rect 35360 21690 35388 22471
rect 35438 22264 35494 22273
rect 35820 22234 35848 22510
rect 35438 22199 35494 22208
rect 35808 22228 35860 22234
rect 35256 21684 35308 21690
rect 35256 21626 35308 21632
rect 35348 21684 35400 21690
rect 35348 21626 35400 21632
rect 34702 21176 34758 21185
rect 35268 21146 35296 21626
rect 34702 21111 34758 21120
rect 35256 21140 35308 21146
rect 35308 21100 35388 21128
rect 35256 21082 35308 21088
rect 35256 20936 35308 20942
rect 35256 20878 35308 20884
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 35268 20482 35296 20878
rect 35360 20602 35388 21100
rect 35348 20596 35400 20602
rect 35348 20538 35400 20544
rect 35176 20454 35296 20482
rect 35176 20262 35204 20454
rect 35164 20256 35216 20262
rect 35164 20198 35216 20204
rect 35176 19825 35204 20198
rect 35162 19816 35218 19825
rect 35162 19751 35218 19760
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 35072 19168 35124 19174
rect 35072 19110 35124 19116
rect 35084 18873 35112 19110
rect 34794 18864 34850 18873
rect 34794 18799 34850 18808
rect 35070 18864 35126 18873
rect 35070 18799 35126 18808
rect 34808 17746 34836 18799
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 34796 17740 34848 17746
rect 34796 17682 34848 17688
rect 35256 17740 35308 17746
rect 35256 17682 35308 17688
rect 34808 16946 34836 17682
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 34716 16918 34836 16946
rect 34716 16726 34744 16918
rect 35268 16794 35296 17682
rect 35452 17626 35480 22199
rect 35808 22170 35860 22176
rect 35820 21486 35848 22170
rect 35716 21480 35768 21486
rect 35716 21422 35768 21428
rect 35808 21480 35860 21486
rect 35808 21422 35860 21428
rect 35624 19848 35676 19854
rect 35624 19790 35676 19796
rect 35636 19242 35664 19790
rect 35624 19236 35676 19242
rect 35624 19178 35676 19184
rect 35530 17776 35586 17785
rect 35530 17711 35532 17720
rect 35584 17711 35586 17720
rect 35532 17682 35584 17688
rect 35452 17598 35572 17626
rect 35438 17096 35494 17105
rect 35438 17031 35494 17040
rect 34796 16788 34848 16794
rect 34796 16730 34848 16736
rect 35256 16788 35308 16794
rect 35256 16730 35308 16736
rect 34704 16720 34756 16726
rect 34704 16662 34756 16668
rect 34808 15586 34836 16730
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 34888 16040 34940 16046
rect 34886 16008 34888 16017
rect 34940 16008 34942 16017
rect 34886 15943 34942 15952
rect 34716 15570 34836 15586
rect 34716 15564 34848 15570
rect 34716 15558 34796 15564
rect 34716 15162 34744 15558
rect 34796 15506 34848 15512
rect 34796 15428 34848 15434
rect 34796 15370 34848 15376
rect 34704 15156 34756 15162
rect 34704 15098 34756 15104
rect 34610 9480 34666 9489
rect 34610 9415 34666 9424
rect 34702 7576 34758 7585
rect 34702 7511 34758 7520
rect 34518 6896 34574 6905
rect 34518 6831 34574 6840
rect 34610 4992 34666 5001
rect 34610 4927 34666 4936
rect 34058 1456 34114 1465
rect 34058 1391 34114 1400
rect 34242 1456 34298 1465
rect 34624 1442 34652 4927
rect 34242 1391 34298 1400
rect 34532 1414 34652 1442
rect 34716 1442 34744 7511
rect 34808 4185 34836 15370
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 35348 11008 35400 11014
rect 35348 10950 35400 10956
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 35256 10124 35308 10130
rect 35256 10066 35308 10072
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 35268 9654 35296 10066
rect 35360 10062 35388 10950
rect 35348 10056 35400 10062
rect 35348 9998 35400 10004
rect 35256 9648 35308 9654
rect 35070 9616 35126 9625
rect 35070 9551 35072 9560
rect 35124 9551 35126 9560
rect 35254 9616 35256 9625
rect 35308 9616 35310 9625
rect 35360 9586 35388 9998
rect 35254 9551 35310 9560
rect 35348 9580 35400 9586
rect 35072 9522 35124 9528
rect 35348 9522 35400 9528
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 35254 6352 35310 6361
rect 35254 6287 35310 6296
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 34794 4176 34850 4185
rect 34794 4111 34850 4120
rect 35268 3505 35296 6287
rect 35452 5545 35480 17031
rect 35544 13705 35572 17598
rect 35728 14385 35756 21422
rect 35900 19916 35952 19922
rect 35900 19858 35952 19864
rect 35912 19174 35940 19858
rect 35900 19168 35952 19174
rect 35900 19110 35952 19116
rect 35714 14376 35770 14385
rect 35714 14311 35770 14320
rect 35530 13696 35586 13705
rect 35530 13631 35586 13640
rect 35808 12776 35860 12782
rect 35808 12718 35860 12724
rect 35820 12102 35848 12718
rect 35900 12436 35952 12442
rect 35900 12378 35952 12384
rect 35808 12096 35860 12102
rect 35808 12038 35860 12044
rect 35820 11694 35848 12038
rect 35808 11688 35860 11694
rect 35808 11630 35860 11636
rect 35820 11014 35848 11630
rect 35808 11008 35860 11014
rect 35808 10950 35860 10956
rect 35438 5536 35494 5545
rect 35438 5471 35494 5480
rect 35254 3496 35310 3505
rect 35254 3431 35310 3440
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 35820 2990 35848 3334
rect 35808 2984 35860 2990
rect 35808 2926 35860 2932
rect 35624 2848 35676 2854
rect 35622 2816 35624 2825
rect 35676 2816 35678 2825
rect 35622 2751 35678 2760
rect 35162 2680 35218 2689
rect 35162 2615 35164 2624
rect 35216 2615 35218 2624
rect 35164 2586 35216 2592
rect 35176 2446 35204 2586
rect 35820 2514 35848 2926
rect 35808 2508 35860 2514
rect 35808 2450 35860 2456
rect 35164 2440 35216 2446
rect 35164 2382 35216 2388
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 34716 1414 35020 1442
rect 34072 800 34100 1391
rect 34532 800 34560 1414
rect 34992 800 35020 1414
rect 35912 800 35940 12378
rect 36004 4049 36032 27406
rect 36096 26586 36124 27542
rect 36266 27503 36322 27512
rect 37188 27532 37240 27538
rect 36280 27130 36308 27503
rect 37188 27474 37240 27480
rect 36268 27124 36320 27130
rect 36268 27066 36320 27072
rect 36176 26920 36228 26926
rect 36176 26862 36228 26868
rect 36084 26580 36136 26586
rect 36084 26522 36136 26528
rect 36084 25832 36136 25838
rect 36084 25774 36136 25780
rect 36096 25265 36124 25774
rect 36082 25256 36138 25265
rect 36082 25191 36138 25200
rect 36084 24608 36136 24614
rect 36084 24550 36136 24556
rect 36096 23730 36124 24550
rect 36084 23724 36136 23730
rect 36084 23666 36136 23672
rect 36084 22568 36136 22574
rect 36082 22536 36084 22545
rect 36136 22536 36138 22545
rect 36082 22471 36138 22480
rect 36084 19848 36136 19854
rect 36084 19790 36136 19796
rect 36096 19378 36124 19790
rect 36084 19372 36136 19378
rect 36084 19314 36136 19320
rect 36188 12442 36216 26862
rect 37200 26790 37228 27474
rect 37188 26784 37240 26790
rect 37240 26732 37320 26738
rect 37188 26726 37320 26732
rect 37200 26710 37320 26726
rect 37292 26042 37320 26710
rect 37280 26036 37332 26042
rect 37280 25978 37332 25984
rect 37188 24812 37240 24818
rect 37384 24800 37412 27814
rect 37240 24772 37412 24800
rect 37188 24754 37240 24760
rect 37372 23520 37424 23526
rect 37372 23462 37424 23468
rect 37384 23225 37412 23462
rect 37370 23216 37426 23225
rect 37370 23151 37426 23160
rect 37278 22672 37334 22681
rect 37278 22607 37280 22616
rect 37332 22607 37334 22616
rect 37280 22578 37332 22584
rect 36266 21992 36322 22001
rect 36266 21927 36322 21936
rect 36280 21146 36308 21927
rect 37476 21321 37504 36314
rect 37462 21312 37518 21321
rect 37462 21247 37518 21256
rect 36268 21140 36320 21146
rect 36268 21082 36320 21088
rect 37280 12844 37332 12850
rect 37280 12786 37332 12792
rect 37188 12776 37240 12782
rect 37292 12753 37320 12786
rect 37188 12718 37240 12724
rect 37278 12744 37334 12753
rect 37200 12594 37228 12718
rect 37278 12679 37334 12688
rect 37200 12566 37320 12594
rect 36176 12436 36228 12442
rect 36176 12378 36228 12384
rect 37292 11898 37320 12566
rect 37280 11892 37332 11898
rect 37280 11834 37332 11840
rect 36084 11688 36136 11694
rect 36084 11630 36136 11636
rect 36096 10266 36124 11630
rect 36084 10260 36136 10266
rect 36084 10202 36136 10208
rect 37370 5536 37426 5545
rect 37370 5471 37426 5480
rect 35990 4040 36046 4049
rect 35990 3975 36046 3984
rect 37384 3194 37412 5471
rect 37738 4040 37794 4049
rect 37738 3975 37794 3984
rect 37372 3188 37424 3194
rect 37372 3130 37424 3136
rect 36360 2304 36412 2310
rect 36360 2246 36412 2252
rect 36372 800 36400 2246
rect 37280 2100 37332 2106
rect 37280 2042 37332 2048
rect 37292 800 37320 2042
rect 37752 800 37780 3975
rect 39578 3904 39634 3913
rect 39578 3839 39634 3848
rect 39118 3088 39174 3097
rect 39118 3023 39174 3032
rect 38198 2544 38254 2553
rect 38198 2479 38254 2488
rect 38212 800 38240 2479
rect 39132 800 39160 3023
rect 39592 800 39620 3839
rect 33230 96 33286 105
rect 33230 31 33286 40
rect 34058 0 34114 800
rect 34518 0 34574 800
rect 34978 0 35034 800
rect 35898 0 35954 800
rect 36358 0 36414 800
rect 37278 0 37334 800
rect 37738 0 37794 800
rect 38198 0 38254 800
rect 39118 0 39174 800
rect 39578 0 39634 800
<< via2 >>
rect 3238 41520 3294 41576
rect 938 38528 994 38584
rect 1398 37712 1454 37768
rect 18 35128 74 35184
rect 2962 40840 3018 40896
rect 35622 41520 35678 41576
rect 3422 40196 3424 40216
rect 3424 40196 3476 40216
rect 3476 40196 3478 40216
rect 3422 40160 3478 40196
rect 3422 38664 3478 38720
rect 2778 38120 2834 38176
rect 1766 37304 1822 37360
rect 2318 37168 2374 37224
rect 1582 34176 1638 34232
rect 1398 29280 1454 29336
rect 1582 23860 1638 23896
rect 1582 23840 1584 23860
rect 1584 23840 1636 23860
rect 1636 23840 1638 23860
rect 1674 21120 1730 21176
rect 3422 34040 3478 34096
rect 3422 33224 3478 33280
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4246 39194
rect 4246 39142 4276 39194
rect 4300 39142 4310 39194
rect 4310 39142 4356 39194
rect 4380 39142 4426 39194
rect 4426 39142 4436 39194
rect 4460 39142 4490 39194
rect 4490 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4066 36760 4122 36816
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4066 35400 4122 35456
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 6182 33360 6238 33416
rect 5998 32816 6054 32872
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 2962 28464 3018 28520
rect 3422 30096 3478 30152
rect 3146 28600 3202 28656
rect 2778 27920 2834 27976
rect 2778 26560 2834 26616
rect 3054 27512 3110 27568
rect 3054 27412 3056 27432
rect 3056 27412 3108 27432
rect 3108 27412 3110 27432
rect 3054 27376 3110 27412
rect 2962 25200 3018 25256
rect 1950 23160 2006 23216
rect 2410 21800 2466 21856
rect 2594 20440 2650 20496
rect 1766 19080 1822 19136
rect 1950 17756 1952 17776
rect 1952 17756 2004 17776
rect 2004 17756 2006 17776
rect 1950 17720 2006 17756
rect 1674 16360 1730 16416
rect 1582 13776 1638 13832
rect 1582 12980 1638 13016
rect 1582 12960 1584 12980
rect 1584 12960 1636 12980
rect 1636 12960 1638 12980
rect 18 5072 74 5128
rect 938 3712 994 3768
rect 478 3032 534 3088
rect 1490 11056 1546 11112
rect 1582 10240 1638 10296
rect 2870 11056 2926 11112
rect 2410 9560 2466 9616
rect 1490 6976 1546 7032
rect 1858 6704 1914 6760
rect 1766 6160 1822 6216
rect 2410 8880 2466 8936
rect 2686 8200 2742 8256
rect 2778 7248 2834 7304
rect 3054 23588 3110 23624
rect 3054 23568 3056 23588
rect 3056 23568 3108 23588
rect 3108 23568 3110 23588
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4066 30932 4122 30968
rect 4066 30912 4068 30932
rect 4068 30912 4120 30932
rect 4120 30912 4122 30932
rect 4066 30504 4122 30560
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4986 30912 5042 30968
rect 4894 30232 4950 30288
rect 4066 29688 4122 29744
rect 3422 23724 3478 23760
rect 3422 23704 3424 23724
rect 3424 23704 3476 23724
rect 3476 23704 3478 23724
rect 3882 26968 3938 27024
rect 3790 24112 3846 24168
rect 3882 23432 3938 23488
rect 3882 23316 3938 23352
rect 3882 23296 3884 23316
rect 3884 23296 3936 23316
rect 3936 23296 3938 23316
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 4710 28872 4766 28928
rect 4710 26968 4766 27024
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 4066 25880 4122 25936
rect 4526 25472 4582 25528
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 3146 19352 3202 19408
rect 3054 18672 3110 18728
rect 3698 22616 3754 22672
rect 3514 21528 3570 21584
rect 3422 19372 3478 19408
rect 3422 19352 3424 19372
rect 3424 19352 3476 19372
rect 3476 19352 3478 19372
rect 3514 19080 3570 19136
rect 3514 15000 3570 15056
rect 3422 14456 3478 14512
rect 3146 12300 3202 12336
rect 3146 12280 3148 12300
rect 3148 12280 3200 12300
rect 3200 12280 3202 12300
rect 3974 23024 4030 23080
rect 4710 24928 4766 24984
rect 5078 26560 5134 26616
rect 4986 26308 5042 26344
rect 4986 26288 4988 26308
rect 4988 26288 5040 26308
rect 5040 26288 5042 26308
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4802 22208 4858 22264
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 3882 21140 3938 21176
rect 3882 21120 3884 21140
rect 3884 21120 3936 21140
rect 3936 21120 3938 21140
rect 3974 20032 4030 20088
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 4618 20440 4674 20496
rect 3882 19216 3938 19272
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4066 19352 4122 19408
rect 4434 18692 4490 18728
rect 4434 18672 4436 18692
rect 4436 18672 4488 18692
rect 4488 18672 4490 18692
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4066 18400 4122 18456
rect 4618 17876 4674 17912
rect 4618 17856 4620 17876
rect 4620 17856 4672 17876
rect 4672 17856 4674 17876
rect 4526 17584 4582 17640
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 3974 16904 4030 16960
rect 3882 16496 3938 16552
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 3882 15408 3938 15464
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4802 18944 4858 19000
rect 4894 18808 4950 18864
rect 5814 26424 5870 26480
rect 5722 26152 5778 26208
rect 5170 22344 5226 22400
rect 5078 21936 5134 21992
rect 5262 21936 5318 21992
rect 5262 20712 5318 20768
rect 5262 19932 5264 19952
rect 5264 19932 5316 19952
rect 5316 19932 5318 19952
rect 5262 19896 5318 19932
rect 3882 14864 3938 14920
rect 3974 14592 4030 14648
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4618 12044 4620 12064
rect 4620 12044 4672 12064
rect 4672 12044 4674 12064
rect 4618 12008 4674 12044
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 3790 11600 3846 11656
rect 5262 18420 5318 18456
rect 5262 18400 5264 18420
rect 5264 18400 5316 18420
rect 5316 18400 5318 18420
rect 5630 19896 5686 19952
rect 6366 30096 6422 30152
rect 6274 25880 6330 25936
rect 6366 24112 6422 24168
rect 5446 16632 5502 16688
rect 4894 14340 4950 14376
rect 4894 14320 4896 14340
rect 4896 14320 4948 14340
rect 4948 14320 4950 14340
rect 5446 15136 5502 15192
rect 5262 14728 5318 14784
rect 5354 14612 5410 14648
rect 5354 14592 5356 14612
rect 5356 14592 5408 14612
rect 5408 14592 5410 14612
rect 6090 20596 6146 20632
rect 6090 20576 6092 20596
rect 6092 20576 6144 20596
rect 6144 20576 6146 20596
rect 6182 20052 6238 20088
rect 6182 20032 6184 20052
rect 6184 20032 6236 20052
rect 6236 20032 6238 20052
rect 5906 17740 5962 17776
rect 5906 17720 5908 17740
rect 5908 17720 5960 17740
rect 5960 17720 5962 17740
rect 5814 14592 5870 14648
rect 5722 13504 5778 13560
rect 5262 13368 5318 13424
rect 4986 13232 5042 13288
rect 4894 12960 4950 13016
rect 5722 13096 5778 13152
rect 6274 17196 6330 17232
rect 6274 17176 6276 17196
rect 6276 17176 6328 17196
rect 6328 17176 6330 17196
rect 6090 15544 6146 15600
rect 5998 12280 6054 12336
rect 6642 23024 6698 23080
rect 6826 37168 6882 37224
rect 6826 36624 6882 36680
rect 6918 33496 6974 33552
rect 7010 33360 7066 33416
rect 7838 38392 7894 38448
rect 7378 37440 7434 37496
rect 6918 33224 6974 33280
rect 7102 33224 7158 33280
rect 8390 35672 8446 35728
rect 10598 38392 10654 38448
rect 9954 37984 10010 38040
rect 9678 37440 9734 37496
rect 9218 37304 9274 37360
rect 10414 37304 10470 37360
rect 11518 37848 11574 37904
rect 13358 38412 13414 38448
rect 13358 38392 13360 38412
rect 13360 38392 13412 38412
rect 13412 38392 13414 38412
rect 13634 37712 13690 37768
rect 10966 36488 11022 36544
rect 9034 34448 9090 34504
rect 7930 31864 7986 31920
rect 7746 31356 7748 31376
rect 7748 31356 7800 31376
rect 7800 31356 7802 31376
rect 7746 31320 7802 31356
rect 6918 30252 6974 30288
rect 6918 30232 6920 30252
rect 6920 30232 6972 30252
rect 6972 30232 6974 30252
rect 7378 30232 7434 30288
rect 7010 26696 7066 26752
rect 7194 26152 7250 26208
rect 7194 25744 7250 25800
rect 7010 24112 7066 24168
rect 7194 23432 7250 23488
rect 7194 22480 7250 22536
rect 7102 22208 7158 22264
rect 7562 24384 7618 24440
rect 7562 23724 7618 23760
rect 7562 23704 7564 23724
rect 7564 23704 7616 23724
rect 7616 23704 7618 23724
rect 7378 20712 7434 20768
rect 7654 23296 7710 23352
rect 7562 22380 7564 22400
rect 7564 22380 7616 22400
rect 7616 22380 7618 22400
rect 7562 22344 7618 22380
rect 8574 30096 8630 30152
rect 8022 29960 8078 30016
rect 8666 28620 8722 28656
rect 8666 28600 8668 28620
rect 8668 28600 8720 28620
rect 8720 28600 8722 28620
rect 10874 32136 10930 32192
rect 9586 30660 9642 30696
rect 9586 30640 9588 30660
rect 9588 30640 9640 30660
rect 9640 30640 9642 30660
rect 9954 30368 10010 30424
rect 9678 30268 9680 30288
rect 9680 30268 9732 30288
rect 9732 30268 9734 30288
rect 9678 30232 9734 30268
rect 8114 27004 8116 27024
rect 8116 27004 8168 27024
rect 8168 27004 8170 27024
rect 8114 26968 8170 27004
rect 9126 26324 9128 26344
rect 9128 26324 9180 26344
rect 9180 26324 9182 26344
rect 9126 26288 9182 26324
rect 8390 26016 8446 26072
rect 8206 25644 8208 25664
rect 8208 25644 8260 25664
rect 8260 25644 8262 25664
rect 8206 25608 8262 25644
rect 7378 20032 7434 20088
rect 7194 19236 7250 19272
rect 7194 19216 7196 19236
rect 7196 19216 7248 19236
rect 7248 19216 7250 19236
rect 6826 16904 6882 16960
rect 6734 15952 6790 16008
rect 7194 18692 7250 18728
rect 7194 18672 7196 18692
rect 7196 18672 7248 18692
rect 7248 18672 7250 18692
rect 7654 19080 7710 19136
rect 7930 21392 7986 21448
rect 7838 21120 7894 21176
rect 8022 21120 8078 21176
rect 7930 19080 7986 19136
rect 7930 18828 7986 18864
rect 7930 18808 7932 18828
rect 7932 18808 7984 18828
rect 7984 18808 7986 18828
rect 7746 18400 7802 18456
rect 7286 17060 7342 17096
rect 7286 17040 7288 17060
rect 7288 17040 7340 17060
rect 7340 17040 7342 17060
rect 7470 16668 7472 16688
rect 7472 16668 7524 16688
rect 7524 16668 7526 16688
rect 6826 14592 6882 14648
rect 6734 14184 6790 14240
rect 7102 15564 7158 15600
rect 7102 15544 7104 15564
rect 7104 15544 7156 15564
rect 7156 15544 7158 15564
rect 7470 16632 7526 16668
rect 7194 15272 7250 15328
rect 6918 12844 6974 12880
rect 6918 12824 6920 12844
rect 6920 12824 6972 12844
rect 6972 12824 6974 12844
rect 6826 12144 6882 12200
rect 6182 11464 6238 11520
rect 3790 9424 3846 9480
rect 3606 8336 3662 8392
rect 3514 7928 3570 7984
rect 3790 7112 3846 7168
rect 3514 4120 3570 4176
rect 3146 3476 3148 3496
rect 3148 3476 3200 3496
rect 3200 3476 3202 3496
rect 3146 3440 3202 3476
rect 3790 2760 3846 2816
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 6642 10784 6698 10840
rect 5538 10124 5594 10160
rect 5538 10104 5540 10124
rect 5540 10104 5592 10124
rect 5592 10104 5594 10124
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 6182 9288 6238 9344
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 5538 7656 5594 7712
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4802 7520 4858 7576
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4066 5480 4122 5536
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4618 4936 4674 4992
rect 4066 4528 4122 4584
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 3974 3576 4030 3632
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4342 2488 4398 2544
rect 4066 2352 4122 2408
rect 3882 1536 3938 1592
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 4066 1400 4122 1456
rect 5998 5888 6054 5944
rect 7470 14900 7472 14920
rect 7472 14900 7524 14920
rect 7524 14900 7526 14920
rect 7470 14864 7526 14900
rect 7378 14728 7434 14784
rect 8206 20440 8262 20496
rect 7930 17856 7986 17912
rect 8022 17584 8078 17640
rect 8298 17992 8354 18048
rect 8298 17856 8354 17912
rect 8942 24928 8998 24984
rect 8850 24268 8906 24304
rect 8850 24248 8852 24268
rect 8852 24248 8904 24268
rect 8904 24248 8906 24268
rect 8942 24112 8998 24168
rect 9310 24792 9366 24848
rect 8942 23588 8998 23624
rect 8942 23568 8944 23588
rect 8944 23568 8996 23588
rect 8996 23568 8998 23588
rect 9126 23568 9182 23624
rect 8942 22752 8998 22808
rect 9218 22616 9274 22672
rect 9218 22344 9274 22400
rect 9218 22208 9274 22264
rect 8574 21836 8576 21856
rect 8576 21836 8628 21856
rect 8628 21836 8630 21856
rect 8574 21800 8630 21836
rect 8666 21528 8722 21584
rect 8666 20576 8722 20632
rect 9218 21936 9274 21992
rect 8850 21292 8852 21312
rect 8852 21292 8904 21312
rect 8904 21292 8906 21312
rect 8850 21256 8906 21292
rect 9770 27104 9826 27160
rect 9586 26288 9642 26344
rect 10322 30232 10378 30288
rect 10414 28872 10470 28928
rect 10138 26732 10140 26752
rect 10140 26732 10192 26752
rect 10192 26732 10194 26752
rect 10138 26696 10194 26732
rect 10322 27920 10378 27976
rect 10046 25644 10048 25664
rect 10048 25644 10100 25664
rect 10100 25644 10102 25664
rect 10046 25608 10102 25644
rect 9586 22072 9642 22128
rect 8850 19488 8906 19544
rect 7930 16496 7986 16552
rect 8022 15136 8078 15192
rect 7838 15020 7894 15056
rect 7838 15000 7840 15020
rect 7840 15000 7892 15020
rect 7892 15000 7894 15020
rect 7654 14456 7710 14512
rect 8390 17620 8392 17640
rect 8392 17620 8444 17640
rect 8444 17620 8446 17640
rect 8390 17584 8446 17620
rect 8666 17856 8722 17912
rect 9218 18536 9274 18592
rect 8850 17176 8906 17232
rect 7562 14184 7618 14240
rect 8482 13640 8538 13696
rect 8206 12300 8262 12336
rect 8206 12280 8208 12300
rect 8208 12280 8260 12300
rect 8260 12280 8262 12300
rect 7470 11872 7526 11928
rect 8482 13368 8538 13424
rect 10230 26424 10286 26480
rect 9954 22072 10010 22128
rect 9954 21392 10010 21448
rect 10138 21256 10194 21312
rect 9862 19080 9918 19136
rect 9678 17992 9734 18048
rect 9586 17484 9588 17504
rect 9588 17484 9640 17504
rect 9640 17484 9642 17504
rect 9586 17448 9642 17484
rect 9678 16632 9734 16688
rect 9402 14764 9404 14784
rect 9404 14764 9456 14784
rect 9456 14764 9458 14784
rect 9402 14728 9458 14764
rect 9310 12960 9366 13016
rect 8666 12144 8722 12200
rect 8390 12008 8446 12064
rect 8206 11212 8262 11248
rect 8206 11192 8208 11212
rect 8208 11192 8260 11212
rect 8260 11192 8262 11212
rect 7930 11092 7932 11112
rect 7932 11092 7984 11112
rect 7984 11092 7986 11112
rect 7930 11056 7986 11092
rect 8666 10920 8722 10976
rect 8482 10804 8538 10840
rect 8482 10784 8484 10804
rect 8484 10784 8536 10804
rect 8536 10784 8538 10804
rect 7286 9444 7342 9480
rect 7286 9424 7288 9444
rect 7288 9424 7340 9444
rect 7340 9424 7342 9444
rect 6274 8900 6330 8936
rect 6274 8880 6276 8900
rect 6276 8880 6328 8900
rect 6328 8880 6330 8900
rect 8206 8472 8262 8528
rect 9586 12960 9642 13016
rect 10230 16108 10286 16144
rect 10230 16088 10232 16108
rect 10232 16088 10284 16108
rect 10284 16088 10286 16108
rect 10046 14864 10102 14920
rect 9862 13132 9864 13152
rect 9864 13132 9916 13152
rect 9916 13132 9918 13152
rect 9862 13096 9918 13132
rect 9494 10784 9550 10840
rect 9402 10648 9458 10704
rect 9310 10240 9366 10296
rect 8758 9988 8814 10024
rect 8758 9968 8760 9988
rect 8760 9968 8812 9988
rect 8812 9968 8814 9988
rect 9494 9460 9496 9480
rect 9496 9460 9548 9480
rect 9548 9460 9550 9480
rect 9494 9424 9550 9460
rect 9586 8608 9642 8664
rect 9034 8472 9090 8528
rect 10230 14476 10286 14512
rect 10230 14456 10232 14476
rect 10232 14456 10284 14476
rect 10284 14456 10286 14476
rect 10322 12860 10324 12880
rect 10324 12860 10376 12880
rect 10376 12860 10378 12880
rect 10322 12824 10378 12860
rect 10138 9288 10194 9344
rect 10138 8472 10194 8528
rect 10046 8336 10102 8392
rect 6918 5480 6974 5536
rect 7378 4664 7434 4720
rect 8482 2488 8538 2544
rect 8298 1572 8300 1592
rect 8300 1572 8352 1592
rect 8352 1572 8354 1592
rect 8298 1536 8354 1572
rect 10230 7148 10232 7168
rect 10232 7148 10284 7168
rect 10284 7148 10286 7168
rect 10230 7112 10286 7148
rect 10138 5480 10194 5536
rect 11058 32000 11114 32056
rect 11242 30368 11298 30424
rect 11518 28600 11574 28656
rect 10598 26560 10654 26616
rect 11518 27784 11574 27840
rect 11058 27532 11114 27568
rect 11058 27512 11060 27532
rect 11060 27512 11112 27532
rect 11112 27512 11114 27532
rect 11702 27512 11758 27568
rect 10506 25200 10562 25256
rect 10506 24928 10562 24984
rect 10966 25780 10968 25800
rect 10968 25780 11020 25800
rect 11020 25780 11022 25800
rect 10966 25744 11022 25780
rect 11058 25472 11114 25528
rect 11058 24248 11114 24304
rect 11610 26288 11666 26344
rect 10782 22616 10838 22672
rect 10506 21020 10508 21040
rect 10508 21020 10560 21040
rect 10560 21020 10562 21040
rect 10506 20984 10562 21020
rect 11242 21664 11298 21720
rect 10782 19352 10838 19408
rect 10690 18944 10746 19000
rect 10506 17176 10562 17232
rect 10506 16496 10562 16552
rect 10506 13096 10562 13152
rect 10506 11736 10562 11792
rect 11794 26324 11796 26344
rect 11796 26324 11848 26344
rect 11848 26324 11850 26344
rect 11794 26288 11850 26324
rect 11794 26036 11850 26072
rect 11794 26016 11796 26036
rect 11796 26016 11848 26036
rect 11848 26016 11850 26036
rect 11794 25880 11850 25936
rect 11886 25336 11942 25392
rect 11702 21936 11758 21992
rect 11334 20576 11390 20632
rect 11886 20576 11942 20632
rect 11610 19932 11612 19952
rect 11612 19932 11664 19952
rect 11664 19932 11666 19952
rect 11610 19896 11666 19932
rect 11794 19896 11850 19952
rect 11334 18284 11390 18320
rect 10782 18148 10838 18184
rect 10782 18128 10784 18148
rect 10784 18128 10836 18148
rect 10836 18128 10838 18148
rect 11334 18264 11336 18284
rect 11336 18264 11388 18284
rect 11388 18264 11390 18284
rect 10690 17584 10746 17640
rect 10782 16768 10838 16824
rect 11150 16904 11206 16960
rect 10966 15680 11022 15736
rect 11702 18672 11758 18728
rect 11518 17876 11574 17912
rect 11518 17856 11520 17876
rect 11520 17856 11572 17876
rect 11572 17856 11574 17876
rect 11426 16360 11482 16416
rect 11058 15156 11114 15192
rect 11058 15136 11060 15156
rect 11060 15136 11112 15156
rect 11112 15136 11114 15156
rect 10966 14864 11022 14920
rect 10782 14184 10838 14240
rect 10506 2932 10508 2952
rect 10508 2932 10560 2952
rect 10560 2932 10562 2952
rect 10506 2896 10562 2932
rect 10322 2508 10378 2544
rect 10322 2488 10324 2508
rect 10324 2488 10376 2508
rect 10376 2488 10378 2508
rect 10782 11092 10784 11112
rect 10784 11092 10836 11112
rect 10836 11092 10838 11112
rect 10782 11056 10838 11092
rect 11242 15036 11244 15056
rect 11244 15036 11296 15056
rect 11296 15036 11298 15056
rect 11242 15000 11298 15036
rect 11610 15680 11666 15736
rect 11610 15408 11666 15464
rect 10966 13504 11022 13560
rect 11242 13232 11298 13288
rect 11058 11212 11114 11248
rect 11058 11192 11060 11212
rect 11060 11192 11112 11212
rect 11112 11192 11114 11212
rect 11334 10412 11336 10432
rect 11336 10412 11388 10432
rect 11388 10412 11390 10432
rect 11334 10376 11390 10412
rect 12622 32852 12624 32872
rect 12624 32852 12676 32872
rect 12676 32852 12678 32872
rect 12622 32816 12678 32852
rect 13358 32172 13360 32192
rect 13360 32172 13412 32192
rect 13412 32172 13414 32192
rect 12622 27784 12678 27840
rect 12254 24556 12256 24576
rect 12256 24556 12308 24576
rect 12308 24556 12310 24576
rect 12254 24520 12310 24556
rect 12438 22616 12494 22672
rect 13358 32136 13414 32172
rect 12990 31184 13046 31240
rect 13358 29960 13414 30016
rect 12990 25336 13046 25392
rect 13174 24828 13176 24848
rect 13176 24828 13228 24848
rect 13228 24828 13230 24848
rect 13174 24792 13230 24828
rect 13726 35944 13782 36000
rect 14278 35944 14334 36000
rect 13634 34992 13690 35048
rect 14094 33224 14150 33280
rect 13910 30368 13966 30424
rect 13634 29552 13690 29608
rect 14738 36896 14794 36952
rect 14554 34468 14610 34504
rect 14554 34448 14556 34468
rect 14556 34448 14608 34468
rect 14608 34448 14610 34468
rect 14462 33496 14518 33552
rect 14370 32544 14426 32600
rect 14186 30232 14242 30288
rect 14094 29280 14150 29336
rect 14094 29044 14096 29064
rect 14096 29044 14148 29064
rect 14148 29044 14150 29064
rect 13726 28600 13782 28656
rect 13450 27240 13506 27296
rect 14094 29008 14150 29044
rect 14646 33360 14702 33416
rect 14278 27104 14334 27160
rect 13174 24384 13230 24440
rect 12622 21392 12678 21448
rect 12254 20032 12310 20088
rect 12622 19252 12624 19272
rect 12624 19252 12676 19272
rect 12676 19252 12678 19272
rect 12622 19216 12678 19252
rect 12898 19252 12900 19272
rect 12900 19252 12952 19272
rect 12952 19252 12954 19272
rect 12898 19216 12954 19252
rect 12346 17040 12402 17096
rect 12806 17720 12862 17776
rect 12714 17448 12770 17504
rect 12898 17448 12954 17504
rect 12714 17040 12770 17096
rect 12162 16360 12218 16416
rect 12622 16088 12678 16144
rect 12162 15408 12218 15464
rect 12530 14320 12586 14376
rect 12254 13368 12310 13424
rect 12070 12688 12126 12744
rect 10874 9968 10930 10024
rect 11426 9424 11482 9480
rect 10874 6840 10930 6896
rect 11242 7112 11298 7168
rect 11150 4256 11206 4312
rect 13266 21836 13268 21856
rect 13268 21836 13320 21856
rect 13320 21836 13322 21856
rect 13266 21800 13322 21836
rect 14370 26968 14426 27024
rect 14094 24520 14150 24576
rect 13910 24268 13966 24304
rect 13910 24248 13912 24268
rect 13912 24248 13964 24268
rect 13964 24248 13966 24268
rect 13358 20884 13360 20904
rect 13360 20884 13412 20904
rect 13412 20884 13414 20904
rect 13358 20848 13414 20884
rect 13266 17992 13322 18048
rect 13082 16632 13138 16688
rect 14094 22344 14150 22400
rect 14094 21292 14096 21312
rect 14096 21292 14148 21312
rect 14148 21292 14150 21312
rect 14094 21256 14150 21292
rect 12990 15544 13046 15600
rect 12806 15408 12862 15464
rect 12990 15272 13046 15328
rect 12714 13640 12770 13696
rect 12622 12960 12678 13016
rect 12714 12824 12770 12880
rect 12622 12552 12678 12608
rect 12438 11056 12494 11112
rect 12714 10784 12770 10840
rect 12898 12552 12954 12608
rect 13266 14048 13322 14104
rect 13082 12552 13138 12608
rect 13450 12416 13506 12472
rect 12990 11056 13046 11112
rect 12898 8880 12954 8936
rect 12162 8744 12218 8800
rect 11518 6568 11574 6624
rect 13266 8880 13322 8936
rect 11978 4392 12034 4448
rect 13634 16768 13690 16824
rect 13818 15000 13874 15056
rect 14186 18944 14242 19000
rect 14002 15272 14058 15328
rect 13634 14320 13690 14376
rect 13726 13776 13782 13832
rect 13726 12552 13782 12608
rect 13634 11212 13690 11248
rect 14002 12552 14058 12608
rect 14094 12316 14096 12336
rect 14096 12316 14148 12336
rect 14148 12316 14150 12336
rect 14094 12280 14150 12316
rect 14370 15136 14426 15192
rect 14370 13640 14426 13696
rect 14278 11736 14334 11792
rect 13634 11192 13636 11212
rect 13636 11192 13688 11212
rect 13688 11192 13690 11212
rect 15566 37848 15622 37904
rect 15658 37304 15714 37360
rect 15750 37168 15806 37224
rect 15290 32816 15346 32872
rect 15382 31184 15438 31240
rect 15658 32852 15660 32872
rect 15660 32852 15712 32872
rect 15712 32852 15714 32872
rect 15658 32816 15714 32852
rect 15750 31900 15752 31920
rect 15752 31900 15804 31920
rect 15804 31900 15806 31920
rect 15750 31864 15806 31900
rect 15474 30912 15530 30968
rect 15198 29552 15254 29608
rect 15014 28056 15070 28112
rect 15474 26988 15530 27024
rect 15474 26968 15476 26988
rect 15476 26968 15528 26988
rect 15528 26968 15530 26988
rect 14646 24112 14702 24168
rect 14738 23568 14794 23624
rect 14646 22092 14702 22128
rect 14646 22072 14648 22092
rect 14648 22072 14700 22092
rect 14700 22072 14702 22092
rect 14646 21020 14648 21040
rect 14648 21020 14700 21040
rect 14700 21020 14702 21040
rect 14646 20984 14702 21020
rect 15290 24812 15346 24848
rect 15290 24792 15292 24812
rect 15292 24792 15344 24812
rect 15344 24792 15346 24812
rect 15382 23840 15438 23896
rect 15290 23024 15346 23080
rect 14646 19352 14702 19408
rect 14646 19080 14702 19136
rect 14738 17992 14794 18048
rect 14738 17620 14740 17640
rect 14740 17620 14792 17640
rect 14792 17620 14794 17640
rect 14738 17584 14794 17620
rect 15198 21256 15254 21312
rect 14554 17076 14556 17096
rect 14556 17076 14608 17096
rect 14608 17076 14610 17096
rect 14554 17040 14610 17076
rect 14554 14320 14610 14376
rect 14554 14048 14610 14104
rect 14554 12552 14610 12608
rect 14738 15308 14740 15328
rect 14740 15308 14792 15328
rect 14792 15308 14794 15328
rect 14738 15272 14794 15308
rect 14738 15000 14794 15056
rect 14738 14456 14794 14512
rect 14922 17040 14978 17096
rect 15474 19116 15476 19136
rect 15476 19116 15528 19136
rect 15528 19116 15530 19136
rect 15474 19080 15530 19116
rect 15198 18264 15254 18320
rect 15198 15680 15254 15736
rect 15014 14728 15070 14784
rect 16210 36624 16266 36680
rect 16302 36352 16358 36408
rect 17314 37748 17316 37768
rect 17316 37748 17368 37768
rect 17368 37748 17370 37768
rect 17314 37712 17370 37748
rect 15750 24792 15806 24848
rect 15566 17856 15622 17912
rect 15658 16496 15714 16552
rect 15198 13096 15254 13152
rect 15106 12844 15162 12880
rect 15106 12824 15108 12844
rect 15108 12824 15160 12844
rect 15160 12824 15162 12844
rect 15198 10240 15254 10296
rect 15014 9016 15070 9072
rect 14370 8780 14372 8800
rect 14372 8780 14424 8800
rect 14424 8780 14426 8800
rect 14370 8744 14426 8780
rect 15382 14068 15438 14104
rect 15382 14048 15384 14068
rect 15384 14048 15436 14068
rect 15436 14048 15438 14068
rect 15566 14184 15622 14240
rect 15382 11636 15384 11656
rect 15384 11636 15436 11656
rect 15436 11636 15438 11656
rect 15382 11600 15438 11636
rect 14646 8356 14702 8392
rect 14646 8336 14648 8356
rect 14648 8336 14700 8356
rect 14700 8336 14702 8356
rect 16394 31356 16396 31376
rect 16396 31356 16448 31376
rect 16448 31356 16450 31376
rect 16394 31320 16450 31356
rect 16394 29960 16450 30016
rect 16394 28464 16450 28520
rect 16118 25880 16174 25936
rect 16118 24112 16174 24168
rect 16302 23060 16304 23080
rect 16304 23060 16356 23080
rect 16356 23060 16358 23080
rect 16302 23024 16358 23060
rect 16118 22480 16174 22536
rect 16026 20440 16082 20496
rect 15842 17176 15898 17232
rect 15934 17040 15990 17096
rect 16302 18944 16358 19000
rect 16210 18808 16266 18864
rect 16026 12824 16082 12880
rect 16210 13504 16266 13560
rect 15842 10140 15844 10160
rect 15844 10140 15896 10160
rect 15896 10140 15898 10160
rect 15842 10104 15898 10140
rect 16026 8608 16082 8664
rect 16118 8472 16174 8528
rect 13910 7112 13966 7168
rect 13542 6704 13598 6760
rect 12898 6568 12954 6624
rect 12530 2644 12586 2680
rect 12530 2624 12532 2644
rect 12532 2624 12584 2644
rect 12584 2624 12586 2644
rect 13818 6740 13820 6760
rect 13820 6740 13872 6760
rect 13872 6740 13874 6760
rect 13818 6704 13874 6740
rect 14002 6432 14058 6488
rect 14554 6296 14610 6352
rect 14370 6160 14426 6216
rect 16210 5208 16266 5264
rect 16118 4256 16174 4312
rect 14278 3304 14334 3360
rect 15658 3052 15714 3088
rect 15658 3032 15660 3052
rect 15660 3032 15712 3052
rect 15712 3032 15714 3052
rect 16578 32272 16634 32328
rect 16670 29008 16726 29064
rect 17130 33260 17132 33280
rect 17132 33260 17184 33280
rect 17184 33260 17186 33280
rect 17130 33224 17186 33260
rect 16486 22616 16542 22672
rect 16578 22480 16634 22536
rect 16486 22344 16542 22400
rect 16762 22752 16818 22808
rect 17038 27104 17094 27160
rect 17774 35556 17830 35592
rect 17774 35536 17776 35556
rect 17776 35536 17828 35556
rect 17828 35536 17830 35556
rect 17774 34040 17830 34096
rect 17038 24792 17094 24848
rect 17038 21936 17094 21992
rect 16946 20884 16948 20904
rect 16948 20884 17000 20904
rect 17000 20884 17002 20904
rect 16946 20848 17002 20884
rect 16670 20440 16726 20496
rect 16946 19252 16948 19272
rect 16948 19252 17000 19272
rect 17000 19252 17002 19272
rect 16946 19216 17002 19252
rect 16946 18808 17002 18864
rect 16670 18128 16726 18184
rect 16578 15136 16634 15192
rect 16946 17040 17002 17096
rect 16946 14184 17002 14240
rect 16578 13912 16634 13968
rect 16670 13640 16726 13696
rect 16578 12824 16634 12880
rect 16486 10920 16542 10976
rect 16854 13368 16910 13424
rect 16946 12960 17002 13016
rect 16670 11464 16726 11520
rect 16670 10684 16672 10704
rect 16672 10684 16724 10704
rect 16724 10684 16726 10704
rect 16670 10648 16726 10684
rect 16670 8372 16672 8392
rect 16672 8372 16724 8392
rect 16724 8372 16726 8392
rect 16670 8336 16726 8372
rect 16854 8492 16910 8528
rect 16854 8472 16856 8492
rect 16856 8472 16908 8492
rect 16908 8472 16910 8492
rect 16854 6860 16910 6896
rect 16854 6840 16856 6860
rect 16856 6840 16908 6860
rect 16908 6840 16910 6860
rect 16670 5616 16726 5672
rect 17406 25744 17462 25800
rect 18418 38392 18474 38448
rect 18050 36116 18052 36136
rect 18052 36116 18104 36136
rect 18104 36116 18106 36136
rect 18050 36080 18106 36116
rect 17958 34856 18014 34912
rect 17958 34060 18014 34096
rect 17958 34040 17960 34060
rect 17960 34040 18012 34060
rect 18012 34040 18014 34060
rect 17866 30912 17922 30968
rect 17498 24928 17554 24984
rect 17958 21664 18014 21720
rect 17314 20032 17370 20088
rect 17222 19624 17278 19680
rect 17130 19216 17186 19272
rect 17222 18536 17278 18592
rect 17590 19216 17646 19272
rect 17774 20712 17830 20768
rect 17314 17448 17370 17504
rect 17222 16496 17278 16552
rect 17774 18128 17830 18184
rect 17498 16496 17554 16552
rect 17498 16224 17554 16280
rect 17498 12552 17554 12608
rect 17314 12280 17370 12336
rect 17130 4936 17186 4992
rect 17774 14864 17830 14920
rect 17682 12824 17738 12880
rect 17958 17992 18014 18048
rect 18970 38120 19026 38176
rect 18878 37576 18934 37632
rect 18326 37304 18382 37360
rect 18602 37324 18658 37360
rect 18602 37304 18604 37324
rect 18604 37304 18656 37324
rect 18656 37304 18658 37324
rect 18234 30912 18290 30968
rect 18786 36488 18842 36544
rect 18326 30660 18382 30696
rect 18326 30640 18328 30660
rect 18328 30640 18380 30660
rect 18380 30640 18382 30660
rect 18234 26016 18290 26072
rect 18510 26288 18566 26344
rect 18510 25200 18566 25256
rect 18142 21292 18144 21312
rect 18144 21292 18196 21312
rect 18196 21292 18198 21312
rect 18142 21256 18198 21292
rect 18142 18808 18198 18864
rect 18142 17720 18198 17776
rect 17958 14048 18014 14104
rect 17682 11872 17738 11928
rect 17406 10240 17462 10296
rect 17590 10648 17646 10704
rect 17498 5888 17554 5944
rect 17222 4664 17278 4720
rect 17222 4256 17278 4312
rect 17130 4120 17186 4176
rect 17866 10260 17922 10296
rect 17866 10240 17868 10260
rect 17868 10240 17920 10260
rect 17920 10240 17922 10260
rect 18050 11620 18106 11656
rect 18050 11600 18052 11620
rect 18052 11600 18104 11620
rect 18104 11600 18106 11620
rect 18142 9868 18144 9888
rect 18144 9868 18196 9888
rect 18196 9868 18198 9888
rect 18142 9832 18198 9868
rect 18418 18944 18474 19000
rect 18694 23044 18750 23080
rect 18694 23024 18696 23044
rect 18696 23024 18748 23044
rect 18748 23024 18750 23044
rect 19062 33360 19118 33416
rect 19580 38650 19636 38652
rect 19660 38650 19716 38652
rect 19740 38650 19796 38652
rect 19820 38650 19876 38652
rect 19580 38598 19606 38650
rect 19606 38598 19636 38650
rect 19660 38598 19670 38650
rect 19670 38598 19716 38650
rect 19740 38598 19786 38650
rect 19786 38598 19796 38650
rect 19820 38598 19850 38650
rect 19850 38598 19876 38650
rect 19580 38596 19636 38598
rect 19660 38596 19716 38598
rect 19740 38596 19796 38598
rect 19820 38596 19876 38598
rect 19430 38548 19486 38584
rect 19430 38528 19432 38548
rect 19432 38528 19484 38548
rect 19484 38528 19486 38548
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 19338 37032 19394 37088
rect 19890 36624 19946 36680
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 19338 33224 19394 33280
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 18878 27920 18934 27976
rect 18878 24656 18934 24712
rect 18602 19352 18658 19408
rect 18602 19080 18658 19136
rect 18602 18128 18658 18184
rect 18786 16632 18842 16688
rect 18602 12724 18604 12744
rect 18604 12724 18656 12744
rect 18656 12724 18658 12744
rect 18602 12688 18658 12724
rect 18510 12552 18566 12608
rect 18510 12280 18566 12336
rect 17958 7520 18014 7576
rect 19062 32000 19118 32056
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 19062 30232 19118 30288
rect 19338 30776 19394 30832
rect 19338 30640 19394 30696
rect 19338 29996 19340 30016
rect 19340 29996 19392 30016
rect 19392 29996 19394 30016
rect 19338 29960 19394 29996
rect 19062 27920 19118 27976
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 19798 28192 19854 28248
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 19154 24928 19210 24984
rect 19062 21428 19064 21448
rect 19064 21428 19116 21448
rect 19116 21428 19118 21448
rect 19062 21392 19118 21428
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 19338 26288 19394 26344
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 19890 23588 19946 23624
rect 19890 23568 19892 23588
rect 19892 23568 19944 23588
rect 19944 23568 19946 23588
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 19246 19896 19302 19952
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 20534 35672 20590 35728
rect 20074 35400 20130 35456
rect 20442 33516 20498 33552
rect 20442 33496 20444 33516
rect 20444 33496 20496 33516
rect 20496 33496 20498 33516
rect 20258 25744 20314 25800
rect 20258 22752 20314 22808
rect 19430 18028 19432 18048
rect 19432 18028 19484 18048
rect 19484 18028 19486 18048
rect 19430 17992 19486 18028
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 19798 16668 19800 16688
rect 19800 16668 19852 16688
rect 19852 16668 19854 16688
rect 19798 16632 19854 16668
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 19338 15272 19394 15328
rect 18970 14048 19026 14104
rect 19890 15136 19946 15192
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 18602 9036 18658 9072
rect 18602 9016 18604 9036
rect 18604 9016 18656 9036
rect 18656 9016 18658 9036
rect 18694 7792 18750 7848
rect 18510 7384 18566 7440
rect 18510 6432 18566 6488
rect 17866 4020 17868 4040
rect 17868 4020 17920 4040
rect 17920 4020 17922 4040
rect 17866 3984 17922 4020
rect 18050 2372 18106 2408
rect 18050 2352 18052 2372
rect 18052 2352 18104 2372
rect 18104 2352 18106 2372
rect 17866 1572 17868 1592
rect 17868 1572 17920 1592
rect 17920 1572 17922 1592
rect 17866 1536 17922 1572
rect 19338 13912 19394 13968
rect 19522 14320 19578 14376
rect 19890 14320 19946 14376
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 19338 12688 19394 12744
rect 19154 11192 19210 11248
rect 19338 12280 19394 12336
rect 20258 20576 20314 20632
rect 20166 17584 20222 17640
rect 20166 14900 20168 14920
rect 20168 14900 20220 14920
rect 20220 14900 20222 14920
rect 20166 14864 20222 14900
rect 20074 12960 20130 13016
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 20534 27920 20590 27976
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 19154 10376 19210 10432
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 20994 33632 21050 33688
rect 22742 38392 22798 38448
rect 22558 37848 22614 37904
rect 22742 35264 22798 35320
rect 22374 34856 22430 34912
rect 21914 33768 21970 33824
rect 21178 33224 21234 33280
rect 21822 33360 21878 33416
rect 21086 31592 21142 31648
rect 20994 30368 21050 30424
rect 21546 31728 21602 31784
rect 21270 30504 21326 30560
rect 21178 29280 21234 29336
rect 20902 21664 20958 21720
rect 20626 20304 20682 20360
rect 20810 15816 20866 15872
rect 20718 15136 20774 15192
rect 19246 9424 19302 9480
rect 18970 9016 19026 9072
rect 18786 7520 18842 7576
rect 18786 5752 18842 5808
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19706 7656 19762 7712
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19430 6840 19486 6896
rect 20350 7404 20406 7440
rect 20350 7384 20352 7404
rect 20352 7384 20404 7404
rect 20404 7384 20406 7404
rect 19062 6296 19118 6352
rect 17958 856 18014 912
rect 18694 856 18750 912
rect 19982 6024 20038 6080
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 19430 5616 19486 5672
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 20718 12688 20774 12744
rect 20810 9560 20866 9616
rect 20810 8880 20866 8936
rect 23478 38528 23534 38584
rect 23202 38412 23258 38448
rect 23202 38392 23204 38412
rect 23204 38392 23256 38412
rect 23256 38392 23258 38412
rect 24398 38392 24454 38448
rect 24582 38392 24638 38448
rect 23570 37440 23626 37496
rect 22466 33532 22468 33552
rect 22468 33532 22520 33552
rect 22520 33532 22522 33552
rect 22466 33496 22522 33532
rect 22098 33088 22154 33144
rect 21638 28056 21694 28112
rect 21362 25336 21418 25392
rect 22282 30132 22284 30152
rect 22284 30132 22336 30152
rect 22336 30132 22338 30152
rect 22282 30096 22338 30132
rect 22374 29960 22430 30016
rect 22190 28620 22246 28656
rect 22190 28600 22192 28620
rect 22192 28600 22244 28620
rect 22244 28600 22246 28620
rect 21178 20576 21234 20632
rect 21362 20712 21418 20768
rect 21270 19488 21326 19544
rect 21546 21664 21602 21720
rect 21178 9832 21234 9888
rect 20902 6296 20958 6352
rect 20442 5888 20498 5944
rect 19982 4528 20038 4584
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 20166 2932 20168 2952
rect 20168 2932 20220 2952
rect 20220 2932 20222 2952
rect 19430 2796 19432 2816
rect 19432 2796 19484 2816
rect 19484 2796 19486 2816
rect 19430 2760 19486 2796
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 20166 2896 20222 2932
rect 21638 20884 21640 20904
rect 21640 20884 21692 20904
rect 21692 20884 21694 20904
rect 21638 20848 21694 20884
rect 22558 29708 22614 29744
rect 22558 29688 22560 29708
rect 22560 29688 22612 29708
rect 22612 29688 22614 29708
rect 23018 30796 23074 30832
rect 23018 30776 23020 30796
rect 23020 30776 23072 30796
rect 23072 30776 23074 30796
rect 23294 34856 23350 34912
rect 23478 29688 23534 29744
rect 22926 28620 22982 28656
rect 22926 28600 22928 28620
rect 22928 28600 22980 28620
rect 22980 28600 22982 28620
rect 22834 26424 22890 26480
rect 21730 17584 21786 17640
rect 21822 15156 21878 15192
rect 21822 15136 21824 15156
rect 21824 15136 21876 15156
rect 21876 15136 21878 15156
rect 21822 11328 21878 11384
rect 22466 16496 22522 16552
rect 22374 15952 22430 16008
rect 22558 15272 22614 15328
rect 22558 12960 22614 13016
rect 22466 12860 22468 12880
rect 22468 12860 22520 12880
rect 22520 12860 22522 12880
rect 22466 12824 22522 12860
rect 22190 7792 22246 7848
rect 22466 7656 22522 7712
rect 22282 7248 22338 7304
rect 22558 6568 22614 6624
rect 21362 5072 21418 5128
rect 21270 3304 21326 3360
rect 22558 2896 22614 2952
rect 23202 28212 23258 28248
rect 23202 28192 23204 28212
rect 23204 28192 23256 28212
rect 23256 28192 23258 28212
rect 23294 20576 23350 20632
rect 23110 17740 23166 17776
rect 23110 17720 23112 17740
rect 23112 17720 23164 17740
rect 23164 17720 23166 17740
rect 23110 10920 23166 10976
rect 23294 9152 23350 9208
rect 23202 4392 23258 4448
rect 24858 37440 24914 37496
rect 24306 37304 24362 37360
rect 25134 36780 25190 36816
rect 25134 36760 25136 36780
rect 25136 36760 25188 36780
rect 25188 36760 25190 36780
rect 24030 36488 24086 36544
rect 23846 34992 23902 35048
rect 23662 33088 23718 33144
rect 23662 31628 23664 31648
rect 23664 31628 23716 31648
rect 23716 31628 23718 31648
rect 23662 31592 23718 31628
rect 23754 31320 23810 31376
rect 23938 33224 23994 33280
rect 24950 35828 25006 35864
rect 24950 35808 24952 35828
rect 24952 35808 25004 35828
rect 25004 35808 25006 35828
rect 25134 34892 25136 34912
rect 25136 34892 25188 34912
rect 25188 34892 25190 34912
rect 25134 34856 25190 34892
rect 24582 34584 24638 34640
rect 24398 32680 24454 32736
rect 25502 33632 25558 33688
rect 24674 31884 24730 31920
rect 24674 31864 24676 31884
rect 24676 31864 24728 31884
rect 24728 31864 24730 31884
rect 24950 31864 25006 31920
rect 24030 27512 24086 27568
rect 23662 26560 23718 26616
rect 23662 24928 23718 24984
rect 23570 19896 23626 19952
rect 23938 25336 23994 25392
rect 24490 27376 24546 27432
rect 24306 24656 24362 24712
rect 23846 21548 23902 21584
rect 23846 21528 23848 21548
rect 23848 21528 23900 21548
rect 23900 21528 23902 21548
rect 23938 19508 23994 19544
rect 23938 19488 23940 19508
rect 23940 19488 23992 19508
rect 23992 19488 23994 19508
rect 24398 23296 24454 23352
rect 24490 20204 24492 20224
rect 24492 20204 24544 20224
rect 24544 20204 24546 20224
rect 24490 20168 24546 20204
rect 24306 19252 24308 19272
rect 24308 19252 24360 19272
rect 24360 19252 24362 19272
rect 24306 19216 24362 19252
rect 24306 18808 24362 18864
rect 23938 18128 23994 18184
rect 23570 10104 23626 10160
rect 24214 17604 24270 17640
rect 24214 17584 24216 17604
rect 24216 17584 24268 17604
rect 24268 17584 24270 17604
rect 23754 16360 23810 16416
rect 23754 15816 23810 15872
rect 23846 14220 23848 14240
rect 23848 14220 23900 14240
rect 23900 14220 23902 14240
rect 23846 14184 23902 14220
rect 24490 15156 24546 15192
rect 24490 15136 24492 15156
rect 24492 15136 24544 15156
rect 24544 15136 24546 15156
rect 23662 7928 23718 7984
rect 23386 2624 23442 2680
rect 24674 27532 24730 27568
rect 24674 27512 24676 27532
rect 24676 27512 24728 27532
rect 24728 27512 24730 27532
rect 24858 27920 24914 27976
rect 24766 26968 24822 27024
rect 25502 32000 25558 32056
rect 26790 38528 26846 38584
rect 25778 31728 25834 31784
rect 26238 29688 26294 29744
rect 26146 29452 26148 29472
rect 26148 29452 26200 29472
rect 26200 29452 26202 29472
rect 26146 29416 26202 29452
rect 25410 28872 25466 28928
rect 25318 28192 25374 28248
rect 25502 27376 25558 27432
rect 25318 27240 25374 27296
rect 25778 25744 25834 25800
rect 25042 25200 25098 25256
rect 25502 24268 25558 24304
rect 25502 24248 25504 24268
rect 25504 24248 25556 24268
rect 25556 24248 25558 24268
rect 24858 23740 24860 23760
rect 24860 23740 24912 23760
rect 24912 23740 24914 23760
rect 24858 23704 24914 23740
rect 25318 23568 25374 23624
rect 25226 20168 25282 20224
rect 24766 19896 24822 19952
rect 25410 19624 25466 19680
rect 24674 9288 24730 9344
rect 25594 20576 25650 20632
rect 27618 35128 27674 35184
rect 27342 34584 27398 34640
rect 26146 26560 26202 26616
rect 26238 26460 26240 26480
rect 26240 26460 26292 26480
rect 26292 26460 26294 26480
rect 26238 26424 26294 26460
rect 26514 25880 26570 25936
rect 26238 23316 26294 23352
rect 26238 23296 26240 23316
rect 26240 23296 26292 23316
rect 26292 23296 26294 23316
rect 25962 22516 25964 22536
rect 25964 22516 26016 22536
rect 26016 22516 26018 22536
rect 25962 22480 26018 22516
rect 26054 21528 26110 21584
rect 25962 20476 25964 20496
rect 25964 20476 26016 20496
rect 26016 20476 26018 20496
rect 25962 20440 26018 20476
rect 25962 19896 26018 19952
rect 25502 17448 25558 17504
rect 25410 15544 25466 15600
rect 25134 15136 25190 15192
rect 25318 14184 25374 14240
rect 25594 12300 25650 12336
rect 25594 12280 25596 12300
rect 25596 12280 25648 12300
rect 25648 12280 25650 12300
rect 26238 19216 26294 19272
rect 26238 17312 26294 17368
rect 26514 17312 26570 17368
rect 27618 34448 27674 34504
rect 27986 31864 28042 31920
rect 30838 38120 30894 38176
rect 30562 37032 30618 37088
rect 30378 34448 30434 34504
rect 30654 34620 30656 34640
rect 30656 34620 30708 34640
rect 30708 34620 30710 34640
rect 30654 34584 30710 34620
rect 30286 34176 30342 34232
rect 30194 33396 30196 33416
rect 30196 33396 30248 33416
rect 30248 33396 30250 33416
rect 29826 32952 29882 33008
rect 28722 32816 28778 32872
rect 27066 26152 27122 26208
rect 27066 23704 27122 23760
rect 26698 20712 26754 20768
rect 26238 16360 26294 16416
rect 25778 9696 25834 9752
rect 25778 9596 25780 9616
rect 25780 9596 25832 9616
rect 25832 9596 25834 9616
rect 25778 9560 25834 9596
rect 25962 9560 26018 9616
rect 26146 9152 26202 9208
rect 24582 5616 24638 5672
rect 24950 6160 25006 6216
rect 24582 3576 24638 3632
rect 24398 2760 24454 2816
rect 26238 5752 26294 5808
rect 26698 14456 26754 14512
rect 26790 12008 26846 12064
rect 26790 4276 26846 4312
rect 26790 4256 26792 4276
rect 26792 4256 26844 4276
rect 26844 4256 26846 4276
rect 27158 22344 27214 22400
rect 27342 21800 27398 21856
rect 27066 19660 27068 19680
rect 27068 19660 27120 19680
rect 27120 19660 27122 19680
rect 27066 19624 27122 19660
rect 26974 18964 27030 19000
rect 26974 18944 26976 18964
rect 26976 18944 27028 18964
rect 27028 18944 27030 18964
rect 27434 17584 27490 17640
rect 27250 16668 27252 16688
rect 27252 16668 27304 16688
rect 27304 16668 27306 16688
rect 27250 16632 27306 16668
rect 27066 16360 27122 16416
rect 27342 9560 27398 9616
rect 27066 6060 27068 6080
rect 27068 6060 27120 6080
rect 27120 6060 27122 6080
rect 27066 6024 27122 6060
rect 26974 5480 27030 5536
rect 27710 29688 27766 29744
rect 27618 26424 27674 26480
rect 28538 31728 28594 31784
rect 28262 29708 28318 29744
rect 28262 29688 28264 29708
rect 28264 29688 28316 29708
rect 28316 29688 28318 29708
rect 27986 28056 28042 28112
rect 27894 20440 27950 20496
rect 27802 18400 27858 18456
rect 27710 17720 27766 17776
rect 27802 15544 27858 15600
rect 27710 15136 27766 15192
rect 28354 26152 28410 26208
rect 28078 22208 28134 22264
rect 28078 20576 28134 20632
rect 28078 18284 28134 18320
rect 28078 18264 28080 18284
rect 28080 18264 28132 18284
rect 28132 18264 28134 18284
rect 27986 12144 28042 12200
rect 29182 32816 29238 32872
rect 29182 31728 29238 31784
rect 28998 30232 29054 30288
rect 30194 33360 30250 33396
rect 30010 31340 30066 31376
rect 30010 31320 30012 31340
rect 30012 31320 30064 31340
rect 30064 31320 30066 31340
rect 30010 30796 30066 30832
rect 30010 30776 30012 30796
rect 30012 30776 30064 30796
rect 30064 30776 30066 30796
rect 29550 30096 29606 30152
rect 28722 27004 28724 27024
rect 28724 27004 28776 27024
rect 28776 27004 28778 27024
rect 28722 26968 28778 27004
rect 28538 25744 28594 25800
rect 28722 25644 28724 25664
rect 28724 25644 28776 25664
rect 28776 25644 28778 25664
rect 28722 25608 28778 25644
rect 28446 24268 28502 24304
rect 28446 24248 28448 24268
rect 28448 24248 28500 24268
rect 28500 24248 28502 24268
rect 28722 11600 28778 11656
rect 28538 11328 28594 11384
rect 28722 6860 28778 6896
rect 28722 6840 28724 6860
rect 28724 6840 28776 6860
rect 28776 6840 28778 6860
rect 28078 5888 28134 5944
rect 27526 3168 27582 3224
rect 27342 2760 27398 2816
rect 29090 27376 29146 27432
rect 29090 26308 29146 26344
rect 29090 26288 29092 26308
rect 29092 26288 29144 26308
rect 29144 26288 29146 26308
rect 29274 28872 29330 28928
rect 29734 29960 29790 30016
rect 29826 29552 29882 29608
rect 29366 25880 29422 25936
rect 30470 29708 30526 29744
rect 30470 29688 30472 29708
rect 30472 29688 30524 29708
rect 30524 29688 30526 29708
rect 30562 28056 30618 28112
rect 29642 21936 29698 21992
rect 29550 20168 29606 20224
rect 28998 17992 29054 18048
rect 29090 17720 29146 17776
rect 29642 18400 29698 18456
rect 29550 17584 29606 17640
rect 29550 16496 29606 16552
rect 30470 25608 30526 25664
rect 30194 23160 30250 23216
rect 30378 22344 30434 22400
rect 30838 27276 30840 27296
rect 30840 27276 30892 27296
rect 30892 27276 30894 27296
rect 30838 27240 30894 27276
rect 30470 21800 30526 21856
rect 30194 20848 30250 20904
rect 30470 20576 30526 20632
rect 29918 17484 29920 17504
rect 29920 17484 29972 17504
rect 29972 17484 29974 17504
rect 29918 17448 29974 17484
rect 30286 19216 30342 19272
rect 30378 17756 30380 17776
rect 30380 17756 30432 17776
rect 30432 17756 30434 17776
rect 30378 17720 30434 17756
rect 30654 18264 30710 18320
rect 31206 36896 31262 36952
rect 31482 38392 31538 38448
rect 31390 38004 31446 38040
rect 31390 37984 31392 38004
rect 31392 37984 31444 38004
rect 31444 37984 31446 38004
rect 31206 26444 31262 26480
rect 31206 26424 31208 26444
rect 31208 26424 31260 26444
rect 31260 26424 31262 26444
rect 32402 38256 32458 38312
rect 34426 39480 34482 39536
rect 33230 37984 33286 38040
rect 35254 40160 35310 40216
rect 34940 39194 34996 39196
rect 35020 39194 35076 39196
rect 35100 39194 35156 39196
rect 35180 39194 35236 39196
rect 34940 39142 34966 39194
rect 34966 39142 34996 39194
rect 35020 39142 35030 39194
rect 35030 39142 35076 39194
rect 35100 39142 35146 39194
rect 35146 39142 35156 39194
rect 35180 39142 35210 39194
rect 35210 39142 35236 39194
rect 34940 39140 34996 39142
rect 35020 39140 35076 39142
rect 35100 39140 35156 39142
rect 35180 39140 35236 39142
rect 35254 38800 35310 38856
rect 34940 38106 34996 38108
rect 35020 38106 35076 38108
rect 35100 38106 35156 38108
rect 35180 38106 35236 38108
rect 34940 38054 34966 38106
rect 34966 38054 34996 38106
rect 35020 38054 35030 38106
rect 35030 38054 35076 38106
rect 35100 38054 35146 38106
rect 35146 38054 35156 38106
rect 35180 38054 35210 38106
rect 35210 38054 35236 38106
rect 34940 38052 34996 38054
rect 35020 38052 35076 38054
rect 35100 38052 35156 38054
rect 35180 38052 35236 38054
rect 34794 37712 34850 37768
rect 32678 36624 32734 36680
rect 31942 35264 31998 35320
rect 31574 24520 31630 24576
rect 30746 16652 30802 16688
rect 30746 16632 30748 16652
rect 30748 16632 30800 16652
rect 30800 16632 30802 16652
rect 30470 15272 30526 15328
rect 30378 13096 30434 13152
rect 29642 12300 29698 12336
rect 29642 12280 29644 12300
rect 29644 12280 29696 12300
rect 29696 12280 29698 12300
rect 29458 11328 29514 11384
rect 29550 10784 29606 10840
rect 29458 5480 29514 5536
rect 29274 4392 29330 4448
rect 29366 2760 29422 2816
rect 31206 18964 31262 19000
rect 31206 18944 31208 18964
rect 31208 18944 31260 18964
rect 31260 18944 31262 18964
rect 31482 20712 31538 20768
rect 31390 17856 31446 17912
rect 31390 17312 31446 17368
rect 31390 15136 31446 15192
rect 31666 20440 31722 20496
rect 32770 32000 32826 32056
rect 32126 29416 32182 29472
rect 32034 26016 32090 26072
rect 32678 27376 32734 27432
rect 31942 16496 31998 16552
rect 31942 15952 31998 16008
rect 30930 12960 30986 13016
rect 31850 13132 31852 13152
rect 31852 13132 31904 13152
rect 31904 13132 31906 13152
rect 31850 13096 31906 13132
rect 30930 12008 30986 12064
rect 32126 14476 32182 14512
rect 32126 14456 32128 14476
rect 32128 14456 32180 14476
rect 32180 14456 32182 14476
rect 32034 10648 32090 10704
rect 30838 6840 30894 6896
rect 32494 15564 32550 15600
rect 32494 15544 32496 15564
rect 32496 15544 32548 15564
rect 32548 15544 32550 15564
rect 32218 7792 32274 7848
rect 31390 4936 31446 4992
rect 32954 22652 32956 22672
rect 32956 22652 33008 22672
rect 33008 22652 33010 22672
rect 32954 22616 33010 22652
rect 34610 33904 34666 33960
rect 33598 31864 33654 31920
rect 33138 26968 33194 27024
rect 33046 19488 33102 19544
rect 30838 2760 30894 2816
rect 33138 5208 33194 5264
rect 33046 4392 33102 4448
rect 32770 3188 32826 3224
rect 32770 3168 32772 3188
rect 32772 3168 32824 3188
rect 32824 3168 32826 3188
rect 1398 720 1454 776
rect 33322 21256 33378 21312
rect 34334 29588 34336 29608
rect 34336 29588 34388 29608
rect 34388 29588 34390 29608
rect 34334 29552 34390 29588
rect 33690 27376 33746 27432
rect 34150 27376 34206 27432
rect 33506 24556 33508 24576
rect 33508 24556 33560 24576
rect 33560 24556 33562 24576
rect 33506 24520 33562 24556
rect 33874 24520 33930 24576
rect 34518 23704 34574 23760
rect 33874 23568 33930 23624
rect 33874 20576 33930 20632
rect 34058 20304 34114 20360
rect 33506 19252 33508 19272
rect 33508 19252 33560 19272
rect 33560 19252 33562 19272
rect 33506 19216 33562 19252
rect 34058 19080 34114 19136
rect 33782 17448 33838 17504
rect 33414 10240 33470 10296
rect 34058 16532 34060 16552
rect 34060 16532 34112 16552
rect 34112 16532 34114 16552
rect 34058 16496 34114 16532
rect 34518 17856 34574 17912
rect 33966 9016 34022 9072
rect 33506 7656 33562 7712
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 35346 34720 35402 34776
rect 35438 34176 35494 34232
rect 35346 34040 35402 34096
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 35254 30640 35310 30696
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 35254 29960 35310 30016
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 36358 38256 36414 38312
rect 35898 37848 35954 37904
rect 36082 37868 36138 37904
rect 36082 37848 36084 37868
rect 36084 37848 36136 37868
rect 36136 37848 36138 37868
rect 35806 37440 35862 37496
rect 38198 37848 38254 37904
rect 36818 36488 36874 36544
rect 39578 37168 39634 37224
rect 36082 35808 36138 35864
rect 37370 35400 37426 35456
rect 35622 31320 35678 31376
rect 35806 31320 35862 31376
rect 35438 29280 35494 29336
rect 34702 27920 34758 27976
rect 35346 27920 35402 27976
rect 37278 29552 37334 29608
rect 37370 28736 37426 28792
rect 36082 28600 36138 28656
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 34886 26560 34942 26616
rect 35254 26560 35310 26616
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 35254 25336 35310 25392
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34702 23024 34758 23080
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 35346 22480 35402 22536
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 35438 22208 35494 22264
rect 34702 21120 34758 21176
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 35162 19760 35218 19816
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 34794 18808 34850 18864
rect 35070 18808 35126 18864
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 35530 17740 35586 17776
rect 35530 17720 35532 17740
rect 35532 17720 35584 17740
rect 35584 17720 35586 17740
rect 35438 17040 35494 17096
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 34886 15988 34888 16008
rect 34888 15988 34940 16008
rect 34940 15988 34942 16008
rect 34886 15952 34942 15988
rect 34610 9424 34666 9480
rect 34702 7520 34758 7576
rect 34518 6840 34574 6896
rect 34610 4936 34666 4992
rect 34058 1400 34114 1456
rect 34242 1400 34298 1456
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 35070 9580 35126 9616
rect 35070 9560 35072 9580
rect 35072 9560 35124 9580
rect 35124 9560 35126 9580
rect 35254 9596 35256 9616
rect 35256 9596 35308 9616
rect 35308 9596 35310 9616
rect 35254 9560 35310 9596
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 35254 6296 35310 6352
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 34794 4120 34850 4176
rect 35714 14320 35770 14376
rect 35530 13640 35586 13696
rect 35438 5480 35494 5536
rect 35254 3440 35310 3496
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 35622 2796 35624 2816
rect 35624 2796 35676 2816
rect 35676 2796 35678 2816
rect 35622 2760 35678 2796
rect 35162 2644 35218 2680
rect 35162 2624 35164 2644
rect 35164 2624 35216 2644
rect 35216 2624 35218 2644
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 36266 27512 36322 27568
rect 36082 25200 36138 25256
rect 36082 22516 36084 22536
rect 36084 22516 36136 22536
rect 36136 22516 36138 22536
rect 36082 22480 36138 22516
rect 37370 23160 37426 23216
rect 37278 22636 37334 22672
rect 37278 22616 37280 22636
rect 37280 22616 37332 22636
rect 37332 22616 37334 22636
rect 36266 21936 36322 21992
rect 37462 21256 37518 21312
rect 37278 12688 37334 12744
rect 37370 5480 37426 5536
rect 35990 3984 36046 4040
rect 37738 3984 37794 4040
rect 39578 3848 39634 3904
rect 39118 3032 39174 3088
rect 38198 2488 38254 2544
rect 33230 40 33286 96
<< metal3 >>
rect 0 41578 800 41608
rect 3233 41578 3299 41581
rect 0 41576 3299 41578
rect 0 41520 3238 41576
rect 3294 41520 3299 41576
rect 0 41518 3299 41520
rect 0 41488 800 41518
rect 3233 41515 3299 41518
rect 35617 41578 35683 41581
rect 38852 41578 39652 41608
rect 35617 41576 39652 41578
rect 35617 41520 35622 41576
rect 35678 41520 39652 41576
rect 35617 41518 39652 41520
rect 35617 41515 35683 41518
rect 38852 41488 39652 41518
rect 0 40898 800 40928
rect 2957 40898 3023 40901
rect 0 40896 3023 40898
rect 0 40840 2962 40896
rect 3018 40840 3023 40896
rect 0 40838 3023 40840
rect 0 40808 800 40838
rect 2957 40835 3023 40838
rect 0 40218 800 40248
rect 3417 40218 3483 40221
rect 0 40216 3483 40218
rect 0 40160 3422 40216
rect 3478 40160 3483 40216
rect 0 40158 3483 40160
rect 0 40128 800 40158
rect 3417 40155 3483 40158
rect 35249 40218 35315 40221
rect 38852 40218 39652 40248
rect 35249 40216 39652 40218
rect 35249 40160 35254 40216
rect 35310 40160 39652 40216
rect 35249 40158 39652 40160
rect 35249 40155 35315 40158
rect 38852 40128 39652 40158
rect 34421 39538 34487 39541
rect 38852 39538 39652 39568
rect 34421 39536 39652 39538
rect 34421 39480 34426 39536
rect 34482 39480 39652 39536
rect 34421 39478 39652 39480
rect 34421 39475 34487 39478
rect 38852 39448 39652 39478
rect 4208 39200 4528 39201
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 34928 39200 35248 39201
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 39135 35248 39136
rect 0 38858 800 38888
rect 35249 38858 35315 38861
rect 38852 38858 39652 38888
rect 0 38798 3434 38858
rect 0 38768 800 38798
rect 3374 38725 3434 38798
rect 35249 38856 39652 38858
rect 35249 38800 35254 38856
rect 35310 38800 39652 38856
rect 35249 38798 39652 38800
rect 35249 38795 35315 38798
rect 38852 38768 39652 38798
rect 3374 38720 3483 38725
rect 3374 38664 3422 38720
rect 3478 38664 3483 38720
rect 3374 38662 3483 38664
rect 3417 38659 3483 38662
rect 19568 38656 19888 38657
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 38591 19888 38592
rect 933 38586 999 38589
rect 17534 38586 17540 38588
rect 933 38584 17540 38586
rect 933 38528 938 38584
rect 994 38528 17540 38584
rect 933 38526 17540 38528
rect 933 38523 999 38526
rect 17534 38524 17540 38526
rect 17604 38524 17610 38588
rect 19425 38586 19491 38589
rect 17726 38584 19491 38586
rect 17726 38528 19430 38584
rect 19486 38528 19491 38584
rect 17726 38526 19491 38528
rect 7833 38450 7899 38453
rect 10174 38450 10180 38452
rect 7833 38448 10180 38450
rect 7833 38392 7838 38448
rect 7894 38392 10180 38448
rect 7833 38390 10180 38392
rect 7833 38387 7899 38390
rect 10174 38388 10180 38390
rect 10244 38388 10250 38452
rect 10593 38450 10659 38453
rect 10910 38450 10916 38452
rect 10593 38448 10916 38450
rect 10593 38392 10598 38448
rect 10654 38392 10916 38448
rect 10593 38390 10916 38392
rect 10593 38387 10659 38390
rect 10910 38388 10916 38390
rect 10980 38388 10986 38452
rect 13353 38450 13419 38453
rect 17726 38450 17786 38526
rect 19425 38523 19491 38526
rect 23473 38586 23539 38589
rect 26785 38586 26851 38589
rect 23473 38584 26851 38586
rect 23473 38528 23478 38584
rect 23534 38528 26790 38584
rect 26846 38528 26851 38584
rect 23473 38526 26851 38528
rect 23473 38523 23539 38526
rect 26785 38523 26851 38526
rect 13353 38448 17786 38450
rect 13353 38392 13358 38448
rect 13414 38392 17786 38448
rect 13353 38390 17786 38392
rect 18413 38450 18479 38453
rect 22737 38450 22803 38453
rect 18413 38448 22803 38450
rect 18413 38392 18418 38448
rect 18474 38392 22742 38448
rect 22798 38392 22803 38448
rect 18413 38390 22803 38392
rect 13353 38387 13419 38390
rect 18413 38387 18479 38390
rect 22737 38387 22803 38390
rect 23197 38450 23263 38453
rect 24393 38450 24459 38453
rect 23197 38448 24459 38450
rect 23197 38392 23202 38448
rect 23258 38392 24398 38448
rect 24454 38392 24459 38448
rect 23197 38390 24459 38392
rect 23197 38387 23263 38390
rect 24393 38387 24459 38390
rect 24577 38450 24643 38453
rect 31477 38450 31543 38453
rect 24577 38448 31543 38450
rect 24577 38392 24582 38448
rect 24638 38392 31482 38448
rect 31538 38392 31543 38448
rect 24577 38390 31543 38392
rect 24577 38387 24643 38390
rect 31477 38387 31543 38390
rect 32397 38314 32463 38317
rect 36353 38314 36419 38317
rect 32397 38312 36419 38314
rect 32397 38256 32402 38312
rect 32458 38256 36358 38312
rect 36414 38256 36419 38312
rect 32397 38254 36419 38256
rect 32397 38251 32463 38254
rect 36353 38251 36419 38254
rect 0 38178 800 38208
rect 2773 38178 2839 38181
rect 0 38176 2839 38178
rect 0 38120 2778 38176
rect 2834 38120 2839 38176
rect 0 38118 2839 38120
rect 0 38088 800 38118
rect 2773 38115 2839 38118
rect 18965 38178 19031 38181
rect 30833 38178 30899 38181
rect 18965 38176 30899 38178
rect 18965 38120 18970 38176
rect 19026 38120 30838 38176
rect 30894 38120 30899 38176
rect 18965 38118 30899 38120
rect 18965 38115 19031 38118
rect 30833 38115 30899 38118
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 34928 38112 35248 38113
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 38047 35248 38048
rect 9949 38042 10015 38045
rect 31385 38042 31451 38045
rect 33225 38042 33291 38045
rect 9949 38040 26986 38042
rect 9949 37984 9954 38040
rect 10010 37984 26986 38040
rect 9949 37982 26986 37984
rect 9949 37979 10015 37982
rect 11513 37906 11579 37909
rect 15561 37906 15627 37909
rect 22553 37906 22619 37909
rect 11513 37904 15440 37906
rect 11513 37848 11518 37904
rect 11574 37848 15440 37904
rect 11513 37846 15440 37848
rect 11513 37843 11579 37846
rect 1393 37770 1459 37773
rect 13629 37770 13695 37773
rect 1393 37768 13695 37770
rect 1393 37712 1398 37768
rect 1454 37712 13634 37768
rect 13690 37712 13695 37768
rect 1393 37710 13695 37712
rect 1393 37707 1459 37710
rect 13629 37707 13695 37710
rect 15380 37634 15440 37846
rect 15561 37904 22619 37906
rect 15561 37848 15566 37904
rect 15622 37848 22558 37904
rect 22614 37848 22619 37904
rect 15561 37846 22619 37848
rect 26926 37906 26986 37982
rect 31385 38040 33291 38042
rect 31385 37984 31390 38040
rect 31446 37984 33230 38040
rect 33286 37984 33291 38040
rect 31385 37982 33291 37984
rect 31385 37979 31451 37982
rect 33225 37979 33291 37982
rect 35893 37906 35959 37909
rect 26926 37904 35959 37906
rect 26926 37848 35898 37904
rect 35954 37848 35959 37904
rect 26926 37846 35959 37848
rect 15561 37843 15627 37846
rect 22553 37843 22619 37846
rect 35893 37843 35959 37846
rect 36077 37906 36143 37909
rect 38193 37906 38259 37909
rect 36077 37904 38259 37906
rect 36077 37848 36082 37904
rect 36138 37848 38198 37904
rect 38254 37848 38259 37904
rect 36077 37846 38259 37848
rect 36077 37843 36143 37846
rect 38193 37843 38259 37846
rect 17309 37770 17375 37773
rect 34789 37770 34855 37773
rect 17309 37768 34855 37770
rect 17309 37712 17314 37768
rect 17370 37712 34794 37768
rect 34850 37712 34855 37768
rect 17309 37710 34855 37712
rect 17309 37707 17375 37710
rect 34789 37707 34855 37710
rect 18873 37634 18939 37637
rect 15380 37632 18939 37634
rect 15380 37576 18878 37632
rect 18934 37576 18939 37632
rect 15380 37574 18939 37576
rect 18873 37571 18939 37574
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 7373 37498 7439 37501
rect 9673 37498 9739 37501
rect 7373 37496 9739 37498
rect 7373 37440 7378 37496
rect 7434 37440 9678 37496
rect 9734 37440 9739 37496
rect 7373 37438 9739 37440
rect 7373 37435 7439 37438
rect 9673 37435 9739 37438
rect 23565 37498 23631 37501
rect 24853 37498 24919 37501
rect 23565 37496 24919 37498
rect 23565 37440 23570 37496
rect 23626 37440 24858 37496
rect 24914 37440 24919 37496
rect 23565 37438 24919 37440
rect 23565 37435 23631 37438
rect 24853 37435 24919 37438
rect 35801 37498 35867 37501
rect 38852 37498 39652 37528
rect 35801 37496 39652 37498
rect 35801 37440 35806 37496
rect 35862 37440 39652 37496
rect 35801 37438 39652 37440
rect 35801 37435 35867 37438
rect 38852 37408 39652 37438
rect 1761 37362 1827 37365
rect 9213 37362 9279 37365
rect 10409 37362 10475 37365
rect 1761 37360 10475 37362
rect 1761 37304 1766 37360
rect 1822 37304 9218 37360
rect 9274 37304 10414 37360
rect 10470 37304 10475 37360
rect 1761 37302 10475 37304
rect 1761 37299 1827 37302
rect 9213 37299 9279 37302
rect 10409 37299 10475 37302
rect 15653 37362 15719 37365
rect 18321 37362 18387 37365
rect 15653 37360 18387 37362
rect 15653 37304 15658 37360
rect 15714 37304 18326 37360
rect 18382 37304 18387 37360
rect 15653 37302 18387 37304
rect 15653 37299 15719 37302
rect 18321 37299 18387 37302
rect 18597 37362 18663 37365
rect 24301 37362 24367 37365
rect 18597 37360 24367 37362
rect 18597 37304 18602 37360
rect 18658 37304 24306 37360
rect 24362 37304 24367 37360
rect 18597 37302 24367 37304
rect 18597 37299 18663 37302
rect 24301 37299 24367 37302
rect 2313 37226 2379 37229
rect 6821 37226 6887 37229
rect 2313 37224 6887 37226
rect 2313 37168 2318 37224
rect 2374 37168 6826 37224
rect 6882 37168 6887 37224
rect 2313 37166 6887 37168
rect 2313 37163 2379 37166
rect 6821 37163 6887 37166
rect 15745 37226 15811 37229
rect 39573 37226 39639 37229
rect 15745 37224 39639 37226
rect 15745 37168 15750 37224
rect 15806 37168 39578 37224
rect 39634 37168 39639 37224
rect 15745 37166 39639 37168
rect 15745 37163 15811 37166
rect 39573 37163 39639 37166
rect 19333 37090 19399 37093
rect 30557 37090 30623 37093
rect 19333 37088 30623 37090
rect 19333 37032 19338 37088
rect 19394 37032 30562 37088
rect 30618 37032 30623 37088
rect 19333 37030 30623 37032
rect 19333 37027 19399 37030
rect 30557 37027 30623 37030
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 14733 36954 14799 36957
rect 31201 36954 31267 36957
rect 14733 36952 31267 36954
rect 14733 36896 14738 36952
rect 14794 36896 31206 36952
rect 31262 36896 31267 36952
rect 14733 36894 31267 36896
rect 14733 36891 14799 36894
rect 31201 36891 31267 36894
rect 0 36818 800 36848
rect 4061 36818 4127 36821
rect 25129 36818 25195 36821
rect 38852 36818 39652 36848
rect 0 36758 1962 36818
rect 0 36728 800 36758
rect 1902 36274 1962 36758
rect 4061 36816 25195 36818
rect 4061 36760 4066 36816
rect 4122 36760 25134 36816
rect 25190 36760 25195 36816
rect 4061 36758 25195 36760
rect 4061 36755 4127 36758
rect 25129 36755 25195 36758
rect 37046 36758 39652 36818
rect 6821 36682 6887 36685
rect 16205 36682 16271 36685
rect 19885 36682 19951 36685
rect 32673 36682 32739 36685
rect 6821 36680 10978 36682
rect 6821 36624 6826 36680
rect 6882 36624 10978 36680
rect 6821 36622 10978 36624
rect 6821 36619 6887 36622
rect 10918 36549 10978 36622
rect 16205 36680 19951 36682
rect 16205 36624 16210 36680
rect 16266 36624 19890 36680
rect 19946 36624 19951 36680
rect 16205 36622 19951 36624
rect 16205 36619 16271 36622
rect 19885 36619 19951 36622
rect 22694 36680 32739 36682
rect 22694 36624 32678 36680
rect 32734 36624 32739 36680
rect 22694 36622 32739 36624
rect 10918 36546 11027 36549
rect 18781 36546 18847 36549
rect 10918 36544 18847 36546
rect 10918 36488 10966 36544
rect 11022 36488 18786 36544
rect 18842 36488 18847 36544
rect 10918 36486 18847 36488
rect 10961 36483 11027 36486
rect 18781 36483 18847 36486
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 16297 36410 16363 36413
rect 22694 36410 22754 36622
rect 32673 36619 32739 36622
rect 24025 36546 24091 36549
rect 36813 36546 36879 36549
rect 24025 36544 36879 36546
rect 24025 36488 24030 36544
rect 24086 36488 36818 36544
rect 36874 36488 36879 36544
rect 24025 36486 36879 36488
rect 24025 36483 24091 36486
rect 36813 36483 36879 36486
rect 37046 36410 37106 36758
rect 38852 36728 39652 36758
rect 16297 36408 18108 36410
rect 16297 36352 16302 36408
rect 16358 36352 18108 36408
rect 16297 36350 18108 36352
rect 16297 36347 16363 36350
rect 18048 36274 18108 36350
rect 20118 36350 22754 36410
rect 35206 36350 37106 36410
rect 20118 36274 20178 36350
rect 1902 36214 17970 36274
rect 18048 36214 20178 36274
rect 0 36138 800 36168
rect 0 36078 3986 36138
rect 0 36048 800 36078
rect 3926 35594 3986 36078
rect 13721 36002 13787 36005
rect 14273 36002 14339 36005
rect 13721 36000 14339 36002
rect 13721 35944 13726 36000
rect 13782 35944 14278 36000
rect 14334 35944 14339 36000
rect 13721 35942 14339 35944
rect 13721 35939 13787 35942
rect 14273 35939 14339 35942
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 17910 35866 17970 36214
rect 18045 36138 18111 36141
rect 35206 36138 35266 36350
rect 38852 36138 39652 36168
rect 18045 36136 35266 36138
rect 18045 36080 18050 36136
rect 18106 36080 35266 36136
rect 18045 36078 35266 36080
rect 36126 36078 39652 36138
rect 18045 36075 18111 36078
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 36126 35869 36186 36078
rect 38852 36048 39652 36078
rect 24945 35866 25011 35869
rect 17910 35864 25011 35866
rect 17910 35808 24950 35864
rect 25006 35808 25011 35864
rect 17910 35806 25011 35808
rect 24945 35803 25011 35806
rect 36077 35864 36186 35869
rect 36077 35808 36082 35864
rect 36138 35808 36186 35864
rect 36077 35806 36186 35808
rect 36077 35803 36143 35806
rect 8385 35730 8451 35733
rect 20529 35730 20595 35733
rect 8385 35728 20595 35730
rect 8385 35672 8390 35728
rect 8446 35672 20534 35728
rect 20590 35672 20595 35728
rect 8385 35670 20595 35672
rect 8385 35667 8451 35670
rect 20529 35667 20595 35670
rect 17769 35594 17835 35597
rect 3926 35592 17835 35594
rect 3926 35536 17774 35592
rect 17830 35536 17835 35592
rect 3926 35534 17835 35536
rect 17769 35531 17835 35534
rect 0 35458 800 35488
rect 4061 35458 4127 35461
rect 0 35456 4127 35458
rect 0 35400 4066 35456
rect 4122 35400 4127 35456
rect 0 35398 4127 35400
rect 0 35368 800 35398
rect 4061 35395 4127 35398
rect 20069 35458 20135 35461
rect 37365 35458 37431 35461
rect 20069 35456 37431 35458
rect 20069 35400 20074 35456
rect 20130 35400 37370 35456
rect 37426 35400 37431 35456
rect 20069 35398 37431 35400
rect 20069 35395 20135 35398
rect 37365 35395 37431 35398
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 22737 35322 22803 35325
rect 31937 35322 32003 35325
rect 22737 35320 32003 35322
rect 22737 35264 22742 35320
rect 22798 35264 31942 35320
rect 31998 35264 32003 35320
rect 22737 35262 32003 35264
rect 22737 35259 22803 35262
rect 31937 35259 32003 35262
rect 13 35186 79 35189
rect 27613 35186 27679 35189
rect 13 35184 27679 35186
rect 13 35128 18 35184
rect 74 35128 27618 35184
rect 27674 35128 27679 35184
rect 13 35126 27679 35128
rect 13 35123 79 35126
rect 27613 35123 27679 35126
rect 13629 35050 13695 35053
rect 23841 35050 23907 35053
rect 13629 35048 23907 35050
rect 13629 34992 13634 35048
rect 13690 34992 23846 35048
rect 23902 34992 23907 35048
rect 13629 34990 23907 34992
rect 13629 34987 13695 34990
rect 23841 34987 23907 34990
rect 17953 34914 18019 34917
rect 22369 34914 22435 34917
rect 17953 34912 22435 34914
rect 17953 34856 17958 34912
rect 18014 34856 22374 34912
rect 22430 34856 22435 34912
rect 17953 34854 22435 34856
rect 17953 34851 18019 34854
rect 22369 34851 22435 34854
rect 23289 34914 23355 34917
rect 25129 34914 25195 34917
rect 23289 34912 25195 34914
rect 23289 34856 23294 34912
rect 23350 34856 25134 34912
rect 25190 34856 25195 34912
rect 23289 34854 25195 34856
rect 23289 34851 23355 34854
rect 25129 34851 25195 34854
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 35341 34778 35407 34781
rect 38852 34778 39652 34808
rect 35341 34776 39652 34778
rect 35341 34720 35346 34776
rect 35402 34720 39652 34776
rect 35341 34718 39652 34720
rect 35341 34715 35407 34718
rect 38852 34688 39652 34718
rect 24577 34642 24643 34645
rect 27337 34642 27403 34645
rect 30649 34642 30715 34645
rect 24577 34640 30715 34642
rect 24577 34584 24582 34640
rect 24638 34584 27342 34640
rect 27398 34584 30654 34640
rect 30710 34584 30715 34640
rect 24577 34582 30715 34584
rect 24577 34579 24643 34582
rect 27337 34579 27403 34582
rect 30649 34579 30715 34582
rect 9029 34506 9095 34509
rect 14549 34506 14615 34509
rect 9029 34504 14615 34506
rect 9029 34448 9034 34504
rect 9090 34448 14554 34504
rect 14610 34448 14615 34504
rect 9029 34446 14615 34448
rect 9029 34443 9095 34446
rect 14549 34443 14615 34446
rect 27613 34506 27679 34509
rect 30373 34506 30439 34509
rect 27613 34504 30439 34506
rect 27613 34448 27618 34504
rect 27674 34448 30378 34504
rect 30434 34448 30439 34504
rect 27613 34446 30439 34448
rect 27613 34443 27679 34446
rect 30373 34443 30439 34446
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 1577 34234 1643 34237
rect 30281 34234 30347 34237
rect 35433 34234 35499 34237
rect 1577 34232 3618 34234
rect 1577 34176 1582 34232
rect 1638 34176 3618 34232
rect 1577 34174 3618 34176
rect 1577 34171 1643 34174
rect 0 34098 800 34128
rect 3417 34098 3483 34101
rect 0 34096 3483 34098
rect 0 34040 3422 34096
rect 3478 34040 3483 34096
rect 0 34038 3483 34040
rect 3558 34098 3618 34174
rect 30281 34232 35499 34234
rect 30281 34176 30286 34232
rect 30342 34176 35438 34232
rect 35494 34176 35499 34232
rect 30281 34174 35499 34176
rect 30281 34171 30347 34174
rect 35433 34171 35499 34174
rect 17769 34098 17835 34101
rect 3558 34096 17835 34098
rect 3558 34040 17774 34096
rect 17830 34040 17835 34096
rect 3558 34038 17835 34040
rect 0 34008 800 34038
rect 3417 34035 3483 34038
rect 17769 34035 17835 34038
rect 17953 34098 18019 34101
rect 35341 34098 35407 34101
rect 38852 34098 39652 34128
rect 17953 34096 35407 34098
rect 17953 34040 17958 34096
rect 18014 34040 35346 34096
rect 35402 34040 35407 34096
rect 17953 34038 35407 34040
rect 17953 34035 18019 34038
rect 35341 34035 35407 34038
rect 35574 34038 39652 34098
rect 34605 33962 34671 33965
rect 35574 33962 35634 34038
rect 38852 34008 39652 34038
rect 34605 33960 35634 33962
rect 34605 33904 34610 33960
rect 34666 33904 35634 33960
rect 34605 33902 35634 33904
rect 34605 33899 34671 33902
rect 21909 33826 21975 33829
rect 20118 33824 21975 33826
rect 20118 33768 21914 33824
rect 21970 33768 21975 33824
rect 20118 33766 21975 33768
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 20118 33690 20178 33766
rect 21909 33763 21975 33766
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 4662 33630 20178 33690
rect 20989 33690 21055 33693
rect 25497 33690 25563 33693
rect 20989 33688 25563 33690
rect 20989 33632 20994 33688
rect 21050 33632 25502 33688
rect 25558 33632 25563 33688
rect 20989 33630 25563 33632
rect 0 33418 800 33448
rect 4662 33418 4722 33630
rect 20989 33627 21055 33630
rect 25497 33627 25563 33630
rect 6913 33554 6979 33557
rect 14457 33554 14523 33557
rect 6913 33552 14523 33554
rect 6913 33496 6918 33552
rect 6974 33496 14462 33552
rect 14518 33496 14523 33552
rect 6913 33494 14523 33496
rect 6913 33491 6979 33494
rect 14457 33491 14523 33494
rect 20437 33554 20503 33557
rect 22461 33554 22527 33557
rect 20437 33552 22527 33554
rect 20437 33496 20442 33552
rect 20498 33496 22466 33552
rect 22522 33496 22527 33552
rect 20437 33494 22527 33496
rect 20437 33491 20503 33494
rect 22461 33491 22527 33494
rect 0 33358 4722 33418
rect 6177 33418 6243 33421
rect 7005 33418 7071 33421
rect 6177 33416 7071 33418
rect 6177 33360 6182 33416
rect 6238 33360 7010 33416
rect 7066 33360 7071 33416
rect 6177 33358 7071 33360
rect 0 33328 800 33358
rect 6177 33355 6243 33358
rect 7005 33355 7071 33358
rect 14641 33418 14707 33421
rect 19057 33418 19123 33421
rect 14641 33416 19123 33418
rect 14641 33360 14646 33416
rect 14702 33360 19062 33416
rect 19118 33360 19123 33416
rect 14641 33358 19123 33360
rect 14641 33355 14707 33358
rect 19057 33355 19123 33358
rect 21817 33418 21883 33421
rect 30189 33418 30255 33421
rect 21817 33416 30255 33418
rect 21817 33360 21822 33416
rect 21878 33360 30194 33416
rect 30250 33360 30255 33416
rect 21817 33358 30255 33360
rect 21817 33355 21883 33358
rect 30189 33355 30255 33358
rect 3417 33282 3483 33285
rect 6913 33282 6979 33285
rect 3417 33280 6979 33282
rect 3417 33224 3422 33280
rect 3478 33224 6918 33280
rect 6974 33224 6979 33280
rect 3417 33222 6979 33224
rect 3417 33219 3483 33222
rect 6913 33219 6979 33222
rect 7097 33282 7163 33285
rect 14089 33282 14155 33285
rect 7097 33280 14155 33282
rect 7097 33224 7102 33280
rect 7158 33224 14094 33280
rect 14150 33224 14155 33280
rect 7097 33222 14155 33224
rect 7097 33219 7163 33222
rect 14089 33219 14155 33222
rect 17125 33282 17191 33285
rect 19333 33282 19399 33285
rect 17125 33280 19399 33282
rect 17125 33224 17130 33280
rect 17186 33224 19338 33280
rect 19394 33224 19399 33280
rect 17125 33222 19399 33224
rect 17125 33219 17191 33222
rect 19333 33219 19399 33222
rect 21173 33282 21239 33285
rect 23933 33282 23999 33285
rect 21173 33280 23999 33282
rect 21173 33224 21178 33280
rect 21234 33224 23938 33280
rect 23994 33224 23999 33280
rect 21173 33222 23999 33224
rect 21173 33219 21239 33222
rect 23933 33219 23999 33222
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 22093 33146 22159 33149
rect 23657 33146 23723 33149
rect 22093 33144 23723 33146
rect 22093 33088 22098 33144
rect 22154 33088 23662 33144
rect 23718 33088 23723 33144
rect 22093 33086 23723 33088
rect 22093 33083 22159 33086
rect 23657 33083 23723 33086
rect 23660 33010 23720 33083
rect 29821 33010 29887 33013
rect 23660 33008 29887 33010
rect 23660 32952 29826 33008
rect 29882 32952 29887 33008
rect 23660 32950 29887 32952
rect 29821 32947 29887 32950
rect 5993 32874 6059 32877
rect 3926 32872 6059 32874
rect 3926 32816 5998 32872
rect 6054 32816 6059 32872
rect 3926 32814 6059 32816
rect 0 32738 800 32768
rect 3926 32738 3986 32814
rect 5993 32811 6059 32814
rect 12617 32874 12683 32877
rect 15285 32874 15351 32877
rect 15653 32874 15719 32877
rect 12617 32872 15719 32874
rect 12617 32816 12622 32872
rect 12678 32816 15290 32872
rect 15346 32816 15658 32872
rect 15714 32816 15719 32872
rect 12617 32814 15719 32816
rect 12617 32811 12683 32814
rect 15285 32811 15351 32814
rect 15653 32811 15719 32814
rect 28717 32874 28783 32877
rect 29177 32874 29243 32877
rect 28717 32872 29243 32874
rect 28717 32816 28722 32872
rect 28778 32816 29182 32872
rect 29238 32816 29243 32872
rect 28717 32814 29243 32816
rect 28717 32811 28783 32814
rect 29177 32811 29243 32814
rect 24393 32738 24459 32741
rect 38852 32738 39652 32768
rect 0 32678 3986 32738
rect 21774 32736 24459 32738
rect 21774 32680 24398 32736
rect 24454 32680 24459 32736
rect 21774 32678 24459 32680
rect 0 32648 800 32678
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 14365 32602 14431 32605
rect 21774 32602 21834 32678
rect 24393 32675 24459 32678
rect 35390 32678 39652 32738
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 14365 32600 21834 32602
rect 14365 32544 14370 32600
rect 14426 32544 21834 32600
rect 14365 32542 21834 32544
rect 14365 32539 14431 32542
rect 16573 32330 16639 32333
rect 16573 32328 20178 32330
rect 16573 32272 16578 32328
rect 16634 32272 20178 32328
rect 16573 32270 20178 32272
rect 16573 32267 16639 32270
rect 10869 32194 10935 32197
rect 13353 32194 13419 32197
rect 10869 32192 13419 32194
rect 10869 32136 10874 32192
rect 10930 32136 13358 32192
rect 13414 32136 13419 32192
rect 10869 32134 13419 32136
rect 20118 32194 20178 32270
rect 35390 32194 35450 32678
rect 38852 32648 39652 32678
rect 20118 32134 35450 32194
rect 10869 32131 10935 32134
rect 13353 32131 13419 32134
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 11053 32058 11119 32061
rect 19057 32058 19123 32061
rect 11053 32056 19123 32058
rect 11053 32000 11058 32056
rect 11114 32000 19062 32056
rect 19118 32000 19123 32056
rect 11053 31998 19123 32000
rect 11053 31995 11119 31998
rect 19057 31995 19123 31998
rect 25497 32058 25563 32061
rect 32765 32058 32831 32061
rect 38852 32058 39652 32088
rect 25497 32056 32690 32058
rect 25497 32000 25502 32056
rect 25558 32000 32690 32056
rect 25497 31998 32690 32000
rect 25497 31995 25563 31998
rect 7925 31922 7991 31925
rect 15745 31922 15811 31925
rect 24669 31922 24735 31925
rect 7925 31920 15811 31922
rect 7925 31864 7930 31920
rect 7986 31864 15750 31920
rect 15806 31864 15811 31920
rect 7925 31862 15811 31864
rect 7925 31859 7991 31862
rect 15745 31859 15811 31862
rect 15886 31920 24735 31922
rect 15886 31864 24674 31920
rect 24730 31864 24735 31920
rect 15886 31862 24735 31864
rect 15886 31786 15946 31862
rect 24669 31859 24735 31862
rect 24945 31922 25011 31925
rect 27981 31922 28047 31925
rect 24945 31920 28047 31922
rect 24945 31864 24950 31920
rect 25006 31864 27986 31920
rect 28042 31864 28047 31920
rect 24945 31862 28047 31864
rect 32630 31922 32690 31998
rect 32765 32056 39652 32058
rect 32765 32000 32770 32056
rect 32826 32000 39652 32056
rect 32765 31998 39652 32000
rect 32765 31995 32831 31998
rect 38852 31968 39652 31998
rect 33593 31922 33659 31925
rect 32630 31920 33659 31922
rect 32630 31864 33598 31920
rect 33654 31864 33659 31920
rect 32630 31862 33659 31864
rect 24945 31859 25011 31862
rect 27981 31859 28047 31862
rect 33593 31859 33659 31862
rect 13862 31726 15946 31786
rect 21541 31786 21607 31789
rect 25773 31786 25839 31789
rect 21541 31784 25839 31786
rect 21541 31728 21546 31784
rect 21602 31728 25778 31784
rect 25834 31728 25839 31784
rect 21541 31726 25839 31728
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 13862 31514 13922 31726
rect 21541 31723 21607 31726
rect 25773 31723 25839 31726
rect 28533 31786 28599 31789
rect 29177 31786 29243 31789
rect 28533 31784 29243 31786
rect 28533 31728 28538 31784
rect 28594 31728 29182 31784
rect 29238 31728 29243 31784
rect 28533 31726 29243 31728
rect 28533 31723 28599 31726
rect 29177 31723 29243 31726
rect 21081 31650 21147 31653
rect 23657 31650 23723 31653
rect 21081 31648 23723 31650
rect 21081 31592 21086 31648
rect 21142 31592 23662 31648
rect 23718 31592 23723 31648
rect 21081 31590 23723 31592
rect 21081 31587 21147 31590
rect 23657 31587 23723 31590
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 7606 31454 13922 31514
rect 0 31378 800 31408
rect 7606 31378 7666 31454
rect 0 31318 7666 31378
rect 7741 31378 7807 31381
rect 16389 31378 16455 31381
rect 7741 31376 9506 31378
rect 7741 31320 7746 31376
rect 7802 31344 9506 31376
rect 9814 31376 16455 31378
rect 9814 31344 16394 31376
rect 7802 31320 16394 31344
rect 16450 31320 16455 31376
rect 7741 31318 16455 31320
rect 0 31288 800 31318
rect 7741 31315 7807 31318
rect 9446 31284 9874 31318
rect 16389 31315 16455 31318
rect 23749 31378 23815 31381
rect 30005 31378 30071 31381
rect 35617 31378 35683 31381
rect 23749 31376 35683 31378
rect 23749 31320 23754 31376
rect 23810 31320 30010 31376
rect 30066 31320 35622 31376
rect 35678 31320 35683 31376
rect 23749 31318 35683 31320
rect 23749 31315 23815 31318
rect 30005 31315 30071 31318
rect 35617 31315 35683 31318
rect 35801 31378 35867 31381
rect 38852 31378 39652 31408
rect 35801 31376 39652 31378
rect 35801 31320 35806 31376
rect 35862 31320 39652 31376
rect 35801 31318 39652 31320
rect 35801 31315 35867 31318
rect 38852 31288 39652 31318
rect 12985 31242 13051 31245
rect 15377 31242 15443 31245
rect 12985 31240 15443 31242
rect 12985 31184 12990 31240
rect 13046 31184 15382 31240
rect 15438 31184 15443 31240
rect 12985 31182 15443 31184
rect 12985 31179 13051 31182
rect 15377 31179 15443 31182
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 4061 30970 4127 30973
rect 4981 30970 5047 30973
rect 15469 30970 15535 30973
rect 4061 30968 15535 30970
rect 4061 30912 4066 30968
rect 4122 30912 4986 30968
rect 5042 30912 15474 30968
rect 15530 30912 15535 30968
rect 4061 30910 15535 30912
rect 4061 30907 4127 30910
rect 4981 30907 5047 30910
rect 15469 30907 15535 30910
rect 17861 30970 17927 30973
rect 18229 30970 18295 30973
rect 17861 30968 18295 30970
rect 17861 30912 17866 30968
rect 17922 30912 18234 30968
rect 18290 30912 18295 30968
rect 17861 30910 18295 30912
rect 17861 30907 17927 30910
rect 18229 30907 18295 30910
rect 19333 30834 19399 30837
rect 23013 30834 23079 30837
rect 30005 30834 30071 30837
rect 19333 30832 19810 30834
rect 19333 30776 19338 30832
rect 19394 30776 19810 30832
rect 19333 30774 19810 30776
rect 19333 30771 19399 30774
rect 0 30698 800 30728
rect 9581 30698 9647 30701
rect 18321 30698 18387 30701
rect 19333 30698 19399 30701
rect 0 30608 858 30698
rect 9581 30696 14474 30698
rect 9581 30640 9586 30696
rect 9642 30640 14474 30696
rect 9581 30638 14474 30640
rect 9581 30635 9647 30638
rect 798 30562 858 30608
rect 4061 30562 4127 30565
rect 798 30560 4127 30562
rect 798 30504 4066 30560
rect 4122 30504 4127 30560
rect 798 30502 4127 30504
rect 14414 30562 14474 30638
rect 18321 30696 19399 30698
rect 18321 30640 18326 30696
rect 18382 30640 19338 30696
rect 19394 30640 19399 30696
rect 18321 30638 19399 30640
rect 19750 30698 19810 30774
rect 23013 30832 30071 30834
rect 23013 30776 23018 30832
rect 23074 30776 30010 30832
rect 30066 30776 30071 30832
rect 23013 30774 30071 30776
rect 23013 30771 23079 30774
rect 30005 30771 30071 30774
rect 35249 30698 35315 30701
rect 19750 30696 35315 30698
rect 19750 30640 35254 30696
rect 35310 30640 35315 30696
rect 19750 30638 35315 30640
rect 18321 30635 18387 30638
rect 19333 30635 19399 30638
rect 35249 30635 35315 30638
rect 21265 30562 21331 30565
rect 14414 30560 21331 30562
rect 14414 30504 21270 30560
rect 21326 30504 21331 30560
rect 14414 30502 21331 30504
rect 4061 30499 4127 30502
rect 21265 30499 21331 30502
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 9949 30426 10015 30429
rect 11237 30426 11303 30429
rect 9949 30424 11303 30426
rect 9949 30368 9954 30424
rect 10010 30368 11242 30424
rect 11298 30368 11303 30424
rect 9949 30366 11303 30368
rect 9949 30363 10015 30366
rect 11237 30363 11303 30366
rect 13905 30426 13971 30429
rect 20989 30426 21055 30429
rect 13905 30424 21055 30426
rect 13905 30368 13910 30424
rect 13966 30368 20994 30424
rect 21050 30368 21055 30424
rect 13905 30366 21055 30368
rect 13905 30363 13971 30366
rect 20989 30363 21055 30366
rect 4889 30290 4955 30293
rect 6913 30290 6979 30293
rect 4889 30288 6979 30290
rect 4889 30232 4894 30288
rect 4950 30232 6918 30288
rect 6974 30232 6979 30288
rect 4889 30230 6979 30232
rect 4889 30227 4955 30230
rect 6913 30227 6979 30230
rect 7373 30290 7439 30293
rect 9673 30290 9739 30293
rect 7373 30288 9739 30290
rect 7373 30232 7378 30288
rect 7434 30232 9678 30288
rect 9734 30232 9739 30288
rect 7373 30230 9739 30232
rect 7373 30227 7439 30230
rect 9673 30227 9739 30230
rect 10317 30290 10383 30293
rect 14181 30290 14247 30293
rect 10317 30288 14247 30290
rect 10317 30232 10322 30288
rect 10378 30232 14186 30288
rect 14242 30232 14247 30288
rect 10317 30230 14247 30232
rect 10317 30227 10383 30230
rect 14181 30227 14247 30230
rect 19057 30290 19123 30293
rect 28993 30290 29059 30293
rect 19057 30288 29059 30290
rect 19057 30232 19062 30288
rect 19118 30232 28998 30288
rect 29054 30232 29059 30288
rect 19057 30230 29059 30232
rect 19057 30227 19123 30230
rect 28993 30227 29059 30230
rect 3417 30154 3483 30157
rect 6361 30154 6427 30157
rect 8569 30154 8635 30157
rect 3417 30152 8635 30154
rect 3417 30096 3422 30152
rect 3478 30096 6366 30152
rect 6422 30096 8574 30152
rect 8630 30096 8635 30152
rect 3417 30094 8635 30096
rect 3417 30091 3483 30094
rect 6361 30091 6427 30094
rect 8569 30091 8635 30094
rect 22277 30154 22343 30157
rect 29545 30154 29611 30157
rect 22277 30152 29611 30154
rect 22277 30096 22282 30152
rect 22338 30096 29550 30152
rect 29606 30096 29611 30152
rect 22277 30094 29611 30096
rect 22277 30091 22343 30094
rect 29545 30091 29611 30094
rect 8017 30018 8083 30021
rect 13353 30018 13419 30021
rect 8017 30016 13419 30018
rect 8017 29960 8022 30016
rect 8078 29960 13358 30016
rect 13414 29960 13419 30016
rect 8017 29958 13419 29960
rect 8017 29955 8083 29958
rect 13353 29955 13419 29958
rect 16389 30018 16455 30021
rect 19333 30018 19399 30021
rect 16389 30016 19399 30018
rect 16389 29960 16394 30016
rect 16450 29960 19338 30016
rect 19394 29960 19399 30016
rect 16389 29958 19399 29960
rect 16389 29955 16455 29958
rect 19333 29955 19399 29958
rect 22369 30018 22435 30021
rect 29729 30018 29795 30021
rect 22369 30016 29795 30018
rect 22369 29960 22374 30016
rect 22430 29960 29734 30016
rect 29790 29960 29795 30016
rect 22369 29958 29795 29960
rect 22369 29955 22435 29958
rect 29729 29955 29795 29958
rect 35249 30018 35315 30021
rect 38852 30018 39652 30048
rect 35249 30016 39652 30018
rect 35249 29960 35254 30016
rect 35310 29960 39652 30016
rect 35249 29958 39652 29960
rect 35249 29955 35315 29958
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 38852 29928 39652 29958
rect 19568 29887 19888 29888
rect 4061 29746 4127 29749
rect 22553 29746 22619 29749
rect 4061 29744 22619 29746
rect 4061 29688 4066 29744
rect 4122 29688 22558 29744
rect 22614 29688 22619 29744
rect 4061 29686 22619 29688
rect 4061 29683 4127 29686
rect 22553 29683 22619 29686
rect 23473 29746 23539 29749
rect 26233 29746 26299 29749
rect 27705 29746 27771 29749
rect 23473 29744 27771 29746
rect 23473 29688 23478 29744
rect 23534 29688 26238 29744
rect 26294 29688 27710 29744
rect 27766 29688 27771 29744
rect 23473 29686 27771 29688
rect 23473 29683 23539 29686
rect 26233 29683 26299 29686
rect 27705 29683 27771 29686
rect 28257 29746 28323 29749
rect 30465 29746 30531 29749
rect 28257 29744 30531 29746
rect 28257 29688 28262 29744
rect 28318 29688 30470 29744
rect 30526 29688 30531 29744
rect 28257 29686 30531 29688
rect 28257 29683 28323 29686
rect 30465 29683 30531 29686
rect 13629 29610 13695 29613
rect 15193 29610 15259 29613
rect 13629 29608 15259 29610
rect 13629 29552 13634 29608
rect 13690 29552 15198 29608
rect 15254 29552 15259 29608
rect 13629 29550 15259 29552
rect 13629 29547 13695 29550
rect 15193 29547 15259 29550
rect 29821 29610 29887 29613
rect 34329 29610 34395 29613
rect 37273 29610 37339 29613
rect 29821 29608 34395 29610
rect 29821 29552 29826 29608
rect 29882 29552 34334 29608
rect 34390 29552 34395 29608
rect 29821 29550 34395 29552
rect 29821 29547 29887 29550
rect 34329 29547 34395 29550
rect 34470 29608 37339 29610
rect 34470 29552 37278 29608
rect 37334 29552 37339 29608
rect 34470 29550 37339 29552
rect 26141 29474 26207 29477
rect 32121 29474 32187 29477
rect 34470 29474 34530 29550
rect 37273 29547 37339 29550
rect 26141 29472 34530 29474
rect 26141 29416 26146 29472
rect 26202 29416 32126 29472
rect 32182 29416 34530 29472
rect 26141 29414 34530 29416
rect 26141 29411 26207 29414
rect 32121 29411 32187 29414
rect 4208 29408 4528 29409
rect 0 29338 800 29368
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 1393 29338 1459 29341
rect 0 29336 1459 29338
rect 0 29280 1398 29336
rect 1454 29280 1459 29336
rect 0 29278 1459 29280
rect 0 29248 800 29278
rect 1393 29275 1459 29278
rect 14089 29338 14155 29341
rect 21173 29338 21239 29341
rect 14089 29336 21239 29338
rect 14089 29280 14094 29336
rect 14150 29280 21178 29336
rect 21234 29280 21239 29336
rect 14089 29278 21239 29280
rect 14089 29275 14155 29278
rect 21173 29275 21239 29278
rect 35433 29338 35499 29341
rect 38852 29338 39652 29368
rect 35433 29336 39652 29338
rect 35433 29280 35438 29336
rect 35494 29280 39652 29336
rect 35433 29278 39652 29280
rect 35433 29275 35499 29278
rect 38852 29248 39652 29278
rect 14089 29066 14155 29069
rect 16665 29066 16731 29069
rect 14089 29064 16731 29066
rect 14089 29008 14094 29064
rect 14150 29008 16670 29064
rect 16726 29008 16731 29064
rect 14089 29006 16731 29008
rect 14089 29003 14155 29006
rect 16665 29003 16731 29006
rect 4705 28930 4771 28933
rect 10409 28930 10475 28933
rect 4705 28928 10475 28930
rect 4705 28872 4710 28928
rect 4766 28872 10414 28928
rect 10470 28872 10475 28928
rect 4705 28870 10475 28872
rect 4705 28867 4771 28870
rect 10409 28867 10475 28870
rect 25405 28930 25471 28933
rect 29269 28930 29335 28933
rect 25405 28928 29335 28930
rect 25405 28872 25410 28928
rect 25466 28872 29274 28928
rect 29330 28872 29335 28928
rect 25405 28870 29335 28872
rect 25405 28867 25471 28870
rect 29269 28867 29335 28870
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 37365 28794 37431 28797
rect 34470 28792 37431 28794
rect 34470 28736 37370 28792
rect 37426 28736 37431 28792
rect 34470 28734 37431 28736
rect 0 28658 800 28688
rect 3141 28658 3207 28661
rect 0 28656 3207 28658
rect 0 28600 3146 28656
rect 3202 28600 3207 28656
rect 0 28598 3207 28600
rect 0 28568 800 28598
rect 3141 28595 3207 28598
rect 8661 28658 8727 28661
rect 11513 28658 11579 28661
rect 8661 28656 11579 28658
rect 8661 28600 8666 28656
rect 8722 28600 11518 28656
rect 11574 28600 11579 28656
rect 8661 28598 11579 28600
rect 8661 28595 8727 28598
rect 11513 28595 11579 28598
rect 13721 28658 13787 28661
rect 22185 28658 22251 28661
rect 13721 28656 22251 28658
rect 13721 28600 13726 28656
rect 13782 28600 22190 28656
rect 22246 28600 22251 28656
rect 13721 28598 22251 28600
rect 13721 28595 13787 28598
rect 22185 28595 22251 28598
rect 22921 28658 22987 28661
rect 34470 28658 34530 28734
rect 37365 28731 37431 28734
rect 22921 28656 34530 28658
rect 22921 28600 22926 28656
rect 22982 28600 34530 28656
rect 22921 28598 34530 28600
rect 36077 28658 36143 28661
rect 38852 28658 39652 28688
rect 36077 28656 39652 28658
rect 36077 28600 36082 28656
rect 36138 28600 39652 28656
rect 36077 28598 39652 28600
rect 22921 28595 22987 28598
rect 36077 28595 36143 28598
rect 38852 28568 39652 28598
rect 2957 28522 3023 28525
rect 16389 28522 16455 28525
rect 2957 28520 16455 28522
rect 2957 28464 2962 28520
rect 3018 28464 16394 28520
rect 16450 28464 16455 28520
rect 2957 28462 16455 28464
rect 2957 28459 3023 28462
rect 16389 28459 16455 28462
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 19793 28250 19859 28253
rect 23197 28250 23263 28253
rect 25313 28250 25379 28253
rect 19793 28248 25379 28250
rect 19793 28192 19798 28248
rect 19854 28192 23202 28248
rect 23258 28192 25318 28248
rect 25374 28192 25379 28248
rect 19793 28190 25379 28192
rect 19793 28187 19859 28190
rect 23197 28187 23263 28190
rect 25313 28187 25379 28190
rect 15009 28114 15075 28117
rect 21633 28114 21699 28117
rect 15009 28112 21699 28114
rect 15009 28056 15014 28112
rect 15070 28056 21638 28112
rect 21694 28056 21699 28112
rect 15009 28054 21699 28056
rect 15009 28051 15075 28054
rect 21633 28051 21699 28054
rect 27981 28114 28047 28117
rect 30557 28114 30623 28117
rect 27981 28112 30623 28114
rect 27981 28056 27986 28112
rect 28042 28056 30562 28112
rect 30618 28056 30623 28112
rect 27981 28054 30623 28056
rect 27981 28051 28047 28054
rect 30557 28051 30623 28054
rect 0 27978 800 28008
rect 2773 27978 2839 27981
rect 0 27976 2839 27978
rect 0 27920 2778 27976
rect 2834 27920 2839 27976
rect 0 27918 2839 27920
rect 0 27888 800 27918
rect 2773 27915 2839 27918
rect 10317 27978 10383 27981
rect 18873 27978 18939 27981
rect 10317 27976 18939 27978
rect 10317 27920 10322 27976
rect 10378 27920 18878 27976
rect 18934 27920 18939 27976
rect 10317 27918 18939 27920
rect 10317 27915 10383 27918
rect 18873 27915 18939 27918
rect 19057 27978 19123 27981
rect 20529 27978 20595 27981
rect 19057 27976 20595 27978
rect 19057 27920 19062 27976
rect 19118 27920 20534 27976
rect 20590 27920 20595 27976
rect 19057 27918 20595 27920
rect 19057 27915 19123 27918
rect 20529 27915 20595 27918
rect 24853 27978 24919 27981
rect 34697 27978 34763 27981
rect 35341 27978 35407 27981
rect 24853 27976 35407 27978
rect 24853 27920 24858 27976
rect 24914 27920 34702 27976
rect 34758 27920 35346 27976
rect 35402 27920 35407 27976
rect 24853 27918 35407 27920
rect 24853 27915 24919 27918
rect 31664 27884 31770 27918
rect 34697 27915 34763 27918
rect 35341 27915 35407 27918
rect 11513 27842 11579 27845
rect 12617 27842 12683 27845
rect 11513 27840 12683 27842
rect 11513 27784 11518 27840
rect 11574 27784 12622 27840
rect 12678 27784 12683 27840
rect 11513 27782 12683 27784
rect 11513 27779 11579 27782
rect 12617 27779 12683 27782
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 3049 27570 3115 27573
rect 11053 27570 11119 27573
rect 3049 27568 11119 27570
rect 3049 27512 3054 27568
rect 3110 27512 11058 27568
rect 11114 27512 11119 27568
rect 3049 27510 11119 27512
rect 3049 27507 3115 27510
rect 11053 27507 11119 27510
rect 11697 27570 11763 27573
rect 24025 27570 24091 27573
rect 11697 27568 24091 27570
rect 11697 27512 11702 27568
rect 11758 27512 24030 27568
rect 24086 27512 24091 27568
rect 11697 27510 24091 27512
rect 11697 27507 11763 27510
rect 24025 27507 24091 27510
rect 24669 27570 24735 27573
rect 36261 27570 36327 27573
rect 24669 27568 36327 27570
rect 24669 27512 24674 27568
rect 24730 27512 36266 27568
rect 36322 27512 36327 27568
rect 24669 27510 36327 27512
rect 24669 27507 24735 27510
rect 36261 27507 36327 27510
rect 3049 27434 3115 27437
rect 24485 27434 24551 27437
rect 3049 27432 24551 27434
rect 3049 27376 3054 27432
rect 3110 27376 24490 27432
rect 24546 27376 24551 27432
rect 3049 27374 24551 27376
rect 3049 27371 3115 27374
rect 24485 27371 24551 27374
rect 25497 27434 25563 27437
rect 29085 27434 29151 27437
rect 32673 27434 32739 27437
rect 33685 27434 33751 27437
rect 25497 27432 29151 27434
rect 25497 27376 25502 27432
rect 25558 27376 29090 27432
rect 29146 27376 29151 27432
rect 25497 27374 29151 27376
rect 25497 27371 25563 27374
rect 29085 27371 29151 27374
rect 32630 27432 33751 27434
rect 32630 27376 32678 27432
rect 32734 27376 33690 27432
rect 33746 27376 33751 27432
rect 32630 27374 33751 27376
rect 32630 27371 32739 27374
rect 33685 27371 33751 27374
rect 34145 27434 34211 27437
rect 34145 27432 35450 27434
rect 34145 27376 34150 27432
rect 34206 27376 35450 27432
rect 34145 27374 35450 27376
rect 34145 27371 34211 27374
rect 13445 27298 13511 27301
rect 25313 27298 25379 27301
rect 13445 27296 25379 27298
rect 13445 27240 13450 27296
rect 13506 27240 25318 27296
rect 25374 27240 25379 27296
rect 13445 27238 25379 27240
rect 13445 27235 13511 27238
rect 25313 27235 25379 27238
rect 30833 27298 30899 27301
rect 32630 27298 32690 27371
rect 30833 27296 32690 27298
rect 30833 27240 30838 27296
rect 30894 27240 32690 27296
rect 30833 27238 32690 27240
rect 35390 27298 35450 27374
rect 38852 27298 39652 27328
rect 35390 27238 39652 27298
rect 30833 27235 30899 27238
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 38852 27208 39652 27238
rect 34928 27167 35248 27168
rect 9765 27162 9831 27165
rect 14273 27162 14339 27165
rect 17033 27164 17099 27165
rect 16982 27162 16988 27164
rect 4662 27160 14339 27162
rect 4662 27104 9770 27160
rect 9826 27104 14278 27160
rect 14334 27104 14339 27160
rect 4662 27102 14339 27104
rect 16942 27102 16988 27162
rect 17052 27160 17099 27164
rect 17094 27104 17099 27160
rect 4662 27029 4722 27102
rect 9765 27099 9831 27102
rect 14273 27099 14339 27102
rect 16982 27100 16988 27102
rect 17052 27100 17099 27104
rect 17033 27099 17099 27100
rect 3877 27026 3943 27029
rect 4662 27026 4771 27029
rect 8109 27026 8175 27029
rect 14365 27026 14431 27029
rect 15469 27026 15535 27029
rect 3877 27024 4852 27026
rect 3877 26968 3882 27024
rect 3938 26968 4710 27024
rect 4766 26968 4852 27024
rect 3877 26966 4852 26968
rect 8109 27024 15535 27026
rect 8109 26968 8114 27024
rect 8170 26968 14370 27024
rect 14426 26968 15474 27024
rect 15530 26968 15535 27024
rect 8109 26966 15535 26968
rect 3877 26963 3943 26966
rect 4705 26963 4771 26966
rect 8109 26963 8175 26966
rect 14365 26963 14431 26966
rect 15469 26963 15535 26966
rect 24761 27026 24827 27029
rect 28717 27026 28783 27029
rect 33133 27026 33199 27029
rect 24761 27024 33199 27026
rect 24761 26968 24766 27024
rect 24822 26968 28722 27024
rect 28778 26968 33138 27024
rect 33194 26968 33199 27024
rect 24761 26966 33199 26968
rect 24761 26963 24827 26966
rect 28717 26963 28783 26966
rect 33133 26963 33199 26966
rect 7005 26754 7071 26757
rect 10133 26754 10199 26757
rect 7005 26752 10199 26754
rect 7005 26696 7010 26752
rect 7066 26696 10138 26752
rect 10194 26696 10199 26752
rect 7005 26694 10199 26696
rect 7005 26691 7071 26694
rect 10133 26691 10199 26694
rect 19568 26688 19888 26689
rect 0 26618 800 26648
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 2773 26618 2839 26621
rect 0 26616 2839 26618
rect 0 26560 2778 26616
rect 2834 26560 2839 26616
rect 0 26558 2839 26560
rect 0 26528 800 26558
rect 2773 26555 2839 26558
rect 5073 26618 5139 26621
rect 10593 26618 10659 26621
rect 5073 26616 10659 26618
rect 5073 26560 5078 26616
rect 5134 26560 10598 26616
rect 10654 26560 10659 26616
rect 5073 26558 10659 26560
rect 5073 26555 5139 26558
rect 10593 26555 10659 26558
rect 23657 26618 23723 26621
rect 26141 26618 26207 26621
rect 34881 26618 34947 26621
rect 23657 26616 34947 26618
rect 23657 26560 23662 26616
rect 23718 26560 26146 26616
rect 26202 26560 34886 26616
rect 34942 26560 34947 26616
rect 23657 26558 34947 26560
rect 23657 26555 23723 26558
rect 26141 26555 26207 26558
rect 34881 26555 34947 26558
rect 35249 26618 35315 26621
rect 38852 26618 39652 26648
rect 35249 26616 39652 26618
rect 35249 26560 35254 26616
rect 35310 26560 39652 26616
rect 35249 26558 39652 26560
rect 35249 26555 35315 26558
rect 38852 26528 39652 26558
rect 5809 26482 5875 26485
rect 10225 26482 10291 26485
rect 5809 26480 10291 26482
rect 5809 26424 5814 26480
rect 5870 26424 10230 26480
rect 10286 26424 10291 26480
rect 5809 26422 10291 26424
rect 5809 26419 5875 26422
rect 10225 26419 10291 26422
rect 22829 26482 22895 26485
rect 26233 26482 26299 26485
rect 27613 26482 27679 26485
rect 31201 26482 31267 26485
rect 22829 26480 26434 26482
rect 22829 26424 22834 26480
rect 22890 26424 26238 26480
rect 26294 26424 26434 26480
rect 22829 26422 26434 26424
rect 22829 26419 22895 26422
rect 26233 26419 26299 26422
rect 4981 26346 5047 26349
rect 9121 26346 9187 26349
rect 4981 26344 9187 26346
rect 4981 26288 4986 26344
rect 5042 26288 9126 26344
rect 9182 26288 9187 26344
rect 4981 26286 9187 26288
rect 4981 26283 5047 26286
rect 9121 26283 9187 26286
rect 9438 26284 9444 26348
rect 9508 26346 9514 26348
rect 9581 26346 9647 26349
rect 11605 26346 11671 26349
rect 9508 26344 11671 26346
rect 9508 26288 9586 26344
rect 9642 26288 11610 26344
rect 11666 26288 11671 26344
rect 9508 26286 11671 26288
rect 9508 26284 9514 26286
rect 9581 26283 9647 26286
rect 11605 26283 11671 26286
rect 11789 26346 11855 26349
rect 18505 26346 18571 26349
rect 19333 26346 19399 26349
rect 11789 26344 19399 26346
rect 11789 26288 11794 26344
rect 11850 26288 18510 26344
rect 18566 26288 19338 26344
rect 19394 26288 19399 26344
rect 11789 26286 19399 26288
rect 26374 26346 26434 26422
rect 27613 26480 31267 26482
rect 27613 26424 27618 26480
rect 27674 26424 31206 26480
rect 31262 26424 31267 26480
rect 27613 26422 31267 26424
rect 27613 26419 27679 26422
rect 31201 26419 31267 26422
rect 29085 26346 29151 26349
rect 26374 26344 29151 26346
rect 26374 26288 29090 26344
rect 29146 26288 29151 26344
rect 26374 26286 29151 26288
rect 11789 26283 11855 26286
rect 18505 26283 18571 26286
rect 19333 26283 19399 26286
rect 29085 26283 29151 26286
rect 5717 26210 5783 26213
rect 7189 26210 7255 26213
rect 5717 26208 7255 26210
rect 5717 26152 5722 26208
rect 5778 26152 7194 26208
rect 7250 26152 7255 26208
rect 5717 26150 7255 26152
rect 5717 26147 5783 26150
rect 7189 26147 7255 26150
rect 27061 26210 27127 26213
rect 28349 26210 28415 26213
rect 27061 26208 28415 26210
rect 27061 26152 27066 26208
rect 27122 26152 28354 26208
rect 28410 26152 28415 26208
rect 27061 26150 28415 26152
rect 27061 26147 27127 26150
rect 28349 26147 28415 26150
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 8385 26074 8451 26077
rect 11789 26074 11855 26077
rect 8385 26072 11855 26074
rect 8385 26016 8390 26072
rect 8446 26016 11794 26072
rect 11850 26016 11855 26072
rect 8385 26014 11855 26016
rect 8385 26011 8451 26014
rect 11789 26011 11855 26014
rect 18229 26074 18295 26077
rect 32029 26074 32095 26077
rect 18229 26072 32095 26074
rect 18229 26016 18234 26072
rect 18290 26016 32034 26072
rect 32090 26016 32095 26072
rect 18229 26014 32095 26016
rect 18229 26011 18295 26014
rect 32029 26011 32095 26014
rect 0 25938 800 25968
rect 4061 25938 4127 25941
rect 0 25936 4127 25938
rect 0 25880 4066 25936
rect 4122 25880 4127 25936
rect 0 25878 4127 25880
rect 0 25848 800 25878
rect 4061 25875 4127 25878
rect 6269 25938 6335 25941
rect 11789 25938 11855 25941
rect 6269 25936 11855 25938
rect 6269 25880 6274 25936
rect 6330 25880 11794 25936
rect 11850 25880 11855 25936
rect 6269 25878 11855 25880
rect 6269 25875 6335 25878
rect 11789 25875 11855 25878
rect 16113 25938 16179 25941
rect 26509 25938 26575 25941
rect 16113 25936 26575 25938
rect 16113 25880 16118 25936
rect 16174 25880 26514 25936
rect 26570 25880 26575 25936
rect 16113 25878 26575 25880
rect 16113 25875 16179 25878
rect 26509 25875 26575 25878
rect 29126 25876 29132 25940
rect 29196 25938 29202 25940
rect 29361 25938 29427 25941
rect 29196 25936 29427 25938
rect 29196 25880 29366 25936
rect 29422 25880 29427 25936
rect 29196 25878 29427 25880
rect 29196 25876 29202 25878
rect 29361 25875 29427 25878
rect 7189 25802 7255 25805
rect 10961 25802 11027 25805
rect 7189 25800 11027 25802
rect 7189 25744 7194 25800
rect 7250 25744 10966 25800
rect 11022 25744 11027 25800
rect 7189 25742 11027 25744
rect 7189 25739 7255 25742
rect 10961 25739 11027 25742
rect 17401 25802 17467 25805
rect 20253 25802 20319 25805
rect 17401 25800 20319 25802
rect 17401 25744 17406 25800
rect 17462 25744 20258 25800
rect 20314 25744 20319 25800
rect 17401 25742 20319 25744
rect 17401 25739 17467 25742
rect 20253 25739 20319 25742
rect 25773 25802 25839 25805
rect 28533 25802 28599 25805
rect 25773 25800 28599 25802
rect 25773 25744 25778 25800
rect 25834 25744 28538 25800
rect 28594 25744 28599 25800
rect 25773 25742 28599 25744
rect 25773 25739 25839 25742
rect 28533 25739 28599 25742
rect 8201 25666 8267 25669
rect 10041 25666 10107 25669
rect 8201 25664 10107 25666
rect 8201 25608 8206 25664
rect 8262 25608 10046 25664
rect 10102 25608 10107 25664
rect 8201 25606 10107 25608
rect 8201 25603 8267 25606
rect 10041 25603 10107 25606
rect 28717 25666 28783 25669
rect 30465 25666 30531 25669
rect 28717 25664 30531 25666
rect 28717 25608 28722 25664
rect 28778 25608 30470 25664
rect 30526 25608 30531 25664
rect 28717 25606 30531 25608
rect 28717 25603 28783 25606
rect 30465 25603 30531 25606
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 4521 25530 4587 25533
rect 11053 25530 11119 25533
rect 4521 25528 11119 25530
rect 4521 25472 4526 25528
rect 4582 25472 11058 25528
rect 11114 25472 11119 25528
rect 4521 25470 11119 25472
rect 4521 25467 4587 25470
rect 11053 25467 11119 25470
rect 11881 25394 11947 25397
rect 12985 25394 13051 25397
rect 21357 25394 21423 25397
rect 11881 25392 21423 25394
rect 11881 25336 11886 25392
rect 11942 25336 12990 25392
rect 13046 25336 21362 25392
rect 21418 25336 21423 25392
rect 11881 25334 21423 25336
rect 11881 25331 11947 25334
rect 12985 25331 13051 25334
rect 21357 25331 21423 25334
rect 23933 25394 23999 25397
rect 35249 25394 35315 25397
rect 23933 25392 35315 25394
rect 23933 25336 23938 25392
rect 23994 25336 35254 25392
rect 35310 25336 35315 25392
rect 23933 25334 35315 25336
rect 23933 25331 23999 25334
rect 35249 25331 35315 25334
rect 0 25258 800 25288
rect 2957 25258 3023 25261
rect 0 25256 3023 25258
rect 0 25200 2962 25256
rect 3018 25200 3023 25256
rect 0 25198 3023 25200
rect 0 25168 800 25198
rect 2957 25195 3023 25198
rect 10501 25258 10567 25261
rect 18505 25258 18571 25261
rect 25037 25258 25103 25261
rect 10501 25256 25103 25258
rect 10501 25200 10506 25256
rect 10562 25200 18510 25256
rect 18566 25200 25042 25256
rect 25098 25200 25103 25256
rect 10501 25198 25103 25200
rect 10501 25195 10567 25198
rect 18505 25195 18571 25198
rect 25037 25195 25103 25198
rect 36077 25258 36143 25261
rect 38852 25258 39652 25288
rect 36077 25256 39652 25258
rect 36077 25200 36082 25256
rect 36138 25200 39652 25256
rect 36077 25198 39652 25200
rect 36077 25195 36143 25198
rect 38852 25168 39652 25198
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 4705 24986 4771 24989
rect 8937 24986 9003 24989
rect 4705 24984 9003 24986
rect 4705 24928 4710 24984
rect 4766 24928 8942 24984
rect 8998 24928 9003 24984
rect 4705 24926 9003 24928
rect 4705 24923 4771 24926
rect 8937 24923 9003 24926
rect 10501 24986 10567 24989
rect 17493 24986 17559 24989
rect 10501 24984 17559 24986
rect 10501 24928 10506 24984
rect 10562 24928 17498 24984
rect 17554 24928 17559 24984
rect 10501 24926 17559 24928
rect 10501 24923 10567 24926
rect 17493 24923 17559 24926
rect 19149 24986 19215 24989
rect 23657 24986 23723 24989
rect 19149 24984 23723 24986
rect 19149 24928 19154 24984
rect 19210 24928 23662 24984
rect 23718 24928 23723 24984
rect 19149 24926 23723 24928
rect 19149 24923 19215 24926
rect 23657 24923 23723 24926
rect 9305 24850 9371 24853
rect 10504 24850 10564 24923
rect 9305 24848 10564 24850
rect 9305 24792 9310 24848
rect 9366 24792 10564 24848
rect 9305 24790 10564 24792
rect 13169 24850 13235 24853
rect 15285 24850 15351 24853
rect 13169 24848 15351 24850
rect 13169 24792 13174 24848
rect 13230 24792 15290 24848
rect 15346 24792 15351 24848
rect 13169 24790 15351 24792
rect 9305 24787 9371 24790
rect 13169 24787 13235 24790
rect 15285 24787 15351 24790
rect 15745 24850 15811 24853
rect 17033 24850 17099 24853
rect 15745 24848 17099 24850
rect 15745 24792 15750 24848
rect 15806 24792 17038 24848
rect 17094 24792 17099 24848
rect 15745 24790 17099 24792
rect 15745 24787 15811 24790
rect 17033 24787 17099 24790
rect 18873 24714 18939 24717
rect 24301 24714 24367 24717
rect 18873 24712 24367 24714
rect 18873 24656 18878 24712
rect 18934 24656 24306 24712
rect 24362 24656 24367 24712
rect 18873 24654 24367 24656
rect 18873 24651 18939 24654
rect 24301 24651 24367 24654
rect 12249 24578 12315 24581
rect 14089 24578 14155 24581
rect 12249 24576 14155 24578
rect 12249 24520 12254 24576
rect 12310 24520 14094 24576
rect 14150 24520 14155 24576
rect 12249 24518 14155 24520
rect 12249 24515 12315 24518
rect 14089 24515 14155 24518
rect 31569 24578 31635 24581
rect 33501 24578 33567 24581
rect 31569 24576 33567 24578
rect 31569 24520 31574 24576
rect 31630 24520 33506 24576
rect 33562 24520 33567 24576
rect 31569 24518 33567 24520
rect 31569 24515 31635 24518
rect 33501 24515 33567 24518
rect 33869 24578 33935 24581
rect 38852 24578 39652 24608
rect 33869 24576 39652 24578
rect 33869 24520 33874 24576
rect 33930 24520 39652 24576
rect 33869 24518 39652 24520
rect 33869 24515 33935 24518
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 38852 24488 39652 24518
rect 19568 24447 19888 24448
rect 7557 24442 7623 24445
rect 13169 24442 13235 24445
rect 7557 24440 13235 24442
rect 7557 24384 7562 24440
rect 7618 24384 13174 24440
rect 13230 24384 13235 24440
rect 7557 24382 13235 24384
rect 7557 24379 7623 24382
rect 13169 24379 13235 24382
rect 8845 24306 8911 24309
rect 11053 24306 11119 24309
rect 13905 24306 13971 24309
rect 8845 24304 13971 24306
rect 8845 24248 8850 24304
rect 8906 24248 11058 24304
rect 11114 24248 13910 24304
rect 13966 24248 13971 24304
rect 8845 24246 13971 24248
rect 8845 24243 8911 24246
rect 11053 24243 11119 24246
rect 13905 24243 13971 24246
rect 25497 24306 25563 24309
rect 28441 24306 28507 24309
rect 25497 24304 28507 24306
rect 25497 24248 25502 24304
rect 25558 24248 28446 24304
rect 28502 24248 28507 24304
rect 25497 24246 28507 24248
rect 25497 24243 25563 24246
rect 28441 24243 28507 24246
rect 3785 24170 3851 24173
rect 6361 24170 6427 24173
rect 7005 24170 7071 24173
rect 3785 24168 7071 24170
rect 3785 24112 3790 24168
rect 3846 24112 6366 24168
rect 6422 24112 7010 24168
rect 7066 24112 7071 24168
rect 3785 24110 7071 24112
rect 3785 24107 3851 24110
rect 6361 24107 6427 24110
rect 7005 24107 7071 24110
rect 8937 24170 9003 24173
rect 14641 24170 14707 24173
rect 16113 24170 16179 24173
rect 8937 24168 16179 24170
rect 8937 24112 8942 24168
rect 8998 24112 14646 24168
rect 14702 24112 16118 24168
rect 16174 24112 16179 24168
rect 8937 24110 16179 24112
rect 8937 24107 9003 24110
rect 14641 24107 14707 24110
rect 16113 24107 16179 24110
rect 4208 23968 4528 23969
rect 0 23898 800 23928
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 1577 23898 1643 23901
rect 0 23896 1643 23898
rect 0 23840 1582 23896
rect 1638 23840 1643 23896
rect 0 23838 1643 23840
rect 0 23808 800 23838
rect 1577 23835 1643 23838
rect 15377 23898 15443 23901
rect 38852 23898 39652 23928
rect 15377 23896 16866 23898
rect 15377 23840 15382 23896
rect 15438 23840 16866 23896
rect 15377 23838 16866 23840
rect 15377 23835 15443 23838
rect 3417 23762 3483 23765
rect 7557 23762 7623 23765
rect 16806 23764 16866 23838
rect 35390 23838 39652 23898
rect 3417 23760 7623 23762
rect 3417 23704 3422 23760
rect 3478 23704 7562 23760
rect 7618 23704 7623 23760
rect 3417 23702 7623 23704
rect 3417 23699 3483 23702
rect 7557 23699 7623 23702
rect 16798 23700 16804 23764
rect 16868 23762 16874 23764
rect 24853 23762 24919 23765
rect 27061 23762 27127 23765
rect 16868 23760 27127 23762
rect 16868 23704 24858 23760
rect 24914 23704 27066 23760
rect 27122 23704 27127 23760
rect 16868 23702 27127 23704
rect 16868 23700 16874 23702
rect 24853 23699 24919 23702
rect 27061 23699 27127 23702
rect 34513 23762 34579 23765
rect 35390 23762 35450 23838
rect 38852 23808 39652 23838
rect 34513 23760 35450 23762
rect 34513 23704 34518 23760
rect 34574 23704 35450 23760
rect 34513 23702 35450 23704
rect 34513 23699 34579 23702
rect 3049 23626 3115 23629
rect 8937 23626 9003 23629
rect 3049 23624 9003 23626
rect 3049 23568 3054 23624
rect 3110 23568 8942 23624
rect 8998 23568 9003 23624
rect 3049 23566 9003 23568
rect 3049 23563 3115 23566
rect 8937 23563 9003 23566
rect 9121 23626 9187 23629
rect 14733 23626 14799 23629
rect 19885 23626 19951 23629
rect 9121 23624 19951 23626
rect 9121 23568 9126 23624
rect 9182 23568 14738 23624
rect 14794 23568 19890 23624
rect 19946 23568 19951 23624
rect 9121 23566 19951 23568
rect 9121 23563 9187 23566
rect 14733 23563 14799 23566
rect 19885 23563 19951 23566
rect 25313 23626 25379 23629
rect 33869 23626 33935 23629
rect 25313 23624 33935 23626
rect 25313 23568 25318 23624
rect 25374 23568 33874 23624
rect 33930 23568 33935 23624
rect 25313 23566 33935 23568
rect 25313 23563 25379 23566
rect 33869 23563 33935 23566
rect 3877 23490 3943 23493
rect 7189 23490 7255 23493
rect 3877 23488 7255 23490
rect 3877 23432 3882 23488
rect 3938 23432 7194 23488
rect 7250 23432 7255 23488
rect 3877 23430 7255 23432
rect 3877 23427 3943 23430
rect 7189 23427 7255 23430
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 3877 23354 3943 23357
rect 7649 23354 7715 23357
rect 3877 23352 7715 23354
rect 3877 23296 3882 23352
rect 3938 23296 7654 23352
rect 7710 23296 7715 23352
rect 3877 23294 7715 23296
rect 3877 23291 3943 23294
rect 7649 23291 7715 23294
rect 24393 23354 24459 23357
rect 26233 23354 26299 23357
rect 24393 23352 26299 23354
rect 24393 23296 24398 23352
rect 24454 23296 26238 23352
rect 26294 23296 26299 23352
rect 24393 23294 26299 23296
rect 24393 23291 24459 23294
rect 26233 23291 26299 23294
rect 0 23218 800 23248
rect 1945 23218 2011 23221
rect 0 23216 2011 23218
rect 0 23160 1950 23216
rect 2006 23160 2011 23216
rect 0 23158 2011 23160
rect 0 23128 800 23158
rect 1945 23155 2011 23158
rect 30189 23218 30255 23221
rect 37365 23218 37431 23221
rect 30189 23216 37431 23218
rect 30189 23160 30194 23216
rect 30250 23160 37370 23216
rect 37426 23160 37431 23216
rect 30189 23158 37431 23160
rect 30189 23155 30255 23158
rect 37365 23155 37431 23158
rect 3969 23082 4035 23085
rect 6637 23082 6703 23085
rect 15285 23082 15351 23085
rect 16297 23082 16363 23085
rect 3969 23080 16363 23082
rect 3969 23024 3974 23080
rect 4030 23024 6642 23080
rect 6698 23024 15290 23080
rect 15346 23024 16302 23080
rect 16358 23024 16363 23080
rect 3969 23022 16363 23024
rect 3969 23019 4035 23022
rect 6637 23019 6703 23022
rect 15285 23019 15351 23022
rect 16297 23019 16363 23022
rect 18689 23082 18755 23085
rect 34697 23082 34763 23085
rect 18689 23080 34763 23082
rect 18689 23024 18694 23080
rect 18750 23024 34702 23080
rect 34758 23024 34763 23080
rect 18689 23022 34763 23024
rect 18689 23019 18755 23022
rect 34697 23019 34763 23022
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 8937 22810 9003 22813
rect 16757 22810 16823 22813
rect 20253 22810 20319 22813
rect 8937 22808 20319 22810
rect 8937 22752 8942 22808
rect 8998 22752 16762 22808
rect 16818 22752 20258 22808
rect 20314 22752 20319 22808
rect 8937 22750 20319 22752
rect 8937 22747 9003 22750
rect 16757 22747 16823 22750
rect 20253 22747 20319 22750
rect 3693 22674 3759 22677
rect 9213 22674 9279 22677
rect 3693 22672 9279 22674
rect 3693 22616 3698 22672
rect 3754 22616 9218 22672
rect 9274 22616 9279 22672
rect 3693 22614 9279 22616
rect 3693 22611 3759 22614
rect 9213 22611 9279 22614
rect 10777 22674 10843 22677
rect 12433 22674 12499 22677
rect 10777 22672 12499 22674
rect 10777 22616 10782 22672
rect 10838 22616 12438 22672
rect 12494 22616 12499 22672
rect 10777 22614 12499 22616
rect 10777 22611 10843 22614
rect 12433 22611 12499 22614
rect 16062 22612 16068 22676
rect 16132 22674 16138 22676
rect 16481 22674 16547 22677
rect 16132 22672 16547 22674
rect 16132 22616 16486 22672
rect 16542 22616 16547 22672
rect 16132 22614 16547 22616
rect 16132 22612 16138 22614
rect 16481 22611 16547 22614
rect 32949 22674 33015 22677
rect 37273 22674 37339 22677
rect 32949 22672 37339 22674
rect 32949 22616 32954 22672
rect 33010 22616 37278 22672
rect 37334 22616 37339 22672
rect 32949 22614 37339 22616
rect 32949 22611 33015 22614
rect 37273 22611 37339 22614
rect 7189 22538 7255 22541
rect 16113 22538 16179 22541
rect 16573 22538 16639 22541
rect 7189 22536 16639 22538
rect 7189 22480 7194 22536
rect 7250 22480 16118 22536
rect 16174 22480 16578 22536
rect 16634 22480 16639 22536
rect 7189 22478 16639 22480
rect 7189 22475 7255 22478
rect 16113 22475 16179 22478
rect 16573 22475 16639 22478
rect 25957 22538 26023 22541
rect 35341 22538 35407 22541
rect 25957 22536 35407 22538
rect 25957 22480 25962 22536
rect 26018 22480 35346 22536
rect 35402 22480 35407 22536
rect 25957 22478 35407 22480
rect 25957 22475 26023 22478
rect 35341 22475 35407 22478
rect 36077 22538 36143 22541
rect 38852 22538 39652 22568
rect 36077 22536 39652 22538
rect 36077 22480 36082 22536
rect 36138 22480 39652 22536
rect 36077 22478 39652 22480
rect 36077 22475 36143 22478
rect 38852 22448 39652 22478
rect 5165 22402 5231 22405
rect 7557 22402 7623 22405
rect 5165 22400 7623 22402
rect 5165 22344 5170 22400
rect 5226 22344 7562 22400
rect 7618 22344 7623 22400
rect 5165 22342 7623 22344
rect 5165 22339 5231 22342
rect 7557 22339 7623 22342
rect 9213 22402 9279 22405
rect 14089 22402 14155 22405
rect 9213 22400 14155 22402
rect 9213 22344 9218 22400
rect 9274 22344 14094 22400
rect 14150 22344 14155 22400
rect 9213 22342 14155 22344
rect 9213 22339 9279 22342
rect 14089 22339 14155 22342
rect 16481 22402 16547 22405
rect 16982 22402 16988 22404
rect 16481 22400 16988 22402
rect 16481 22344 16486 22400
rect 16542 22344 16988 22400
rect 16481 22342 16988 22344
rect 16481 22339 16547 22342
rect 16982 22340 16988 22342
rect 17052 22340 17058 22404
rect 27153 22402 27219 22405
rect 30373 22402 30439 22405
rect 27153 22400 30439 22402
rect 27153 22344 27158 22400
rect 27214 22344 30378 22400
rect 30434 22344 30439 22400
rect 27153 22342 30439 22344
rect 27153 22339 27219 22342
rect 30373 22339 30439 22342
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 4797 22266 4863 22269
rect 7097 22266 7163 22269
rect 9213 22266 9279 22269
rect 4797 22264 9279 22266
rect 4797 22208 4802 22264
rect 4858 22208 7102 22264
rect 7158 22208 9218 22264
rect 9274 22208 9279 22264
rect 4797 22206 9279 22208
rect 4797 22203 4863 22206
rect 7097 22203 7163 22206
rect 9213 22203 9279 22206
rect 28073 22266 28139 22269
rect 35433 22266 35499 22269
rect 28073 22264 35499 22266
rect 28073 22208 28078 22264
rect 28134 22208 35438 22264
rect 35494 22208 35499 22264
rect 28073 22206 35499 22208
rect 28073 22203 28139 22206
rect 35433 22203 35499 22206
rect 9581 22130 9647 22133
rect 9949 22130 10015 22133
rect 14641 22130 14707 22133
rect 9581 22128 14707 22130
rect 9581 22072 9586 22128
rect 9642 22072 9954 22128
rect 10010 22072 14646 22128
rect 14702 22072 14707 22128
rect 9581 22070 14707 22072
rect 9581 22067 9647 22070
rect 9949 22067 10015 22070
rect 14641 22067 14707 22070
rect 5073 21994 5139 21997
rect 5257 21994 5323 21997
rect 5073 21992 5323 21994
rect 5073 21936 5078 21992
rect 5134 21936 5262 21992
rect 5318 21936 5323 21992
rect 5073 21934 5323 21936
rect 5073 21931 5139 21934
rect 5257 21931 5323 21934
rect 9213 21994 9279 21997
rect 11697 21994 11763 21997
rect 9213 21992 11763 21994
rect 9213 21936 9218 21992
rect 9274 21936 11702 21992
rect 11758 21936 11763 21992
rect 9213 21934 11763 21936
rect 9213 21931 9279 21934
rect 11697 21931 11763 21934
rect 16798 21932 16804 21996
rect 16868 21994 16874 21996
rect 17033 21994 17099 21997
rect 16868 21992 17099 21994
rect 16868 21936 17038 21992
rect 17094 21936 17099 21992
rect 16868 21934 17099 21936
rect 16868 21932 16874 21934
rect 17033 21931 17099 21934
rect 29637 21994 29703 21997
rect 36261 21994 36327 21997
rect 29637 21992 36327 21994
rect 29637 21936 29642 21992
rect 29698 21936 36266 21992
rect 36322 21936 36327 21992
rect 29637 21934 36327 21936
rect 29637 21931 29703 21934
rect 36261 21931 36327 21934
rect 0 21858 800 21888
rect 2405 21858 2471 21861
rect 0 21856 2471 21858
rect 0 21800 2410 21856
rect 2466 21800 2471 21856
rect 0 21798 2471 21800
rect 0 21768 800 21798
rect 2405 21795 2471 21798
rect 8569 21858 8635 21861
rect 13261 21858 13327 21861
rect 8569 21856 13327 21858
rect 8569 21800 8574 21856
rect 8630 21800 13266 21856
rect 13322 21800 13327 21856
rect 8569 21798 13327 21800
rect 8569 21795 8635 21798
rect 13261 21795 13327 21798
rect 27337 21858 27403 21861
rect 30465 21858 30531 21861
rect 38852 21858 39652 21888
rect 27337 21856 30531 21858
rect 27337 21800 27342 21856
rect 27398 21800 30470 21856
rect 30526 21800 30531 21856
rect 27337 21798 30531 21800
rect 27337 21795 27403 21798
rect 30465 21795 30531 21798
rect 35390 21798 39652 21858
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 11237 21722 11303 21725
rect 17953 21722 18019 21725
rect 20897 21722 20963 21725
rect 21541 21722 21607 21725
rect 11237 21720 21607 21722
rect 11237 21664 11242 21720
rect 11298 21664 17958 21720
rect 18014 21664 20902 21720
rect 20958 21664 21546 21720
rect 21602 21664 21607 21720
rect 11237 21662 21607 21664
rect 11237 21659 11303 21662
rect 17953 21659 18019 21662
rect 20897 21659 20963 21662
rect 21541 21659 21607 21662
rect 3509 21586 3575 21589
rect 8661 21586 8727 21589
rect 3509 21584 8727 21586
rect 3509 21528 3514 21584
rect 3570 21528 8666 21584
rect 8722 21528 8727 21584
rect 3509 21526 8727 21528
rect 3509 21523 3575 21526
rect 8661 21523 8727 21526
rect 23841 21586 23907 21589
rect 26049 21586 26115 21589
rect 23841 21584 26115 21586
rect 23841 21528 23846 21584
rect 23902 21528 26054 21584
rect 26110 21528 26115 21584
rect 23841 21526 26115 21528
rect 23841 21523 23907 21526
rect 26049 21523 26115 21526
rect 7925 21450 7991 21453
rect 9949 21450 10015 21453
rect 12617 21450 12683 21453
rect 7925 21448 12683 21450
rect 7925 21392 7930 21448
rect 7986 21392 9954 21448
rect 10010 21392 12622 21448
rect 12678 21392 12683 21448
rect 7925 21390 12683 21392
rect 7925 21387 7991 21390
rect 9949 21387 10015 21390
rect 12617 21387 12683 21390
rect 19057 21450 19123 21453
rect 35390 21450 35450 21798
rect 38852 21768 39652 21798
rect 19057 21448 35450 21450
rect 19057 21392 19062 21448
rect 19118 21392 35450 21448
rect 19057 21390 35450 21392
rect 19057 21387 19123 21390
rect 8845 21314 8911 21317
rect 10133 21314 10199 21317
rect 14089 21314 14155 21317
rect 8845 21312 10199 21314
rect 8845 21256 8850 21312
rect 8906 21256 10138 21312
rect 10194 21256 10199 21312
rect 8845 21254 10199 21256
rect 8845 21251 8911 21254
rect 10133 21251 10199 21254
rect 10366 21312 14155 21314
rect 10366 21256 14094 21312
rect 14150 21256 14155 21312
rect 10366 21254 14155 21256
rect 0 21178 800 21208
rect 1669 21178 1735 21181
rect 0 21176 1735 21178
rect 0 21120 1674 21176
rect 1730 21120 1735 21176
rect 0 21118 1735 21120
rect 0 21088 800 21118
rect 1669 21115 1735 21118
rect 3877 21178 3943 21181
rect 7833 21178 7899 21181
rect 3877 21176 7899 21178
rect 3877 21120 3882 21176
rect 3938 21120 7838 21176
rect 7894 21120 7899 21176
rect 3877 21118 7899 21120
rect 3877 21115 3943 21118
rect 7833 21115 7899 21118
rect 8017 21178 8083 21181
rect 10366 21178 10426 21254
rect 14089 21251 14155 21254
rect 15193 21314 15259 21317
rect 18137 21314 18203 21317
rect 15193 21312 18203 21314
rect 15193 21256 15198 21312
rect 15254 21256 18142 21312
rect 18198 21256 18203 21312
rect 15193 21254 18203 21256
rect 15193 21251 15259 21254
rect 18137 21251 18203 21254
rect 33317 21314 33383 21317
rect 37457 21314 37523 21317
rect 33317 21312 37523 21314
rect 33317 21256 33322 21312
rect 33378 21256 37462 21312
rect 37518 21256 37523 21312
rect 33317 21254 37523 21256
rect 33317 21251 33383 21254
rect 37457 21251 37523 21254
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 8017 21176 10426 21178
rect 8017 21120 8022 21176
rect 8078 21120 10426 21176
rect 8017 21118 10426 21120
rect 34697 21178 34763 21181
rect 38852 21178 39652 21208
rect 34697 21176 39652 21178
rect 34697 21120 34702 21176
rect 34758 21120 39652 21176
rect 34697 21118 39652 21120
rect 8017 21115 8083 21118
rect 34697 21115 34763 21118
rect 38852 21088 39652 21118
rect 10501 21042 10567 21045
rect 14641 21042 14707 21045
rect 10501 21040 14707 21042
rect 10501 20984 10506 21040
rect 10562 20984 14646 21040
rect 14702 20984 14707 21040
rect 10501 20982 14707 20984
rect 10501 20979 10567 20982
rect 14641 20979 14707 20982
rect 13353 20906 13419 20909
rect 16941 20906 17007 20909
rect 13353 20904 17007 20906
rect 13353 20848 13358 20904
rect 13414 20848 16946 20904
rect 17002 20848 17007 20904
rect 13353 20846 17007 20848
rect 13353 20843 13419 20846
rect 16941 20843 17007 20846
rect 21633 20906 21699 20909
rect 30189 20906 30255 20909
rect 21633 20904 30255 20906
rect 21633 20848 21638 20904
rect 21694 20848 30194 20904
rect 30250 20848 30255 20904
rect 21633 20846 30255 20848
rect 21633 20843 21699 20846
rect 30189 20843 30255 20846
rect 5257 20770 5323 20773
rect 7373 20770 7439 20773
rect 5257 20768 7439 20770
rect 5257 20712 5262 20768
rect 5318 20712 7378 20768
rect 7434 20712 7439 20768
rect 5257 20710 7439 20712
rect 5257 20707 5323 20710
rect 7373 20707 7439 20710
rect 17769 20770 17835 20773
rect 21357 20770 21423 20773
rect 17769 20768 21423 20770
rect 17769 20712 17774 20768
rect 17830 20712 21362 20768
rect 21418 20712 21423 20768
rect 17769 20710 21423 20712
rect 17769 20707 17835 20710
rect 21357 20707 21423 20710
rect 26693 20770 26759 20773
rect 31477 20770 31543 20773
rect 26693 20768 31543 20770
rect 26693 20712 26698 20768
rect 26754 20712 31482 20768
rect 31538 20712 31543 20768
rect 26693 20710 31543 20712
rect 26693 20707 26759 20710
rect 31477 20707 31543 20710
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 6085 20634 6151 20637
rect 8661 20634 8727 20637
rect 11329 20634 11395 20637
rect 6085 20632 11395 20634
rect 6085 20576 6090 20632
rect 6146 20576 8666 20632
rect 8722 20576 11334 20632
rect 11390 20576 11395 20632
rect 6085 20574 11395 20576
rect 6085 20571 6151 20574
rect 8661 20571 8727 20574
rect 11329 20571 11395 20574
rect 11881 20634 11947 20637
rect 20253 20634 20319 20637
rect 21173 20634 21239 20637
rect 11881 20632 21239 20634
rect 11881 20576 11886 20632
rect 11942 20576 20258 20632
rect 20314 20576 21178 20632
rect 21234 20576 21239 20632
rect 11881 20574 21239 20576
rect 11881 20571 11947 20574
rect 20253 20571 20319 20574
rect 21173 20571 21239 20574
rect 23289 20634 23355 20637
rect 25589 20634 25655 20637
rect 23289 20632 25655 20634
rect 23289 20576 23294 20632
rect 23350 20576 25594 20632
rect 25650 20576 25655 20632
rect 23289 20574 25655 20576
rect 23289 20571 23355 20574
rect 25589 20571 25655 20574
rect 28073 20634 28139 20637
rect 30465 20634 30531 20637
rect 33869 20634 33935 20637
rect 28073 20632 33935 20634
rect 28073 20576 28078 20632
rect 28134 20576 30470 20632
rect 30526 20576 33874 20632
rect 33930 20576 33935 20632
rect 28073 20574 33935 20576
rect 28073 20571 28139 20574
rect 30465 20571 30531 20574
rect 33869 20571 33935 20574
rect 0 20498 800 20528
rect 2589 20498 2655 20501
rect 0 20496 2655 20498
rect 0 20440 2594 20496
rect 2650 20440 2655 20496
rect 0 20438 2655 20440
rect 0 20408 800 20438
rect 2589 20435 2655 20438
rect 4613 20498 4679 20501
rect 8201 20498 8267 20501
rect 16021 20498 16087 20501
rect 4613 20496 16087 20498
rect 4613 20440 4618 20496
rect 4674 20440 8206 20496
rect 8262 20440 16026 20496
rect 16082 20440 16087 20496
rect 4613 20438 16087 20440
rect 4613 20435 4679 20438
rect 8201 20435 8267 20438
rect 16021 20435 16087 20438
rect 16665 20498 16731 20501
rect 25957 20498 26023 20501
rect 16665 20496 26023 20498
rect 16665 20440 16670 20496
rect 16726 20440 25962 20496
rect 26018 20440 26023 20496
rect 16665 20438 26023 20440
rect 16665 20435 16731 20438
rect 25957 20435 26023 20438
rect 27889 20498 27955 20501
rect 31661 20498 31727 20501
rect 27889 20496 31727 20498
rect 27889 20440 27894 20496
rect 27950 20440 31666 20496
rect 31722 20440 31727 20496
rect 27889 20438 31727 20440
rect 27889 20435 27955 20438
rect 31661 20435 31727 20438
rect 20621 20362 20687 20365
rect 34053 20362 34119 20365
rect 20621 20360 34119 20362
rect 20621 20304 20626 20360
rect 20682 20304 34058 20360
rect 34114 20304 34119 20360
rect 20621 20302 34119 20304
rect 20621 20299 20687 20302
rect 34053 20299 34119 20302
rect 24485 20226 24551 20229
rect 25221 20226 25287 20229
rect 29545 20226 29611 20229
rect 24485 20224 29611 20226
rect 24485 20168 24490 20224
rect 24546 20168 25226 20224
rect 25282 20168 29550 20224
rect 29606 20168 29611 20224
rect 24485 20166 29611 20168
rect 24485 20163 24551 20166
rect 25221 20163 25287 20166
rect 29545 20163 29611 20166
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 3969 20090 4035 20093
rect 6177 20090 6243 20093
rect 3969 20088 6243 20090
rect 3969 20032 3974 20088
rect 4030 20032 6182 20088
rect 6238 20032 6243 20088
rect 3969 20030 6243 20032
rect 3969 20027 4035 20030
rect 6177 20027 6243 20030
rect 7373 20090 7439 20093
rect 9438 20090 9444 20092
rect 7373 20088 9444 20090
rect 7373 20032 7378 20088
rect 7434 20032 9444 20088
rect 7373 20030 9444 20032
rect 7373 20027 7439 20030
rect 9438 20028 9444 20030
rect 9508 20090 9514 20092
rect 12249 20090 12315 20093
rect 17309 20090 17375 20093
rect 9508 20030 11852 20090
rect 9508 20028 9514 20030
rect 11792 19957 11852 20030
rect 12249 20088 17375 20090
rect 12249 20032 12254 20088
rect 12310 20032 17314 20088
rect 17370 20032 17375 20088
rect 12249 20030 17375 20032
rect 12249 20027 12315 20030
rect 17309 20027 17375 20030
rect 5257 19954 5323 19957
rect 5625 19954 5691 19957
rect 11605 19954 11671 19957
rect 5257 19952 11671 19954
rect 5257 19896 5262 19952
rect 5318 19896 5630 19952
rect 5686 19896 11610 19952
rect 11666 19896 11671 19952
rect 5257 19894 11671 19896
rect 5257 19891 5323 19894
rect 5625 19891 5691 19894
rect 11605 19891 11671 19894
rect 11789 19952 11855 19957
rect 11789 19896 11794 19952
rect 11850 19896 11855 19952
rect 11789 19891 11855 19896
rect 19241 19954 19307 19957
rect 23565 19954 23631 19957
rect 19241 19952 23631 19954
rect 19241 19896 19246 19952
rect 19302 19896 23570 19952
rect 23626 19896 23631 19952
rect 19241 19894 23631 19896
rect 19241 19891 19307 19894
rect 23565 19891 23631 19894
rect 24761 19954 24827 19957
rect 25957 19954 26023 19957
rect 24761 19952 26023 19954
rect 24761 19896 24766 19952
rect 24822 19896 25962 19952
rect 26018 19896 26023 19952
rect 24761 19894 26023 19896
rect 24761 19891 24827 19894
rect 25957 19891 26023 19894
rect 35157 19818 35223 19821
rect 38852 19818 39652 19848
rect 35157 19816 39652 19818
rect 35157 19760 35162 19816
rect 35218 19760 39652 19816
rect 35157 19758 39652 19760
rect 35157 19755 35223 19758
rect 38852 19728 39652 19758
rect 16982 19620 16988 19684
rect 17052 19682 17058 19684
rect 17217 19682 17283 19685
rect 17052 19680 17283 19682
rect 17052 19624 17222 19680
rect 17278 19624 17283 19680
rect 17052 19622 17283 19624
rect 17052 19620 17058 19622
rect 17217 19619 17283 19622
rect 25405 19682 25471 19685
rect 27061 19682 27127 19685
rect 25405 19680 27127 19682
rect 25405 19624 25410 19680
rect 25466 19624 27066 19680
rect 27122 19624 27127 19680
rect 25405 19622 27127 19624
rect 25405 19619 25471 19622
rect 27061 19619 27127 19622
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 8845 19546 8911 19549
rect 21265 19546 21331 19549
rect 8845 19544 21331 19546
rect 8845 19488 8850 19544
rect 8906 19488 21270 19544
rect 21326 19488 21331 19544
rect 8845 19486 21331 19488
rect 8845 19483 8911 19486
rect 21265 19483 21331 19486
rect 23933 19546 23999 19549
rect 33041 19546 33107 19549
rect 23933 19544 33107 19546
rect 23933 19488 23938 19544
rect 23994 19488 33046 19544
rect 33102 19488 33107 19544
rect 23933 19486 33107 19488
rect 23933 19483 23999 19486
rect 33041 19483 33107 19486
rect 3141 19410 3207 19413
rect 3417 19410 3483 19413
rect 3141 19408 3483 19410
rect 3141 19352 3146 19408
rect 3202 19352 3422 19408
rect 3478 19352 3483 19408
rect 3141 19350 3483 19352
rect 3141 19347 3207 19350
rect 3417 19347 3483 19350
rect 4061 19410 4127 19413
rect 7598 19410 7604 19412
rect 4061 19408 7604 19410
rect 4061 19352 4066 19408
rect 4122 19352 7604 19408
rect 4061 19350 7604 19352
rect 4061 19347 4127 19350
rect 7598 19348 7604 19350
rect 7668 19348 7674 19412
rect 10777 19410 10843 19413
rect 14641 19410 14707 19413
rect 10777 19408 14707 19410
rect 10777 19352 10782 19408
rect 10838 19352 14646 19408
rect 14702 19352 14707 19408
rect 10777 19350 14707 19352
rect 10777 19347 10843 19350
rect 14641 19347 14707 19350
rect 16430 19348 16436 19412
rect 16500 19410 16506 19412
rect 18597 19410 18663 19413
rect 16500 19408 18663 19410
rect 16500 19352 18602 19408
rect 18658 19352 18663 19408
rect 16500 19350 18663 19352
rect 16500 19348 16506 19350
rect 18597 19347 18663 19350
rect 3877 19274 3943 19277
rect 7189 19274 7255 19277
rect 12617 19274 12683 19277
rect 3877 19272 12683 19274
rect 3877 19216 3882 19272
rect 3938 19216 7194 19272
rect 7250 19216 12622 19272
rect 12678 19216 12683 19272
rect 3877 19214 12683 19216
rect 3877 19211 3943 19214
rect 7189 19211 7255 19214
rect 12617 19211 12683 19214
rect 12893 19274 12959 19277
rect 16941 19276 17007 19277
rect 16941 19274 16988 19276
rect 12893 19272 14842 19274
rect 12893 19216 12898 19272
rect 12954 19216 14842 19272
rect 12893 19214 14842 19216
rect 16896 19272 16988 19274
rect 16896 19216 16946 19272
rect 16896 19214 16988 19216
rect 12893 19211 12959 19214
rect 0 19138 800 19168
rect 1761 19138 1827 19141
rect 0 19136 1827 19138
rect 0 19080 1766 19136
rect 1822 19080 1827 19136
rect 0 19078 1827 19080
rect 0 19048 800 19078
rect 1761 19075 1827 19078
rect 3509 19138 3575 19141
rect 7649 19138 7715 19141
rect 7925 19138 7991 19141
rect 3509 19136 7991 19138
rect 3509 19080 3514 19136
rect 3570 19080 7654 19136
rect 7710 19080 7930 19136
rect 7986 19080 7991 19136
rect 3509 19078 7991 19080
rect 3509 19075 3575 19078
rect 7649 19075 7715 19078
rect 7925 19075 7991 19078
rect 9857 19138 9923 19141
rect 14641 19138 14707 19141
rect 9857 19136 14707 19138
rect 9857 19080 9862 19136
rect 9918 19080 14646 19136
rect 14702 19080 14707 19136
rect 9857 19078 14707 19080
rect 14782 19138 14842 19214
rect 16941 19212 16988 19214
rect 17052 19212 17058 19276
rect 17125 19274 17191 19277
rect 17585 19274 17651 19277
rect 17125 19272 17651 19274
rect 17125 19216 17130 19272
rect 17186 19216 17590 19272
rect 17646 19216 17651 19272
rect 17125 19214 17651 19216
rect 16941 19211 17007 19212
rect 17125 19211 17191 19214
rect 17585 19211 17651 19214
rect 24301 19274 24367 19277
rect 26233 19274 26299 19277
rect 24301 19272 26299 19274
rect 24301 19216 24306 19272
rect 24362 19216 26238 19272
rect 26294 19216 26299 19272
rect 24301 19214 26299 19216
rect 24301 19211 24367 19214
rect 26233 19211 26299 19214
rect 30281 19274 30347 19277
rect 33501 19274 33567 19277
rect 30281 19272 33567 19274
rect 30281 19216 30286 19272
rect 30342 19216 33506 19272
rect 33562 19216 33567 19272
rect 30281 19214 33567 19216
rect 30281 19211 30347 19214
rect 33501 19211 33567 19214
rect 15469 19138 15535 19141
rect 18597 19138 18663 19141
rect 14782 19136 18663 19138
rect 14782 19080 15474 19136
rect 15530 19080 18602 19136
rect 18658 19080 18663 19136
rect 14782 19078 18663 19080
rect 9857 19075 9923 19078
rect 14641 19075 14707 19078
rect 15469 19075 15535 19078
rect 18597 19075 18663 19078
rect 34053 19138 34119 19141
rect 38852 19138 39652 19168
rect 34053 19136 39652 19138
rect 34053 19080 34058 19136
rect 34114 19080 39652 19136
rect 34053 19078 39652 19080
rect 34053 19075 34119 19078
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 38852 19048 39652 19078
rect 19568 19007 19888 19008
rect 4797 19002 4863 19005
rect 10685 19002 10751 19005
rect 4797 19000 10751 19002
rect 4797 18944 4802 19000
rect 4858 18944 10690 19000
rect 10746 18944 10751 19000
rect 4797 18942 10751 18944
rect 4797 18939 4863 18942
rect 10685 18939 10751 18942
rect 14181 19002 14247 19005
rect 16297 19002 16363 19005
rect 18413 19002 18479 19005
rect 14181 19000 18479 19002
rect 14181 18944 14186 19000
rect 14242 18944 16302 19000
rect 16358 18944 18418 19000
rect 18474 18944 18479 19000
rect 14181 18942 18479 18944
rect 14181 18939 14247 18942
rect 16297 18939 16363 18942
rect 18413 18939 18479 18942
rect 26969 19002 27035 19005
rect 31201 19002 31267 19005
rect 26969 19000 31267 19002
rect 26969 18944 26974 19000
rect 27030 18944 31206 19000
rect 31262 18944 31267 19000
rect 26969 18942 31267 18944
rect 26969 18939 27035 18942
rect 31201 18939 31267 18942
rect 4889 18866 4955 18869
rect 7925 18866 7991 18869
rect 16205 18866 16271 18869
rect 4889 18864 16271 18866
rect 4889 18808 4894 18864
rect 4950 18808 7930 18864
rect 7986 18808 16210 18864
rect 16266 18808 16271 18864
rect 4889 18806 16271 18808
rect 4889 18803 4955 18806
rect 7925 18803 7991 18806
rect 16205 18803 16271 18806
rect 16941 18866 17007 18869
rect 18137 18866 18203 18869
rect 18454 18866 18460 18868
rect 16941 18864 18460 18866
rect 16941 18808 16946 18864
rect 17002 18808 18142 18864
rect 18198 18808 18460 18864
rect 16941 18806 18460 18808
rect 16941 18803 17007 18806
rect 18137 18803 18203 18806
rect 18454 18804 18460 18806
rect 18524 18804 18530 18868
rect 24301 18866 24367 18869
rect 34789 18866 34855 18869
rect 35065 18866 35131 18869
rect 24301 18864 35131 18866
rect 24301 18808 24306 18864
rect 24362 18808 34794 18864
rect 34850 18808 35070 18864
rect 35126 18808 35131 18864
rect 24301 18806 35131 18808
rect 24301 18803 24367 18806
rect 34789 18803 34855 18806
rect 35065 18803 35131 18806
rect 3049 18730 3115 18733
rect 4429 18730 4495 18733
rect 7189 18730 7255 18733
rect 11697 18730 11763 18733
rect 3049 18728 7114 18730
rect 3049 18672 3054 18728
rect 3110 18672 4434 18728
rect 4490 18672 7114 18728
rect 3049 18670 7114 18672
rect 3049 18667 3115 18670
rect 4429 18667 4495 18670
rect 7054 18594 7114 18670
rect 7189 18728 11763 18730
rect 7189 18672 7194 18728
rect 7250 18672 11702 18728
rect 11758 18672 11763 18728
rect 7189 18670 11763 18672
rect 7189 18667 7255 18670
rect 11697 18667 11763 18670
rect 9213 18594 9279 18597
rect 17217 18594 17283 18597
rect 7054 18592 17283 18594
rect 7054 18536 9218 18592
rect 9274 18536 17222 18592
rect 17278 18536 17283 18592
rect 7054 18534 17283 18536
rect 9213 18531 9279 18534
rect 17217 18531 17283 18534
rect 4208 18528 4528 18529
rect 0 18458 800 18488
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 4061 18458 4127 18461
rect 0 18456 4127 18458
rect 0 18400 4066 18456
rect 4122 18400 4127 18456
rect 0 18398 4127 18400
rect 0 18368 800 18398
rect 4061 18395 4127 18398
rect 5257 18458 5323 18461
rect 7741 18458 7807 18461
rect 5257 18456 7807 18458
rect 5257 18400 5262 18456
rect 5318 18400 7746 18456
rect 7802 18400 7807 18456
rect 5257 18398 7807 18400
rect 5257 18395 5323 18398
rect 7741 18395 7807 18398
rect 27797 18458 27863 18461
rect 29637 18458 29703 18461
rect 27797 18456 29703 18458
rect 27797 18400 27802 18456
rect 27858 18400 29642 18456
rect 29698 18400 29703 18456
rect 27797 18398 29703 18400
rect 27797 18395 27863 18398
rect 29637 18395 29703 18398
rect 11329 18322 11395 18325
rect 15193 18322 15259 18325
rect 11329 18320 15259 18322
rect 11329 18264 11334 18320
rect 11390 18264 15198 18320
rect 15254 18264 15259 18320
rect 11329 18262 15259 18264
rect 11329 18259 11395 18262
rect 15193 18259 15259 18262
rect 28073 18322 28139 18325
rect 30649 18322 30715 18325
rect 28073 18320 30715 18322
rect 28073 18264 28078 18320
rect 28134 18264 30654 18320
rect 30710 18264 30715 18320
rect 28073 18262 30715 18264
rect 28073 18259 28139 18262
rect 30649 18259 30715 18262
rect 10777 18186 10843 18189
rect 16665 18186 16731 18189
rect 10777 18184 16731 18186
rect 10777 18128 10782 18184
rect 10838 18128 16670 18184
rect 16726 18128 16731 18184
rect 10777 18126 16731 18128
rect 10777 18123 10843 18126
rect 16665 18123 16731 18126
rect 17350 18124 17356 18188
rect 17420 18186 17426 18188
rect 17769 18186 17835 18189
rect 17420 18184 17835 18186
rect 17420 18128 17774 18184
rect 17830 18128 17835 18184
rect 17420 18126 17835 18128
rect 17420 18124 17426 18126
rect 17769 18123 17835 18126
rect 18597 18186 18663 18189
rect 23933 18186 23999 18189
rect 18597 18184 23999 18186
rect 18597 18128 18602 18184
rect 18658 18128 23938 18184
rect 23994 18128 23999 18184
rect 18597 18126 23999 18128
rect 18597 18123 18663 18126
rect 23933 18123 23999 18126
rect 8293 18050 8359 18053
rect 9673 18050 9739 18053
rect 13261 18050 13327 18053
rect 8293 18048 8724 18050
rect 8293 17992 8298 18048
rect 8354 17992 8724 18048
rect 8293 17990 8724 17992
rect 8293 17987 8359 17990
rect 8664 17917 8724 17990
rect 9673 18048 13327 18050
rect 9673 17992 9678 18048
rect 9734 17992 13266 18048
rect 13322 17992 13327 18048
rect 9673 17990 13327 17992
rect 9673 17987 9739 17990
rect 13261 17987 13327 17990
rect 14733 18050 14799 18053
rect 17953 18050 18019 18053
rect 19425 18050 19491 18053
rect 14733 18048 19491 18050
rect 14733 17992 14738 18048
rect 14794 17992 17958 18048
rect 18014 17992 19430 18048
rect 19486 17992 19491 18048
rect 14733 17990 19491 17992
rect 14733 17987 14799 17990
rect 17953 17987 18019 17990
rect 19425 17987 19491 17990
rect 28993 18050 29059 18053
rect 29126 18050 29132 18052
rect 28993 18048 29132 18050
rect 28993 17992 28998 18048
rect 29054 17992 29132 18048
rect 28993 17990 29132 17992
rect 28993 17987 29059 17990
rect 29126 17988 29132 17990
rect 29196 17988 29202 18052
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 4613 17914 4679 17917
rect 7925 17914 7991 17917
rect 8293 17914 8359 17917
rect 4613 17912 8359 17914
rect 4613 17856 4618 17912
rect 4674 17856 7930 17912
rect 7986 17856 8298 17912
rect 8354 17856 8359 17912
rect 4613 17854 8359 17856
rect 4613 17851 4679 17854
rect 7925 17851 7991 17854
rect 8293 17851 8359 17854
rect 8661 17912 8727 17917
rect 8661 17856 8666 17912
rect 8722 17856 8727 17912
rect 8661 17851 8727 17856
rect 11513 17914 11579 17917
rect 15561 17914 15627 17917
rect 31385 17914 31451 17917
rect 34513 17914 34579 17917
rect 11513 17912 18200 17914
rect 11513 17856 11518 17912
rect 11574 17856 15566 17912
rect 15622 17856 18200 17912
rect 11513 17854 18200 17856
rect 11513 17851 11579 17854
rect 15561 17851 15627 17854
rect 0 17778 800 17808
rect 18140 17781 18200 17854
rect 31385 17912 34579 17914
rect 31385 17856 31390 17912
rect 31446 17856 34518 17912
rect 34574 17856 34579 17912
rect 31385 17854 34579 17856
rect 31385 17851 31451 17854
rect 34513 17851 34579 17854
rect 1945 17778 2011 17781
rect 0 17776 2011 17778
rect 0 17720 1950 17776
rect 2006 17720 2011 17776
rect 0 17718 2011 17720
rect 0 17688 800 17718
rect 1945 17715 2011 17718
rect 5901 17778 5967 17781
rect 12801 17778 12867 17781
rect 5901 17776 12867 17778
rect 5901 17720 5906 17776
rect 5962 17720 12806 17776
rect 12862 17720 12867 17776
rect 5901 17718 12867 17720
rect 5901 17715 5967 17718
rect 12801 17715 12867 17718
rect 18137 17776 18203 17781
rect 18137 17720 18142 17776
rect 18198 17720 18203 17776
rect 18137 17715 18203 17720
rect 23105 17778 23171 17781
rect 27705 17778 27771 17781
rect 23105 17776 27771 17778
rect 23105 17720 23110 17776
rect 23166 17720 27710 17776
rect 27766 17720 27771 17776
rect 23105 17718 27771 17720
rect 23105 17715 23171 17718
rect 27705 17715 27771 17718
rect 29085 17778 29151 17781
rect 30373 17778 30439 17781
rect 29085 17776 30439 17778
rect 29085 17720 29090 17776
rect 29146 17720 30378 17776
rect 30434 17720 30439 17776
rect 29085 17718 30439 17720
rect 29085 17715 29151 17718
rect 30373 17715 30439 17718
rect 35525 17778 35591 17781
rect 38852 17778 39652 17808
rect 35525 17776 39652 17778
rect 35525 17720 35530 17776
rect 35586 17720 39652 17776
rect 35525 17718 39652 17720
rect 35525 17715 35591 17718
rect 38852 17688 39652 17718
rect 4521 17642 4587 17645
rect 8017 17642 8083 17645
rect 4521 17640 8083 17642
rect 4521 17584 4526 17640
rect 4582 17584 8022 17640
rect 8078 17584 8083 17640
rect 4521 17582 8083 17584
rect 4521 17579 4587 17582
rect 8017 17579 8083 17582
rect 8385 17642 8451 17645
rect 10685 17642 10751 17645
rect 8385 17640 10751 17642
rect 8385 17584 8390 17640
rect 8446 17584 10690 17640
rect 10746 17584 10751 17640
rect 8385 17582 10751 17584
rect 8385 17579 8451 17582
rect 10685 17579 10751 17582
rect 14733 17642 14799 17645
rect 20161 17642 20227 17645
rect 14733 17640 20227 17642
rect 14733 17584 14738 17640
rect 14794 17584 20166 17640
rect 20222 17584 20227 17640
rect 14733 17582 20227 17584
rect 14733 17579 14799 17582
rect 20161 17579 20227 17582
rect 21725 17642 21791 17645
rect 24209 17642 24275 17645
rect 21725 17640 24275 17642
rect 21725 17584 21730 17640
rect 21786 17584 24214 17640
rect 24270 17584 24275 17640
rect 21725 17582 24275 17584
rect 21725 17579 21791 17582
rect 24209 17579 24275 17582
rect 27429 17642 27495 17645
rect 29545 17642 29611 17645
rect 27429 17640 29611 17642
rect 27429 17584 27434 17640
rect 27490 17584 29550 17640
rect 29606 17584 29611 17640
rect 27429 17582 29611 17584
rect 27429 17579 27495 17582
rect 29545 17579 29611 17582
rect 9581 17506 9647 17509
rect 12709 17506 12775 17509
rect 9581 17504 12775 17506
rect 9581 17448 9586 17504
rect 9642 17448 12714 17504
rect 12770 17448 12775 17504
rect 9581 17446 12775 17448
rect 9581 17443 9647 17446
rect 12709 17443 12775 17446
rect 12893 17506 12959 17509
rect 17309 17506 17375 17509
rect 12893 17504 17375 17506
rect 12893 17448 12898 17504
rect 12954 17448 17314 17504
rect 17370 17448 17375 17504
rect 12893 17446 17375 17448
rect 12893 17443 12959 17446
rect 17309 17443 17375 17446
rect 25497 17506 25563 17509
rect 29913 17506 29979 17509
rect 33777 17506 33843 17509
rect 25497 17504 33843 17506
rect 25497 17448 25502 17504
rect 25558 17448 29918 17504
rect 29974 17448 33782 17504
rect 33838 17448 33843 17504
rect 25497 17446 33843 17448
rect 25497 17443 25563 17446
rect 29913 17443 29979 17446
rect 33777 17443 33843 17446
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 26233 17370 26299 17373
rect 26509 17370 26575 17373
rect 31385 17370 31451 17373
rect 26233 17368 31451 17370
rect 26233 17312 26238 17368
rect 26294 17312 26514 17368
rect 26570 17312 31390 17368
rect 31446 17312 31451 17368
rect 26233 17310 31451 17312
rect 26233 17307 26299 17310
rect 26509 17307 26575 17310
rect 31385 17307 31451 17310
rect 6269 17234 6335 17237
rect 8845 17234 8911 17237
rect 6269 17232 8911 17234
rect 6269 17176 6274 17232
rect 6330 17176 8850 17232
rect 8906 17176 8911 17232
rect 6269 17174 8911 17176
rect 6269 17171 6335 17174
rect 8845 17171 8911 17174
rect 10501 17234 10567 17237
rect 15837 17234 15903 17237
rect 10501 17232 15903 17234
rect 10501 17176 10506 17232
rect 10562 17176 15842 17232
rect 15898 17176 15903 17232
rect 10501 17174 15903 17176
rect 10501 17171 10567 17174
rect 15837 17171 15903 17174
rect 7281 17098 7347 17101
rect 12341 17098 12407 17101
rect 7281 17096 12407 17098
rect 7281 17040 7286 17096
rect 7342 17040 12346 17096
rect 12402 17040 12407 17096
rect 7281 17038 12407 17040
rect 7281 17035 7347 17038
rect 12341 17035 12407 17038
rect 12709 17098 12775 17101
rect 14549 17098 14615 17101
rect 12709 17096 14615 17098
rect 12709 17040 12714 17096
rect 12770 17040 14554 17096
rect 14610 17040 14615 17096
rect 12709 17038 14615 17040
rect 12709 17035 12775 17038
rect 14549 17035 14615 17038
rect 14917 17098 14983 17101
rect 15929 17098 15995 17101
rect 16941 17098 17007 17101
rect 14917 17096 17007 17098
rect 14917 17040 14922 17096
rect 14978 17040 15934 17096
rect 15990 17040 16946 17096
rect 17002 17040 17007 17096
rect 14917 17038 17007 17040
rect 14917 17035 14983 17038
rect 15929 17035 15995 17038
rect 16941 17035 17007 17038
rect 35433 17098 35499 17101
rect 38852 17098 39652 17128
rect 35433 17096 39652 17098
rect 35433 17040 35438 17096
rect 35494 17040 39652 17096
rect 35433 17038 39652 17040
rect 35433 17035 35499 17038
rect 38852 17008 39652 17038
rect 3969 16962 4035 16965
rect 6821 16962 6887 16965
rect 11145 16962 11211 16965
rect 3969 16960 6887 16962
rect 3969 16904 3974 16960
rect 4030 16904 6826 16960
rect 6882 16904 6887 16960
rect 3969 16902 6887 16904
rect 3969 16899 4035 16902
rect 6821 16899 6887 16902
rect 9446 16960 11211 16962
rect 9446 16904 11150 16960
rect 11206 16904 11211 16960
rect 9446 16902 11211 16904
rect 5441 16690 5507 16693
rect 7465 16690 7531 16693
rect 9446 16690 9506 16902
rect 11145 16899 11211 16902
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 10777 16826 10843 16829
rect 13629 16826 13695 16829
rect 10777 16824 13695 16826
rect 10777 16768 10782 16824
rect 10838 16768 13634 16824
rect 13690 16768 13695 16824
rect 10777 16766 13695 16768
rect 10777 16763 10843 16766
rect 13629 16763 13695 16766
rect 5441 16688 7531 16690
rect 5441 16632 5446 16688
rect 5502 16632 7470 16688
rect 7526 16632 7531 16688
rect 5441 16630 7531 16632
rect 5441 16627 5507 16630
rect 7465 16627 7531 16630
rect 7790 16630 9506 16690
rect 9673 16690 9739 16693
rect 13077 16690 13143 16693
rect 9673 16688 13143 16690
rect 9673 16632 9678 16688
rect 9734 16632 13082 16688
rect 13138 16632 13143 16688
rect 9673 16630 13143 16632
rect 3877 16554 3943 16557
rect 7790 16554 7850 16630
rect 9673 16627 9739 16630
rect 13077 16627 13143 16630
rect 18781 16690 18847 16693
rect 19793 16690 19859 16693
rect 18781 16688 19859 16690
rect 18781 16632 18786 16688
rect 18842 16632 19798 16688
rect 19854 16632 19859 16688
rect 18781 16630 19859 16632
rect 18781 16627 18847 16630
rect 19793 16627 19859 16630
rect 27245 16690 27311 16693
rect 30741 16690 30807 16693
rect 27245 16688 30807 16690
rect 27245 16632 27250 16688
rect 27306 16632 30746 16688
rect 30802 16632 30807 16688
rect 27245 16630 30807 16632
rect 27245 16627 27311 16630
rect 30741 16627 30807 16630
rect 3877 16552 7850 16554
rect 3877 16496 3882 16552
rect 3938 16496 7850 16552
rect 3877 16494 7850 16496
rect 7925 16554 7991 16557
rect 10501 16554 10567 16557
rect 7925 16552 10567 16554
rect 7925 16496 7930 16552
rect 7986 16496 10506 16552
rect 10562 16496 10567 16552
rect 7925 16494 10567 16496
rect 3877 16491 3943 16494
rect 7925 16491 7991 16494
rect 10501 16491 10567 16494
rect 13486 16492 13492 16556
rect 13556 16554 13562 16556
rect 15653 16554 15719 16557
rect 17217 16554 17283 16557
rect 13556 16552 17283 16554
rect 13556 16496 15658 16552
rect 15714 16496 17222 16552
rect 17278 16496 17283 16552
rect 13556 16494 17283 16496
rect 13556 16492 13562 16494
rect 15653 16491 15719 16494
rect 17217 16491 17283 16494
rect 17493 16554 17559 16557
rect 22461 16554 22527 16557
rect 17493 16552 22527 16554
rect 17493 16496 17498 16552
rect 17554 16496 22466 16552
rect 22522 16496 22527 16552
rect 17493 16494 22527 16496
rect 17493 16491 17559 16494
rect 22461 16491 22527 16494
rect 29545 16554 29611 16557
rect 31937 16554 32003 16557
rect 29545 16552 32003 16554
rect 29545 16496 29550 16552
rect 29606 16496 31942 16552
rect 31998 16496 32003 16552
rect 29545 16494 32003 16496
rect 29545 16491 29611 16494
rect 31937 16491 32003 16494
rect 34053 16554 34119 16557
rect 34053 16552 36370 16554
rect 34053 16496 34058 16552
rect 34114 16496 36370 16552
rect 34053 16494 36370 16496
rect 34053 16491 34119 16494
rect 0 16418 800 16448
rect 1669 16418 1735 16421
rect 0 16416 1735 16418
rect 0 16360 1674 16416
rect 1730 16360 1735 16416
rect 0 16358 1735 16360
rect 0 16328 800 16358
rect 1669 16355 1735 16358
rect 11421 16418 11487 16421
rect 12157 16418 12223 16421
rect 11421 16416 12223 16418
rect 11421 16360 11426 16416
rect 11482 16360 12162 16416
rect 12218 16360 12223 16416
rect 11421 16358 12223 16360
rect 11421 16355 11487 16358
rect 12157 16355 12223 16358
rect 23749 16418 23815 16421
rect 26233 16418 26299 16421
rect 27061 16418 27127 16421
rect 23749 16416 27127 16418
rect 23749 16360 23754 16416
rect 23810 16360 26238 16416
rect 26294 16360 27066 16416
rect 27122 16360 27127 16416
rect 23749 16358 27127 16360
rect 36310 16418 36370 16494
rect 38852 16418 39652 16448
rect 36310 16358 39652 16418
rect 23749 16355 23815 16358
rect 26233 16355 26299 16358
rect 27061 16355 27127 16358
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 38852 16328 39652 16358
rect 34928 16287 35248 16288
rect 17493 16282 17559 16285
rect 4846 16280 17559 16282
rect 4846 16224 17498 16280
rect 17554 16224 17559 16280
rect 4846 16222 17559 16224
rect 0 15738 800 15768
rect 4846 15738 4906 16222
rect 17493 16219 17559 16222
rect 10225 16146 10291 16149
rect 12617 16146 12683 16149
rect 10225 16144 12683 16146
rect 10225 16088 10230 16144
rect 10286 16088 12622 16144
rect 12678 16088 12683 16144
rect 10225 16086 12683 16088
rect 10225 16083 10291 16086
rect 12617 16083 12683 16086
rect 6729 16010 6795 16013
rect 22369 16010 22435 16013
rect 6729 16008 22435 16010
rect 6729 15952 6734 16008
rect 6790 15952 22374 16008
rect 22430 15952 22435 16008
rect 6729 15950 22435 15952
rect 6729 15947 6795 15950
rect 22369 15947 22435 15950
rect 31937 16010 32003 16013
rect 34881 16010 34947 16013
rect 31937 16008 34947 16010
rect 31937 15952 31942 16008
rect 31998 15952 34886 16008
rect 34942 15952 34947 16008
rect 31937 15950 34947 15952
rect 31937 15947 32003 15950
rect 34881 15947 34947 15950
rect 20805 15874 20871 15877
rect 23749 15874 23815 15877
rect 20805 15872 23815 15874
rect 20805 15816 20810 15872
rect 20866 15816 23754 15872
rect 23810 15816 23815 15872
rect 20805 15814 23815 15816
rect 20805 15811 20871 15814
rect 23749 15811 23815 15814
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 0 15678 4906 15738
rect 10961 15738 11027 15741
rect 11605 15738 11671 15741
rect 15193 15738 15259 15741
rect 10961 15736 15259 15738
rect 10961 15680 10966 15736
rect 11022 15680 11610 15736
rect 11666 15680 15198 15736
rect 15254 15680 15259 15736
rect 10961 15678 15259 15680
rect 0 15648 800 15678
rect 10961 15675 11027 15678
rect 11605 15675 11671 15678
rect 15193 15675 15259 15678
rect 6085 15602 6151 15605
rect 7097 15602 7163 15605
rect 12985 15602 13051 15605
rect 6085 15600 13051 15602
rect 6085 15544 6090 15600
rect 6146 15544 7102 15600
rect 7158 15544 12990 15600
rect 13046 15544 13051 15600
rect 6085 15542 13051 15544
rect 6085 15539 6151 15542
rect 7097 15539 7163 15542
rect 12985 15539 13051 15542
rect 25405 15602 25471 15605
rect 27797 15602 27863 15605
rect 32489 15602 32555 15605
rect 25405 15600 32555 15602
rect 25405 15544 25410 15600
rect 25466 15544 27802 15600
rect 27858 15544 32494 15600
rect 32550 15544 32555 15600
rect 25405 15542 32555 15544
rect 25405 15539 25471 15542
rect 27797 15539 27863 15542
rect 32489 15539 32555 15542
rect 3877 15466 3943 15469
rect 11605 15466 11671 15469
rect 12157 15466 12223 15469
rect 12801 15466 12867 15469
rect 3877 15464 12867 15466
rect 3877 15408 3882 15464
rect 3938 15408 11610 15464
rect 11666 15408 12162 15464
rect 12218 15408 12806 15464
rect 12862 15408 12867 15464
rect 3877 15406 12867 15408
rect 3877 15403 3943 15406
rect 11605 15403 11671 15406
rect 12157 15403 12223 15406
rect 12801 15403 12867 15406
rect 7189 15330 7255 15333
rect 12985 15330 13051 15333
rect 13997 15330 14063 15333
rect 7189 15328 14063 15330
rect 7189 15272 7194 15328
rect 7250 15272 12990 15328
rect 13046 15272 14002 15328
rect 14058 15272 14063 15328
rect 7189 15270 14063 15272
rect 7189 15267 7255 15270
rect 12985 15267 13051 15270
rect 13997 15267 14063 15270
rect 14733 15330 14799 15333
rect 19333 15330 19399 15333
rect 14733 15328 19399 15330
rect 14733 15272 14738 15328
rect 14794 15272 19338 15328
rect 19394 15272 19399 15328
rect 14733 15270 19399 15272
rect 14733 15267 14799 15270
rect 19333 15267 19399 15270
rect 22553 15330 22619 15333
rect 30465 15330 30531 15333
rect 22553 15328 30531 15330
rect 22553 15272 22558 15328
rect 22614 15272 30470 15328
rect 30526 15272 30531 15328
rect 22553 15270 30531 15272
rect 22553 15267 22619 15270
rect 30465 15267 30531 15270
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 5441 15194 5507 15197
rect 8017 15194 8083 15197
rect 11053 15194 11119 15197
rect 14365 15194 14431 15197
rect 5441 15192 8218 15194
rect 5441 15136 5446 15192
rect 5502 15136 8022 15192
rect 8078 15136 8218 15192
rect 5441 15134 8218 15136
rect 5441 15131 5507 15134
rect 8017 15131 8083 15134
rect 3509 15058 3575 15061
rect 7833 15058 7899 15061
rect 3509 15056 7899 15058
rect 3509 15000 3514 15056
rect 3570 15000 7838 15056
rect 7894 15000 7899 15056
rect 3509 14998 7899 15000
rect 8158 15058 8218 15134
rect 11053 15192 14431 15194
rect 11053 15136 11058 15192
rect 11114 15136 14370 15192
rect 14426 15136 14431 15192
rect 11053 15134 14431 15136
rect 11053 15131 11119 15134
rect 14365 15131 14431 15134
rect 16573 15194 16639 15197
rect 19885 15194 19951 15197
rect 20713 15194 20779 15197
rect 16573 15192 20779 15194
rect 16573 15136 16578 15192
rect 16634 15136 19890 15192
rect 19946 15136 20718 15192
rect 20774 15136 20779 15192
rect 16573 15134 20779 15136
rect 16573 15131 16639 15134
rect 19885 15131 19951 15134
rect 20713 15131 20779 15134
rect 21817 15194 21883 15197
rect 24485 15194 24551 15197
rect 21817 15192 24551 15194
rect 21817 15136 21822 15192
rect 21878 15136 24490 15192
rect 24546 15136 24551 15192
rect 21817 15134 24551 15136
rect 21817 15131 21883 15134
rect 24485 15131 24551 15134
rect 25129 15194 25195 15197
rect 27705 15194 27771 15197
rect 31385 15194 31451 15197
rect 25129 15192 31451 15194
rect 25129 15136 25134 15192
rect 25190 15136 27710 15192
rect 27766 15136 31390 15192
rect 31446 15136 31451 15192
rect 25129 15134 31451 15136
rect 25129 15131 25195 15134
rect 27705 15131 27771 15134
rect 31385 15131 31451 15134
rect 11237 15058 11303 15061
rect 8158 15056 11303 15058
rect 8158 15000 11242 15056
rect 11298 15000 11303 15056
rect 8158 14998 11303 15000
rect 3509 14995 3575 14998
rect 7833 14995 7899 14998
rect 11237 14995 11303 14998
rect 13813 15058 13879 15061
rect 14733 15058 14799 15061
rect 13813 15056 14799 15058
rect 13813 15000 13818 15056
rect 13874 15000 14738 15056
rect 14794 15000 14799 15056
rect 13813 14998 14799 15000
rect 13813 14995 13879 14998
rect 14733 14995 14799 14998
rect 35566 14996 35572 15060
rect 35636 15058 35642 15060
rect 38852 15058 39652 15088
rect 35636 14998 39652 15058
rect 35636 14996 35642 14998
rect 38852 14968 39652 14998
rect 3877 14922 3943 14925
rect 7465 14922 7531 14925
rect 3877 14920 7531 14922
rect 3877 14864 3882 14920
rect 3938 14864 7470 14920
rect 7526 14864 7531 14920
rect 3877 14862 7531 14864
rect 3877 14859 3943 14862
rect 7465 14859 7531 14862
rect 10041 14922 10107 14925
rect 10961 14922 11027 14925
rect 10041 14920 11027 14922
rect 10041 14864 10046 14920
rect 10102 14864 10966 14920
rect 11022 14864 11027 14920
rect 10041 14862 11027 14864
rect 10041 14859 10107 14862
rect 10961 14859 11027 14862
rect 17769 14922 17835 14925
rect 17902 14922 17908 14924
rect 17769 14920 17908 14922
rect 17769 14864 17774 14920
rect 17830 14864 17908 14920
rect 17769 14862 17908 14864
rect 17769 14859 17835 14862
rect 17902 14860 17908 14862
rect 17972 14922 17978 14924
rect 20161 14922 20227 14925
rect 17972 14920 20227 14922
rect 17972 14864 20166 14920
rect 20222 14864 20227 14920
rect 17972 14862 20227 14864
rect 17972 14860 17978 14862
rect 20161 14859 20227 14862
rect 5257 14786 5323 14789
rect 7373 14786 7439 14789
rect 5257 14784 7439 14786
rect 5257 14728 5262 14784
rect 5318 14728 7378 14784
rect 7434 14728 7439 14784
rect 5257 14726 7439 14728
rect 5257 14723 5323 14726
rect 7373 14723 7439 14726
rect 9397 14786 9463 14789
rect 15009 14786 15075 14789
rect 9397 14784 15075 14786
rect 9397 14728 9402 14784
rect 9458 14728 15014 14784
rect 15070 14728 15075 14784
rect 9397 14726 15075 14728
rect 9397 14723 9463 14726
rect 15009 14723 15075 14726
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 3969 14652 4035 14653
rect 3918 14650 3924 14652
rect 3878 14590 3924 14650
rect 3988 14648 4035 14652
rect 4030 14592 4035 14648
rect 3918 14588 3924 14590
rect 3988 14588 4035 14592
rect 3969 14587 4035 14588
rect 5349 14650 5415 14653
rect 5809 14650 5875 14653
rect 6821 14650 6887 14653
rect 5349 14648 6887 14650
rect 5349 14592 5354 14648
rect 5410 14592 5814 14648
rect 5870 14592 6826 14648
rect 6882 14592 6887 14648
rect 5349 14590 6887 14592
rect 5349 14587 5415 14590
rect 5809 14587 5875 14590
rect 6821 14587 6887 14590
rect 3417 14514 3483 14517
rect 7649 14514 7715 14517
rect 3417 14512 7715 14514
rect 3417 14456 3422 14512
rect 3478 14456 7654 14512
rect 7710 14456 7715 14512
rect 3417 14454 7715 14456
rect 3417 14451 3483 14454
rect 7649 14451 7715 14454
rect 10225 14514 10291 14517
rect 14733 14514 14799 14517
rect 10225 14512 14799 14514
rect 10225 14456 10230 14512
rect 10286 14456 14738 14512
rect 14794 14456 14799 14512
rect 10225 14454 14799 14456
rect 10225 14451 10291 14454
rect 14733 14451 14799 14454
rect 26693 14514 26759 14517
rect 32121 14514 32187 14517
rect 26693 14512 32187 14514
rect 26693 14456 26698 14512
rect 26754 14456 32126 14512
rect 32182 14456 32187 14512
rect 26693 14454 32187 14456
rect 26693 14451 26759 14454
rect 32121 14451 32187 14454
rect 0 14378 800 14408
rect 4889 14378 4955 14381
rect 12525 14378 12591 14381
rect 0 14318 4768 14378
rect 0 14288 800 14318
rect 4708 14242 4768 14318
rect 4889 14376 12591 14378
rect 4889 14320 4894 14376
rect 4950 14320 12530 14376
rect 12586 14320 12591 14376
rect 4889 14318 12591 14320
rect 4889 14315 4955 14318
rect 12525 14315 12591 14318
rect 13629 14378 13695 14381
rect 14549 14378 14615 14381
rect 19517 14378 19583 14381
rect 19885 14378 19951 14381
rect 13629 14376 19951 14378
rect 13629 14320 13634 14376
rect 13690 14320 14554 14376
rect 14610 14320 19522 14376
rect 19578 14320 19890 14376
rect 19946 14320 19951 14376
rect 13629 14318 19951 14320
rect 13629 14315 13695 14318
rect 14549 14315 14615 14318
rect 19517 14315 19583 14318
rect 19885 14315 19951 14318
rect 35709 14378 35775 14381
rect 38852 14378 39652 14408
rect 35709 14376 39652 14378
rect 35709 14320 35714 14376
rect 35770 14320 39652 14376
rect 35709 14318 39652 14320
rect 35709 14315 35775 14318
rect 38852 14288 39652 14318
rect 6729 14242 6795 14245
rect 4708 14240 6795 14242
rect 4708 14184 6734 14240
rect 6790 14184 6795 14240
rect 4708 14182 6795 14184
rect 6729 14179 6795 14182
rect 7557 14242 7623 14245
rect 10777 14242 10843 14245
rect 15561 14242 15627 14245
rect 7557 14240 15627 14242
rect 7557 14184 7562 14240
rect 7618 14184 10782 14240
rect 10838 14184 15566 14240
rect 15622 14184 15627 14240
rect 7557 14182 15627 14184
rect 7557 14179 7623 14182
rect 10777 14179 10843 14182
rect 15561 14179 15627 14182
rect 16614 14180 16620 14244
rect 16684 14242 16690 14244
rect 16941 14242 17007 14245
rect 16684 14240 17007 14242
rect 16684 14184 16946 14240
rect 17002 14184 17007 14240
rect 16684 14182 17007 14184
rect 16684 14180 16690 14182
rect 16941 14179 17007 14182
rect 23841 14242 23907 14245
rect 25313 14242 25379 14245
rect 23841 14240 25379 14242
rect 23841 14184 23846 14240
rect 23902 14184 25318 14240
rect 25374 14184 25379 14240
rect 23841 14182 25379 14184
rect 23841 14179 23907 14182
rect 25313 14179 25379 14182
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 13261 14106 13327 14109
rect 14549 14106 14615 14109
rect 15377 14106 15443 14109
rect 13261 14104 15443 14106
rect 13261 14048 13266 14104
rect 13322 14048 14554 14104
rect 14610 14048 15382 14104
rect 15438 14048 15443 14104
rect 13261 14046 15443 14048
rect 15564 14106 15624 14179
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 17953 14106 18019 14109
rect 18965 14106 19031 14109
rect 15564 14104 19031 14106
rect 15564 14048 17958 14104
rect 18014 14048 18970 14104
rect 19026 14048 19031 14104
rect 15564 14046 19031 14048
rect 13261 14043 13327 14046
rect 14549 14043 14615 14046
rect 15377 14043 15443 14046
rect 17953 14043 18019 14046
rect 18965 14043 19031 14046
rect 16573 13970 16639 13973
rect 19333 13970 19399 13973
rect 16573 13968 19399 13970
rect 16573 13912 16578 13968
rect 16634 13912 19338 13968
rect 19394 13912 19399 13968
rect 16573 13910 19399 13912
rect 16573 13907 16639 13910
rect 19333 13907 19399 13910
rect 1577 13834 1643 13837
rect 1534 13832 1643 13834
rect 1534 13776 1582 13832
rect 1638 13776 1643 13832
rect 1534 13771 1643 13776
rect 13721 13834 13787 13837
rect 17902 13834 17908 13836
rect 13721 13832 17908 13834
rect 13721 13776 13726 13832
rect 13782 13776 17908 13832
rect 13721 13774 17908 13776
rect 13721 13771 13787 13774
rect 17902 13772 17908 13774
rect 17972 13772 17978 13836
rect 0 13698 800 13728
rect 1534 13698 1594 13771
rect 0 13638 1594 13698
rect 8477 13698 8543 13701
rect 12709 13698 12775 13701
rect 8477 13696 12775 13698
rect 8477 13640 8482 13696
rect 8538 13640 12714 13696
rect 12770 13640 12775 13696
rect 8477 13638 12775 13640
rect 0 13608 800 13638
rect 8477 13635 8543 13638
rect 12709 13635 12775 13638
rect 14365 13698 14431 13701
rect 16665 13698 16731 13701
rect 14365 13696 16731 13698
rect 14365 13640 14370 13696
rect 14426 13640 16670 13696
rect 16726 13640 16731 13696
rect 14365 13638 16731 13640
rect 14365 13635 14431 13638
rect 16665 13635 16731 13638
rect 35525 13698 35591 13701
rect 38852 13698 39652 13728
rect 35525 13696 39652 13698
rect 35525 13640 35530 13696
rect 35586 13640 39652 13696
rect 35525 13638 39652 13640
rect 35525 13635 35591 13638
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 38852 13608 39652 13638
rect 19568 13567 19888 13568
rect 5717 13562 5783 13565
rect 10961 13562 11027 13565
rect 5717 13560 11027 13562
rect 5717 13504 5722 13560
rect 5778 13504 10966 13560
rect 11022 13504 11027 13560
rect 5717 13502 11027 13504
rect 5717 13499 5783 13502
rect 10961 13499 11027 13502
rect 16062 13500 16068 13564
rect 16132 13562 16138 13564
rect 16205 13562 16271 13565
rect 16132 13560 16271 13562
rect 16132 13504 16210 13560
rect 16266 13504 16271 13560
rect 16132 13502 16271 13504
rect 16132 13500 16138 13502
rect 16205 13499 16271 13502
rect 5257 13426 5323 13429
rect 8477 13426 8543 13429
rect 5257 13424 8543 13426
rect 5257 13368 5262 13424
rect 5318 13368 8482 13424
rect 8538 13368 8543 13424
rect 5257 13366 8543 13368
rect 5257 13363 5323 13366
rect 8477 13363 8543 13366
rect 12249 13426 12315 13429
rect 16849 13426 16915 13429
rect 12249 13424 16915 13426
rect 12249 13368 12254 13424
rect 12310 13368 16854 13424
rect 16910 13368 16915 13424
rect 12249 13366 16915 13368
rect 12249 13363 12315 13366
rect 16849 13363 16915 13366
rect 4981 13290 5047 13293
rect 11237 13290 11303 13293
rect 4981 13288 11303 13290
rect 4981 13232 4986 13288
rect 5042 13232 11242 13288
rect 11298 13232 11303 13288
rect 4981 13230 11303 13232
rect 4981 13227 5047 13230
rect 11237 13227 11303 13230
rect 5717 13154 5783 13157
rect 9857 13154 9923 13157
rect 5717 13152 9923 13154
rect 5717 13096 5722 13152
rect 5778 13096 9862 13152
rect 9918 13096 9923 13152
rect 5717 13094 9923 13096
rect 5717 13091 5783 13094
rect 9857 13091 9923 13094
rect 10501 13154 10567 13157
rect 15193 13154 15259 13157
rect 10501 13152 15259 13154
rect 10501 13096 10506 13152
rect 10562 13096 15198 13152
rect 15254 13096 15259 13152
rect 10501 13094 15259 13096
rect 10501 13091 10567 13094
rect 15193 13091 15259 13094
rect 30373 13154 30439 13157
rect 31845 13154 31911 13157
rect 30373 13152 31911 13154
rect 30373 13096 30378 13152
rect 30434 13096 31850 13152
rect 31906 13096 31911 13152
rect 30373 13094 31911 13096
rect 30373 13091 30439 13094
rect 31845 13091 31911 13094
rect 4208 13088 4528 13089
rect 0 13018 800 13048
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 13023 35248 13024
rect 1577 13018 1643 13021
rect 0 13016 1643 13018
rect 0 12960 1582 13016
rect 1638 12960 1643 13016
rect 0 12958 1643 12960
rect 0 12928 800 12958
rect 1577 12955 1643 12958
rect 4889 13018 4955 13021
rect 9305 13018 9371 13021
rect 4889 13016 9371 13018
rect 4889 12960 4894 13016
rect 4950 12960 9310 13016
rect 9366 12960 9371 13016
rect 4889 12958 9371 12960
rect 4889 12955 4955 12958
rect 9305 12955 9371 12958
rect 9581 13018 9647 13021
rect 12617 13018 12683 13021
rect 9581 13016 12683 13018
rect 9581 12960 9586 13016
rect 9642 12960 12622 13016
rect 12678 12960 12683 13016
rect 9581 12958 12683 12960
rect 9581 12955 9647 12958
rect 12617 12955 12683 12958
rect 16941 13018 17007 13021
rect 20069 13018 20135 13021
rect 16941 13016 20135 13018
rect 16941 12960 16946 13016
rect 17002 12960 20074 13016
rect 20130 12960 20135 13016
rect 16941 12958 20135 12960
rect 16941 12955 17007 12958
rect 20069 12955 20135 12958
rect 22553 13018 22619 13021
rect 30925 13018 30991 13021
rect 22553 13016 30991 13018
rect 22553 12960 22558 13016
rect 22614 12960 30930 13016
rect 30986 12960 30991 13016
rect 22553 12958 30991 12960
rect 22553 12955 22619 12958
rect 30925 12955 30991 12958
rect 6913 12882 6979 12885
rect 10317 12882 10383 12885
rect 12709 12882 12775 12885
rect 6913 12880 12775 12882
rect 6913 12824 6918 12880
rect 6974 12824 10322 12880
rect 10378 12824 12714 12880
rect 12770 12824 12775 12880
rect 6913 12822 12775 12824
rect 6913 12819 6979 12822
rect 10317 12819 10383 12822
rect 12709 12819 12775 12822
rect 15101 12882 15167 12885
rect 16021 12882 16087 12885
rect 15101 12880 16087 12882
rect 15101 12824 15106 12880
rect 15162 12824 16026 12880
rect 16082 12824 16087 12880
rect 15101 12822 16087 12824
rect 15101 12819 15167 12822
rect 16021 12819 16087 12822
rect 16573 12884 16639 12885
rect 16573 12880 16620 12884
rect 16684 12882 16690 12884
rect 17677 12882 17743 12885
rect 22461 12882 22527 12885
rect 16573 12824 16578 12880
rect 16573 12820 16620 12824
rect 16684 12822 16730 12882
rect 17677 12880 22527 12882
rect 17677 12824 17682 12880
rect 17738 12824 22466 12880
rect 22522 12824 22527 12880
rect 17677 12822 22527 12824
rect 16684 12820 16690 12822
rect 16573 12819 16639 12820
rect 17677 12819 17743 12822
rect 22461 12819 22527 12822
rect 12065 12746 12131 12749
rect 18597 12746 18663 12749
rect 12065 12744 18663 12746
rect 12065 12688 12070 12744
rect 12126 12688 18602 12744
rect 18658 12688 18663 12744
rect 12065 12686 18663 12688
rect 12065 12683 12131 12686
rect 18597 12683 18663 12686
rect 19333 12744 19399 12749
rect 19333 12688 19338 12744
rect 19394 12688 19399 12744
rect 19333 12683 19399 12688
rect 20713 12746 20779 12749
rect 37273 12746 37339 12749
rect 20713 12744 37339 12746
rect 20713 12688 20718 12744
rect 20774 12688 37278 12744
rect 37334 12688 37339 12744
rect 20713 12686 37339 12688
rect 20713 12683 20779 12686
rect 37273 12683 37339 12686
rect 12617 12610 12683 12613
rect 12893 12610 12959 12613
rect 12617 12608 12959 12610
rect 12617 12552 12622 12608
rect 12678 12552 12898 12608
rect 12954 12552 12959 12608
rect 12617 12550 12959 12552
rect 12617 12547 12683 12550
rect 12893 12547 12959 12550
rect 13077 12610 13143 12613
rect 13721 12610 13787 12613
rect 13077 12608 13787 12610
rect 13077 12552 13082 12608
rect 13138 12552 13726 12608
rect 13782 12552 13787 12608
rect 13077 12550 13787 12552
rect 13077 12547 13143 12550
rect 13721 12547 13787 12550
rect 13997 12610 14063 12613
rect 14549 12610 14615 12613
rect 17493 12610 17559 12613
rect 18505 12610 18571 12613
rect 13997 12608 18571 12610
rect 13997 12552 14002 12608
rect 14058 12552 14554 12608
rect 14610 12552 17498 12608
rect 17554 12552 18510 12608
rect 18566 12552 18571 12608
rect 13997 12550 18571 12552
rect 13997 12547 14063 12550
rect 14549 12547 14615 12550
rect 17493 12547 17559 12550
rect 18505 12547 18571 12550
rect 13445 12476 13511 12477
rect 13445 12474 13492 12476
rect 13400 12472 13492 12474
rect 13400 12416 13450 12472
rect 13400 12414 13492 12416
rect 13445 12412 13492 12414
rect 13556 12412 13562 12476
rect 13445 12411 13511 12412
rect 19336 12341 19396 12683
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 3141 12338 3207 12341
rect 5993 12338 6059 12341
rect 3141 12336 6059 12338
rect 3141 12280 3146 12336
rect 3202 12280 5998 12336
rect 6054 12280 6059 12336
rect 3141 12278 6059 12280
rect 3141 12275 3207 12278
rect 5993 12275 6059 12278
rect 8201 12338 8267 12341
rect 14089 12338 14155 12341
rect 17309 12340 17375 12341
rect 18505 12340 18571 12341
rect 17309 12338 17356 12340
rect 8201 12336 14155 12338
rect 8201 12280 8206 12336
rect 8262 12280 14094 12336
rect 14150 12280 14155 12336
rect 8201 12278 14155 12280
rect 17264 12336 17356 12338
rect 17264 12280 17314 12336
rect 17264 12278 17356 12280
rect 8201 12275 8267 12278
rect 14089 12275 14155 12278
rect 17309 12276 17356 12278
rect 17420 12276 17426 12340
rect 18454 12338 18460 12340
rect 18414 12278 18460 12338
rect 18524 12336 18571 12340
rect 18566 12280 18571 12336
rect 18454 12276 18460 12278
rect 18524 12276 18571 12280
rect 17309 12275 17375 12276
rect 18505 12275 18571 12276
rect 19333 12336 19399 12341
rect 19333 12280 19338 12336
rect 19394 12280 19399 12336
rect 19333 12275 19399 12280
rect 25589 12338 25655 12341
rect 29637 12338 29703 12341
rect 38852 12338 39652 12368
rect 25589 12336 29703 12338
rect 25589 12280 25594 12336
rect 25650 12280 29642 12336
rect 29698 12280 29703 12336
rect 25589 12278 29703 12280
rect 25589 12275 25655 12278
rect 29637 12275 29703 12278
rect 38702 12278 39652 12338
rect 6821 12202 6887 12205
rect 8661 12202 8727 12205
rect 6821 12200 8727 12202
rect 6821 12144 6826 12200
rect 6882 12144 8666 12200
rect 8722 12144 8727 12200
rect 6821 12142 8727 12144
rect 6821 12139 6887 12142
rect 8661 12139 8727 12142
rect 27981 12202 28047 12205
rect 38702 12202 38762 12278
rect 38852 12248 39652 12278
rect 27981 12200 38762 12202
rect 27981 12144 27986 12200
rect 28042 12144 38762 12200
rect 27981 12142 38762 12144
rect 27981 12139 28047 12142
rect 4613 12066 4679 12069
rect 8385 12066 8451 12069
rect 4613 12064 8451 12066
rect 4613 12008 4618 12064
rect 4674 12008 8390 12064
rect 8446 12008 8451 12064
rect 4613 12006 8451 12008
rect 4613 12003 4679 12006
rect 8385 12003 8451 12006
rect 26785 12066 26851 12069
rect 30925 12066 30991 12069
rect 26785 12064 30991 12066
rect 26785 12008 26790 12064
rect 26846 12008 30930 12064
rect 30986 12008 30991 12064
rect 26785 12006 30991 12008
rect 26785 12003 26851 12006
rect 30925 12003 30991 12006
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 7465 11930 7531 11933
rect 17677 11930 17743 11933
rect 7465 11928 17743 11930
rect 7465 11872 7470 11928
rect 7526 11872 17682 11928
rect 17738 11872 17743 11928
rect 7465 11870 17743 11872
rect 7465 11867 7531 11870
rect 17677 11867 17743 11870
rect 10501 11794 10567 11797
rect 14273 11794 14339 11797
rect 10501 11792 14339 11794
rect 10501 11736 10506 11792
rect 10562 11736 14278 11792
rect 14334 11736 14339 11792
rect 10501 11734 14339 11736
rect 10501 11731 10567 11734
rect 14273 11731 14339 11734
rect 0 11658 800 11688
rect 3785 11658 3851 11661
rect 0 11656 3851 11658
rect 0 11600 3790 11656
rect 3846 11600 3851 11656
rect 0 11598 3851 11600
rect 0 11568 800 11598
rect 3785 11595 3851 11598
rect 15377 11658 15443 11661
rect 18045 11658 18111 11661
rect 15377 11656 18111 11658
rect 15377 11600 15382 11656
rect 15438 11600 18050 11656
rect 18106 11600 18111 11656
rect 15377 11598 18111 11600
rect 15377 11595 15443 11598
rect 18045 11595 18111 11598
rect 28717 11658 28783 11661
rect 38852 11658 39652 11688
rect 28717 11656 39652 11658
rect 28717 11600 28722 11656
rect 28778 11600 39652 11656
rect 28717 11598 39652 11600
rect 28717 11595 28783 11598
rect 38852 11568 39652 11598
rect 6177 11522 6243 11525
rect 16665 11522 16731 11525
rect 6177 11520 16731 11522
rect 6177 11464 6182 11520
rect 6238 11464 16670 11520
rect 16726 11464 16731 11520
rect 6177 11462 16731 11464
rect 6177 11459 6243 11462
rect 16665 11459 16731 11462
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 21817 11386 21883 11389
rect 28533 11386 28599 11389
rect 29453 11386 29519 11389
rect 21817 11384 29519 11386
rect 21817 11328 21822 11384
rect 21878 11328 28538 11384
rect 28594 11328 29458 11384
rect 29514 11328 29519 11384
rect 21817 11326 29519 11328
rect 21817 11323 21883 11326
rect 28533 11323 28599 11326
rect 29453 11323 29519 11326
rect 8201 11250 8267 11253
rect 11053 11250 11119 11253
rect 8201 11248 11119 11250
rect 8201 11192 8206 11248
rect 8262 11192 11058 11248
rect 11114 11192 11119 11248
rect 8201 11190 11119 11192
rect 8201 11187 8267 11190
rect 11053 11187 11119 11190
rect 13629 11250 13695 11253
rect 19149 11250 19215 11253
rect 13629 11248 19215 11250
rect 13629 11192 13634 11248
rect 13690 11192 19154 11248
rect 19210 11192 19215 11248
rect 13629 11190 19215 11192
rect 13629 11187 13695 11190
rect 19149 11187 19215 11190
rect 1485 11114 1551 11117
rect 1350 11112 1551 11114
rect 1350 11056 1490 11112
rect 1546 11056 1551 11112
rect 1350 11054 1551 11056
rect 0 10978 800 11008
rect 1350 10978 1410 11054
rect 1485 11051 1551 11054
rect 2865 11114 2931 11117
rect 7925 11114 7991 11117
rect 2865 11112 7991 11114
rect 2865 11056 2870 11112
rect 2926 11056 7930 11112
rect 7986 11056 7991 11112
rect 2865 11054 7991 11056
rect 2865 11051 2931 11054
rect 7925 11051 7991 11054
rect 10777 11114 10843 11117
rect 12433 11114 12499 11117
rect 12985 11114 13051 11117
rect 10777 11112 13051 11114
rect 10777 11056 10782 11112
rect 10838 11056 12438 11112
rect 12494 11056 12990 11112
rect 13046 11056 13051 11112
rect 10777 11054 13051 11056
rect 10777 11051 10843 11054
rect 12433 11051 12499 11054
rect 12985 11051 13051 11054
rect 0 10918 1410 10978
rect 8661 10978 8727 10981
rect 16481 10978 16547 10981
rect 23105 10978 23171 10981
rect 8661 10976 23171 10978
rect 8661 10920 8666 10976
rect 8722 10920 16486 10976
rect 16542 10920 23110 10976
rect 23166 10920 23171 10976
rect 8661 10918 23171 10920
rect 0 10888 800 10918
rect 8661 10915 8727 10918
rect 16481 10915 16547 10918
rect 23105 10915 23171 10918
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 6637 10842 6703 10845
rect 8477 10842 8543 10845
rect 6637 10840 8543 10842
rect 6637 10784 6642 10840
rect 6698 10784 8482 10840
rect 8538 10784 8543 10840
rect 6637 10782 8543 10784
rect 6637 10779 6703 10782
rect 8477 10779 8543 10782
rect 9489 10842 9555 10845
rect 12709 10842 12775 10845
rect 9489 10840 12775 10842
rect 9489 10784 9494 10840
rect 9550 10784 12714 10840
rect 12770 10784 12775 10840
rect 9489 10782 12775 10784
rect 9489 10779 9555 10782
rect 12709 10779 12775 10782
rect 17534 10780 17540 10844
rect 17604 10842 17610 10844
rect 29545 10842 29611 10845
rect 17604 10840 29611 10842
rect 17604 10784 29550 10840
rect 29606 10784 29611 10840
rect 17604 10782 29611 10784
rect 17604 10780 17610 10782
rect 29545 10779 29611 10782
rect 9397 10706 9463 10709
rect 16665 10706 16731 10709
rect 9397 10704 16731 10706
rect 9397 10648 9402 10704
rect 9458 10648 16670 10704
rect 16726 10648 16731 10704
rect 9397 10646 16731 10648
rect 9397 10643 9463 10646
rect 16665 10643 16731 10646
rect 17585 10706 17651 10709
rect 32029 10706 32095 10709
rect 17585 10704 32095 10706
rect 17585 10648 17590 10704
rect 17646 10648 32034 10704
rect 32090 10648 32095 10704
rect 17585 10646 32095 10648
rect 17585 10643 17651 10646
rect 32029 10643 32095 10646
rect 11329 10434 11395 10437
rect 19149 10434 19215 10437
rect 11329 10432 19215 10434
rect 11329 10376 11334 10432
rect 11390 10376 19154 10432
rect 19210 10376 19215 10432
rect 11329 10374 19215 10376
rect 11329 10371 11395 10374
rect 19149 10371 19215 10374
rect 19568 10368 19888 10369
rect 0 10298 800 10328
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 1577 10298 1643 10301
rect 0 10296 1643 10298
rect 0 10240 1582 10296
rect 1638 10240 1643 10296
rect 0 10238 1643 10240
rect 0 10208 800 10238
rect 1577 10235 1643 10238
rect 9305 10298 9371 10301
rect 15193 10298 15259 10301
rect 17401 10298 17467 10301
rect 17861 10300 17927 10301
rect 17861 10298 17908 10300
rect 9305 10296 17467 10298
rect 9305 10240 9310 10296
rect 9366 10240 15198 10296
rect 15254 10240 17406 10296
rect 17462 10240 17467 10296
rect 9305 10238 17467 10240
rect 17816 10296 17908 10298
rect 17816 10240 17866 10296
rect 17816 10238 17908 10240
rect 9305 10235 9371 10238
rect 15193 10235 15259 10238
rect 17401 10235 17467 10238
rect 17861 10236 17908 10238
rect 17972 10236 17978 10300
rect 33409 10298 33475 10301
rect 38852 10298 39652 10328
rect 33409 10296 39652 10298
rect 33409 10240 33414 10296
rect 33470 10240 39652 10296
rect 33409 10238 39652 10240
rect 17861 10235 17927 10236
rect 33409 10235 33475 10238
rect 38852 10208 39652 10238
rect 5533 10162 5599 10165
rect 15837 10162 15903 10165
rect 23565 10162 23631 10165
rect 5533 10160 23631 10162
rect 5533 10104 5538 10160
rect 5594 10104 15842 10160
rect 15898 10104 23570 10160
rect 23626 10104 23631 10160
rect 5533 10102 23631 10104
rect 5533 10099 5599 10102
rect 15837 10099 15903 10102
rect 23565 10099 23631 10102
rect 8753 10026 8819 10029
rect 10869 10026 10935 10029
rect 8753 10024 10935 10026
rect 8753 9968 8758 10024
rect 8814 9968 10874 10024
rect 10930 9968 10935 10024
rect 8753 9966 10935 9968
rect 8753 9963 8819 9966
rect 10869 9963 10935 9966
rect 18137 9890 18203 9893
rect 21173 9890 21239 9893
rect 18137 9888 21239 9890
rect 18137 9832 18142 9888
rect 18198 9832 21178 9888
rect 21234 9832 21239 9888
rect 18137 9830 21239 9832
rect 18137 9827 18203 9830
rect 21173 9827 21239 9830
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 25773 9754 25839 9757
rect 20670 9752 25839 9754
rect 20670 9696 25778 9752
rect 25834 9696 25839 9752
rect 20670 9694 25839 9696
rect 2405 9618 2471 9621
rect 20670 9618 20730 9694
rect 25773 9691 25839 9694
rect 2405 9616 20730 9618
rect 2405 9560 2410 9616
rect 2466 9560 20730 9616
rect 2405 9558 20730 9560
rect 20805 9618 20871 9621
rect 25773 9618 25839 9621
rect 20805 9616 25839 9618
rect 20805 9560 20810 9616
rect 20866 9560 25778 9616
rect 25834 9560 25839 9616
rect 20805 9558 25839 9560
rect 2405 9555 2471 9558
rect 20805 9555 20871 9558
rect 25773 9555 25839 9558
rect 25957 9618 26023 9621
rect 27337 9618 27403 9621
rect 35065 9618 35131 9621
rect 25957 9616 35131 9618
rect 25957 9560 25962 9616
rect 26018 9560 27342 9616
rect 27398 9560 35070 9616
rect 35126 9560 35131 9616
rect 25957 9558 35131 9560
rect 25957 9555 26023 9558
rect 27337 9555 27403 9558
rect 35065 9555 35131 9558
rect 35249 9618 35315 9621
rect 38852 9618 39652 9648
rect 35249 9616 39652 9618
rect 35249 9560 35254 9616
rect 35310 9560 39652 9616
rect 35249 9558 39652 9560
rect 35249 9555 35315 9558
rect 38852 9528 39652 9558
rect 3785 9482 3851 9485
rect 7281 9482 7347 9485
rect 3785 9480 7347 9482
rect 3785 9424 3790 9480
rect 3846 9424 7286 9480
rect 7342 9424 7347 9480
rect 3785 9422 7347 9424
rect 3785 9419 3851 9422
rect 7281 9419 7347 9422
rect 9489 9482 9555 9485
rect 11421 9482 11487 9485
rect 9489 9480 11487 9482
rect 9489 9424 9494 9480
rect 9550 9424 11426 9480
rect 11482 9424 11487 9480
rect 9489 9422 11487 9424
rect 9489 9419 9555 9422
rect 11421 9419 11487 9422
rect 19241 9482 19307 9485
rect 34605 9482 34671 9485
rect 19241 9480 34671 9482
rect 19241 9424 19246 9480
rect 19302 9424 34610 9480
rect 34666 9424 34671 9480
rect 19241 9422 34671 9424
rect 19241 9419 19307 9422
rect 34605 9419 34671 9422
rect 6177 9346 6243 9349
rect 10133 9346 10199 9349
rect 6177 9344 10199 9346
rect 6177 9288 6182 9344
rect 6238 9288 10138 9344
rect 10194 9288 10199 9344
rect 6177 9286 10199 9288
rect 6177 9283 6243 9286
rect 10133 9283 10199 9286
rect 24669 9346 24735 9349
rect 24669 9344 35266 9346
rect 24669 9288 24674 9344
rect 24730 9288 35266 9344
rect 24669 9286 35266 9288
rect 24669 9283 24735 9286
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 23289 9210 23355 9213
rect 26141 9210 26207 9213
rect 23289 9208 26207 9210
rect 23289 9152 23294 9208
rect 23350 9152 26146 9208
rect 26202 9152 26207 9208
rect 23289 9150 26207 9152
rect 23289 9147 23355 9150
rect 26141 9147 26207 9150
rect 15009 9074 15075 9077
rect 18597 9074 18663 9077
rect 15009 9072 18663 9074
rect 15009 9016 15014 9072
rect 15070 9016 18602 9072
rect 18658 9016 18663 9072
rect 15009 9014 18663 9016
rect 15009 9011 15075 9014
rect 18597 9011 18663 9014
rect 18965 9074 19031 9077
rect 33961 9074 34027 9077
rect 18965 9072 34027 9074
rect 18965 9016 18970 9072
rect 19026 9016 33966 9072
rect 34022 9016 34027 9072
rect 18965 9014 34027 9016
rect 18965 9011 19031 9014
rect 33961 9011 34027 9014
rect 0 8938 800 8968
rect 2405 8938 2471 8941
rect 0 8936 2471 8938
rect 0 8880 2410 8936
rect 2466 8880 2471 8936
rect 0 8878 2471 8880
rect 0 8848 800 8878
rect 2405 8875 2471 8878
rect 6269 8938 6335 8941
rect 12893 8938 12959 8941
rect 6269 8936 12959 8938
rect 6269 8880 6274 8936
rect 6330 8880 12898 8936
rect 12954 8880 12959 8936
rect 6269 8878 12959 8880
rect 6269 8875 6335 8878
rect 12893 8875 12959 8878
rect 13261 8938 13327 8941
rect 20805 8938 20871 8941
rect 13261 8936 20871 8938
rect 13261 8880 13266 8936
rect 13322 8880 20810 8936
rect 20866 8880 20871 8936
rect 13261 8878 20871 8880
rect 35206 8938 35266 9286
rect 38852 8938 39652 8968
rect 35206 8878 39652 8938
rect 13261 8875 13327 8878
rect 20805 8875 20871 8878
rect 38852 8848 39652 8878
rect 12157 8802 12223 8805
rect 14365 8802 14431 8805
rect 12157 8800 14431 8802
rect 12157 8744 12162 8800
rect 12218 8744 14370 8800
rect 14426 8744 14431 8800
rect 12157 8742 14431 8744
rect 12157 8739 12223 8742
rect 14365 8739 14431 8742
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 9581 8666 9647 8669
rect 16021 8666 16087 8669
rect 9581 8664 16087 8666
rect 9581 8608 9586 8664
rect 9642 8608 16026 8664
rect 16082 8608 16087 8664
rect 9581 8606 16087 8608
rect 9581 8603 9647 8606
rect 16021 8603 16087 8606
rect 8201 8530 8267 8533
rect 9029 8530 9095 8533
rect 10133 8530 10199 8533
rect 16113 8530 16179 8533
rect 16849 8530 16915 8533
rect 8201 8528 16915 8530
rect 8201 8472 8206 8528
rect 8262 8472 9034 8528
rect 9090 8472 10138 8528
rect 10194 8472 16118 8528
rect 16174 8472 16854 8528
rect 16910 8472 16915 8528
rect 8201 8470 16915 8472
rect 8201 8467 8267 8470
rect 9029 8467 9095 8470
rect 10133 8467 10199 8470
rect 16113 8467 16179 8470
rect 16849 8467 16915 8470
rect 3601 8394 3667 8397
rect 10041 8394 10107 8397
rect 3601 8392 10107 8394
rect 3601 8336 3606 8392
rect 3662 8336 10046 8392
rect 10102 8336 10107 8392
rect 3601 8334 10107 8336
rect 3601 8331 3667 8334
rect 10041 8331 10107 8334
rect 14641 8394 14707 8397
rect 16665 8394 16731 8397
rect 14641 8392 16731 8394
rect 14641 8336 14646 8392
rect 14702 8336 16670 8392
rect 16726 8336 16731 8392
rect 14641 8334 16731 8336
rect 14641 8331 14707 8334
rect 16665 8331 16731 8334
rect 0 8258 800 8288
rect 2681 8258 2747 8261
rect 0 8256 2747 8258
rect 0 8200 2686 8256
rect 2742 8200 2747 8256
rect 0 8198 2747 8200
rect 0 8168 800 8198
rect 2681 8195 2747 8198
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 3509 7986 3575 7989
rect 23657 7986 23723 7989
rect 3509 7984 23723 7986
rect 3509 7928 3514 7984
rect 3570 7928 23662 7984
rect 23718 7928 23723 7984
rect 3509 7926 23723 7928
rect 3509 7923 3575 7926
rect 23657 7923 23723 7926
rect 18689 7850 18755 7853
rect 22185 7850 22251 7853
rect 18689 7848 22251 7850
rect 18689 7792 18694 7848
rect 18750 7792 22190 7848
rect 22246 7792 22251 7848
rect 18689 7790 22251 7792
rect 18689 7787 18755 7790
rect 22185 7787 22251 7790
rect 32213 7850 32279 7853
rect 32213 7848 35450 7850
rect 32213 7792 32218 7848
rect 32274 7792 35450 7848
rect 32213 7790 35450 7792
rect 32213 7787 32279 7790
rect 5533 7714 5599 7717
rect 19701 7714 19767 7717
rect 5533 7712 19767 7714
rect 5533 7656 5538 7712
rect 5594 7656 19706 7712
rect 19762 7656 19767 7712
rect 5533 7654 19767 7656
rect 5533 7651 5599 7654
rect 19701 7651 19767 7654
rect 22461 7714 22527 7717
rect 33501 7714 33567 7717
rect 22461 7712 33567 7714
rect 22461 7656 22466 7712
rect 22522 7656 33506 7712
rect 33562 7656 33567 7712
rect 22461 7654 33567 7656
rect 22461 7651 22527 7654
rect 33501 7651 33567 7654
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 4797 7578 4863 7581
rect 17953 7578 18019 7581
rect 4797 7576 18019 7578
rect 4797 7520 4802 7576
rect 4858 7520 17958 7576
rect 18014 7520 18019 7576
rect 4797 7518 18019 7520
rect 4797 7515 4863 7518
rect 17953 7515 18019 7518
rect 18781 7578 18847 7581
rect 34697 7578 34763 7581
rect 18781 7576 34763 7578
rect 18781 7520 18786 7576
rect 18842 7520 34702 7576
rect 34758 7520 34763 7576
rect 18781 7518 34763 7520
rect 35390 7578 35450 7790
rect 38852 7578 39652 7608
rect 35390 7518 39652 7578
rect 18781 7515 18847 7518
rect 34697 7515 34763 7518
rect 38852 7488 39652 7518
rect 18505 7442 18571 7445
rect 20345 7442 20411 7445
rect 18505 7440 20411 7442
rect 18505 7384 18510 7440
rect 18566 7384 20350 7440
rect 20406 7384 20411 7440
rect 18505 7382 20411 7384
rect 18505 7379 18571 7382
rect 20345 7379 20411 7382
rect 2773 7306 2839 7309
rect 22277 7306 22343 7309
rect 2773 7304 22343 7306
rect 2773 7248 2778 7304
rect 2834 7248 22282 7304
rect 22338 7248 22343 7304
rect 2773 7246 22343 7248
rect 2773 7243 2839 7246
rect 22277 7243 22343 7246
rect 3785 7170 3851 7173
rect 10225 7170 10291 7173
rect 3785 7168 10291 7170
rect 3785 7112 3790 7168
rect 3846 7112 10230 7168
rect 10286 7112 10291 7168
rect 3785 7110 10291 7112
rect 3785 7107 3851 7110
rect 10225 7107 10291 7110
rect 11237 7170 11303 7173
rect 13905 7170 13971 7173
rect 11237 7168 13971 7170
rect 11237 7112 11242 7168
rect 11298 7112 13910 7168
rect 13966 7112 13971 7168
rect 11237 7110 13971 7112
rect 11237 7107 11303 7110
rect 13905 7107 13971 7110
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 1485 7034 1551 7037
rect 798 7032 1551 7034
rect 798 6976 1490 7032
rect 1546 6976 1551 7032
rect 798 6974 1551 6976
rect 798 6928 858 6974
rect 1485 6971 1551 6974
rect 0 6838 858 6928
rect 10869 6898 10935 6901
rect 16849 6898 16915 6901
rect 19425 6898 19491 6901
rect 10869 6896 13738 6898
rect 10869 6840 10874 6896
rect 10930 6840 13738 6896
rect 10869 6838 13738 6840
rect 0 6808 800 6838
rect 10869 6835 10935 6838
rect 1853 6762 1919 6765
rect 13537 6762 13603 6765
rect 1853 6760 13603 6762
rect 1853 6704 1858 6760
rect 1914 6704 13542 6760
rect 13598 6704 13603 6760
rect 1853 6702 13603 6704
rect 13678 6762 13738 6838
rect 16849 6896 19491 6898
rect 16849 6840 16854 6896
rect 16910 6840 19430 6896
rect 19486 6840 19491 6896
rect 16849 6838 19491 6840
rect 16849 6835 16915 6838
rect 19425 6835 19491 6838
rect 28717 6898 28783 6901
rect 30833 6898 30899 6901
rect 28717 6896 30899 6898
rect 28717 6840 28722 6896
rect 28778 6840 30838 6896
rect 30894 6840 30899 6896
rect 28717 6838 30899 6840
rect 28717 6835 28783 6838
rect 30833 6835 30899 6838
rect 34513 6898 34579 6901
rect 38852 6898 39652 6928
rect 34513 6896 39652 6898
rect 34513 6840 34518 6896
rect 34574 6840 39652 6896
rect 34513 6838 39652 6840
rect 34513 6835 34579 6838
rect 38852 6808 39652 6838
rect 13813 6762 13879 6765
rect 13678 6760 13879 6762
rect 13678 6704 13818 6760
rect 13874 6704 13879 6760
rect 13678 6702 13879 6704
rect 1853 6699 1919 6702
rect 13537 6699 13603 6702
rect 13813 6699 13879 6702
rect 10910 6564 10916 6628
rect 10980 6626 10986 6628
rect 11513 6626 11579 6629
rect 10980 6624 11579 6626
rect 10980 6568 11518 6624
rect 11574 6568 11579 6624
rect 10980 6566 11579 6568
rect 10980 6564 10986 6566
rect 11513 6563 11579 6566
rect 12893 6626 12959 6629
rect 22553 6626 22619 6629
rect 12893 6624 22619 6626
rect 12893 6568 12898 6624
rect 12954 6568 22558 6624
rect 22614 6568 22619 6624
rect 12893 6566 22619 6568
rect 12893 6563 12959 6566
rect 22553 6563 22619 6566
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 13997 6490 14063 6493
rect 18505 6490 18571 6493
rect 13997 6488 18571 6490
rect 13997 6432 14002 6488
rect 14058 6432 18510 6488
rect 18566 6432 18571 6488
rect 13997 6430 18571 6432
rect 13997 6427 14063 6430
rect 18505 6427 18571 6430
rect 14549 6354 14615 6357
rect 19057 6354 19123 6357
rect 14549 6352 19123 6354
rect 14549 6296 14554 6352
rect 14610 6296 19062 6352
rect 19118 6296 19123 6352
rect 14549 6294 19123 6296
rect 14549 6291 14615 6294
rect 19057 6291 19123 6294
rect 20897 6354 20963 6357
rect 35249 6354 35315 6357
rect 20897 6352 35315 6354
rect 20897 6296 20902 6352
rect 20958 6296 35254 6352
rect 35310 6296 35315 6352
rect 20897 6294 35315 6296
rect 20897 6291 20963 6294
rect 35249 6291 35315 6294
rect 0 6218 800 6248
rect 1761 6218 1827 6221
rect 0 6216 1827 6218
rect 0 6160 1766 6216
rect 1822 6160 1827 6216
rect 0 6158 1827 6160
rect 0 6128 800 6158
rect 1761 6155 1827 6158
rect 14365 6218 14431 6221
rect 24945 6218 25011 6221
rect 14365 6216 25011 6218
rect 14365 6160 14370 6216
rect 14426 6160 24950 6216
rect 25006 6160 25011 6216
rect 14365 6158 25011 6160
rect 14365 6155 14431 6158
rect 24945 6155 25011 6158
rect 28942 6156 28948 6220
rect 29012 6218 29018 6220
rect 38852 6218 39652 6248
rect 29012 6158 39652 6218
rect 29012 6156 29018 6158
rect 38852 6128 39652 6158
rect 19977 6082 20043 6085
rect 27061 6082 27127 6085
rect 19977 6080 27127 6082
rect 19977 6024 19982 6080
rect 20038 6024 27066 6080
rect 27122 6024 27127 6080
rect 19977 6022 27127 6024
rect 19977 6019 20043 6022
rect 27061 6019 27127 6022
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 5993 5946 6059 5949
rect 17493 5946 17559 5949
rect 5993 5944 17559 5946
rect 5993 5888 5998 5944
rect 6054 5888 17498 5944
rect 17554 5888 17559 5944
rect 5993 5886 17559 5888
rect 5993 5883 6059 5886
rect 17493 5883 17559 5886
rect 20437 5946 20503 5949
rect 28073 5946 28139 5949
rect 20437 5944 28139 5946
rect 20437 5888 20442 5944
rect 20498 5888 28078 5944
rect 28134 5888 28139 5944
rect 20437 5886 28139 5888
rect 20437 5883 20503 5886
rect 28073 5883 28139 5886
rect 18781 5810 18847 5813
rect 26233 5810 26299 5813
rect 18781 5808 26299 5810
rect 18781 5752 18786 5808
rect 18842 5752 26238 5808
rect 26294 5752 26299 5808
rect 18781 5750 26299 5752
rect 18781 5747 18847 5750
rect 26233 5747 26299 5750
rect 16665 5674 16731 5677
rect 19425 5674 19491 5677
rect 16665 5672 19491 5674
rect 16665 5616 16670 5672
rect 16726 5616 19430 5672
rect 19486 5616 19491 5672
rect 16665 5614 19491 5616
rect 16665 5611 16731 5614
rect 19425 5611 19491 5614
rect 24577 5674 24643 5677
rect 28942 5674 28948 5676
rect 24577 5672 28948 5674
rect 24577 5616 24582 5672
rect 24638 5616 28948 5672
rect 24577 5614 28948 5616
rect 24577 5611 24643 5614
rect 28942 5612 28948 5614
rect 29012 5612 29018 5676
rect 0 5538 800 5568
rect 4061 5538 4127 5541
rect 0 5536 4127 5538
rect 0 5480 4066 5536
rect 4122 5480 4127 5536
rect 0 5478 4127 5480
rect 0 5448 800 5478
rect 4061 5475 4127 5478
rect 6913 5538 6979 5541
rect 10133 5538 10199 5541
rect 6913 5536 10199 5538
rect 6913 5480 6918 5536
rect 6974 5480 10138 5536
rect 10194 5480 10199 5536
rect 6913 5478 10199 5480
rect 6913 5475 6979 5478
rect 10133 5475 10199 5478
rect 26969 5538 27035 5541
rect 29453 5538 29519 5541
rect 26969 5536 29519 5538
rect 26969 5480 26974 5536
rect 27030 5480 29458 5536
rect 29514 5480 29519 5536
rect 26969 5478 29519 5480
rect 26969 5475 27035 5478
rect 29453 5475 29519 5478
rect 35433 5538 35499 5541
rect 37365 5538 37431 5541
rect 35433 5536 37431 5538
rect 35433 5480 35438 5536
rect 35494 5480 37370 5536
rect 37426 5480 37431 5536
rect 35433 5478 37431 5480
rect 35433 5475 35499 5478
rect 37365 5475 37431 5478
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 16205 5266 16271 5269
rect 33133 5266 33199 5269
rect 16205 5264 33199 5266
rect 16205 5208 16210 5264
rect 16266 5208 33138 5264
rect 33194 5208 33199 5264
rect 16205 5206 33199 5208
rect 16205 5203 16271 5206
rect 33133 5203 33199 5206
rect 13 5130 79 5133
rect 21357 5130 21423 5133
rect 13 5128 21423 5130
rect 13 5072 18 5128
rect 74 5072 21362 5128
rect 21418 5072 21423 5128
rect 13 5070 21423 5072
rect 13 5067 79 5070
rect 21357 5067 21423 5070
rect 4613 4994 4679 4997
rect 17125 4994 17191 4997
rect 4613 4992 17191 4994
rect 4613 4936 4618 4992
rect 4674 4936 17130 4992
rect 17186 4936 17191 4992
rect 4613 4934 17191 4936
rect 4613 4931 4679 4934
rect 17125 4931 17191 4934
rect 31385 4994 31451 4997
rect 34605 4994 34671 4997
rect 31385 4992 34671 4994
rect 31385 4936 31390 4992
rect 31446 4936 34610 4992
rect 34666 4936 34671 4992
rect 31385 4934 34671 4936
rect 31385 4931 31451 4934
rect 34605 4931 34671 4934
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 38852 4858 39652 4888
rect 26926 4798 39652 4858
rect 7373 4722 7439 4725
rect 17217 4722 17283 4725
rect 7373 4720 17283 4722
rect 7373 4664 7378 4720
rect 7434 4664 17222 4720
rect 17278 4664 17283 4720
rect 7373 4662 17283 4664
rect 7373 4659 7439 4662
rect 17217 4659 17283 4662
rect 4061 4586 4127 4589
rect 19977 4586 20043 4589
rect 4061 4584 20043 4586
rect 4061 4528 4066 4584
rect 4122 4528 19982 4584
rect 20038 4528 20043 4584
rect 4061 4526 20043 4528
rect 4061 4523 4127 4526
rect 19977 4523 20043 4526
rect 11973 4450 12039 4453
rect 23197 4450 23263 4453
rect 11973 4448 23263 4450
rect 11973 4392 11978 4448
rect 12034 4392 23202 4448
rect 23258 4392 23263 4448
rect 11973 4390 23263 4392
rect 11973 4387 12039 4390
rect 23197 4387 23263 4390
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 11145 4314 11211 4317
rect 16113 4314 16179 4317
rect 11145 4312 16179 4314
rect 11145 4256 11150 4312
rect 11206 4256 16118 4312
rect 16174 4256 16179 4312
rect 11145 4254 16179 4256
rect 11145 4251 11211 4254
rect 16113 4251 16179 4254
rect 17217 4314 17283 4317
rect 26785 4314 26851 4317
rect 17217 4312 26851 4314
rect 17217 4256 17222 4312
rect 17278 4256 26790 4312
rect 26846 4256 26851 4312
rect 17217 4254 26851 4256
rect 17217 4251 17283 4254
rect 26785 4251 26851 4254
rect 0 4178 800 4208
rect 3509 4178 3575 4181
rect 0 4176 3575 4178
rect 0 4120 3514 4176
rect 3570 4120 3575 4176
rect 0 4118 3575 4120
rect 0 4088 800 4118
rect 3509 4115 3575 4118
rect 17125 4178 17191 4181
rect 26926 4178 26986 4798
rect 38852 4768 39652 4798
rect 29269 4450 29335 4453
rect 33041 4450 33107 4453
rect 29269 4448 33107 4450
rect 29269 4392 29274 4448
rect 29330 4392 33046 4448
rect 33102 4392 33107 4448
rect 29269 4390 33107 4392
rect 29269 4387 29335 4390
rect 33041 4387 33107 4390
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 17125 4176 26986 4178
rect 17125 4120 17130 4176
rect 17186 4120 26986 4176
rect 17125 4118 26986 4120
rect 34789 4178 34855 4181
rect 38852 4178 39652 4208
rect 34789 4176 39652 4178
rect 34789 4120 34794 4176
rect 34850 4120 39652 4176
rect 34789 4118 39652 4120
rect 17125 4115 17191 4118
rect 34789 4115 34855 4118
rect 38852 4088 39652 4118
rect 17861 4042 17927 4045
rect 35985 4042 36051 4045
rect 37733 4042 37799 4045
rect 17861 4040 24226 4042
rect 17861 3984 17866 4040
rect 17922 3984 24226 4040
rect 17861 3982 24226 3984
rect 17861 3979 17927 3982
rect 24166 3906 24226 3982
rect 35985 4040 37799 4042
rect 35985 3984 35990 4040
rect 36046 3984 37738 4040
rect 37794 3984 37799 4040
rect 35985 3982 37799 3984
rect 35985 3979 36051 3982
rect 37733 3979 37799 3982
rect 39573 3906 39639 3909
rect 24166 3904 39639 3906
rect 24166 3848 39578 3904
rect 39634 3848 39639 3904
rect 24166 3846 39639 3848
rect 39573 3843 39639 3846
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 933 3770 999 3773
rect 933 3768 14474 3770
rect 933 3712 938 3768
rect 994 3712 14474 3768
rect 933 3710 14474 3712
rect 933 3707 999 3710
rect 3969 3634 4035 3637
rect 798 3632 4035 3634
rect 798 3576 3974 3632
rect 4030 3576 4035 3632
rect 798 3574 4035 3576
rect 14414 3634 14474 3710
rect 24577 3634 24643 3637
rect 14414 3632 24643 3634
rect 14414 3576 24582 3632
rect 24638 3576 24643 3632
rect 14414 3574 24643 3576
rect 798 3528 858 3574
rect 3969 3571 4035 3574
rect 24577 3571 24643 3574
rect 0 3438 858 3528
rect 3141 3498 3207 3501
rect 35249 3498 35315 3501
rect 38852 3498 39652 3528
rect 3141 3496 34714 3498
rect 3141 3440 3146 3496
rect 3202 3440 34714 3496
rect 3141 3438 34714 3440
rect 0 3408 800 3438
rect 3141 3435 3207 3438
rect 14273 3362 14339 3365
rect 21265 3362 21331 3365
rect 14273 3360 21331 3362
rect 14273 3304 14278 3360
rect 14334 3304 21270 3360
rect 21326 3304 21331 3360
rect 14273 3302 21331 3304
rect 14273 3299 14339 3302
rect 21265 3299 21331 3302
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 17902 3226 17908 3228
rect 14414 3166 17908 3226
rect 473 3090 539 3093
rect 14414 3090 14474 3166
rect 17902 3164 17908 3166
rect 17972 3164 17978 3228
rect 27521 3226 27587 3229
rect 32765 3226 32831 3229
rect 27521 3224 32831 3226
rect 27521 3168 27526 3224
rect 27582 3168 32770 3224
rect 32826 3168 32831 3224
rect 27521 3166 32831 3168
rect 27521 3163 27587 3166
rect 32765 3163 32831 3166
rect 473 3088 14474 3090
rect 473 3032 478 3088
rect 534 3032 14474 3088
rect 473 3030 14474 3032
rect 15653 3090 15719 3093
rect 28942 3090 28948 3092
rect 15653 3088 28948 3090
rect 15653 3032 15658 3088
rect 15714 3032 28948 3088
rect 15653 3030 28948 3032
rect 473 3027 539 3030
rect 15653 3027 15719 3030
rect 28942 3028 28948 3030
rect 29012 3028 29018 3092
rect 34654 3090 34714 3438
rect 35249 3496 39652 3498
rect 35249 3440 35254 3496
rect 35310 3440 39652 3496
rect 35249 3438 39652 3440
rect 35249 3435 35315 3438
rect 38852 3408 39652 3438
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 39113 3090 39179 3093
rect 34654 3088 39179 3090
rect 34654 3032 39118 3088
rect 39174 3032 39179 3088
rect 34654 3030 39179 3032
rect 39113 3027 39179 3030
rect 10501 2954 10567 2957
rect 20161 2954 20227 2957
rect 22553 2954 22619 2957
rect 10501 2952 20040 2954
rect 10501 2896 10506 2952
rect 10562 2896 20040 2952
rect 10501 2894 20040 2896
rect 10501 2891 10567 2894
rect 0 2818 800 2848
rect 3785 2818 3851 2821
rect 0 2816 3851 2818
rect 0 2760 3790 2816
rect 3846 2760 3851 2816
rect 0 2758 3851 2760
rect 0 2728 800 2758
rect 3785 2755 3851 2758
rect 17902 2756 17908 2820
rect 17972 2818 17978 2820
rect 19425 2818 19491 2821
rect 17972 2816 19491 2818
rect 17972 2760 19430 2816
rect 19486 2760 19491 2816
rect 17972 2758 19491 2760
rect 19980 2818 20040 2894
rect 20161 2952 22619 2954
rect 20161 2896 20166 2952
rect 20222 2896 22558 2952
rect 22614 2896 22619 2952
rect 20161 2894 22619 2896
rect 20161 2891 20227 2894
rect 22553 2891 22619 2894
rect 24393 2818 24459 2821
rect 19980 2816 24459 2818
rect 19980 2760 24398 2816
rect 24454 2760 24459 2816
rect 19980 2758 24459 2760
rect 17972 2756 17978 2758
rect 19425 2755 19491 2758
rect 24393 2755 24459 2758
rect 27337 2818 27403 2821
rect 29361 2818 29427 2821
rect 27337 2816 29427 2818
rect 27337 2760 27342 2816
rect 27398 2760 29366 2816
rect 29422 2760 29427 2816
rect 27337 2758 29427 2760
rect 27337 2755 27403 2758
rect 29361 2755 29427 2758
rect 30833 2818 30899 2821
rect 35617 2818 35683 2821
rect 30833 2816 35683 2818
rect 30833 2760 30838 2816
rect 30894 2760 35622 2816
rect 35678 2760 35683 2816
rect 30833 2758 35683 2760
rect 30833 2755 30899 2758
rect 35617 2755 35683 2758
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 10174 2620 10180 2684
rect 10244 2682 10250 2684
rect 12525 2682 12591 2685
rect 10244 2680 12591 2682
rect 10244 2624 12530 2680
rect 12586 2624 12591 2680
rect 10244 2622 12591 2624
rect 10244 2620 10250 2622
rect 12525 2619 12591 2622
rect 23381 2682 23447 2685
rect 35157 2682 35223 2685
rect 23381 2680 35223 2682
rect 23381 2624 23386 2680
rect 23442 2624 35162 2680
rect 35218 2624 35223 2680
rect 23381 2622 35223 2624
rect 23381 2619 23447 2622
rect 35157 2619 35223 2622
rect 4337 2546 4403 2549
rect 8477 2546 8543 2549
rect 4337 2544 8543 2546
rect 4337 2488 4342 2544
rect 4398 2488 8482 2544
rect 8538 2488 8543 2544
rect 4337 2486 8543 2488
rect 4337 2483 4403 2486
rect 8477 2483 8543 2486
rect 10317 2546 10383 2549
rect 38193 2546 38259 2549
rect 10317 2544 38259 2546
rect 10317 2488 10322 2544
rect 10378 2488 38198 2544
rect 38254 2488 38259 2544
rect 10317 2486 38259 2488
rect 10317 2483 10383 2486
rect 38193 2483 38259 2486
rect 4061 2410 4127 2413
rect 18045 2410 18111 2413
rect 4061 2408 18111 2410
rect 4061 2352 4066 2408
rect 4122 2352 18050 2408
rect 18106 2352 18111 2408
rect 4061 2350 18111 2352
rect 4061 2347 4127 2350
rect 18045 2347 18111 2350
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
rect 38852 2138 39652 2168
rect 35436 2078 39652 2138
rect 17902 1668 17908 1732
rect 17972 1730 17978 1732
rect 17972 1670 19442 1730
rect 17972 1668 17978 1670
rect 3877 1594 3943 1597
rect 8293 1594 8359 1597
rect 3877 1592 8359 1594
rect 3877 1536 3882 1592
rect 3938 1536 8298 1592
rect 8354 1536 8359 1592
rect 3877 1534 8359 1536
rect 3877 1531 3943 1534
rect 8293 1531 8359 1534
rect 17861 1592 17927 1597
rect 17861 1536 17866 1592
rect 17922 1536 17927 1592
rect 17861 1531 17927 1536
rect 19382 1594 19442 1670
rect 35436 1594 35496 2078
rect 38852 2048 39652 2078
rect 19382 1534 35496 1594
rect 0 1458 800 1488
rect 4061 1458 4127 1461
rect 0 1456 4127 1458
rect 0 1400 4066 1456
rect 4122 1400 4127 1456
rect 0 1398 4127 1400
rect 17864 1458 17924 1531
rect 17864 1398 17970 1458
rect 0 1368 800 1398
rect 4061 1395 4127 1398
rect 17910 1324 17970 1398
rect 28942 1396 28948 1460
rect 29012 1458 29018 1460
rect 34053 1458 34119 1461
rect 29012 1456 34119 1458
rect 29012 1400 34058 1456
rect 34114 1400 34119 1456
rect 29012 1398 34119 1400
rect 29012 1396 29018 1398
rect 34053 1395 34119 1398
rect 34237 1458 34303 1461
rect 38852 1458 39652 1488
rect 34237 1456 39652 1458
rect 34237 1400 34242 1456
rect 34298 1400 39652 1456
rect 34237 1398 39652 1400
rect 34237 1395 34303 1398
rect 38852 1368 39652 1398
rect 17902 1260 17908 1324
rect 17972 1260 17978 1324
rect 17953 914 18019 917
rect 18689 914 18755 917
rect 17953 912 18755 914
rect 17953 856 17958 912
rect 18014 856 18694 912
rect 18750 856 18755 912
rect 17953 854 18755 856
rect 17953 851 18019 854
rect 18689 851 18755 854
rect 0 778 800 808
rect 1393 778 1459 781
rect 0 776 1459 778
rect 0 720 1398 776
rect 1454 720 1459 776
rect 0 718 1459 720
rect 0 688 800 718
rect 1393 715 1459 718
rect 33225 98 33291 101
rect 38852 98 39652 128
rect 33225 96 39652 98
rect 33225 40 33230 96
rect 33286 40 39652 96
rect 33225 38 39652 40
rect 33225 35 33291 38
rect 38852 8 39652 38
<< via3 >>
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 34936 39196 35000 39200
rect 34936 39140 34940 39196
rect 34940 39140 34996 39196
rect 34996 39140 35000 39196
rect 34936 39136 35000 39140
rect 35016 39196 35080 39200
rect 35016 39140 35020 39196
rect 35020 39140 35076 39196
rect 35076 39140 35080 39196
rect 35016 39136 35080 39140
rect 35096 39196 35160 39200
rect 35096 39140 35100 39196
rect 35100 39140 35156 39196
rect 35156 39140 35160 39196
rect 35096 39136 35160 39140
rect 35176 39196 35240 39200
rect 35176 39140 35180 39196
rect 35180 39140 35236 39196
rect 35236 39140 35240 39196
rect 35176 39136 35240 39140
rect 19576 38652 19640 38656
rect 19576 38596 19580 38652
rect 19580 38596 19636 38652
rect 19636 38596 19640 38652
rect 19576 38592 19640 38596
rect 19656 38652 19720 38656
rect 19656 38596 19660 38652
rect 19660 38596 19716 38652
rect 19716 38596 19720 38652
rect 19656 38592 19720 38596
rect 19736 38652 19800 38656
rect 19736 38596 19740 38652
rect 19740 38596 19796 38652
rect 19796 38596 19800 38652
rect 19736 38592 19800 38596
rect 19816 38652 19880 38656
rect 19816 38596 19820 38652
rect 19820 38596 19876 38652
rect 19876 38596 19880 38652
rect 19816 38592 19880 38596
rect 17540 38524 17604 38588
rect 10180 38388 10244 38452
rect 10916 38388 10980 38452
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 34936 38108 35000 38112
rect 34936 38052 34940 38108
rect 34940 38052 34996 38108
rect 34996 38052 35000 38108
rect 34936 38048 35000 38052
rect 35016 38108 35080 38112
rect 35016 38052 35020 38108
rect 35020 38052 35076 38108
rect 35076 38052 35080 38108
rect 35016 38048 35080 38052
rect 35096 38108 35160 38112
rect 35096 38052 35100 38108
rect 35100 38052 35156 38108
rect 35156 38052 35160 38108
rect 35096 38048 35160 38052
rect 35176 38108 35240 38112
rect 35176 38052 35180 38108
rect 35180 38052 35236 38108
rect 35236 38052 35240 38108
rect 35176 38048 35240 38052
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 16988 27160 17052 27164
rect 16988 27104 17038 27160
rect 17038 27104 17052 27160
rect 16988 27100 17052 27104
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 9444 26284 9508 26348
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 29132 25876 29196 25940
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 16804 23700 16868 23764
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 16068 22612 16132 22676
rect 16988 22340 17052 22404
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 16804 21932 16868 21996
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 9444 20028 9508 20092
rect 16988 19620 17052 19684
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 7604 19348 7668 19412
rect 16436 19348 16500 19412
rect 16988 19272 17052 19276
rect 16988 19216 17002 19272
rect 17002 19216 17052 19272
rect 16988 19212 17052 19216
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 18460 18804 18524 18868
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 17356 18124 17420 18188
rect 29132 17988 29196 18052
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 13492 16492 13556 16556
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 35572 14996 35636 15060
rect 17908 14860 17972 14924
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 3924 14648 3988 14652
rect 3924 14592 3974 14648
rect 3974 14592 3988 14648
rect 3924 14588 3988 14592
rect 16620 14180 16684 14244
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 17908 13772 17972 13836
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 16068 13500 16132 13564
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 16620 12880 16684 12884
rect 16620 12824 16634 12880
rect 16634 12824 16684 12880
rect 16620 12820 16684 12824
rect 13492 12472 13556 12476
rect 13492 12416 13506 12472
rect 13506 12416 13556 12472
rect 13492 12412 13556 12416
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 17356 12336 17420 12340
rect 17356 12280 17370 12336
rect 17370 12280 17420 12336
rect 17356 12276 17420 12280
rect 18460 12336 18524 12340
rect 18460 12280 18510 12336
rect 18510 12280 18524 12336
rect 18460 12276 18524 12280
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 17540 10780 17604 10844
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 17908 10296 17972 10300
rect 17908 10240 17922 10296
rect 17922 10240 17972 10296
rect 17908 10236 17972 10240
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 10916 6564 10980 6628
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 28948 6156 29012 6220
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 28948 5612 29012 5676
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 17908 3164 17972 3228
rect 28948 3028 29012 3092
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 17908 2756 17972 2820
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 10180 2620 10244 2684
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
rect 17908 1668 17972 1732
rect 28948 1396 29012 1460
rect 17908 1260 17972 1324
<< metal4 >>
rect 4208 39200 4528 39216
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 19568 38656 19888 39216
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 17539 38588 17605 38589
rect 17539 38524 17540 38588
rect 17604 38524 17605 38588
rect 17539 38523 17605 38524
rect 10179 38452 10245 38453
rect 10179 38388 10180 38452
rect 10244 38388 10245 38452
rect 10179 38387 10245 38388
rect 10915 38452 10981 38453
rect 10915 38388 10916 38452
rect 10980 38388 10981 38452
rect 10915 38387 10981 38388
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36212 4528 36960
rect 4208 35976 4250 36212
rect 4486 35976 4528 36212
rect 4208 35936 4528 35976
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 9443 26348 9509 26349
rect 9443 26284 9444 26348
rect 9508 26284 9509 26348
rect 9443 26283 9509 26284
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 9446 20093 9506 26283
rect 9443 20092 9509 20093
rect 9443 20028 9444 20092
rect 9508 20028 9509 20092
rect 9443 20027 9509 20028
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5576 4528 6496
rect 4208 5472 4250 5576
rect 4486 5472 4528 5576
rect 4208 5408 4216 5472
rect 4520 5408 4528 5472
rect 4208 5340 4250 5408
rect 4486 5340 4528 5408
rect 4208 4384 4528 5340
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 10182 2685 10242 38387
rect 10918 6629 10978 38387
rect 16987 27164 17053 27165
rect 16987 27100 16988 27164
rect 17052 27100 17053 27164
rect 16987 27099 17053 27100
rect 16803 23764 16869 23765
rect 16803 23700 16804 23764
rect 16868 23700 16869 23764
rect 16803 23699 16869 23700
rect 16067 22676 16133 22677
rect 16067 22612 16068 22676
rect 16132 22612 16133 22676
rect 16067 22611 16133 22612
rect 13491 16556 13557 16557
rect 13491 16492 13492 16556
rect 13556 16492 13557 16556
rect 13491 16491 13557 16492
rect 13494 12477 13554 16491
rect 16070 13565 16130 22611
rect 16806 21997 16866 23699
rect 16990 22405 17050 27099
rect 16987 22404 17053 22405
rect 16987 22340 16988 22404
rect 17052 22340 17053 22404
rect 16987 22339 17053 22340
rect 16803 21996 16869 21997
rect 16803 21932 16804 21996
rect 16868 21932 16869 21996
rect 16803 21931 16869 21932
rect 16987 19684 17053 19685
rect 16987 19620 16988 19684
rect 17052 19620 17053 19684
rect 16987 19619 17053 19620
rect 16990 19277 17050 19619
rect 16987 19276 17053 19277
rect 16987 19212 16988 19276
rect 17052 19212 17053 19276
rect 16987 19211 17053 19212
rect 17355 18188 17421 18189
rect 17355 18124 17356 18188
rect 17420 18124 17421 18188
rect 17355 18123 17421 18124
rect 16619 14244 16685 14245
rect 16619 14180 16620 14244
rect 16684 14180 16685 14244
rect 16619 14179 16685 14180
rect 16067 13564 16133 13565
rect 16067 13500 16068 13564
rect 16132 13500 16133 13564
rect 16067 13499 16133 13500
rect 16622 12885 16682 14179
rect 16619 12884 16685 12885
rect 16619 12820 16620 12884
rect 16684 12820 16685 12884
rect 16619 12819 16685 12820
rect 13491 12476 13557 12477
rect 13491 12412 13492 12476
rect 13556 12412 13557 12476
rect 13491 12411 13557 12412
rect 17358 12341 17418 18123
rect 17355 12340 17421 12341
rect 17355 12276 17356 12340
rect 17420 12276 17421 12340
rect 17355 12275 17421 12276
rect 17542 10845 17602 38523
rect 19568 37568 19888 38592
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 34928 39200 35248 39216
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 38112 35248 39136
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 37024 35248 38048
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36212 35248 36960
rect 34928 35976 34970 36212
rect 35206 35976 35248 36212
rect 34928 35936 35248 35976
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 29131 25940 29197 25941
rect 29131 25876 29132 25940
rect 29196 25876 29197 25940
rect 29131 25875 29197 25876
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20894 19888 21184
rect 19568 20658 19610 20894
rect 19846 20658 19888 20894
rect 19568 20160 19888 20658
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 18459 18868 18525 18869
rect 18459 18804 18460 18868
rect 18524 18804 18525 18868
rect 18459 18803 18525 18804
rect 17907 14924 17973 14925
rect 17907 14860 17908 14924
rect 17972 14860 17973 14924
rect 17907 14859 17973 14860
rect 17910 13837 17970 14859
rect 17907 13836 17973 13837
rect 17907 13772 17908 13836
rect 17972 13772 17973 13836
rect 17907 13771 17973 13772
rect 17539 10844 17605 10845
rect 17539 10780 17540 10844
rect 17604 10780 17605 10844
rect 17539 10779 17605 10780
rect 17910 10301 17970 13771
rect 18462 12341 18522 18803
rect 19568 17984 19888 19008
rect 29134 18053 29194 25875
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 29131 18052 29197 18053
rect 29131 17988 29132 18052
rect 29196 17988 29197 18052
rect 29131 17987 29197 17988
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 18459 12340 18525 12341
rect 18459 12276 18460 12340
rect 18524 12276 18525 12340
rect 18459 12275 18525 12276
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 17907 10300 17973 10301
rect 17907 10236 17908 10300
rect 17972 10236 17973 10300
rect 17907 10235 17973 10236
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 10915 6628 10981 6629
rect 10915 6564 10916 6628
rect 10980 6564 10981 6628
rect 10915 6563 10981 6564
rect 19568 6016 19888 7040
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 35571 15060 35637 15061
rect 35571 14996 35572 15060
rect 35636 14996 35637 15060
rect 35571 14995 35637 14996
rect 35574 14738 35634 14995
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 28947 6220 29013 6221
rect 28947 6156 28948 6220
rect 29012 6156 29013 6220
rect 28947 6155 29013 6156
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 28950 5677 29010 6155
rect 28947 5676 29013 5677
rect 28947 5612 28948 5676
rect 29012 5612 29013 5676
rect 28947 5611 29013 5612
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 17907 3228 17973 3229
rect 17907 3164 17908 3228
rect 17972 3164 17973 3228
rect 17907 3163 17973 3164
rect 17910 2821 17970 3163
rect 17907 2820 17973 2821
rect 17907 2756 17908 2820
rect 17972 2756 17973 2820
rect 17907 2755 17973 2756
rect 19568 2752 19888 3776
rect 34928 5576 35248 6496
rect 34928 5472 34970 5576
rect 35206 5472 35248 5576
rect 34928 5408 34936 5472
rect 35240 5408 35248 5472
rect 34928 5340 34970 5408
rect 35206 5340 35248 5408
rect 34928 4384 35248 5340
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 28947 3092 29013 3093
rect 28947 3028 28948 3092
rect 29012 3028 29013 3092
rect 28947 3027 29013 3028
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 10179 2684 10245 2685
rect 10179 2620 10180 2684
rect 10244 2620 10245 2684
rect 10179 2619 10245 2620
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 19568 2128 19888 2688
rect 17907 1732 17973 1733
rect 17907 1668 17908 1732
rect 17972 1668 17973 1732
rect 17907 1667 17973 1668
rect 17910 1325 17970 1667
rect 28950 1461 29010 3027
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2128 35248 2144
rect 28947 1460 29013 1461
rect 28947 1396 28948 1460
rect 29012 1396 29013 1460
rect 28947 1395 29013 1396
rect 17907 1324 17973 1325
rect 17907 1260 17908 1324
rect 17972 1260 17973 1324
rect 17907 1259 17973 1260
<< via4 >>
rect 4250 35976 4486 36212
rect 7518 19412 7754 19498
rect 7518 19348 7604 19412
rect 7604 19348 7668 19412
rect 7668 19348 7754 19412
rect 7518 19262 7754 19348
rect 3838 14652 4074 14738
rect 3838 14588 3924 14652
rect 3924 14588 3988 14652
rect 3988 14588 4074 14652
rect 3838 14502 4074 14588
rect 4250 5472 4486 5576
rect 4250 5408 4280 5472
rect 4280 5408 4296 5472
rect 4296 5408 4360 5472
rect 4360 5408 4376 5472
rect 4376 5408 4440 5472
rect 4440 5408 4456 5472
rect 4456 5408 4486 5472
rect 4250 5340 4486 5408
rect 16350 19412 16586 19498
rect 16350 19348 16436 19412
rect 16436 19348 16500 19412
rect 16500 19348 16586 19412
rect 16350 19262 16586 19348
rect 34970 35976 35206 36212
rect 19610 20658 19846 20894
rect 35486 14502 35722 14738
rect 34970 5472 35206 5576
rect 34970 5408 35000 5472
rect 35000 5408 35016 5472
rect 35016 5408 35080 5472
rect 35080 5408 35096 5472
rect 35096 5408 35160 5472
rect 35160 5408 35176 5472
rect 35176 5408 35206 5472
rect 34970 5340 35206 5408
<< metal5 >>
rect 1104 36212 38548 36254
rect 1104 35976 4250 36212
rect 4486 35976 34970 36212
rect 35206 35976 38548 36212
rect 1104 35934 38548 35976
rect 1104 20894 38548 20936
rect 1104 20658 19610 20894
rect 19846 20658 38548 20894
rect 1104 20616 38548 20658
rect 7476 19498 16628 19540
rect 7476 19262 7518 19498
rect 7754 19262 16350 19498
rect 16586 19262 16628 19498
rect 7476 19220 16628 19262
rect 3796 14738 35764 14780
rect 3796 14502 3838 14738
rect 4074 14502 35486 14738
rect 35722 14502 35764 14738
rect 3796 14460 35764 14502
rect 1104 5576 38548 5618
rect 1104 5340 4250 5576
rect 4486 5340 34970 5576
rect 35206 5340 38548 5576
rect 1104 5298 38548 5340
use sky130_fd_sc_hd__decap_3  PHY_0 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 1104 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606120353
transform 1 0 1104 0 1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__D /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 1564 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__CLK
timestamp 1606120353
transform 1 0 1932 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 1380 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 2484 0 -1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 1380 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_1_7
timestamp 1606120353
transform 1 0 1748 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_1_11
timestamp 1606120353
transform 1 0 2116 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_1_31 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 3956 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_1_23
timestamp 1606120353
transform 1 0 3220 0 1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp 1606120353
transform 1 0 4048 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1606120353
transform 1 0 3588 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1606120353
transform 1 0 3220 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__CLK
timestamp 1606120353
transform 1 0 3404 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__D
timestamp 1606120353
transform 1 0 3772 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__D
timestamp 1606120353
transform 1 0 4048 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 3956 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_1_34
timestamp 1606120353
transform 1 0 4232 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__CLK
timestamp 1606120353
transform 1 0 4416 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_1_38
timestamp 1606120353
transform 1 0 4600 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1120_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 4324 0 -1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606120353
transform 1 0 6808 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606120353
transform 1 0 6716 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54
timestamp 1606120353
transform 1 0 6072 0 -1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1606120353
transform 1 0 6900 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_1_50
timestamp 1606120353
transform 1 0 5704 0 1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_1_58
timestamp 1606120353
transform 1 0 6440 0 1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1606120353
transform 1 0 6808 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1119_
timestamp 1606120353
transform 1 0 8464 0 1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__D
timestamp 1606120353
transform 1 0 8280 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__CLK
timestamp 1606120353
transform 1 0 8464 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__CLK
timestamp 1606120353
transform 1 0 9108 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 8004 0 -1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79
timestamp 1606120353
transform 1 0 8372 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_0_82
timestamp 1606120353
transform 1 0 8648 0 -1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86
timestamp 1606120353
transform 1 0 9016 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74
timestamp 1606120353
transform 1 0 7912 0 1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_1_99
timestamp 1606120353
transform 1 0 10212 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94
timestamp 1606120353
transform 1 0 9752 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1606120353
transform 1 0 9292 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__D
timestamp 1606120353
transform 1 0 9476 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606120353
transform 1 0 9660 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_1_103
timestamp 1606120353
transform 1 0 10580 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__CLK
timestamp 1606120353
transform 1 0 10764 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__D
timestamp 1606120353
transform 1 0 10396 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_1_107
timestamp 1606120353
transform 1 0 10948 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1142_
timestamp 1606120353
transform 1 0 10028 0 -1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  FILLER_1_119
timestamp 1606120353
transform 1 0 12052 0 1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1606120353
transform 1 0 12144 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1606120353
transform 1 0 11776 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__CLK
timestamp 1606120353
transform 1 0 11960 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_0_125
timestamp 1606120353
transform 1 0 12604 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__D
timestamp 1606120353
transform 1 0 12328 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606120353
transform 1 0 12328 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606120353
transform 1 0 12512 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1606120353
transform 1 0 12420 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1217_
timestamp 1606120353
transform 1 0 12880 0 -1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__D
timestamp 1606120353
transform 1 0 15180 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__D
timestamp 1606120353
transform 1 0 14812 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__CLK
timestamp 1606120353
transform 1 0 14444 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_0_147
timestamp 1606120353
transform 1 0 14628 0 -1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_1_135
timestamp 1606120353
transform 1 0 13524 0 1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_1_143
timestamp 1606120353
transform 1 0 14260 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_1_147
timestamp 1606120353
transform 1 0 14628 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_1_151
timestamp 1606120353
transform 1 0 14996 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1139_
timestamp 1606120353
transform 1 0 15364 0 1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606120353
transform 1 0 15364 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__CLK
timestamp 1606120353
transform 1 0 15640 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156
timestamp 1606120353
transform 1 0 15456 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_0_160
timestamp 1606120353
transform 1 0 15824 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_0_172
timestamp 1606120353
transform 1 0 16928 0 -1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_1_174
timestamp 1606120353
transform 1 0 17112 0 1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1204_
timestamp 1606120353
transform 1 0 18308 0 -1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606120353
transform 1 0 18216 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606120353
transform 1 0 17940 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__D
timestamp 1606120353
transform 1 0 18032 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__CLK
timestamp 1606120353
transform 1 0 17664 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1606120353
transform 1 0 17848 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1606120353
transform 1 0 17848 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1606120353
transform 1 0 18032 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_1_196 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 19136 0 1 2720
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1215_
timestamp 1606120353
transform 1 0 19872 0 1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606120353
transform 1 0 21068 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__D
timestamp 1606120353
transform 1 0 19688 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__D
timestamp 1606120353
transform 1 0 20884 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__CLK
timestamp 1606120353
transform 1 0 20516 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_0_206
timestamp 1606120353
transform 1 0 20056 0 -1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_0_210
timestamp 1606120353
transform 1 0 20424 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1606120353
transform 1 0 20700 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_0_218
timestamp 1606120353
transform 1 0 21160 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1168_
timestamp 1606120353
transform 1 0 21436 0 -1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__D
timestamp 1606120353
transform 1 0 23092 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_0_240
timestamp 1606120353
transform 1 0 23184 0 -1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_1_223
timestamp 1606120353
transform 1 0 21620 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_1_235
timestamp 1606120353
transform 1 0 22724 0 1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_1_241
timestamp 1606120353
transform 1 0 23276 0 1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_1_249
timestamp 1606120353
transform 1 0 24012 0 1 2720
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_1_245
timestamp 1606120353
transform 1 0 23644 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_0_249
timestamp 1606120353
transform 1 0 24012 0 -1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__CLK
timestamp 1606120353
transform 1 0 23828 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606120353
transform 1 0 23552 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606120353
transform 1 0 23920 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__CLK
timestamp 1606120353
transform 1 0 24748 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__D
timestamp 1606120353
transform 1 0 24564 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_0_259
timestamp 1606120353
transform 1 0 24932 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1175_
timestamp 1606120353
transform 1 0 24748 0 1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1169_
timestamp 1606120353
transform 1 0 27140 0 -1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606120353
transform 1 0 26772 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__D
timestamp 1606120353
transform 1 0 26588 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__CLK
timestamp 1606120353
transform 1 0 26220 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_271
timestamp 1606120353
transform 1 0 26036 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_275
timestamp 1606120353
transform 1 0 26404 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_0_280
timestamp 1606120353
transform 1 0 26864 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_1_276
timestamp 1606120353
transform 1 0 26496 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1206_
timestamp 1606120353
transform 1 0 29256 0 1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606120353
transform 1 0 29164 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__D
timestamp 1606120353
transform 1 0 28980 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__CLK
timestamp 1606120353
transform 1 0 29256 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_0_302
timestamp 1606120353
transform 1 0 28888 0 -1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_0_308
timestamp 1606120353
transform 1 0 29440 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_1_288
timestamp 1606120353
transform 1 0 27600 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_1_300
timestamp 1606120353
transform 1 0 28704 0 1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606120353
transform 1 0 29624 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__CLK
timestamp 1606120353
transform 1 0 31188 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_0_311
timestamp 1606120353
transform 1 0 29716 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_0_323
timestamp 1606120353
transform 1 0 30820 0 -1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_1_325
timestamp 1606120353
transform 1 0 31004 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_1_329
timestamp 1606120353
transform 1 0 31372 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_339
timestamp 1606120353
transform 1 0 32292 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_335
timestamp 1606120353
transform 1 0 31924 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_331
timestamp 1606120353
transform 1 0 31556 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__CLK
timestamp 1606120353
transform 1 0 31740 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__D
timestamp 1606120353
transform 1 0 31556 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__D
timestamp 1606120353
transform 1 0 32108 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606120353
transform 1 0 32476 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_1_352
timestamp 1606120353
transform 1 0 33488 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_0_342
timestamp 1606120353
transform 1 0 32568 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1166_
timestamp 1606120353
transform 1 0 31740 0 1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1214_
timestamp 1606120353
transform 1 0 35420 0 -1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606120353
transform 1 0 35328 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606120353
transform 1 0 34776 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__D
timestamp 1606120353
transform 1 0 35144 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__CLK
timestamp 1606120353
transform 1 0 34776 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_0_354
timestamp 1606120353
transform 1 0 33672 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_0_368
timestamp 1606120353
transform 1 0 34960 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_1_364
timestamp 1606120353
transform 1 0 34592 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_1_367
timestamp 1606120353
transform 1 0 34868 0 1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1212_
timestamp 1606120353
transform 1 0 35788 0 1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__D
timestamp 1606120353
transform 1 0 35604 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_0_392
timestamp 1606120353
transform 1 0 37168 0 -1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_1_396
timestamp 1606120353
transform 1 0 37536 0 1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606120353
transform -1 0 38548 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606120353
transform -1 0 38548 0 1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606120353
transform 1 0 38180 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_0_400
timestamp 1606120353
transform 1 0 37904 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1218_
timestamp 1606120353
transform 1 0 1472 0 -1 3808
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606120353
transform 1 0 1104 0 -1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1606120353
transform 1 0 1380 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1200_
timestamp 1606120353
transform 1 0 4048 0 -1 3808
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606120353
transform 1 0 3956 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_2_23
timestamp 1606120353
transform 1 0 3220 0 -1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_2_51
timestamp 1606120353
transform 1 0 5796 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_63
timestamp 1606120353
transform 1 0 6900 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__CLK
timestamp 1606120353
transform 1 0 8372 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_2_75
timestamp 1606120353
transform 1 0 8004 0 -1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_2_81
timestamp 1606120353
transform 1 0 8556 0 -1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1201_
timestamp 1606120353
transform 1 0 10120 0 -1 3808
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606120353
transform 1 0 9568 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1606120353
transform 1 0 9292 0 -1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_2_93
timestamp 1606120353
transform 1 0 9660 0 -1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_2_97
timestamp 1606120353
transform 1 0 10028 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1606120353
transform 1 0 11868 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1606120353
transform 1 0 12972 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1227_
timestamp 1606120353
transform 1 0 15272 0 -1 3808
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606120353
transform 1 0 15180 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1606120353
transform 1 0 14076 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_173
timestamp 1606120353
transform 1 0 17020 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__CLK
timestamp 1606120353
transform 1 0 19136 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_2_185
timestamp 1606120353
transform 1 0 18124 0 -1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_2_193
timestamp 1606120353
transform 1 0 18860 0 -1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_2_198
timestamp 1606120353
transform 1 0 19320 0 -1 3808
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606120353
transform 1 0 20792 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__CLK
timestamp 1606120353
transform 1 0 19872 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_2_206
timestamp 1606120353
transform 1 0 20056 0 -1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1606120353
transform 1 0 20884 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1211_
timestamp 1606120353
transform 1 0 23092 0 -1 3808
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1606120353
transform 1 0 21988 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__CLK
timestamp 1606120353
transform 1 0 25392 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_2_258
timestamp 1606120353
transform 1 0 24840 0 -1 3808
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606120353
transform 1 0 26404 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__CLK
timestamp 1606120353
transform 1 0 26680 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_2_266
timestamp 1606120353
transform 1 0 25576 0 -1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_2_274
timestamp 1606120353
transform 1 0 26312 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_2_276
timestamp 1606120353
transform 1 0 26496 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_2_280
timestamp 1606120353
transform 1 0 26864 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_292
timestamp 1606120353
transform 1 0 27968 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_304
timestamp 1606120353
transform 1 0 29072 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_316
timestamp 1606120353
transform 1 0 30176 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_2_328
timestamp 1606120353
transform 1 0 31280 0 -1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1202_
timestamp 1606120353
transform 1 0 32108 0 -1 3808
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606120353
transform 1 0 32016 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_2_356
timestamp 1606120353
transform 1 0 33856 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_2_368
timestamp 1606120353
transform 1 0 34960 0 -1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__CLK
timestamp 1606120353
transform 1 0 35788 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_2_376
timestamp 1606120353
transform 1 0 35696 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_2_379
timestamp 1606120353
transform 1 0 35972 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_2_391
timestamp 1606120353
transform 1 0 37076 0 -1 3808
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606120353
transform -1 0 38548 0 -1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606120353
transform 1 0 37628 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_2_398
timestamp 1606120353
transform 1 0 37720 0 -1 3808
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606120353
transform 1 0 1104 0 1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606120353
transform 1 0 1380 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1606120353
transform 1 0 2484 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1606120353
transform 1 0 3588 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1606120353
transform 1 0 4692 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606120353
transform 1 0 6716 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1606120353
transform 1 0 5796 0 1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606120353
transform 1 0 6532 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1606120353
transform 1 0 6808 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1125_
timestamp 1606120353
transform 1 0 8372 0 1 3808
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__D
timestamp 1606120353
transform 1 0 8188 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_3_74
timestamp 1606120353
transform 1 0 7912 0 1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__D
timestamp 1606120353
transform 1 0 10764 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__CLK
timestamp 1606120353
transform 1 0 11132 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_3_98
timestamp 1606120353
transform 1 0 10120 0 1 3808
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_3_104
timestamp 1606120353
transform 1 0 10672 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_3_107
timestamp 1606120353
transform 1 0 10948 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606120353
transform 1 0 12328 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_3_111
timestamp 1606120353
transform 1 0 11316 0 1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1606120353
transform 1 0 12052 0 1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1606120353
transform 1 0 12420 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1606120353
transform 1 0 13524 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1606120353
transform 1 0 14628 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1606120353
transform 1 0 15732 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_3_171
timestamp 1606120353
transform 1 0 16836 0 1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1198_
timestamp 1606120353
transform 1 0 19136 0 1 3808
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606120353
transform 1 0 17940 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__D
timestamp 1606120353
transform 1 0 18952 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__D
timestamp 1606120353
transform 1 0 17756 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__CLK
timestamp 1606120353
transform 1 0 18216 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1606120353
transform 1 0 17572 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_184
timestamp 1606120353
transform 1 0 18032 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_3_188
timestamp 1606120353
transform 1 0 18400 0 1 3808
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_3_215
timestamp 1606120353
transform 1 0 20884 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_227
timestamp 1606120353
transform 1 0 21988 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_3_239
timestamp 1606120353
transform 1 0 23092 0 1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1176_
timestamp 1606120353
transform 1 0 25392 0 1 3808
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606120353
transform 1 0 23552 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__D
timestamp 1606120353
transform 1 0 25208 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_3_243
timestamp 1606120353
transform 1 0 23460 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1606120353
transform 1 0 23644 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_3_257
timestamp 1606120353
transform 1 0 24748 0 1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_3_261
timestamp 1606120353
transform 1 0 25116 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__D
timestamp 1606120353
transform 1 0 27324 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_283
timestamp 1606120353
transform 1 0 27140 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606120353
transform 1 0 29164 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_3_287
timestamp 1606120353
transform 1 0 27508 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_3_299
timestamp 1606120353
transform 1 0 28612 0 1 3808
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_3_306
timestamp 1606120353
transform 1 0 29256 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_318
timestamp 1606120353
transform 1 0 30360 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_3_330
timestamp 1606120353
transform 1 0 31464 0 1 3808
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__D
timestamp 1606120353
transform 1 0 32108 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__CLK
timestamp 1606120353
transform 1 0 32476 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_3_336
timestamp 1606120353
transform 1 0 32016 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_3_339
timestamp 1606120353
transform 1 0 32292 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_3_343
timestamp 1606120353
transform 1 0 32660 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606120353
transform 1 0 34776 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_3_355
timestamp 1606120353
transform 1 0 33764 0 1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_3_363
timestamp 1606120353
transform 1 0 34500 0 1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_3_367
timestamp 1606120353
transform 1 0 34868 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_379
timestamp 1606120353
transform 1 0 35972 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_391
timestamp 1606120353
transform 1 0 37076 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606120353
transform -1 0 38548 0 1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_3_403
timestamp 1606120353
transform 1 0 38180 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606120353
transform 1 0 1104 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606120353
transform 1 0 1380 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1606120353
transform 1 0 2484 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606120353
transform 1 0 3956 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1606120353
transform 1 0 3588 0 -1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1606120353
transform 1 0 4048 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1606120353
transform 1 0 5152 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1606120353
transform 1 0 6256 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__CLK
timestamp 1606120353
transform 1 0 8832 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1606120353
transform 1 0 7360 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1606120353
transform 1 0 8464 0 -1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_4_86
timestamp 1606120353
transform 1 0 9016 0 -1 4896
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1143_
timestamp 1606120353
transform 1 0 10764 0 -1 4896
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606120353
transform 1 0 9568 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1606120353
transform 1 0 9660 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_124
timestamp 1606120353
transform 1 0 12512 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606120353
transform 1 0 15180 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_4_136
timestamp 1606120353
transform 1 0 13616 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1606120353
transform 1 0 14720 0 -1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1606120353
transform 1 0 15088 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1606120353
transform 1 0 15272 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1606120353
transform 1 0 16376 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1135_
timestamp 1606120353
transform 1 0 17756 0 -1 4896
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  FILLER_4_178
timestamp 1606120353
transform 1 0 17480 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606120353
transform 1 0 20792 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_4_200
timestamp 1606120353
transform 1 0 19504 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1606120353
transform 1 0 20608 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1606120353
transform 1 0 20884 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1606120353
transform 1 0 21988 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1606120353
transform 1 0 23092 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1606120353
transform 1 0 24196 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1606120353
transform 1 0 25300 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1220_
timestamp 1606120353
transform 1 0 26496 0 -1 4896
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606120353
transform 1 0 26404 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_4_295
timestamp 1606120353
transform 1 0 28244 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_307
timestamp 1606120353
transform 1 0 29348 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_319
timestamp 1606120353
transform 1 0 30452 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1188_
timestamp 1606120353
transform 1 0 32108 0 -1 4896
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606120353
transform 1 0 32016 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_4_331
timestamp 1606120353
transform 1 0 31556 0 -1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_4_335
timestamp 1606120353
transform 1 0 31924 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_4_356
timestamp 1606120353
transform 1 0 33856 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_368
timestamp 1606120353
transform 1 0 34960 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_380
timestamp 1606120353
transform 1 0 36064 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_4_392
timestamp 1606120353
transform 1 0 37168 0 -1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_4_396
timestamp 1606120353
transform 1 0 37536 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606120353
transform -1 0 38548 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606120353
transform 1 0 37628 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_4_398
timestamp 1606120353
transform 1 0 37720 0 -1 4896
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606120353
transform 1 0 1104 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606120353
transform 1 0 1380 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606120353
transform 1 0 2484 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1606120353
transform 1 0 3588 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1606120353
transform 1 0 4692 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606120353
transform 1 0 6716 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1606120353
transform 1 0 5796 0 1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606120353
transform 1 0 6532 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1606120353
transform 1 0 6808 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1131_
timestamp 1606120353
transform 1 0 8832 0 1 4896
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__D
timestamp 1606120353
transform 1 0 8648 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_5_74
timestamp 1606120353
transform 1 0 7912 0 1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_5_103
timestamp 1606120353
transform 1 0 10580 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606120353
transform 1 0 12328 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__D
timestamp 1606120353
transform 1 0 12696 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__CLK
timestamp 1606120353
transform 1 0 13064 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_5_115
timestamp 1606120353
transform 1 0 11684 0 1 4896
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1606120353
transform 1 0 12236 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_5_123
timestamp 1606120353
transform 1 0 12420 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_5_128
timestamp 1606120353
transform 1 0 12880 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_5_132
timestamp 1606120353
transform 1 0 13248 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_144
timestamp 1606120353
transform 1 0 14352 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__D
timestamp 1606120353
transform 1 0 15640 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__CLK
timestamp 1606120353
transform 1 0 16008 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_156
timestamp 1606120353
transform 1 0 15456 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_160
timestamp 1606120353
transform 1 0 15824 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_5_164
timestamp 1606120353
transform 1 0 16192 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_5_176
timestamp 1606120353
transform 1 0 17296 0 1 4896
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606120353
transform 1 0 17940 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1606120353
transform 1 0 17848 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1606120353
transform 1 0 18032 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1606120353
transform 1 0 19136 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1606120353
transform 1 0 20240 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_5_220
timestamp 1606120353
transform 1 0 21344 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_clk /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 21620 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_clk_A
timestamp 1606120353
transform 1 0 22080 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_226
timestamp 1606120353
transform 1 0 21896 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_5_230
timestamp 1606120353
transform 1 0 22264 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_5_242
timestamp 1606120353
transform 1 0 23368 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606120353
transform 1 0 23552 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_clk
timestamp 1606120353
transform 1 0 25392 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_clk_A
timestamp 1606120353
transform 1 0 23828 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_245
timestamp 1606120353
transform 1 0 23644 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1606120353
transform 1 0 24012 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_5_261
timestamp 1606120353
transform 1 0 25116 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_clk_A
timestamp 1606120353
transform 1 0 25852 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_267
timestamp 1606120353
transform 1 0 25668 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_5_271
timestamp 1606120353
transform 1 0 26036 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_283
timestamp 1606120353
transform 1 0 27140 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606120353
transform 1 0 29164 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_5_295
timestamp 1606120353
transform 1 0 28244 0 1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_5_303
timestamp 1606120353
transform 1 0 28980 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_5_306
timestamp 1606120353
transform 1 0 29256 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_318
timestamp 1606120353
transform 1 0 30360 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_330
timestamp 1606120353
transform 1 0 31464 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_342
timestamp 1606120353
transform 1 0 32568 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606120353
transform 1 0 34776 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_5_354
timestamp 1606120353
transform 1 0 33672 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_367
timestamp 1606120353
transform 1 0 34868 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_379
timestamp 1606120353
transform 1 0 35972 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_391
timestamp 1606120353
transform 1 0 37076 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606120353
transform -1 0 38548 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_5_403
timestamp 1606120353
transform 1 0 38180 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606120353
transform 1 0 1104 0 -1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606120353
transform 1 0 1104 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606120353
transform 1 0 1380 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606120353
transform 1 0 2484 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606120353
transform 1 0 1380 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1606120353
transform 1 0 2484 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606120353
transform 1 0 3956 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606120353
transform 1 0 3588 0 -1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1606120353
transform 1 0 4048 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1606120353
transform 1 0 5152 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1606120353
transform 1 0 3588 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1606120353
transform 1 0 4692 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1606120353
transform 1 0 6716 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1606120353
transform 1 0 6256 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1606120353
transform 1 0 5796 0 1 5984
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606120353
transform 1 0 6532 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_7_62
timestamp 1606120353
transform 1 0 6808 0 1 5984
box 0 -48 736 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_clk
timestamp 1606120353
transform 1 0 7636 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_clk_A
timestamp 1606120353
transform 1 0 8096 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1606120353
transform 1 0 7360 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1606120353
transform 1 0 8464 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_7_70
timestamp 1606120353
transform 1 0 7544 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_7_74
timestamp 1606120353
transform 1 0 7912 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_7_78
timestamp 1606120353
transform 1 0 8280 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_7_96
timestamp 1606120353
transform 1 0 9936 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_7_90
timestamp 1606120353
transform 1 0 9384 0 1 5984
box 0 -48 552 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_clk
timestamp 1606120353
transform 1 0 10028 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606120353
transform 1 0 9568 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_7_108
timestamp 1606120353
transform 1 0 11040 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_7_104
timestamp 1606120353
transform 1 0 10672 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_7_100
timestamp 1606120353
transform 1 0 10304 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__CLK
timestamp 1606120353
transform 1 0 11224 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_clk_A
timestamp 1606120353
transform 1 0 10856 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__D
timestamp 1606120353
transform 1 0 10488 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1606120353
transform 1 0 10764 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1606120353
transform 1 0 9660 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_7_112
timestamp 1606120353
transform 1 0 11408 0 1 5984
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_6_117
timestamp 1606120353
transform 1 0 11868 0 -1 5984
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A2
timestamp 1606120353
transform 1 0 12144 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_7_132
timestamp 1606120353
transform 1 0 13248 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_7_128
timestamp 1606120353
transform 1 0 12880 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_7_123
timestamp 1606120353
transform 1 0 12420 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_6_125
timestamp 1606120353
transform 1 0 12604 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__B2
timestamp 1606120353
transform 1 0 12696 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A1
timestamp 1606120353
transform 1 0 13064 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1606120353
transform 1 0 12328 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1094_
timestamp 1606120353
transform 1 0 12696 0 -1 5984
box 0 -48 1748 592
use sky130_fd_sc_hd__o22a_4  _0789_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 14076 0 1 5984
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606120353
transform 1 0 15180 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A1
timestamp 1606120353
transform 1 0 13892 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__B1
timestamp 1606120353
transform 1 0 13432 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__B2
timestamp 1606120353
transform 1 0 14628 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_6_145
timestamp 1606120353
transform 1 0 14444 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1606120353
transform 1 0 14812 0 -1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_6_154
timestamp 1606120353
transform 1 0 15272 0 -1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_7_136
timestamp 1606120353
transform 1 0 13616 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_7_165
timestamp 1606120353
transform 1 0 16284 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_7_161
timestamp 1606120353
transform 1 0 15916 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_7_155
timestamp 1606120353
transform 1 0 15364 0 1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B1
timestamp 1606120353
transform 1 0 15732 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B2
timestamp 1606120353
transform 1 0 16100 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_7_173
timestamp 1606120353
transform 1 0 17020 0 1 5984
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1606120353
transform 1 0 16652 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A2
timestamp 1606120353
transform 1 0 16836 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A1
timestamp 1606120353
transform 1 0 16468 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1103_
timestamp 1606120353
transform 1 0 15640 0 -1 5984
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_4  FILLER_7_184
timestamp 1606120353
transform 1 0 18032 0 1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__B2
timestamp 1606120353
transform 1 0 17756 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1606120353
transform 1 0 17940 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_7_191
timestamp 1606120353
transform 1 0 18676 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_7_188
timestamp 1606120353
transform 1 0 18400 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_6_195
timestamp 1606120353
transform 1 0 19044 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_6_191
timestamp 1606120353
transform 1 0 18676 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__CLK
timestamp 1606120353
transform 1 0 19228 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A2
timestamp 1606120353
transform 1 0 18860 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__B1
timestamp 1606120353
transform 1 0 18492 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A1
timestamp 1606120353
transform 1 0 18492 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__D
timestamp 1606120353
transform 1 0 18860 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1606120353
transform 1 0 17388 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1133_
timestamp 1606120353
transform 1 0 19044 0 1 5984
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606120353
transform 1 0 20792 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_6_199
timestamp 1606120353
transform 1 0 19412 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_6_211
timestamp 1606120353
transform 1 0 20516 0 -1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1606120353
transform 1 0 20884 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_214
timestamp 1606120353
transform 1 0 20792 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__D
timestamp 1606120353
transform 1 0 22172 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__CLK
timestamp 1606120353
transform 1 0 22540 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1606120353
transform 1 0 21988 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_6_239
timestamp 1606120353
transform 1 0 23092 0 -1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_7_226
timestamp 1606120353
transform 1 0 21896 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_7_231
timestamp 1606120353
transform 1 0 22356 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_7_235
timestamp 1606120353
transform 1 0 22724 0 1 5984
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1606120353
transform 1 0 23552 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_clk
timestamp 1606120353
transform 1 0 23460 0 -1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_6_246
timestamp 1606120353
transform 1 0 23736 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_258
timestamp 1606120353
transform 1 0 24840 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_7_243
timestamp 1606120353
transform 1 0 23460 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1606120353
transform 1 0 23644 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1606120353
transform 1 0 24748 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606120353
transform 1 0 26404 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__D
timestamp 1606120353
transform 1 0 27048 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__CLK
timestamp 1606120353
transform 1 0 27416 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_6_270
timestamp 1606120353
transform 1 0 25944 0 -1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_6_274
timestamp 1606120353
transform 1 0 26312 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_6_276
timestamp 1606120353
transform 1 0 26496 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_269
timestamp 1606120353
transform 1 0 25852 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_7_281
timestamp 1606120353
transform 1 0 26956 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_7_284
timestamp 1606120353
transform 1 0 27232 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1606120353
transform 1 0 29164 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_6_288
timestamp 1606120353
transform 1 0 27600 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_300
timestamp 1606120353
transform 1 0 28704 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_288
timestamp 1606120353
transform 1 0 27600 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_7_300
timestamp 1606120353
transform 1 0 28704 0 1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_7_304
timestamp 1606120353
transform 1 0 29072 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_7_306
timestamp 1606120353
transform 1 0 29256 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_312
timestamp 1606120353
transform 1 0 29808 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_324
timestamp 1606120353
transform 1 0 30912 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_318
timestamp 1606120353
transform 1 0 30360 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_330
timestamp 1606120353
transform 1 0 31464 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606120353
transform 1 0 32016 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_6_337
timestamp 1606120353
transform 1 0 32108 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_349
timestamp 1606120353
transform 1 0 33212 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_342
timestamp 1606120353
transform 1 0 32568 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1606120353
transform 1 0 34776 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_6_361
timestamp 1606120353
transform 1 0 34316 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_373
timestamp 1606120353
transform 1 0 35420 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_354
timestamp 1606120353
transform 1 0 33672 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_367
timestamp 1606120353
transform 1 0 34868 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_385
timestamp 1606120353
transform 1 0 36524 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_379
timestamp 1606120353
transform 1 0 35972 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_391
timestamp 1606120353
transform 1 0 37076 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606120353
transform -1 0 38548 0 -1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606120353
transform -1 0 38548 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606120353
transform 1 0 37628 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_6_398
timestamp 1606120353
transform 1 0 37720 0 -1 5984
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_7_403
timestamp 1606120353
transform 1 0 38180 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606120353
transform 1 0 1104 0 -1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1606120353
transform 1 0 1380 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1606120353
transform 1 0 2484 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1606120353
transform 1 0 3956 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606120353
transform 1 0 3588 0 -1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1606120353
transform 1 0 4048 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1606120353
transform 1 0 5152 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1606120353
transform 1 0 6256 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1606120353
transform 1 0 7360 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_8_80
timestamp 1606120353
transform 1 0 8464 0 -1 7072
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_8_88
timestamp 1606120353
transform 1 0 9200 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1093_
timestamp 1606120353
transform 1 0 10488 0 -1 7072
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1606120353
transform 1 0 9568 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__B1
timestamp 1606120353
transform 1 0 10304 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__A2
timestamp 1606120353
transform 1 0 9936 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__CLK
timestamp 1606120353
transform 1 0 9384 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_8_93
timestamp 1606120353
transform 1 0 9660 0 -1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_8_98
timestamp 1606120353
transform 1 0 10120 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _0794_
timestamp 1606120353
transform 1 0 13064 0 -1 7072
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__D
timestamp 1606120353
transform 1 0 12880 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__CLK
timestamp 1606120353
transform 1 0 12512 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_8_121
timestamp 1606120353
transform 1 0 12236 0 -1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_8_126
timestamp 1606120353
transform 1 0 12696 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1606120353
transform 1 0 15180 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__B1
timestamp 1606120353
transform 1 0 14536 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A2
timestamp 1606120353
transform 1 0 14904 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_144
timestamp 1606120353
transform 1 0 14352 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_148
timestamp 1606120353
transform 1 0 14720 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1606120353
transform 1 0 15088 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_8_154
timestamp 1606120353
transform 1 0 15272 0 -1 7072
box 0 -48 736 592
use sky130_fd_sc_hd__o22a_4  _0807_
timestamp 1606120353
transform 1 0 16100 0 -1 7072
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_1  FILLER_8_162
timestamp 1606120353
transform 1 0 16008 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _0796_
timestamp 1606120353
transform 1 0 18492 0 -1 7072
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1606120353
transform 1 0 17388 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1606120353
transform 1 0 20792 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A1
timestamp 1606120353
transform 1 0 21068 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__D
timestamp 1606120353
transform 1 0 20148 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_8_203
timestamp 1606120353
transform 1 0 19780 0 -1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_8_209
timestamp 1606120353
transform 1 0 20332 0 -1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1606120353
transform 1 0 20700 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_8_215
timestamp 1606120353
transform 1 0 20884 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_219
timestamp 1606120353
transform 1 0 21252 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1144_
timestamp 1606120353
transform 1 0 22172 0 -1 7072
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A2
timestamp 1606120353
transform 1 0 21436 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_8_223
timestamp 1606120353
transform 1 0 21620 0 -1 7072
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_8_248
timestamp 1606120353
transform 1 0 23920 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_260
timestamp 1606120353
transform 1 0 25024 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1167_
timestamp 1606120353
transform 1 0 27048 0 -1 7072
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1606120353
transform 1 0 26404 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_8_272
timestamp 1606120353
transform 1 0 26128 0 -1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_8_276
timestamp 1606120353
transform 1 0 26496 0 -1 7072
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_8_301
timestamp 1606120353
transform 1 0 28796 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_313
timestamp 1606120353
transform 1 0 29900 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_8_325
timestamp 1606120353
transform 1 0 31004 0 -1 7072
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1606120353
transform 1 0 32016 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_8_333
timestamp 1606120353
transform 1 0 31740 0 -1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_8_337
timestamp 1606120353
transform 1 0 32108 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_349
timestamp 1606120353
transform 1 0 33212 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_361
timestamp 1606120353
transform 1 0 34316 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_373
timestamp 1606120353
transform 1 0 35420 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_385
timestamp 1606120353
transform 1 0 36524 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606120353
transform -1 0 38548 0 -1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1606120353
transform 1 0 37628 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_8_398
timestamp 1606120353
transform 1 0 37720 0 -1 7072
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606120353
transform 1 0 1104 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606120353
transform 1 0 1380 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1606120353
transform 1 0 2484 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1606120353
transform 1 0 3588 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1606120353
transform 1 0 4692 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1606120353
transform 1 0 6716 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1606120353
transform 1 0 5796 0 1 7072
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1606120353
transform 1 0 6532 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1606120353
transform 1 0 6808 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_clk
timestamp 1606120353
transform 1 0 8648 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_clk_A
timestamp 1606120353
transform 1 0 8464 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_9_74
timestamp 1606120353
transform 1 0 7912 0 1 7072
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILLER_9_85
timestamp 1606120353
transform 1 0 8924 0 1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__o22a_4  _0786_
timestamp 1606120353
transform 1 0 10304 0 1 7072
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__A1
timestamp 1606120353
transform 1 0 10120 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__B2
timestamp 1606120353
transform 1 0 9752 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__D
timestamp 1606120353
transform 1 0 9384 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_9_89
timestamp 1606120353
transform 1 0 9292 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_9_92
timestamp 1606120353
transform 1 0 9568 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_96
timestamp 1606120353
transform 1 0 9936 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1096_
timestamp 1606120353
transform 1 0 12880 0 1 7072
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1606120353
transform 1 0 12328 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A1
timestamp 1606120353
transform 1 0 12144 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A2
timestamp 1606120353
transform 1 0 12604 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__B1
timestamp 1606120353
transform 1 0 11776 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1606120353
transform 1 0 11592 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1606120353
transform 1 0 11960 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1606120353
transform 1 0 12420 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_9_127
timestamp 1606120353
transform 1 0 12788 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__D
timestamp 1606120353
transform 1 0 15272 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__CLK
timestamp 1606120353
transform 1 0 14904 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_9_147
timestamp 1606120353
transform 1 0 14628 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_9_152
timestamp 1606120353
transform 1 0 15088 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__B2
timestamp 1606120353
transform 1 0 15916 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__B1
timestamp 1606120353
transform 1 0 16284 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_9_156
timestamp 1606120353
transform 1 0 15456 0 1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_9_160
timestamp 1606120353
transform 1 0 15824 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_9_163
timestamp 1606120353
transform 1 0 16100 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_9_167
timestamp 1606120353
transform 1 0 16468 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1606120353
transform 1 0 17940 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__D
timestamp 1606120353
transform 1 0 17756 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__CLK
timestamp 1606120353
transform 1 0 18216 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 1606120353
transform 1 0 17572 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_184
timestamp 1606120353
transform 1 0 18032 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_9_188
timestamp 1606120353
transform 1 0 18400 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1101_
timestamp 1606120353
transform 1 0 20148 0 1 7072
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__B2
timestamp 1606120353
transform 1 0 19964 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_9_200
timestamp 1606120353
transform 1 0 19504 0 1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_9_204
timestamp 1606120353
transform 1 0 19872 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__B1
timestamp 1606120353
transform 1 0 22080 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_clk_A
timestamp 1606120353
transform 1 0 22908 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_226
timestamp 1606120353
transform 1 0 21896 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_9_230
timestamp 1606120353
transform 1 0 22264 0 1 7072
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_9_236
timestamp 1606120353
transform 1 0 22816 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_9_239
timestamp 1606120353
transform 1 0 23092 0 1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1606120353
transform 1 0 23552 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_9_243
timestamp 1606120353
transform 1 0 23460 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1606120353
transform 1 0 23644 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1606120353
transform 1 0 24748 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_269
timestamp 1606120353
transform 1 0 25852 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1606120353
transform 1 0 26956 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1606120353
transform 1 0 29164 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1606120353
transform 1 0 28060 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_306
timestamp 1606120353
transform 1 0 29256 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_318
timestamp 1606120353
transform 1 0 30360 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_330
timestamp 1606120353
transform 1 0 31464 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_342
timestamp 1606120353
transform 1 0 32568 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1606120353
transform 1 0 34776 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_9_354
timestamp 1606120353
transform 1 0 33672 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_367
timestamp 1606120353
transform 1 0 34868 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_379
timestamp 1606120353
transform 1 0 35972 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_391
timestamp 1606120353
transform 1 0 37076 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606120353
transform -1 0 38548 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_9_403
timestamp 1606120353
transform 1 0 38180 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606120353
transform 1 0 1104 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1606120353
transform 1 0 1380 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1606120353
transform 1 0 2484 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1606120353
transform 1 0 3956 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1606120353
transform 1 0 3588 0 -1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1606120353
transform 1 0 4048 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1606120353
transform 1 0 5152 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1606120353
transform 1 0 6256 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A1
timestamp 1606120353
transform 1 0 8924 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1606120353
transform 1 0 7360 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1606120353
transform 1 0 8464 0 -1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_10_84
timestamp 1606120353
transform 1 0 8832 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1606120353
transform 1 0 9108 0 -1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1109_
timestamp 1606120353
transform 1 0 9660 0 -1 8160
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1606120353
transform 1 0 9568 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1606120353
transform 1 0 9476 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__a21o_4  _0784_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 12144 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_10_112
timestamp 1606120353
transform 1 0 11408 0 -1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_10_132
timestamp 1606120353
transform 1 0 13248 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1111_
timestamp 1606120353
transform 1 0 15272 0 -1 8160
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1606120353
transform 1 0 15180 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__A2
timestamp 1606120353
transform 1 0 13432 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__B1
timestamp 1606120353
transform 1 0 13800 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__B1
timestamp 1606120353
transform 1 0 14996 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_10_136
timestamp 1606120353
transform 1 0 13616 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_10_140
timestamp 1606120353
transform 1 0 13984 0 -1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_10_148
timestamp 1606120353
transform 1 0 14720 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_10_173
timestamp 1606120353
transform 1 0 17020 0 -1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1097_
timestamp 1606120353
transform 1 0 17756 0 -1 8160
box 0 -48 1748 592
use sky130_fd_sc_hd__o22a_4  _0804_
timestamp 1606120353
transform 1 0 20884 0 -1 8160
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1606120353
transform 1 0 20792 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__CLK
timestamp 1606120353
transform 1 0 20148 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_10_200
timestamp 1606120353
transform 1 0 19504 0 -1 8160
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_10_206
timestamp 1606120353
transform 1 0 20056 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_10_209
timestamp 1606120353
transform 1 0 20332 0 -1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1606120353
transform 1 0 20700 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_clk
timestamp 1606120353
transform 1 0 22908 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_10_229
timestamp 1606120353
transform 1 0 22172 0 -1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_10_240
timestamp 1606120353
transform 1 0 23184 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_252
timestamp 1606120353
transform 1 0 24288 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_10_264
timestamp 1606120353
transform 1 0 25392 0 -1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1606120353
transform 1 0 26404 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_10_272
timestamp 1606120353
transform 1 0 26128 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_10_276
timestamp 1606120353
transform 1 0 26496 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_288
timestamp 1606120353
transform 1 0 27600 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_300
timestamp 1606120353
transform 1 0 28704 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_312
timestamp 1606120353
transform 1 0 29808 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_324
timestamp 1606120353
transform 1 0 30912 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1606120353
transform 1 0 32016 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_10_337
timestamp 1606120353
transform 1 0 32108 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_349
timestamp 1606120353
transform 1 0 33212 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_361
timestamp 1606120353
transform 1 0 34316 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_373
timestamp 1606120353
transform 1 0 35420 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_385
timestamp 1606120353
transform 1 0 36524 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606120353
transform -1 0 38548 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1606120353
transform 1 0 37628 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_10_398
timestamp 1606120353
transform 1 0 37720 0 -1 8160
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606120353
transform 1 0 1104 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1606120353
transform 1 0 1380 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1606120353
transform 1 0 2484 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1606120353
transform 1 0 3588 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1606120353
transform 1 0 4692 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1606120353
transform 1 0 6716 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__D
timestamp 1606120353
transform 1 0 7084 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__A
timestamp 1606120353
transform 1 0 6072 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_11_51
timestamp 1606120353
transform 1 0 5796 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_11_56
timestamp 1606120353
transform 1 0 6256 0 1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1606120353
transform 1 0 6624 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_11_62
timestamp 1606120353
transform 1 0 6808 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__o22a_4  _0816_
timestamp 1606120353
transform 1 0 8924 0 1 8160
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__B1
timestamp 1606120353
transform 1 0 8740 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__B2
timestamp 1606120353
transform 1 0 8372 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__CLK
timestamp 1606120353
transform 1 0 7452 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_67
timestamp 1606120353
transform 1 0 7268 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_11_71
timestamp 1606120353
transform 1 0 7636 0 1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_11_81
timestamp 1606120353
transform 1 0 8556 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A1_N
timestamp 1606120353
transform 1 0 10856 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__B1
timestamp 1606120353
transform 1 0 11224 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A2_N
timestamp 1606120353
transform 1 0 10488 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_11_99
timestamp 1606120353
transform 1 0 10212 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_11_104
timestamp 1606120353
transform 1 0 10672 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_108
timestamp 1606120353
transform 1 0 11040 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_11_116
timestamp 1606120353
transform 1 0 11776 0 1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_11_112
timestamp 1606120353
transform 1 0 11408 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A
timestamp 1606120353
transform 1 0 12144 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__B2
timestamp 1606120353
transform 1 0 11592 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_128
timestamp 1606120353
transform 1 0 12880 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_11_123
timestamp 1606120353
transform 1 0 12420 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__A1
timestamp 1606120353
transform 1 0 12696 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__B
timestamp 1606120353
transform 1 0 13064 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1606120353
transform 1 0 12328 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__a21o_4  _0793_
timestamp 1606120353
transform 1 0 13248 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__A1_N
timestamp 1606120353
transform 1 0 15272 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__A2_N
timestamp 1606120353
transform 1 0 14904 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A2
timestamp 1606120353
transform 1 0 14536 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_144
timestamp 1606120353
transform 1 0 14352 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_148
timestamp 1606120353
transform 1 0 14720 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_152
timestamp 1606120353
transform 1 0 15088 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _0818_
timestamp 1606120353
transform 1 0 15916 0 1 8160
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__B2
timestamp 1606120353
transform 1 0 15640 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_156
timestamp 1606120353
transform 1 0 15456 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_11_160
timestamp 1606120353
transform 1 0 15824 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_11_175
timestamp 1606120353
transform 1 0 17204 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_187
timestamp 1606120353
transform 1 0 18308 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_179
timestamp 1606120353
transform 1 0 17572 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__CLK
timestamp 1606120353
transform 1 0 17756 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A1
timestamp 1606120353
transform 1 0 17388 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1606120353
transform 1 0 17940 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0662_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 18032 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_11_191
timestamp 1606120353
transform 1 0 18676 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__D
timestamp 1606120353
transform 1 0 18860 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0662__A
timestamp 1606120353
transform 1 0 18492 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_11_195
timestamp 1606120353
transform 1 0 19044 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_207
timestamp 1606120353
transform 1 0 20148 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_219
timestamp 1606120353
transform 1 0 21252 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_231
timestamp 1606120353
transform 1 0 22356 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1606120353
transform 1 0 23552 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_11_243
timestamp 1606120353
transform 1 0 23460 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1606120353
transform 1 0 23644 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1606120353
transform 1 0 24748 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_clk_A
timestamp 1606120353
transform 1 0 25944 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_11_269
timestamp 1606120353
transform 1 0 25852 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_11_272
timestamp 1606120353
transform 1 0 26128 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_284
timestamp 1606120353
transform 1 0 27232 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1606120353
transform 1 0 29164 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_11_296
timestamp 1606120353
transform 1 0 28336 0 1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_11_304
timestamp 1606120353
transform 1 0 29072 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_11_306
timestamp 1606120353
transform 1 0 29256 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_318
timestamp 1606120353
transform 1 0 30360 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_330
timestamp 1606120353
transform 1 0 31464 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_342
timestamp 1606120353
transform 1 0 32568 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1606120353
transform 1 0 34776 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_11_354
timestamp 1606120353
transform 1 0 33672 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_367
timestamp 1606120353
transform 1 0 34868 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_379
timestamp 1606120353
transform 1 0 35972 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_391
timestamp 1606120353
transform 1 0 37076 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606120353
transform -1 0 38548 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_11_403
timestamp 1606120353
transform 1 0 38180 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606120353
transform 1 0 1104 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__CLK
timestamp 1606120353
transform 1 0 1932 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1606120353
transform 1 0 1380 0 -1 9248
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_12_11
timestamp 1606120353
transform 1 0 2116 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1606120353
transform 1 0 3956 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_12_23
timestamp 1606120353
transform 1 0 3220 0 -1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1606120353
transform 1 0 4048 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_12_44
timestamp 1606120353
transform 1 0 5152 0 -1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _0678_
timestamp 1606120353
transform 1 0 6072 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1110_
timestamp 1606120353
transform 1 0 7084 0 -1 9248
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_2  FILLER_12_52
timestamp 1606120353
transform 1 0 5888 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_12_57
timestamp 1606120353
transform 1 0 6348 0 -1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A2
timestamp 1606120353
transform 1 0 9016 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_84
timestamp 1606120353
transform 1 0 8832 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1606120353
transform 1 0 9200 0 -1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _0637_
timestamp 1606120353
transform 1 0 9844 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__a2bb2o_4  _0788_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 10856 0 -1 9248
box 0 -48 1472 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1606120353
transform 1 0 9568 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__A
timestamp 1606120353
transform 1 0 10304 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1606120353
transform 1 0 9660 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_98
timestamp 1606120353
transform 1 0 10120 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_12_102
timestamp 1606120353
transform 1 0 10488 0 -1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _0783_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 13064 0 -1 9248
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__A
timestamp 1606120353
transform 1 0 12604 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_12_122
timestamp 1606120353
transform 1 0 12328 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_12_127
timestamp 1606120353
transform 1 0 12788 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__a2bb2o_4  _0795_
timestamp 1606120353
transform 1 0 15272 0 -1 9248
box 0 -48 1472 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1606120353
transform 1 0 15180 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A1_N
timestamp 1606120353
transform 1 0 13892 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B1
timestamp 1606120353
transform 1 0 14260 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__B
timestamp 1606120353
transform 1 0 14628 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_137
timestamp 1606120353
transform 1 0 13708 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1606120353
transform 1 0 14076 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_145
timestamp 1606120353
transform 1 0 14444 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1606120353
transform 1 0 14812 0 -1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_12_170
timestamp 1606120353
transform 1 0 16744 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1095_
timestamp 1606120353
transform 1 0 18308 0 -1 9248
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_4  FILLER_12_182
timestamp 1606120353
transform 1 0 17848 0 -1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_12_186
timestamp 1606120353
transform 1 0 18216 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1606120353
transform 1 0 20792 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_12_206
timestamp 1606120353
transform 1 0 20056 0 -1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1606120353
transform 1 0 20884 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1606120353
transform 1 0 21988 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1606120353
transform 1 0 23092 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A
timestamp 1606120353
transform 1 0 25392 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__CLK
timestamp 1606120353
transform 1 0 24380 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_251
timestamp 1606120353
transform 1 0 24196 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_12_255
timestamp 1606120353
transform 1 0 24564 0 -1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_12_263
timestamp 1606120353
transform 1 0 25300 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1606120353
transform 1 0 26404 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_clk
timestamp 1606120353
transform 1 0 25944 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_12_266
timestamp 1606120353
transform 1 0 25576 0 -1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_12_273
timestamp 1606120353
transform 1 0 26220 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_12_276
timestamp 1606120353
transform 1 0 26496 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_288
timestamp 1606120353
transform 1 0 27600 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_300
timestamp 1606120353
transform 1 0 28704 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_312
timestamp 1606120353
transform 1 0 29808 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_324
timestamp 1606120353
transform 1 0 30912 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1606120353
transform 1 0 32016 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_12_337
timestamp 1606120353
transform 1 0 32108 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_349
timestamp 1606120353
transform 1 0 33212 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_361
timestamp 1606120353
transform 1 0 34316 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_373
timestamp 1606120353
transform 1 0 35420 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_385
timestamp 1606120353
transform 1 0 36524 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606120353
transform -1 0 38548 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1606120353
transform 1 0 37628 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_12_398
timestamp 1606120353
transform 1 0 37720 0 -1 9248
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1137_
timestamp 1606120353
transform 1 0 1932 0 1 9248
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606120353
transform 1 0 1104 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606120353
transform 1 0 1104 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__D
timestamp 1606120353
transform 1 0 1748 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1606120353
transform 1 0 1380 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1606120353
transform 1 0 1380 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1606120353
transform 1 0 2484 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1606120353
transform 1 0 4048 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1606120353
transform 1 0 3588 0 -1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1606120353
transform 1 0 3956 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_14_44
timestamp 1606120353
transform 1 0 5152 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_14_40
timestamp 1606120353
transform 1 0 4784 0 -1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_14_36
timestamp 1606120353
transform 1 0 4416 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_13_44
timestamp 1606120353
transform 1 0 5152 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_13_40
timestamp 1606120353
transform 1 0 4784 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_clk_A
timestamp 1606120353
transform 1 0 4600 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A2
timestamp 1606120353
transform 1 0 4232 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_13_28
timestamp 1606120353
transform 1 0 3680 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1606120353
transform 1 0 5796 0 1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_13_47
timestamp 1606120353
transform 1 0 5428 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__CLK
timestamp 1606120353
transform 1 0 5612 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__D
timestamp 1606120353
transform 1 0 5244 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_14_64
timestamp 1606120353
transform 1 0 6992 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_13_62
timestamp 1606120353
transform 1 0 6808 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__B2
timestamp 1606120353
transform 1 0 6532 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__B1
timestamp 1606120353
transform 1 0 7084 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1606120353
transform 1 0 6716 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1112_
timestamp 1606120353
transform 1 0 5244 0 -1 10336
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_6  FILLER_14_73
timestamp 1606120353
transform 1 0 7820 0 -1 10336
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_14_69
timestamp 1606120353
transform 1 0 7452 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A2
timestamp 1606120353
transform 1 0 7636 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A1
timestamp 1606120353
transform 1 0 7268 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1606120353
transform 1 0 9200 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_84
timestamp 1606120353
transform 1 0 8832 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1606120353
transform 1 0 8556 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_clk_A
timestamp 1606120353
transform 1 0 8372 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__A
timestamp 1606120353
transform 1 0 8740 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__A1_N
timestamp 1606120353
transform 1 0 9016 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0691_
timestamp 1606120353
transform 1 0 8556 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_13_85
timestamp 1606120353
transform 1 0 8924 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__o22a_4  _0817_
timestamp 1606120353
transform 1 0 7268 0 1 9248
box 0 -48 1288 592
use sky130_fd_sc_hd__inv_8  _0554_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 10948 0 -1 10336
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1606120353
transform 1 0 9568 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0554__A
timestamp 1606120353
transform 1 0 10948 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__B1
timestamp 1606120353
transform 1 0 9384 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_13_97
timestamp 1606120353
transform 1 0 10028 0 1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_13_105
timestamp 1606120353
transform 1 0 10764 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_13_109
timestamp 1606120353
transform 1 0 11132 0 1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1606120353
transform 1 0 9660 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_14_105
timestamp 1606120353
transform 1 0 10764 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_116
timestamp 1606120353
transform 1 0 11776 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_13_119
timestamp 1606120353
transform 1 0 12052 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0503__A
timestamp 1606120353
transform 1 0 11868 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__D
timestamp 1606120353
transform 1 0 11960 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_120
timestamp 1606120353
transform 1 0 12144 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__D
timestamp 1606120353
transform 1 0 12328 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1606120353
transform 1 0 12328 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_14_124
timestamp 1606120353
transform 1 0 12512 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_123
timestamp 1606120353
transform 1 0 12420 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__A
timestamp 1606120353
transform 1 0 12604 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_128
timestamp 1606120353
transform 1 0 12880 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_127
timestamp 1606120353
transform 1 0 12788 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__D
timestamp 1606120353
transform 1 0 12696 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_131
timestamp 1606120353
transform 1 0 13156 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B2
timestamp 1606120353
transform 1 0 12972 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0568__B1
timestamp 1606120353
transform 1 0 13064 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_14_132
timestamp 1606120353
transform 1 0 13248 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_14_140
timestamp 1606120353
transform 1 0 13984 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_135
timestamp 1606120353
transform 1 0 13524 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A2_N
timestamp 1606120353
transform 1 0 14168 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__B
timestamp 1606120353
transform 1 0 13340 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0792_
timestamp 1606120353
transform 1 0 13340 0 -1 10336
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILLER_14_150
timestamp 1606120353
transform 1 0 14904 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_14_144
timestamp 1606120353
transform 1 0 14352 0 -1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_13_153
timestamp 1606120353
transform 1 0 15180 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__A2_N
timestamp 1606120353
transform 1 0 14720 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1606120353
transform 1 0 15180 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0787_
timestamp 1606120353
transform 1 0 15272 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__a2bb2o_4  _0790_
timestamp 1606120353
transform 1 0 13708 0 1 9248
box 0 -48 1472 592
use sky130_fd_sc_hd__fill_2  FILLER_14_157
timestamp 1606120353
transform 1 0 15548 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_13_157
timestamp 1606120353
transform 1 0 15548 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__A
timestamp 1606120353
transform 1 0 15364 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_14_161
timestamp 1606120353
transform 1 0 15916 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__B1
timestamp 1606120353
transform 1 0 15732 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0813_
timestamp 1606120353
transform 1 0 15916 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_14_166
timestamp 1606120353
transform 1 0 16376 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_164
timestamp 1606120353
transform 1 0 16192 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__A
timestamp 1606120353
transform 1 0 16192 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A
timestamp 1606120353
transform 1 0 16376 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_170
timestamp 1606120353
transform 1 0 16744 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_13_168
timestamp 1606120353
transform 1 0 16560 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_clk_A
timestamp 1606120353
transform 1 0 16560 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0806_
timestamp 1606120353
transform 1 0 16928 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0785_
timestamp 1606120353
transform 1 0 16928 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_14_175
timestamp 1606120353
transform 1 0 17204 0 -1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1606120353
transform 1 0 17204 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__A
timestamp 1606120353
transform 1 0 17388 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__A
timestamp 1606120353
transform 1 0 17756 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__B
timestamp 1606120353
transform 1 0 17572 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1606120353
transform 1 0 17572 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_181
timestamp 1606120353
transform 1 0 17756 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0799_
timestamp 1606120353
transform 1 0 17940 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1606120353
transform 1 0 17940 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A
timestamp 1606120353
transform 1 0 18216 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1606120353
transform 1 0 18032 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_14_186
timestamp 1606120353
transform 1 0 18216 0 -1 10336
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1606120353
transform 1 0 19228 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_13_188
timestamp 1606120353
transform 1 0 18400 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__A2
timestamp 1606120353
transform 1 0 18768 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0557__A
timestamp 1606120353
transform 1 0 18768 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0557_
timestamp 1606120353
transform 1 0 18952 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__o22a_4  _0791_
timestamp 1606120353
transform 1 0 18952 0 1 9248
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_8  FILLER_14_205
timestamp 1606120353
transform 1 0 19964 0 -1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_14_201
timestamp 1606120353
transform 1 0 19596 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_208
timestamp 1606120353
transform 1 0 20240 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__B1
timestamp 1606120353
transform 1 0 19780 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__A1
timestamp 1606120353
transform 1 0 19412 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1606120353
transform 1 0 20884 0 -1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1606120353
transform 1 0 20700 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__B2
timestamp 1606120353
transform 1 0 20424 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1606120353
transform 1 0 20792 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_13_212
timestamp 1606120353
transform 1 0 20608 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_14_227
timestamp 1606120353
transform 1 0 21988 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_14_223
timestamp 1606120353
transform 1 0 21620 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_13_226
timestamp 1606120353
transform 1 0 21896 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_clk_A
timestamp 1606120353
transform 1 0 21712 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__D
timestamp 1606120353
transform 1 0 22264 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_clk
timestamp 1606120353
transform 1 0 21712 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_13_240
timestamp 1606120353
transform 1 0 23184 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_13_236
timestamp 1606120353
transform 1 0 22816 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_13_232
timestamp 1606120353
transform 1 0 22448 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__CLK
timestamp 1606120353
transform 1 0 22632 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_clk
timestamp 1606120353
transform 1 0 23276 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1208_
timestamp 1606120353
transform 1 0 22264 0 -1 10336
box 0 -48 1748 592
use sky130_fd_sc_hd__buf_1  _0963_
timestamp 1606120353
transform 1 0 25392 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1118_
timestamp 1606120353
transform 1 0 24380 0 1 9248
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1606120353
transform 1 0 23552 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__D
timestamp 1606120353
transform 1 0 24196 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_clk_A
timestamp 1606120353
transform 1 0 23828 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_245
timestamp 1606120353
transform 1 0 23644 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_249
timestamp 1606120353
transform 1 0 24012 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_14_249
timestamp 1606120353
transform 1 0 24012 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_14_261
timestamp 1606120353
transform 1 0 25116 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_14_267
timestamp 1606120353
transform 1 0 25668 0 -1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__decap_6  FILLER_13_272
timestamp 1606120353
transform 1 0 26128 0 1 9248
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILLER_14_276
timestamp 1606120353
transform 1 0 26496 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_13_278
timestamp 1606120353
transform 1 0 26680 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A
timestamp 1606120353
transform 1 0 26772 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1606120353
transform 1 0 26404 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0954_
timestamp 1606120353
transform 1 0 26772 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_14_286
timestamp 1606120353
transform 1 0 27416 0 -1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_14_282
timestamp 1606120353
transform 1 0 27048 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_13_281
timestamp 1606120353
transform 1 0 26956 0 1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__CLK
timestamp 1606120353
transform 1 0 27232 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0957_
timestamp 1606120353
transform 1 0 27784 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1606120353
transform 1 0 29164 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__A
timestamp 1606120353
transform 1 0 27784 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_13_289
timestamp 1606120353
transform 1 0 27692 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_13_292
timestamp 1606120353
transform 1 0 27968 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_13_304
timestamp 1606120353
transform 1 0 29072 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_13_306
timestamp 1606120353
transform 1 0 29256 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_14_293
timestamp 1606120353
transform 1 0 28060 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_14_305
timestamp 1606120353
transform 1 0 29164 0 -1 10336
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_14_318
timestamp 1606120353
transform 1 0 30360 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_314
timestamp 1606120353
transform 1 0 29992 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_14_311
timestamp 1606120353
transform 1 0 29716 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__C1
timestamp 1606120353
transform 1 0 29808 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__A2
timestamp 1606120353
transform 1 0 30176 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_14_326
timestamp 1606120353
transform 1 0 31096 0 -1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_14_322
timestamp 1606120353
transform 1 0 30728 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__B1
timestamp 1606120353
transform 1 0 30912 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__B1
timestamp 1606120353
transform 1 0 30544 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_13_330
timestamp 1606120353
transform 1 0 31464 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_13_318
timestamp 1606120353
transform 1 0 30360 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1606120353
transform 1 0 32016 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_13_342
timestamp 1606120353
transform 1 0 32568 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_14_334
timestamp 1606120353
transform 1 0 31832 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_14_337
timestamp 1606120353
transform 1 0 32108 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_14_349
timestamp 1606120353
transform 1 0 33212 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1223_
timestamp 1606120353
transform 1 0 35144 0 -1 10336
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1606120353
transform 1 0 34776 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__D
timestamp 1606120353
transform 1 0 35144 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__CLK
timestamp 1606120353
transform 1 0 35512 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_13_354
timestamp 1606120353
transform 1 0 33672 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_13_367
timestamp 1606120353
transform 1 0 34868 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_13_372
timestamp 1606120353
transform 1 0 35328 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_14_361
timestamp 1606120353
transform 1 0 34316 0 -1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_14_369
timestamp 1606120353
transform 1 0 35052 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_13_376
timestamp 1606120353
transform 1 0 35696 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_13_388
timestamp 1606120353
transform 1 0 36800 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_14_389
timestamp 1606120353
transform 1 0 36892 0 -1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606120353
transform -1 0 38548 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606120353
transform -1 0 38548 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1606120353
transform 1 0 37628 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_13_400
timestamp 1606120353
transform 1 0 37904 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_14_398
timestamp 1606120353
transform 1 0 37720 0 -1 10336
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606120353
transform 1 0 1104 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__D
timestamp 1606120353
transform 1 0 1564 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__CLK
timestamp 1606120353
transform 1 0 1932 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1606120353
transform 1 0 1380 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_7
timestamp 1606120353
transform 1 0 1748 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_15_11
timestamp 1606120353
transform 1 0 2116 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_clk
timestamp 1606120353
transform 1 0 4600 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__B1
timestamp 1606120353
transform 1 0 4048 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__B2
timestamp 1606120353
transform 1 0 4416 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A1
timestamp 1606120353
transform 1 0 3680 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_15_23
timestamp 1606120353
transform 1 0 3220 0 1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_15_27
timestamp 1606120353
transform 1 0 3588 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_15_30
timestamp 1606120353
transform 1 0 3864 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_34
timestamp 1606120353
transform 1 0 4232 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_15_41
timestamp 1606120353
transform 1 0 4876 0 1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_15_52
timestamp 1606120353
transform 1 0 5888 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp 1606120353
transform 1 0 5520 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_15_45
timestamp 1606120353
transform 1 0 5244 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A2
timestamp 1606120353
transform 1 0 5336 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__B2
timestamp 1606120353
transform 1 0 5704 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1606120353
transform 1 0 6624 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_15_56
timestamp 1606120353
transform 1 0 6256 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A1
timestamp 1606120353
transform 1 0 6440 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__B1
timestamp 1606120353
transform 1 0 6072 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_15_62
timestamp 1606120353
transform 1 0 6808 0 1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1606120353
transform 1 0 6716 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__a2bb2o_4  _0605_
timestamp 1606120353
transform 1 0 8740 0 1 10336
box 0 -48 1472 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_clk
timestamp 1606120353
transform 1 0 8464 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__B
timestamp 1606120353
transform 1 0 8096 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__A
timestamp 1606120353
transform 1 0 7728 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_70
timestamp 1606120353
transform 1 0 7544 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_74
timestamp 1606120353
transform 1 0 7912 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1606120353
transform 1 0 8280 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__A1_N
timestamp 1606120353
transform 1 0 10856 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__A2_N
timestamp 1606120353
transform 1 0 11224 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__B1
timestamp 1606120353
transform 1 0 10488 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_15_99
timestamp 1606120353
transform 1 0 10212 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_15_104
timestamp 1606120353
transform 1 0 10672 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_108
timestamp 1606120353
transform 1 0 11040 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0560_
timestamp 1606120353
transform 1 0 12880 0 1 10336
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1606120353
transform 1 0 12328 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__B2
timestamp 1606120353
transform 1 0 11592 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0568__A2
timestamp 1606120353
transform 1 0 12696 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__A
timestamp 1606120353
transform 1 0 12144 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_112
timestamp 1606120353
transform 1 0 11408 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_15_116
timestamp 1606120353
transform 1 0 11776 0 1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_15_123
timestamp 1606120353
transform 1 0 12420 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0667_
timestamp 1606120353
transform 1 0 14444 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__A
timestamp 1606120353
transform 1 0 14904 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__B2
timestamp 1606120353
transform 1 0 15272 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0568__A1
timestamp 1606120353
transform 1 0 13892 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__A1_N
timestamp 1606120353
transform 1 0 14260 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_137
timestamp 1606120353
transform 1 0 13708 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_141
timestamp 1606120353
transform 1 0 14076 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_148
timestamp 1606120353
transform 1 0 14720 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_152
timestamp 1606120353
transform 1 0 15088 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0603_
timestamp 1606120353
transform 1 0 16192 0 1 10336
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__A2_N
timestamp 1606120353
transform 1 0 15640 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__A1_N
timestamp 1606120353
transform 1 0 16008 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_156
timestamp 1606120353
transform 1 0 15456 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_160
timestamp 1606120353
transform 1 0 15824 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_15_173
timestamp 1606120353
transform 1 0 17020 0 1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _0661_
timestamp 1606120353
transform 1 0 18308 0 1 10336
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1606120353
transform 1 0 17940 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__A
timestamp 1606120353
transform 1 0 17756 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__A
timestamp 1606120353
transform 1 0 19320 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0614__A
timestamp 1606120353
transform 1 0 17388 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1606120353
transform 1 0 17572 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_15_184
timestamp 1606120353
transform 1 0 18032 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_15_196
timestamp 1606120353
transform 1 0 19136 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0713_
timestamp 1606120353
transform 1 0 19872 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__A
timestamp 1606120353
transform 1 0 20332 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_15_200
timestamp 1606120353
transform 1 0 19504 0 1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_15_207
timestamp 1606120353
transform 1 0 20148 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_15_211
timestamp 1606120353
transform 1 0 20516 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_15_223
timestamp 1606120353
transform 1 0 21620 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_15_235
timestamp 1606120353
transform 1 0 22724 0 1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_15_245
timestamp 1606120353
transform 1 0 23644 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_15_243
timestamp 1606120353
transform 1 0 23460 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1606120353
transform 1 0 23552 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A
timestamp 1606120353
transform 1 0 23828 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_15_249
timestamp 1606120353
transform 1 0 24012 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0962_
timestamp 1606120353
transform 1 0 24104 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_15_253
timestamp 1606120353
transform 1 0 24380 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_257
timestamp 1606120353
transform 1 0 24748 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A
timestamp 1606120353
transform 1 0 24564 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A
timestamp 1606120353
transform 1 0 24932 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0981_
timestamp 1606120353
transform 1 0 25116 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1606120353
transform 1 0 25392 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1210_
timestamp 1606120353
transform 1 0 26680 0 1 10336
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__D
timestamp 1606120353
transform 1 0 26496 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A
timestamp 1606120353
transform 1 0 26128 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A
timestamp 1606120353
transform 1 0 25576 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_15_268
timestamp 1606120353
transform 1 0 25760 0 1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_15_274
timestamp 1606120353
transform 1 0 26312 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1606120353
transform 1 0 29164 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A
timestamp 1606120353
transform 1 0 28612 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_297
timestamp 1606120353
transform 1 0 28428 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_15_301
timestamp 1606120353
transform 1 0 28796 0 1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_15_306
timestamp 1606120353
transform 1 0 29256 0 1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__a211o_4  _0961_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 30176 0 1 10336
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__A1
timestamp 1606120353
transform 1 0 29992 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A1
timestamp 1606120353
transform 1 0 29624 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_312
timestamp 1606120353
transform 1 0 29808 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_330
timestamp 1606120353
transform 1 0 31464 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__C1
timestamp 1606120353
transform 1 0 31648 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_15_334
timestamp 1606120353
transform 1 0 31832 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_15_346
timestamp 1606120353
transform 1 0 32936 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1606120353
transform 1 0 34776 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_15_358
timestamp 1606120353
transform 1 0 34040 0 1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_15_367
timestamp 1606120353
transform 1 0 34868 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_15_379
timestamp 1606120353
transform 1 0 35972 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_15_391
timestamp 1606120353
transform 1 0 37076 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606120353
transform -1 0 38548 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_15_403
timestamp 1606120353
transform 1 0 38180 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1140_
timestamp 1606120353
transform 1 0 1380 0 -1 11424
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606120353
transform 1 0 1104 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_16_22
timestamp 1606120353
transform 1 0 3128 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__o22a_4  _0814_
timestamp 1606120353
transform 1 0 4048 0 -1 11424
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1606120353
transform 1 0 3956 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__CLK
timestamp 1606120353
transform 1 0 3404 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1606120353
transform 1 0 3588 0 -1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__o22a_4  _0819_
timestamp 1606120353
transform 1 0 6072 0 -1 11424
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_clk_A
timestamp 1606120353
transform 1 0 5888 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_clk_A
timestamp 1606120353
transform 1 0 5520 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_46
timestamp 1606120353
transform 1 0 5336 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_50
timestamp 1606120353
transform 1 0 5704 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0692_
timestamp 1606120353
transform 1 0 8096 0 -1 11424
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__A2_N
timestamp 1606120353
transform 1 0 8924 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__A
timestamp 1606120353
transform 1 0 7912 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__D
timestamp 1606120353
transform 1 0 7544 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_68
timestamp 1606120353
transform 1 0 7360 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_72
timestamp 1606120353
transform 1 0 7728 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_83
timestamp 1606120353
transform 1 0 8740 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_87
timestamp 1606120353
transform 1 0 9108 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_97
timestamp 1606120353
transform 1 0 10028 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1606120353
transform 1 0 9660 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1606120353
transform 1 0 9476 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__D
timestamp 1606120353
transform 1 0 10212 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__D
timestamp 1606120353
transform 1 0 9844 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__B2
timestamp 1606120353
transform 1 0 9292 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1606120353
transform 1 0 9568 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_16_101
timestamp 1606120353
transform 1 0 10396 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__D
timestamp 1606120353
transform 1 0 10672 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__a2bb2o_4  _0559_
timestamp 1606120353
transform 1 0 10856 0 -1 11424
box 0 -48 1472 592
use sky130_fd_sc_hd__o21ai_4  _0568_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 13064 0 -1 11424
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__B
timestamp 1606120353
transform 1 0 12512 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__C
timestamp 1606120353
transform 1 0 12880 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_122
timestamp 1606120353
transform 1 0 12328 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_126
timestamp 1606120353
transform 1 0 12696 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__a2bb2o_4  _0615_
timestamp 1606120353
transform 1 0 15272 0 -1 11424
box 0 -48 1472 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1606120353
transform 1 0 15180 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__B1
timestamp 1606120353
transform 1 0 14720 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_16_143
timestamp 1606120353
transform 1 0 14260 0 -1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_16_147
timestamp 1606120353
transform 1 0 14628 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1606120353
transform 1 0 14904 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__B2
timestamp 1606120353
transform 1 0 16928 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__A1
timestamp 1606120353
transform 1 0 17296 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1606120353
transform 1 0 16744 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1606120353
transform 1 0 17112 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0562_
timestamp 1606120353
transform 1 0 19044 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _0614_
timestamp 1606120353
transform 1 0 17480 0 -1 11424
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__A
timestamp 1606120353
transform 1 0 18492 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__D
timestamp 1606120353
transform 1 0 18860 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_187
timestamp 1606120353
transform 1 0 18308 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_191
timestamp 1606120353
transform 1 0 18676 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_198
timestamp 1606120353
transform 1 0 19320 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1606120353
transform 1 0 20792 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__C
timestamp 1606120353
transform 1 0 19504 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__C
timestamp 1606120353
transform 1 0 19872 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0516__A
timestamp 1606120353
transform 1 0 20240 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0504__A
timestamp 1606120353
transform 1 0 20608 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_202
timestamp 1606120353
transform 1 0 19688 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_206
timestamp 1606120353
transform 1 0 20056 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_210
timestamp 1606120353
transform 1 0 20424 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_16_215
timestamp 1606120353
transform 1 0 20884 0 -1 11424
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A2
timestamp 1606120353
transform 1 0 21620 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__B1
timestamp 1606120353
transform 1 0 21988 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_225
timestamp 1606120353
transform 1 0 21804 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_16_229
timestamp 1606120353
transform 1 0 22172 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_16_241
timestamp 1606120353
transform 1 0 23276 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0947_
timestamp 1606120353
transform 1 0 24472 0 -1 11424
box 0 -48 828 592
use sky130_fd_sc_hd__buf_1  _0956_
timestamp 1606120353
transform 1 0 23460 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__A
timestamp 1606120353
transform 1 0 23920 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_246
timestamp 1606120353
transform 1 0 23736 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_16_250
timestamp 1606120353
transform 1 0 24104 0 -1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_16_263
timestamp 1606120353
transform 1 0 25300 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_16_267
timestamp 1606120353
transform 1 0 25668 0 -1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__D
timestamp 1606120353
transform 1 0 25484 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__D
timestamp 1606120353
transform 1 0 26036 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1606120353
transform 1 0 26496 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_16_273
timestamp 1606120353
transform 1 0 26220 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1606120353
transform 1 0 26404 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_16_280
timestamp 1606120353
transform 1 0 26864 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0951_
timestamp 1606120353
transform 1 0 26588 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_16_284
timestamp 1606120353
transform 1 0 27232 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__B
timestamp 1606120353
transform 1 0 27048 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__D
timestamp 1606120353
transform 1 0 27416 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0945_
timestamp 1606120353
transform 1 0 28428 0 -1 11424
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILLER_16_288
timestamp 1606120353
transform 1 0 27600 0 -1 11424
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_16_296
timestamp 1606120353
transform 1 0 28336 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_16_306
timestamp 1606120353
transform 1 0 29256 0 -1 11424
box 0 -48 552 592
use sky130_fd_sc_hd__a211o_4  _0967_
timestamp 1606120353
transform 1 0 29992 0 -1 11424
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A2
timestamp 1606120353
transform 1 0 29808 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_16_328
timestamp 1606120353
transform 1 0 31280 0 -1 11424
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1606120353
transform 1 0 32016 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_16_337
timestamp 1606120353
transform 1 0 32108 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_16_349
timestamp 1606120353
transform 1 0 33212 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_16_361
timestamp 1606120353
transform 1 0 34316 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_16_373
timestamp 1606120353
transform 1 0 35420 0 -1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__CLK
timestamp 1606120353
transform 1 0 35788 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_16_379
timestamp 1606120353
transform 1 0 35972 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_16_391
timestamp 1606120353
transform 1 0 37076 0 -1 11424
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606120353
transform -1 0 38548 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1606120353
transform 1 0 37628 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_16_398
timestamp 1606120353
transform 1 0 37720 0 -1 11424
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606120353
transform 1 0 1104 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__D
timestamp 1606120353
transform 1 0 1564 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__CLK
timestamp 1606120353
transform 1 0 1932 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1606120353
transform 1 0 1380 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1606120353
transform 1 0 1748 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_17_11
timestamp 1606120353
transform 1 0 2116 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1108_
timestamp 1606120353
transform 1 0 3404 0 1 11424
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__D
timestamp 1606120353
transform 1 0 3220 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_17_44
timestamp 1606120353
transform 1 0 5152 0 1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _0627_
timestamp 1606120353
transform 1 0 6808 0 1 11424
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1606120353
transform 1 0 6716 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_clk
timestamp 1606120353
transform 1 0 6440 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0627__A
timestamp 1606120353
transform 1 0 6256 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A2
timestamp 1606120353
transform 1 0 5888 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A1
timestamp 1606120353
transform 1 0 5520 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_50
timestamp 1606120353
transform 1 0 5704 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1606120353
transform 1 0 6072 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0639_
timestamp 1606120353
transform 1 0 8648 0 1 11424
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0640__A
timestamp 1606120353
transform 1 0 8188 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__B
timestamp 1606120353
transform 1 0 7820 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_71
timestamp 1606120353
transform 1 0 7636 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_75
timestamp 1606120353
transform 1 0 8004 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_17_79
timestamp 1606120353
transform 1 0 8372 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _0604_
timestamp 1606120353
transform 1 0 10028 0 1 11424
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__A
timestamp 1606120353
transform 1 0 9844 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__B
timestamp 1606120353
transform 1 0 11040 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0600__A
timestamp 1606120353
transform 1 0 9476 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_89
timestamp 1606120353
transform 1 0 9292 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_93
timestamp 1606120353
transform 1 0 9660 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_106
timestamp 1606120353
transform 1 0 10856 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1606120353
transform 1 0 11224 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__nor4_4  _0578_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 12420 0 1 11424
box 0 -48 1564 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1606120353
transform 1 0 12328 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__A
timestamp 1606120353
transform 1 0 12144 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0598__A
timestamp 1606120353
transform 1 0 11776 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__A
timestamp 1606120353
transform 1 0 11408 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1606120353
transform 1 0 11592 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1606120353
transform 1 0 11960 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__a2bb2o_4  _0577_
timestamp 1606120353
transform 1 0 14720 0 1 11424
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0518__A
timestamp 1606120353
transform 1 0 14536 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__A
timestamp 1606120353
transform 1 0 14168 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_140
timestamp 1606120353
transform 1 0 13984 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_144
timestamp 1606120353
transform 1 0 14352 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0517_
timestamp 1606120353
transform 1 0 16928 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__A2
timestamp 1606120353
transform 1 0 16652 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1606120353
transform 1 0 16192 0 1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_17_168
timestamp 1606120353
transform 1 0 16560 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_17_171
timestamp 1606120353
transform 1 0 16836 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1606120353
transform 1 0 17204 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0575_
timestamp 1606120353
transform 1 0 18032 0 1 11424
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1606120353
transform 1 0 17940 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0517__A
timestamp 1606120353
transform 1 0 17388 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0572__A
timestamp 1606120353
transform 1 0 19044 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__B1
timestamp 1606120353
transform 1 0 17756 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1606120353
transform 1 0 17572 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1606120353
transform 1 0 18860 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_197
timestamp 1606120353
transform 1 0 19228 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0516_
timestamp 1606120353
transform 1 0 19872 0 1 11424
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0571__A
timestamp 1606120353
transform 1 0 20884 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__D
timestamp 1606120353
transform 1 0 19412 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_17_201
timestamp 1606120353
transform 1 0 19596 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_17_213
timestamp 1606120353
transform 1 0 20700 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_17_217
timestamp 1606120353
transform 1 0 21068 0 1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__o21ai_4  _1038_
timestamp 1606120353
transform 1 0 21620 0 1 11424
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A1
timestamp 1606120353
transform 1 0 21436 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A
timestamp 1606120353
transform 1 0 23000 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A
timestamp 1606120353
transform 1 0 23368 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1606120353
transform 1 0 22816 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1606120353
transform 1 0 23184 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _1003_
timestamp 1606120353
transform 1 0 23736 0 1 11424
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1606120353
transform 1 0 23552 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__B
timestamp 1606120353
transform 1 0 24840 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A
timestamp 1606120353
transform 1 0 25208 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_17_245
timestamp 1606120353
transform 1 0 23644 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_17_255
timestamp 1606120353
transform 1 0 24564 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_17_260
timestamp 1606120353
transform 1 0 25024 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1606120353
transform 1 0 25392 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0953_
timestamp 1606120353
transform 1 0 26220 0 1 11424
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A
timestamp 1606120353
transform 1 0 27232 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__A
timestamp 1606120353
transform 1 0 26036 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__C
timestamp 1606120353
transform 1 0 25576 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_17_268
timestamp 1606120353
transform 1 0 25760 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_17_282
timestamp 1606120353
transform 1 0 27048 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_286
timestamp 1606120353
transform 1 0 27416 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1008_
timestamp 1606120353
transform 1 0 27784 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1606120353
transform 1 0 29164 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A
timestamp 1606120353
transform 1 0 28612 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1606120353
transform 1 0 28244 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__C
timestamp 1606120353
transform 1 0 27600 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_293
timestamp 1606120353
transform 1 0 28060 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_297
timestamp 1606120353
transform 1 0 28428 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_17_301
timestamp 1606120353
transform 1 0 28796 0 1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_17_306
timestamp 1606120353
transform 1 0 29256 0 1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _0942_
timestamp 1606120353
transform 1 0 30084 0 1 11424
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__A
timestamp 1606120353
transform 1 0 29624 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__B
timestamp 1606120353
transform 1 0 31464 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A
timestamp 1606120353
transform 1 0 31096 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_17_312
timestamp 1606120353
transform 1 0 29808 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_17_324
timestamp 1606120353
transform 1 0 30912 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_328
timestamp 1606120353
transform 1 0 31280 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0946_
timestamp 1606120353
transform 1 0 31648 0 1 11424
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A
timestamp 1606120353
transform 1 0 32476 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A
timestamp 1606120353
transform 1 0 32844 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_339
timestamp 1606120353
transform 1 0 32292 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_343
timestamp 1606120353
transform 1 0 32660 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_17_347
timestamp 1606120353
transform 1 0 33028 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1606120353
transform 1 0 34776 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_17_359
timestamp 1606120353
transform 1 0 34132 0 1 11424
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_17_365
timestamp 1606120353
transform 1 0 34684 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_17_367
timestamp 1606120353
transform 1 0 34868 0 1 11424
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1160_
timestamp 1606120353
transform 1 0 35788 0 1 11424
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__D
timestamp 1606120353
transform 1 0 35604 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_17_396
timestamp 1606120353
transform 1 0 37536 0 1 11424
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606120353
transform -1 0 38548 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1219_
timestamp 1606120353
transform 1 0 1472 0 -1 12512
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606120353
transform 1 0 1104 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1606120353
transform 1 0 1380 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0670_
timestamp 1606120353
transform 1 0 4140 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1606120353
transform 1 0 3956 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__A
timestamp 1606120353
transform 1 0 4600 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__D
timestamp 1606120353
transform 1 0 5152 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_18_23
timestamp 1606120353
transform 1 0 3220 0 -1 12512
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_18_32
timestamp 1606120353
transform 1 0 4048 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_18_36
timestamp 1606120353
transform 1 0 4416 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_18_40
timestamp 1606120353
transform 1 0 4784 0 -1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__a21o_4  _0693_
timestamp 1606120353
transform 1 0 6348 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_clk
timestamp 1606120353
transform 1 0 5704 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__B1
timestamp 1606120353
transform 1 0 6164 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__D
timestamp 1606120353
transform 1 0 5520 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_46
timestamp 1606120353
transform 1 0 5336 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_53
timestamp 1606120353
transform 1 0 5980 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_69
timestamp 1606120353
transform 1 0 7452 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__C
timestamp 1606120353
transform 1 0 7636 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_73
timestamp 1606120353
transform 1 0 7820 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__A
timestamp 1606120353
transform 1 0 8004 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0640_
timestamp 1606120353
transform 1 0 8188 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_18_80
timestamp 1606120353
transform 1 0 8464 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_84
timestamp 1606120353
transform 1 0 8832 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__A
timestamp 1606120353
transform 1 0 8648 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__B
timestamp 1606120353
transform 1 0 9016 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_88
timestamp 1606120353
transform 1 0 9200 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0600_
timestamp 1606120353
transform 1 0 9660 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__and2_4  _0638_
timestamp 1606120353
transform 1 0 10672 0 -1 12512
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1606120353
transform 1 0 9568 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__C
timestamp 1606120353
transform 1 0 9384 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__A
timestamp 1606120353
transform 1 0 10488 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__B
timestamp 1606120353
transform 1 0 10120 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_96
timestamp 1606120353
transform 1 0 9936 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_100
timestamp 1606120353
transform 1 0 10304 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_111
timestamp 1606120353
transform 1 0 11316 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__C
timestamp 1606120353
transform 1 0 11500 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_115
timestamp 1606120353
transform 1 0 11684 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__B
timestamp 1606120353
transform 1 0 11868 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0598_
timestamp 1606120353
transform 1 0 12052 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_18_122
timestamp 1606120353
transform 1 0 12328 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__C
timestamp 1606120353
transform 1 0 12512 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_126
timestamp 1606120353
transform 1 0 12696 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__D
timestamp 1606120353
transform 1 0 12880 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_130
timestamp 1606120353
transform 1 0 13064 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__D
timestamp 1606120353
transform 1 0 13248 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_134
timestamp 1606120353
transform 1 0 13432 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1606120353
transform 1 0 13800 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__A
timestamp 1606120353
transform 1 0 13616 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__B
timestamp 1606120353
transform 1 0 13984 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0593_
timestamp 1606120353
transform 1 0 14168 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_18_145
timestamp 1606120353
transform 1 0 14444 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_18_150
timestamp 1606120353
transform 1 0 14904 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__B2
timestamp 1606120353
transform 1 0 14720 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1606120353
transform 1 0 15180 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0518_
timestamp 1606120353
transform 1 0 15272 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__o22a_4  _0625_
timestamp 1606120353
transform 1 0 16652 0 -1 12512
box 0 -48 1288 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk
timestamp 1606120353
transform 1 0 16376 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__A
timestamp 1606120353
transform 1 0 15916 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_18_157
timestamp 1606120353
transform 1 0 15548 0 -1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_18_163
timestamp 1606120353
transform 1 0 16100 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _0572_
timestamp 1606120353
transform 1 0 18676 0 -1 12512
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__B
timestamp 1606120353
transform 1 0 18124 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__C
timestamp 1606120353
transform 1 0 18492 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_183
timestamp 1606120353
transform 1 0 17940 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_187
timestamp 1606120353
transform 1 0 18308 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0571_
timestamp 1606120353
transform 1 0 20884 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1606120353
transform 1 0 20792 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__D
timestamp 1606120353
transform 1 0 19688 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0570__B
timestamp 1606120353
transform 1 0 20240 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0522__A
timestamp 1606120353
transform 1 0 20608 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_200
timestamp 1606120353
transform 1 0 19504 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_18_204
timestamp 1606120353
transform 1 0 19872 0 -1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_18_210
timestamp 1606120353
transform 1 0 20424 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_18_218
timestamp 1606120353
transform 1 0 21160 0 -1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_18_222
timestamp 1606120353
transform 1 0 21528 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__B1
timestamp 1606120353
transform 1 0 21620 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_225
timestamp 1606120353
transform 1 0 21804 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A2
timestamp 1606120353
transform 1 0 21988 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_229
timestamp 1606120353
transform 1 0 22172 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0948_
timestamp 1606120353
transform 1 0 22356 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_18_234
timestamp 1606120353
transform 1 0 22632 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__A
timestamp 1606120353
transform 1 0 22816 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_18_238
timestamp 1606120353
transform 1 0 23000 0 -1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _1035_
timestamp 1606120353
transform 1 0 23368 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__or4_4  _0940_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 24840 0 -1 12512
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__A
timestamp 1606120353
transform 1 0 23828 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__B
timestamp 1606120353
transform 1 0 24196 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__C
timestamp 1606120353
transform 1 0 24564 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_245
timestamp 1606120353
transform 1 0 23644 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_249
timestamp 1606120353
transform 1 0 24012 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1606120353
transform 1 0 24380 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_18_257
timestamp 1606120353
transform 1 0 24748 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__or4_4  _0994_
timestamp 1606120353
transform 1 0 27048 0 -1 12512
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1606120353
transform 1 0 26404 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__B
timestamp 1606120353
transform 1 0 26036 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__C
timestamp 1606120353
transform 1 0 26680 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_18_267
timestamp 1606120353
transform 1 0 25668 0 -1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_18_273
timestamp 1606120353
transform 1 0 26220 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_276
timestamp 1606120353
transform 1 0 26496 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_280
timestamp 1606120353
transform 1 0 26864 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0949_
timestamp 1606120353
transform 1 0 28612 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__B
timestamp 1606120353
transform 1 0 28152 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A
timestamp 1606120353
transform 1 0 29348 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_18_291
timestamp 1606120353
transform 1 0 27876 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_18_296
timestamp 1606120353
transform 1 0 28336 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_18_302
timestamp 1606120353
transform 1 0 28888 0 -1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_18_306
timestamp 1606120353
transform 1 0 29256 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_18_309
timestamp 1606120353
transform 1 0 29532 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0941_
timestamp 1606120353
transform 1 0 29624 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_18_313
timestamp 1606120353
transform 1 0 29900 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_317
timestamp 1606120353
transform 1 0 30268 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A
timestamp 1606120353
transform 1 0 30084 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__C
timestamp 1606120353
transform 1 0 30452 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_321
timestamp 1606120353
transform 1 0 30636 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__B
timestamp 1606120353
transform 1 0 30820 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0965_
timestamp 1606120353
transform 1 0 31004 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_18_328
timestamp 1606120353
transform 1 0 31280 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A2
timestamp 1606120353
transform 1 0 31464 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0966_
timestamp 1606120353
transform 1 0 32108 0 -1 12512
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1606120353
transform 1 0 32016 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_18_332
timestamp 1606120353
transform 1 0 31648 0 -1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_18_346
timestamp 1606120353
transform 1 0 32936 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_18_358
timestamp 1606120353
transform 1 0 34040 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_18_370
timestamp 1606120353
transform 1 0 35144 0 -1 12512
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__CLK
timestamp 1606120353
transform 1 0 35788 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_18_376
timestamp 1606120353
transform 1 0 35696 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_18_379
timestamp 1606120353
transform 1 0 35972 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_18_391
timestamp 1606120353
transform 1 0 37076 0 -1 12512
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606120353
transform -1 0 38548 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1606120353
transform 1 0 37628 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_18_398
timestamp 1606120353
transform 1 0 37720 0 -1 12512
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1129_
timestamp 1606120353
transform 1 0 1380 0 -1 13600
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606120353
transform 1 0 1104 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606120353
transform 1 0 1104 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__D
timestamp 1606120353
transform 1 0 1564 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__CLK
timestamp 1606120353
transform 1 0 1932 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1606120353
transform 1 0 1380 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 1606120353
transform 1 0 1748 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_19_11
timestamp 1606120353
transform 1 0 2116 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_20_22
timestamp 1606120353
transform 1 0 3128 0 -1 13600
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1606120353
transform 1 0 4048 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1606120353
transform 1 0 3864 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1606120353
transform 1 0 3956 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_20_42
timestamp 1606120353
transform 1 0 4968 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_20_36
timestamp 1606120353
transform 1 0 4416 0 -1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_19_44
timestamp 1606120353
transform 1 0 5152 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_19_41
timestamp 1606120353
transform 1 0 4876 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_19_35
timestamp 1606120353
transform 1 0 4324 0 1 12512
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__D
timestamp 1606120353
transform 1 0 4784 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0543__A
timestamp 1606120353
transform 1 0 4232 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__D
timestamp 1606120353
transform 1 0 5152 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__C
timestamp 1606120353
transform 1 0 4968 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_19_23
timestamp 1606120353
transform 1 0 3220 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_19_52
timestamp 1606120353
transform 1 0 5888 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_19_48
timestamp 1606120353
transform 1 0 5520 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__B
timestamp 1606120353
transform 1 0 5704 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__B
timestamp 1606120353
transform 1 0 6164 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__A
timestamp 1606120353
transform 1 0 5336 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_20_65
timestamp 1606120353
transform 1 0 7084 0 -1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_20_59
timestamp 1606120353
transform 1 0 6532 0 -1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_19_62
timestamp 1606120353
transform 1 0 6808 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1606120353
transform 1 0 6348 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__C
timestamp 1606120353
transform 1 0 6900 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__A
timestamp 1606120353
transform 1 0 6532 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1606120353
transform 1 0 6716 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0599_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 6900 0 1 12512
box 0 -48 828 592
use sky130_fd_sc_hd__nor3_4  _0626_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 5336 0 -1 13600
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_20_71
timestamp 1606120353
transform 1 0 7636 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_19_77
timestamp 1606120353
transform 1 0 8188 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_19_72
timestamp 1606120353
transform 1 0 7728 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__B
timestamp 1606120353
transform 1 0 7452 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__C
timestamp 1606120353
transform 1 0 7820 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__B
timestamp 1606120353
transform 1 0 8004 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0602_
timestamp 1606120353
transform 1 0 8004 0 -1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_20_88
timestamp 1606120353
transform 1 0 9200 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1606120353
transform 1 0 8832 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__B
timestamp 1606120353
transform 1 0 9016 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__nor4_4  _0612_
timestamp 1606120353
transform 1 0 8464 0 1 12512
box 0 -48 1564 592
use sky130_fd_sc_hd__fill_2  FILLER_20_96
timestamp 1606120353
transform 1 0 9936 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_97
timestamp 1606120353
transform 1 0 10028 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__D
timestamp 1606120353
transform 1 0 9384 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1606120353
transform 1 0 9568 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0519_
timestamp 1606120353
transform 1 0 9660 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_20_104
timestamp 1606120353
transform 1 0 10672 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_100
timestamp 1606120353
transform 1 0 10304 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1606120353
transform 1 0 10396 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__A
timestamp 1606120353
transform 1 0 10580 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__A
timestamp 1606120353
transform 1 0 10488 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__B
timestamp 1606120353
transform 1 0 10120 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0519__A
timestamp 1606120353
transform 1 0 10212 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0647_
timestamp 1606120353
transform 1 0 10764 0 1 12512
box 0 -48 828 592
use sky130_fd_sc_hd__and4_4  _0641_
timestamp 1606120353
transform 1 0 10856 0 -1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_20_119
timestamp 1606120353
transform 1 0 12052 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_115
timestamp 1606120353
transform 1 0 11684 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1606120353
transform 1 0 11960 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1606120353
transform 1 0 11592 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__D
timestamp 1606120353
transform 1 0 12236 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__C
timestamp 1606120353
transform 1 0 11868 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__A
timestamp 1606120353
transform 1 0 11776 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__B
timestamp 1606120353
transform 1 0 12144 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_19_130
timestamp 1606120353
transform 1 0 13064 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_19_126
timestamp 1606120353
transform 1 0 12696 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__A
timestamp 1606120353
transform 1 0 12880 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1606120353
transform 1 0 12328 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0601_
timestamp 1606120353
transform 1 0 12420 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__nor3_4  _0574_
timestamp 1606120353
transform 1 0 12420 0 -1 13600
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_3  FILLER_20_140
timestamp 1606120353
transform 1 0 13984 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_20_136
timestamp 1606120353
transform 1 0 13616 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__B
timestamp 1606120353
transform 1 0 14260 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__A
timestamp 1606120353
transform 1 0 13800 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__C
timestamp 1606120353
transform 1 0 13432 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_149
timestamp 1606120353
transform 1 0 14812 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_145
timestamp 1606120353
transform 1 0 14444 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_153
timestamp 1606120353
transform 1 0 15180 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__A
timestamp 1606120353
transform 1 0 14628 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__B
timestamp 1606120353
transform 1 0 14996 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1606120353
transform 1 0 15180 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0563_
timestamp 1606120353
transform 1 0 15272 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__nand4_4  _0567_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 13616 0 1 12512
box 0 -48 1564 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1606120353
transform 1 0 16100 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_20_157
timestamp 1606120353
transform 1 0 15548 0 -1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_19_157
timestamp 1606120353
transform 1 0 15548 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__C
timestamp 1606120353
transform 1 0 15916 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0563__A
timestamp 1606120353
transform 1 0 15364 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__D
timestamp 1606120353
transform 1 0 15732 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0576_
timestamp 1606120353
transform 1 0 15916 0 1 12512
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_19_170
timestamp 1606120353
transform 1 0 16744 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__A
timestamp 1606120353
transform 1 0 16928 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0643_
timestamp 1606120353
transform 1 0 16284 0 -1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_20_174
timestamp 1606120353
transform 1 0 17112 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_174
timestamp 1606120353
transform 1 0 17112 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__B
timestamp 1606120353
transform 1 0 17296 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__C
timestamp 1606120353
transform 1 0 17296 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_178
timestamp 1606120353
transform 1 0 17480 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_19_184
timestamp 1606120353
transform 1 0 18032 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_19_178
timestamp 1606120353
transform 1 0 17480 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__C
timestamp 1606120353
transform 1 0 17664 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__A
timestamp 1606120353
transform 1 0 17756 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1606120353
transform 1 0 17940 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0642_
timestamp 1606120353
transform 1 0 17848 0 -1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILLER_20_191
timestamp 1606120353
transform 1 0 18676 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_19_188
timestamp 1606120353
transform 1 0 18400 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__A
timestamp 1606120353
transform 1 0 18952 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__A
timestamp 1606120353
transform 1 0 18492 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0561_
timestamp 1606120353
transform 1 0 18676 0 1 12512
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILLER_20_196
timestamp 1606120353
transform 1 0 19136 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_20_206
timestamp 1606120353
transform 1 0 20056 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_202
timestamp 1606120353
transform 1 0 19688 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_204
timestamp 1606120353
transform 1 0 19872 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_200
timestamp 1606120353
transform 1 0 19504 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__C
timestamp 1606120353
transform 1 0 19872 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__B
timestamp 1606120353
transform 1 0 20056 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__A
timestamp 1606120353
transform 1 0 19688 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0564_
timestamp 1606120353
transform 1 0 19412 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1606120353
transform 1 0 20424 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_215
timestamp 1606120353
transform 1 0 20884 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__D
timestamp 1606120353
transform 1 0 20608 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__D
timestamp 1606120353
transform 1 0 20240 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1606120353
transform 1 0 20792 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _0570_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 20240 0 1 12512
box 0 -48 644 592
use sky130_fd_sc_hd__inv_8  _0522_
timestamp 1606120353
transform 1 0 20884 0 -1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_19_219
timestamp 1606120353
transform 1 0 21252 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0570__A
timestamp 1606120353
transform 1 0 21068 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_228
timestamp 1606120353
transform 1 0 22080 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_224
timestamp 1606120353
transform 1 0 21712 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__B1
timestamp 1606120353
transform 1 0 22264 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A
timestamp 1606120353
transform 1 0 21896 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A1
timestamp 1606120353
transform 1 0 21436 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_241
timestamp 1606120353
transform 1 0 23276 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_237
timestamp 1606120353
transform 1 0 22908 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_232
timestamp 1606120353
transform 1 0 22448 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_240
timestamp 1606120353
transform 1 0 23184 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_236
timestamp 1606120353
transform 1 0 22816 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__D
timestamp 1606120353
transform 1 0 23092 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__B
timestamp 1606120353
transform 1 0 23000 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__A
timestamp 1606120353
transform 1 0 23368 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1040_
timestamp 1606120353
transform 1 0 22632 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _1041_
timestamp 1606120353
transform 1 0 21620 0 1 12512
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_19_245
timestamp 1606120353
transform 1 0 23644 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__D
timestamp 1606120353
transform 1 0 23460 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1606120353
transform 1 0 23552 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__or4_4  _1039_
timestamp 1606120353
transform 1 0 23644 0 -1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__or4_4  _1034_
timestamp 1606120353
transform 1 0 23828 0 1 12512
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_20_258
timestamp 1606120353
transform 1 0 24840 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_254
timestamp 1606120353
transform 1 0 24472 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_260
timestamp 1606120353
transform 1 0 25024 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_256
timestamp 1606120353
transform 1 0 24656 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A
timestamp 1606120353
transform 1 0 25024 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__D
timestamp 1606120353
transform 1 0 24656 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__C
timestamp 1606120353
transform 1 0 24840 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_19_264
timestamp 1606120353
transform 1 0 25392 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__A
timestamp 1606120353
transform 1 0 25208 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0969_
timestamp 1606120353
transform 1 0 25208 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_20_272
timestamp 1606120353
transform 1 0 26128 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_20_269
timestamp 1606120353
transform 1 0 25852 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_20_265
timestamp 1606120353
transform 1 0 25484 0 -1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_19_268
timestamp 1606120353
transform 1 0 25760 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__A
timestamp 1606120353
transform 1 0 25944 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__A
timestamp 1606120353
transform 1 0 25852 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0964_
timestamp 1606120353
transform 1 0 26036 0 1 12512
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_20_279
timestamp 1606120353
transform 1 0 26772 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_280
timestamp 1606120353
transform 1 0 26864 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A
timestamp 1606120353
transform 1 0 26956 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__B
timestamp 1606120353
transform 1 0 27048 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1606120353
transform 1 0 26404 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0972_
timestamp 1606120353
transform 1 0 26496 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_20_283
timestamp 1606120353
transform 1 0 27140 0 -1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_19_284
timestamp 1606120353
transform 1 0 27232 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__D
timestamp 1606120353
transform 1 0 27416 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_290
timestamp 1606120353
transform 1 0 27784 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_20_287
timestamp 1606120353
transform 1 0 27508 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__A
timestamp 1606120353
transform 1 0 27968 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__C
timestamp 1606120353
transform 1 0 27600 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _1027_
timestamp 1606120353
transform 1 0 27600 0 1 12512
box 0 -48 828 592
use sky130_fd_sc_hd__and3_4  _1010_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 28152 0 -1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILLER_20_303
timestamp 1606120353
transform 1 0 28980 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_19_301
timestamp 1606120353
transform 1 0 28796 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_297
timestamp 1606120353
transform 1 0 28428 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A
timestamp 1606120353
transform 1 0 28980 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__C
timestamp 1606120353
transform 1 0 28612 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_20_308
timestamp 1606120353
transform 1 0 29440 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_19_306
timestamp 1606120353
transform 1 0 29256 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A
timestamp 1606120353
transform 1 0 29256 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1606120353
transform 1 0 29164 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _1028_
timestamp 1606120353
transform 1 0 29348 0 1 12512
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_19_318
timestamp 1606120353
transform 1 0 30360 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_314
timestamp 1606120353
transform 1 0 29992 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__A
timestamp 1606120353
transform 1 0 30176 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__or3_4  _0960_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 29716 0 -1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_20_328
timestamp 1606120353
transform 1 0 31280 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_324
timestamp 1606120353
transform 1 0 30912 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_320
timestamp 1606120353
transform 1 0 30544 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_322
timestamp 1606120353
transform 1 0 30728 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__B
timestamp 1606120353
transform 1 0 30728 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A1
timestamp 1606120353
transform 1 0 31464 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__B1
timestamp 1606120353
transform 1 0 31096 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__B
timestamp 1606120353
transform 1 0 30544 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A1
timestamp 1606120353
transform 1 0 30912 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__a21oi_4  _0975_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 31096 0 1 12512
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_20_332
timestamp 1606120353
transform 1 0 31648 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_339
timestamp 1606120353
transform 1 0 32292 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__C
timestamp 1606120353
transform 1 0 31832 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__A
timestamp 1606120353
transform 1 0 32476 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1606120353
transform 1 0 32016 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__nor2_4  _1036_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 32108 0 -1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_20_350
timestamp 1606120353
transform 1 0 33304 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_346
timestamp 1606120353
transform 1 0 32936 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_343
timestamp 1606120353
transform 1 0 32660 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__B
timestamp 1606120353
transform 1 0 32844 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__B1
timestamp 1606120353
transform 1 0 33488 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A2
timestamp 1606120353
transform 1 0 33120 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_19_347
timestamp 1606120353
transform 1 0 33028 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1606120353
transform 1 0 34776 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__A1
timestamp 1606120353
transform 1 0 33856 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_19_359
timestamp 1606120353
transform 1 0 34132 0 1 12512
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_19_365
timestamp 1606120353
transform 1 0 34684 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_19_367
timestamp 1606120353
transform 1 0 34868 0 1 12512
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_20_354
timestamp 1606120353
transform 1 0 33672 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_20_358
timestamp 1606120353
transform 1 0 34040 0 -1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_20_370
timestamp 1606120353
transform 1 0 35144 0 -1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1152_
timestamp 1606120353
transform 1 0 35788 0 1 12512
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__D
timestamp 1606120353
transform 1 0 35604 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_19_396
timestamp 1606120353
transform 1 0 37536 0 1 12512
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_20_382
timestamp 1606120353
transform 1 0 36248 0 -1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_20_394
timestamp 1606120353
transform 1 0 37352 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606120353
transform -1 0 38548 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606120353
transform -1 0 38548 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1606120353
transform 1 0 37628 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_20_398
timestamp 1606120353
transform 1 0 37720 0 -1 13600
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606120353
transform 1 0 1104 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__D
timestamp 1606120353
transform 1 0 3036 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__CLK
timestamp 1606120353
transform 1 0 2668 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1606120353
transform 1 0 1380 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_21_15
timestamp 1606120353
transform 1 0 2484 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_19
timestamp 1606120353
transform 1 0 2852 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1107_
timestamp 1606120353
transform 1 0 3220 0 1 13600
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__C
timestamp 1606120353
transform 1 0 5152 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_42
timestamp 1606120353
transform 1 0 4968 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0624_
timestamp 1606120353
transform 1 0 5704 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__and2_4  _0628_
timestamp 1606120353
transform 1 0 6808 0 1 13600
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1606120353
transform 1 0 6716 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__A
timestamp 1606120353
transform 1 0 6532 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0624__A
timestamp 1606120353
transform 1 0 6164 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__A
timestamp 1606120353
transform 1 0 5520 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_46
timestamp 1606120353
transform 1 0 5336 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1606120353
transform 1 0 5980 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1606120353
transform 1 0 6348 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0613_
timestamp 1606120353
transform 1 0 8464 0 1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__B
timestamp 1606120353
transform 1 0 7636 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__C
timestamp 1606120353
transform 1 0 8280 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_69
timestamp 1606120353
transform 1 0 7452 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_21_73
timestamp 1606120353
transform 1 0 7820 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_21_77
timestamp 1606120353
transform 1 0 8188 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0696_
timestamp 1606120353
transform 1 0 10028 0 1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__A
timestamp 1606120353
transform 1 0 9844 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__C
timestamp 1606120353
transform 1 0 9476 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__C
timestamp 1606120353
transform 1 0 11040 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_89
timestamp 1606120353
transform 1 0 9292 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_93
timestamp 1606120353
transform 1 0 9660 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_106
timestamp 1606120353
transform 1 0 10856 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1606120353
transform 1 0 11224 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__B
timestamp 1606120353
transform 1 0 11408 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1606120353
transform 1 0 11592 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__D
timestamp 1606120353
transform 1 0 11776 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1606120353
transform 1 0 11960 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__C
timestamp 1606120353
transform 1 0 12144 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1606120353
transform 1 0 12328 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1606120353
transform 1 0 12420 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0569_
timestamp 1606120353
transform 1 0 12604 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_21_128
timestamp 1606120353
transform 1 0 12880 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__A
timestamp 1606120353
transform 1 0 13064 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1606120353
transform 1 0 13248 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0558_
timestamp 1606120353
transform 1 0 13616 0 1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__buf_1  _0566_
timestamp 1606120353
transform 1 0 15180 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__D
timestamp 1606120353
transform 1 0 13432 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__A
timestamp 1606120353
transform 1 0 14996 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__B
timestamp 1606120353
transform 1 0 14628 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_145
timestamp 1606120353
transform 1 0 14444 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_149
timestamp 1606120353
transform 1 0 14812 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0646_
timestamp 1606120353
transform 1 0 16376 0 1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__C
timestamp 1606120353
transform 1 0 15916 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_21_156
timestamp 1606120353
transform 1 0 15456 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_21_160
timestamp 1606120353
transform 1 0 15824 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_21_163
timestamp 1606120353
transform 1 0 16100 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_21_175
timestamp 1606120353
transform 1 0 17204 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__or4_4  _0556_
timestamp 1606120353
transform 1 0 18952 0 1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1606120353
transform 1 0 17940 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__B
timestamp 1606120353
transform 1 0 18768 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__A
timestamp 1606120353
transform 1 0 17572 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__B
timestamp 1606120353
transform 1 0 18400 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1606120353
transform 1 0 17756 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_21_184
timestamp 1606120353
transform 1 0 18032 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_21_190
timestamp 1606120353
transform 1 0 18584 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0504_
timestamp 1606120353
transform 1 0 20516 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__A
timestamp 1606120353
transform 1 0 19964 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0523__A
timestamp 1606120353
transform 1 0 20976 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__C
timestamp 1606120353
transform 1 0 20332 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A1
timestamp 1606120353
transform 1 0 21344 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_203
timestamp 1606120353
transform 1 0 19780 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_207
timestamp 1606120353
transform 1 0 20148 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_214
timestamp 1606120353
transform 1 0 20792 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_218
timestamp 1606120353
transform 1 0 21160 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1030_
timestamp 1606120353
transform 1 0 21528 0 1 13600
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__B
timestamp 1606120353
transform 1 0 23368 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__C
timestamp 1606120353
transform 1 0 23000 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_21_235
timestamp 1606120353
transform 1 0 22724 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1606120353
transform 1 0 23184 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0950_
timestamp 1606120353
transform 1 0 24380 0 1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1606120353
transform 1 0 23552 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A
timestamp 1606120353
transform 1 0 23920 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__D
timestamp 1606120353
transform 1 0 25392 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_21_245
timestamp 1606120353
transform 1 0 23644 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_21_250
timestamp 1606120353
transform 1 0 24104 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_21_262
timestamp 1606120353
transform 1 0 25208 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _1000_
timestamp 1606120353
transform 1 0 25944 0 1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__B
timestamp 1606120353
transform 1 0 25760 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A
timestamp 1606120353
transform 1 0 26956 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A
timestamp 1606120353
transform 1 0 27324 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_266
timestamp 1606120353
transform 1 0 25576 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_279
timestamp 1606120353
transform 1 0 26772 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_283
timestamp 1606120353
transform 1 0 27140 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0955_
timestamp 1606120353
transform 1 0 29256 0 1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__buf_1  _0995_
timestamp 1606120353
transform 1 0 27508 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1606120353
transform 1 0 29164 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__D
timestamp 1606120353
transform 1 0 28980 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__C
timestamp 1606120353
transform 1 0 28428 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A
timestamp 1606120353
transform 1 0 28060 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_21_290
timestamp 1606120353
transform 1 0 27784 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_21_295
timestamp 1606120353
transform 1 0 28244 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_21_299
timestamp 1606120353
transform 1 0 28612 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__o21a_4  _1037_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 30912 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__C
timestamp 1606120353
transform 1 0 30268 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__A
timestamp 1606120353
transform 1 0 30636 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_315
timestamp 1606120353
transform 1 0 30084 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_319
timestamp 1606120353
transform 1 0 30452 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_21_323
timestamp 1606120353
transform 1 0 30820 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__o21ai_4  _0997_
timestamp 1606120353
transform 1 0 32752 0 1 13600
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A1
timestamp 1606120353
transform 1 0 32568 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A
timestamp 1606120353
transform 1 0 32200 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_336
timestamp 1606120353
transform 1 0 32016 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_340
timestamp 1606120353
transform 1 0 32384 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1606120353
transform 1 0 34776 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__B1
timestamp 1606120353
transform 1 0 34132 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__A2
timestamp 1606120353
transform 1 0 34500 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_357
timestamp 1606120353
transform 1 0 33948 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_361
timestamp 1606120353
transform 1 0 34316 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_21_365
timestamp 1606120353
transform 1 0 34684 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_21_367
timestamp 1606120353
transform 1 0 34868 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_21_379
timestamp 1606120353
transform 1 0 35972 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_21_391
timestamp 1606120353
transform 1 0 37076 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606120353
transform -1 0 38548 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_21_403
timestamp 1606120353
transform 1 0 38180 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606120353
transform 1 0 1104 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__D
timestamp 1606120353
transform 1 0 1564 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__B2
timestamp 1606120353
transform 1 0 3036 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__CLK
timestamp 1606120353
transform 1 0 1932 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1606120353
transform 1 0 1380 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_7
timestamp 1606120353
transform 1 0 1748 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_22_11
timestamp 1606120353
transform 1 0 2116 0 -1 14688
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_22_19
timestamp 1606120353
transform 1 0 2852 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1606120353
transform 1 0 3220 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__D
timestamp 1606120353
transform 1 0 3404 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1606120353
transform 1 0 3588 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__C
timestamp 1606120353
transform 1 0 3772 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_22_32
timestamp 1606120353
transform 1 0 4048 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1606120353
transform 1 0 3956 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0543_
timestamp 1606120353
transform 1 0 4140 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_22_36
timestamp 1606120353
transform 1 0 4416 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__A
timestamp 1606120353
transform 1 0 4600 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_22_40
timestamp 1606120353
transform 1 0 4784 0 -1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_22_44
timestamp 1606120353
transform 1 0 5152 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_22_47
timestamp 1606120353
transform 1 0 5428 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__B
timestamp 1606120353
transform 1 0 5244 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__B1
timestamp 1606120353
transform 1 0 5612 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_51
timestamp 1606120353
transform 1 0 5796 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__B2
timestamp 1606120353
transform 1 0 5980 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_22_55
timestamp 1606120353
transform 1 0 6164 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0629_
timestamp 1606120353
transform 1 0 6440 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_22_61
timestamp 1606120353
transform 1 0 6716 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__A
timestamp 1606120353
transform 1 0 6992 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_66
timestamp 1606120353
transform 1 0 7176 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0702_
timestamp 1606120353
transform 1 0 7912 0 -1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__B
timestamp 1606120353
transform 1 0 8924 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A
timestamp 1606120353
transform 1 0 7728 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__C
timestamp 1606120353
transform 1 0 7360 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_70
timestamp 1606120353
transform 1 0 7544 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_83
timestamp 1606120353
transform 1 0 8740 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_87
timestamp 1606120353
transform 1 0 9108 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0698_
timestamp 1606120353
transform 1 0 9936 0 -1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1606120353
transform 1 0 9568 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__A
timestamp 1606120353
transform 1 0 10948 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__A
timestamp 1606120353
transform 1 0 9292 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1606120353
transform 1 0 9476 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1606120353
transform 1 0 9660 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_22_105
timestamp 1606120353
transform 1 0 10764 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_109
timestamp 1606120353
transform 1 0 11132 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0503_
timestamp 1606120353
transform 1 0 11868 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__and4_4  _0580_
timestamp 1606120353
transform 1 0 13064 0 -1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__B
timestamp 1606120353
transform 1 0 12880 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__B
timestamp 1606120353
transform 1 0 12420 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__B
timestamp 1606120353
transform 1 0 11316 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__A
timestamp 1606120353
transform 1 0 11684 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_113
timestamp 1606120353
transform 1 0 11500 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_22_120
timestamp 1606120353
transform 1 0 12144 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_22_125
timestamp 1606120353
transform 1 0 12604 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1606120353
transform 1 0 15180 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__C
timestamp 1606120353
transform 1 0 14076 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0566__A
timestamp 1606120353
transform 1 0 14996 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__B2
timestamp 1606120353
transform 1 0 14444 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_139
timestamp 1606120353
transform 1 0 13892 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_143
timestamp 1606120353
transform 1 0 14260 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_22_147
timestamp 1606120353
transform 1 0 14628 0 -1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_22_154
timestamp 1606120353
transform 1 0 15272 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0645_
timestamp 1606120353
transform 1 0 15916 0 -1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0553__A
timestamp 1606120353
transform 1 0 15456 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__B
timestamp 1606120353
transform 1 0 16928 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_22_158
timestamp 1606120353
transform 1 0 15640 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_22_170
timestamp 1606120353
transform 1 0 16744 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_22_174
timestamp 1606120353
transform 1 0 17112 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__and4_4  _0586_
timestamp 1606120353
transform 1 0 19136 0 -1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__and4_4  _0587_
timestamp 1606120353
transform 1 0 17572 0 -1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__D
timestamp 1606120353
transform 1 0 18952 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__A
timestamp 1606120353
transform 1 0 18584 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__C
timestamp 1606120353
transform 1 0 17388 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_188
timestamp 1606120353
transform 1 0 18400 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_192
timestamp 1606120353
transform 1 0 18768 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0523_
timestamp 1606120353
transform 1 0 20884 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1606120353
transform 1 0 20792 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__D
timestamp 1606120353
transform 1 0 20148 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__D
timestamp 1606120353
transform 1 0 20516 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_205
timestamp 1606120353
transform 1 0 19964 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_209
timestamp 1606120353
transform 1 0 20332 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_22_213
timestamp 1606120353
transform 1 0 20700 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_22_218
timestamp 1606120353
transform 1 0 21160 0 -1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A2
timestamp 1606120353
transform 1 0 21528 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_224
timestamp 1606120353
transform 1 0 21712 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1004_
timestamp 1606120353
transform 1 0 21896 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_22_229
timestamp 1606120353
transform 1 0 22172 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__A
timestamp 1606120353
transform 1 0 22356 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_233
timestamp 1606120353
transform 1 0 22540 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A
timestamp 1606120353
transform 1 0 22724 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1032_
timestamp 1606120353
transform 1 0 22908 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_22_240
timestamp 1606120353
transform 1 0 23184 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__C
timestamp 1606120353
transform 1 0 23368 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _1031_
timestamp 1606120353
transform 1 0 23920 0 -1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A
timestamp 1606120353
transform 1 0 23736 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__C
timestamp 1606120353
transform 1 0 25208 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_244
timestamp 1606120353
transform 1 0 23552 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_22_257
timestamp 1606120353
transform 1 0 24748 0 -1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_22_261
timestamp 1606120353
transform 1 0 25116 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_22_264
timestamp 1606120353
transform 1 0 25392 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__C
timestamp 1606120353
transform 1 0 25576 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_268
timestamp 1606120353
transform 1 0 25760 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A
timestamp 1606120353
transform 1 0 25944 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_22_272
timestamp 1606120353
transform 1 0 26128 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1606120353
transform 1 0 26404 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0999_
timestamp 1606120353
transform 1 0 26496 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_22_279
timestamp 1606120353
transform 1 0 26772 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__D
timestamp 1606120353
transform 1 0 26956 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_283
timestamp 1606120353
transform 1 0 27140 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A
timestamp 1606120353
transform 1 0 27324 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _0952_
timestamp 1606120353
transform 1 0 28428 0 -1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__B
timestamp 1606120353
transform 1 0 29440 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__B
timestamp 1606120353
transform 1 0 28244 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A
timestamp 1606120353
transform 1 0 27876 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_22_287
timestamp 1606120353
transform 1 0 27508 0 -1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_22_293
timestamp 1606120353
transform 1 0 28060 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1606120353
transform 1 0 29256 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__nor3_4  _1029_
timestamp 1606120353
transform 1 0 30084 0 -1 14688
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__C
timestamp 1606120353
transform 1 0 29808 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A2
timestamp 1606120353
transform 1 0 31464 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_310
timestamp 1606120353
transform 1 0 29624 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_22_314
timestamp 1606120353
transform 1 0 29992 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_22_328
timestamp 1606120353
transform 1 0 31280 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_340
timestamp 1606120353
transform 1 0 32384 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_332
timestamp 1606120353
transform 1 0 31648 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__B1
timestamp 1606120353
transform 1 0 31832 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1606120353
transform 1 0 32016 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0979_
timestamp 1606120353
transform 1 0 32108 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_22_348
timestamp 1606120353
transform 1 0 33120 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_22_344
timestamp 1606120353
transform 1 0 32752 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__B1
timestamp 1606120353
transform 1 0 32936 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A1
timestamp 1606120353
transform 1 0 32568 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1002_
timestamp 1606120353
transform 1 0 33396 0 -1 14688
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILLER_22_364
timestamp 1606120353
transform 1 0 34592 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_22_376
timestamp 1606120353
transform 1 0 35696 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_22_388
timestamp 1606120353
transform 1 0 36800 0 -1 14688
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_22_396
timestamp 1606120353
transform 1 0 37536 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606120353
transform -1 0 38548 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1606120353
transform 1 0 37628 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_22_398
timestamp 1606120353
transform 1 0 37720 0 -1 14688
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1136_
timestamp 1606120353
transform 1 0 1380 0 1 14688
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606120353
transform 1 0 1104 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_23_22
timestamp 1606120353
transform 1 0 3128 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _0812_
timestamp 1606120353
transform 1 0 3864 0 1 14688
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__B1
timestamp 1606120353
transform 1 0 3680 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__B
timestamp 1606120353
transform 1 0 3312 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_26
timestamp 1606120353
transform 1 0 3496 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_44
timestamp 1606120353
transform 1 0 5152 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_23_48
timestamp 1606120353
transform 1 0 5520 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_23_51
timestamp 1606120353
transform 1 0 5796 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__A3
timestamp 1606120353
transform 1 0 5612 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_55
timestamp 1606120353
transform 1 0 6164 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__A1
timestamp 1606120353
transform 1 0 5980 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1606120353
transform 1 0 6532 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__A2
timestamp 1606120353
transform 1 0 6348 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_62
timestamp 1606120353
transform 1 0 6808 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1606120353
transform 1 0 6716 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__A
timestamp 1606120353
transform 1 0 7176 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0701_
timestamp 1606120353
transform 1 0 8924 0 1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__or4_4  _0703_
timestamp 1606120353
transform 1 0 7360 0 1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__C
timestamp 1606120353
transform 1 0 8740 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__D
timestamp 1606120353
transform 1 0 8372 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_77
timestamp 1606120353
transform 1 0 8188 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_81
timestamp 1606120353
transform 1 0 8556 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0699_
timestamp 1606120353
transform 1 0 10764 0 1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__C
timestamp 1606120353
transform 1 0 10580 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0606__A
timestamp 1606120353
transform 1 0 9936 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_94
timestamp 1606120353
transform 1 0 9752 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_98
timestamp 1606120353
transform 1 0 10120 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_23_102
timestamp 1606120353
transform 1 0 10488 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0583_
timestamp 1606120353
transform 1 0 12420 0 1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1606120353
transform 1 0 12328 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__A
timestamp 1606120353
transform 1 0 12144 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__C
timestamp 1606120353
transform 1 0 11776 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_114
timestamp 1606120353
transform 1 0 11592 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1606120353
transform 1 0 11960 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_132
timestamp 1606120353
transform 1 0 13248 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__a22oi_4  _0573_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 14444 0 1 14688
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__A2
timestamp 1606120353
transform 1 0 14260 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__A
timestamp 1606120353
transform 1 0 13432 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__B
timestamp 1606120353
transform 1 0 13800 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_136
timestamp 1606120353
transform 1 0 13616 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_23_140
timestamp 1606120353
transform 1 0 13984 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0565_
timestamp 1606120353
transform 1 0 16744 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__A
timestamp 1606120353
transform 1 0 16468 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0565__A
timestamp 1606120353
transform 1 0 17204 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_162
timestamp 1606120353
transform 1 0 16008 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_23_166
timestamp 1606120353
transform 1 0 16376 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_23_169
timestamp 1606120353
transform 1 0 16652 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_23_173
timestamp 1606120353
transform 1 0 17020 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0588_
timestamp 1606120353
transform 1 0 18308 0 1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1606120353
transform 1 0 17940 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__A
timestamp 1606120353
transform 1 0 19320 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__C
timestamp 1606120353
transform 1 0 17572 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_177
timestamp 1606120353
transform 1 0 17388 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1606120353
transform 1 0 17756 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_23_184
timestamp 1606120353
transform 1 0 18032 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_23_196
timestamp 1606120353
transform 1 0 19136 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0555_
timestamp 1606120353
transform 1 0 19872 0 1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__B
timestamp 1606120353
transform 1 0 19688 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__A
timestamp 1606120353
transform 1 0 21068 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_200
timestamp 1606120353
transform 1 0 19504 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_213
timestamp 1606120353
transform 1 0 20700 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_23_219
timestamp 1606120353
transform 1 0 21252 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1033_
timestamp 1606120353
transform 1 0 21620 0 1 14688
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A1
timestamp 1606120353
transform 1 0 21436 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__B
timestamp 1606120353
transform 1 0 23368 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__C
timestamp 1606120353
transform 1 0 23000 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_236
timestamp 1606120353
transform 1 0 22816 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1606120353
transform 1 0 23184 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _1024_
timestamp 1606120353
transform 1 0 24012 0 1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1606120353
transform 1 0 23552 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A
timestamp 1606120353
transform 1 0 25392 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__B
timestamp 1606120353
transform 1 0 23828 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__D
timestamp 1606120353
transform 1 0 25024 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_245
timestamp 1606120353
transform 1 0 23644 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_258
timestamp 1606120353
transform 1 0 24840 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_262
timestamp 1606120353
transform 1 0 25208 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0978_
timestamp 1606120353
transform 1 0 25944 0 1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__B
timestamp 1606120353
transform 1 0 26956 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__B
timestamp 1606120353
transform 1 0 25760 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__C
timestamp 1606120353
transform 1 0 27324 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_266
timestamp 1606120353
transform 1 0 25576 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_279
timestamp 1606120353
transform 1 0 26772 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_283
timestamp 1606120353
transform 1 0 27140 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_290
timestamp 1606120353
transform 1 0 27784 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _1001_
timestamp 1606120353
transform 1 0 27508 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_23_294
timestamp 1606120353
transform 1 0 28152 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_23_297
timestamp 1606120353
transform 1 0 28428 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__C
timestamp 1606120353
transform 1 0 28244 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_301
timestamp 1606120353
transform 1 0 28796 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__D
timestamp 1606120353
transform 1 0 28612 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_306
timestamp 1606120353
transform 1 0 29256 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__B
timestamp 1606120353
transform 1 0 28980 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1606120353
transform 1 0 29164 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A
timestamp 1606120353
transform 1 0 29440 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__nor3_4  _0988_
timestamp 1606120353
transform 1 0 29624 0 1 14688
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__C
timestamp 1606120353
transform 1 0 31004 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__D
timestamp 1606120353
transform 1 0 31372 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_323
timestamp 1606120353
transform 1 0 30820 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_327
timestamp 1606120353
transform 1 0 31188 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0996_
timestamp 1606120353
transform 1 0 32476 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A2
timestamp 1606120353
transform 1 0 32292 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A
timestamp 1606120353
transform 1 0 31924 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_331
timestamp 1606120353
transform 1 0 31556 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1606120353
transform 1 0 32108 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_361
timestamp 1606120353
transform 1 0 34316 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_357
timestamp 1606120353
transform 1 0 33948 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_353
timestamp 1606120353
transform 1 0 33580 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__B1
timestamp 1606120353
transform 1 0 34500 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A1
timestamp 1606120353
transform 1 0 34132 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__B
timestamp 1606120353
transform 1 0 33764 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_367
timestamp 1606120353
transform 1 0 34868 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_23_365
timestamp 1606120353
transform 1 0 34684 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A2
timestamp 1606120353
transform 1 0 35052 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1606120353
transform 1 0 34776 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_23_371
timestamp 1606120353
transform 1 0 35236 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_23_383
timestamp 1606120353
transform 1 0 36340 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_23_395
timestamp 1606120353
transform 1 0 37444 0 1 14688
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606120353
transform -1 0 38548 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_23_403
timestamp 1606120353
transform 1 0 38180 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606120353
transform 1 0 1104 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__D
timestamp 1606120353
transform 1 0 1564 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A2
timestamp 1606120353
transform 1 0 3036 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1606120353
transform 1 0 1380 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_24_7
timestamp 1606120353
transform 1 0 1748 0 -1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_24_19
timestamp 1606120353
transform 1 0 2852 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_23
timestamp 1606120353
transform 1 0 3220 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A1
timestamp 1606120353
transform 1 0 3404 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1606120353
transform 1 0 3588 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A4
timestamp 1606120353
transform 1 0 3772 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1606120353
transform 1 0 3956 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_24_32
timestamp 1606120353
transform 1 0 4048 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_24_37
timestamp 1606120353
transform 1 0 4508 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A2
timestamp 1606120353
transform 1 0 4324 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0592_
timestamp 1606120353
transform 1 0 4600 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_24_41
timestamp 1606120353
transform 1 0 4876 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__A2
timestamp 1606120353
transform 1 0 5060 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__a32o_4  _0590_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 5612 0 -1 15776
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__C1
timestamp 1606120353
transform 1 0 5428 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_45
timestamp 1606120353
transform 1 0 5244 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_66
timestamp 1606120353
transform 1 0 7176 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0704_
timestamp 1606120353
transform 1 0 7912 0 -1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__A
timestamp 1606120353
transform 1 0 8924 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__C
timestamp 1606120353
transform 1 0 7360 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__B
timestamp 1606120353
transform 1 0 7728 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_70
timestamp 1606120353
transform 1 0 7544 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_83
timestamp 1606120353
transform 1 0 8740 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_87
timestamp 1606120353
transform 1 0 9108 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0606_
timestamp 1606120353
transform 1 0 9660 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__and4_4  _0697_
timestamp 1606120353
transform 1 0 10856 0 -1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1606120353
transform 1 0 9568 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__C
timestamp 1606120353
transform 1 0 10672 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__B
timestamp 1606120353
transform 1 0 9292 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__C
timestamp 1606120353
transform 1 0 10120 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1606120353
transform 1 0 9476 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_24_96
timestamp 1606120353
transform 1 0 9936 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_24_100
timestamp 1606120353
transform 1 0 10304 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__nor4_4  _0589_
timestamp 1606120353
transform 1 0 12880 0 -1 15776
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__A
timestamp 1606120353
transform 1 0 12420 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__C
timestamp 1606120353
transform 1 0 12052 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_24_115
timestamp 1606120353
transform 1 0 11684 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_24_121
timestamp 1606120353
transform 1 0 12236 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_24_125
timestamp 1606120353
transform 1 0 12604 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0553_
timestamp 1606120353
transform 1 0 15272 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1606120353
transform 1 0 15180 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__D
timestamp 1606120353
transform 1 0 14628 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__D
timestamp 1606120353
transform 1 0 14996 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_145
timestamp 1606120353
transform 1 0 14444 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_149
timestamp 1606120353
transform 1 0 14812 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0644_
timestamp 1606120353
transform 1 0 16468 0 -1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0538__A
timestamp 1606120353
transform 1 0 16008 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_24_157
timestamp 1606120353
transform 1 0 15548 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_24_161
timestamp 1606120353
transform 1 0 15916 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_24_164
timestamp 1606120353
transform 1 0 16192 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_24_176
timestamp 1606120353
transform 1 0 17296 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__and4_4  _0585_
timestamp 1606120353
transform 1 0 18860 0 -1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__B
timestamp 1606120353
transform 1 0 18032 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__C
timestamp 1606120353
transform 1 0 18676 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__B
timestamp 1606120353
transform 1 0 17664 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_182
timestamp 1606120353
transform 1 0 17848 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_24_186
timestamp 1606120353
transform 1 0 18216 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_24_190
timestamp 1606120353
transform 1 0 18584 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_24_202
timestamp 1606120353
transform 1 0 19688 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1606120353
transform 1 0 20056 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__D
timestamp 1606120353
transform 1 0 19872 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1606120353
transform 1 0 20424 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A
timestamp 1606120353
transform 1 0 20240 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A2
timestamp 1606120353
transform 1 0 20608 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1606120353
transform 1 0 20792 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1606120353
transform 1 0 20884 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__B2
timestamp 1606120353
transform 1 0 21068 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1606120353
transform 1 0 21252 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _1015_
timestamp 1606120353
transform 1 0 22816 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _1025_
timestamp 1606120353
transform 1 0 21804 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__D
timestamp 1606120353
transform 1 0 23276 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B1
timestamp 1606120353
transform 1 0 21620 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A2
timestamp 1606120353
transform 1 0 22264 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__B1
timestamp 1606120353
transform 1 0 22632 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_228
timestamp 1606120353
transform 1 0 22080 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_232
timestamp 1606120353
transform 1 0 22448 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_239
timestamp 1606120353
transform 1 0 23092 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1007_
timestamp 1606120353
transform 1 0 25392 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__or4_4  _1014_
timestamp 1606120353
transform 1 0 23828 0 -1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__B
timestamp 1606120353
transform 1 0 24840 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__C
timestamp 1606120353
transform 1 0 25208 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__A
timestamp 1606120353
transform 1 0 23644 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_243
timestamp 1606120353
transform 1 0 23460 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_256
timestamp 1606120353
transform 1 0 24656 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_260
timestamp 1606120353
transform 1 0 25024 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0991_
timestamp 1606120353
transform 1 0 26496 0 -1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1606120353
transform 1 0 26404 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__B
timestamp 1606120353
transform 1 0 26220 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__D
timestamp 1606120353
transform 1 0 25852 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_267
timestamp 1606120353
transform 1 0 25668 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_271
timestamp 1606120353
transform 1 0 26036 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_285
timestamp 1606120353
transform 1 0 27324 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _1009_
timestamp 1606120353
transform 1 0 28244 0 -1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__C
timestamp 1606120353
transform 1 0 29256 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A
timestamp 1606120353
transform 1 0 27508 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__D
timestamp 1606120353
transform 1 0 27876 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_289
timestamp 1606120353
transform 1 0 27692 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_293
timestamp 1606120353
transform 1 0 28060 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_304
timestamp 1606120353
transform 1 0 29072 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_308
timestamp 1606120353
transform 1 0 29440 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0987_
timestamp 1606120353
transform 1 0 29808 0 -1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A
timestamp 1606120353
transform 1 0 29624 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__B
timestamp 1606120353
transform 1 0 30820 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__B
timestamp 1606120353
transform 1 0 31188 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_321
timestamp 1606120353
transform 1 0 30636 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_325
timestamp 1606120353
transform 1 0 31004 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_24_329
timestamp 1606120353
transform 1 0 31372 0 -1 15776
box 0 -48 552 592
use sky130_fd_sc_hd__nor2_4  _1026_
timestamp 1606120353
transform 1 0 32108 0 -1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1606120353
transform 1 0 32016 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A2
timestamp 1606120353
transform 1 0 33120 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_24_335
timestamp 1606120353
transform 1 0 31924 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_24_346
timestamp 1606120353
transform 1 0 32936 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_24_350
timestamp 1606120353
transform 1 0 33304 0 -1 15776
box 0 -48 552 592
use sky130_fd_sc_hd__o21ai_4  _1016_
timestamp 1606120353
transform 1 0 33948 0 -1 15776
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_1  FILLER_24_356
timestamp 1606120353
transform 1 0 33856 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_24_370
timestamp 1606120353
transform 1 0 35144 0 -1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_24_382
timestamp 1606120353
transform 1 0 36248 0 -1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_24_394
timestamp 1606120353
transform 1 0 37352 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606120353
transform -1 0 38548 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1606120353
transform 1 0 37628 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_24_398
timestamp 1606120353
transform 1 0 37720 0 -1 15776
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1124_
timestamp 1606120353
transform 1 0 1380 0 1 15776
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606120353
transform 1 0 1104 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_25_22
timestamp 1606120353
transform 1 0 3128 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__a211o_4  _0632_
timestamp 1606120353
transform 1 0 4692 0 1 15776
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__A1
timestamp 1606120353
transform 1 0 4508 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A1
timestamp 1606120353
transform 1 0 4140 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__B1
timestamp 1606120353
transform 1 0 3772 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A3
timestamp 1606120353
transform 1 0 3404 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_27
timestamp 1606120353
transform 1 0 3588 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_31
timestamp 1606120353
transform 1 0 3956 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_35
timestamp 1606120353
transform 1 0 4324 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0631_
timestamp 1606120353
transform 1 0 6808 0 1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1606120353
transform 1 0 6716 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__A
timestamp 1606120353
transform 1 0 6532 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0541__A
timestamp 1606120353
transform 1 0 6164 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1606120353
transform 1 0 5980 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1606120353
transform 1 0 6348 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__nor4_4  _0618_
timestamp 1606120353
transform 1 0 8740 0 1 15776
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__C
timestamp 1606120353
transform 1 0 7820 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A
timestamp 1606120353
transform 1 0 8188 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__A
timestamp 1606120353
transform 1 0 8556 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_71
timestamp 1606120353
transform 1 0 7636 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_75
timestamp 1606120353
transform 1 0 8004 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_79
timestamp 1606120353
transform 1 0 8372 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0534_
timestamp 1606120353
transform 1 0 11040 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0513__A
timestamp 1606120353
transform 1 0 10488 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__A
timestamp 1606120353
transform 1 0 10856 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_100
timestamp 1606120353
transform 1 0 10304 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_104
timestamp 1606120353
transform 1 0 10672 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0579_
timestamp 1606120353
transform 1 0 12420 0 1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1606120353
transform 1 0 12328 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__B
timestamp 1606120353
transform 1 0 12144 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0534__A
timestamp 1606120353
transform 1 0 11500 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_111
timestamp 1606120353
transform 1 0 11316 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_25_115
timestamp 1606120353
transform 1 0 11684 0 1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1606120353
transform 1 0 12052 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1606120353
transform 1 0 13248 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _0505_
timestamp 1606120353
transform 1 0 13984 0 1 15776
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0505__A
timestamp 1606120353
transform 1 0 14812 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0505__B
timestamp 1606120353
transform 1 0 13800 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0531__A
timestamp 1606120353
transform 1 0 13432 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__C
timestamp 1606120353
transform 1 0 15180 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_136
timestamp 1606120353
transform 1 0 13616 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_147
timestamp 1606120353
transform 1 0 14628 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_151
timestamp 1606120353
transform 1 0 14996 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_155
timestamp 1606120353
transform 1 0 15364 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0533__A
timestamp 1606120353
transform 1 0 15548 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_25_159
timestamp 1606120353
transform 1 0 15732 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0538_
timestamp 1606120353
transform 1 0 16008 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1606120353
transform 1 0 16284 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__B
timestamp 1606120353
transform 1 0 16560 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_170
timestamp 1606120353
transform 1 0 16744 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__A
timestamp 1606120353
transform 1 0 16928 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_174
timestamp 1606120353
transform 1 0 17112 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__D
timestamp 1606120353
transform 1 0 17296 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0584_
timestamp 1606120353
transform 1 0 18032 0 1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1606120353
transform 1 0 17940 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__B
timestamp 1606120353
transform 1 0 19044 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__A
timestamp 1606120353
transform 1 0 17756 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_25_178
timestamp 1606120353
transform 1 0 17480 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_25_193
timestamp 1606120353
transform 1 0 18860 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_197
timestamp 1606120353
transform 1 0 19228 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0581_
timestamp 1606120353
transform 1 0 19596 0 1 15776
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0581__A
timestamp 1606120353
transform 1 0 20424 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__A
timestamp 1606120353
transform 1 0 19412 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__B1
timestamp 1606120353
transform 1 0 20884 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A1
timestamp 1606120353
transform 1 0 21252 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_208
timestamp 1606120353
transform 1 0 20240 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_25_212
timestamp 1606120353
transform 1 0 20608 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_25_217
timestamp 1606120353
transform 1 0 21068 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1081_
timestamp 1606120353
transform 1 0 21528 0 1 15776
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A1
timestamp 1606120353
transform 1 0 22908 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__D
timestamp 1606120353
transform 1 0 23368 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_25_221
timestamp 1606120353
transform 1 0 21436 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_25_235
timestamp 1606120353
transform 1 0 22724 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_25_239
timestamp 1606120353
transform 1 0 23092 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0977_
timestamp 1606120353
transform 1 0 23644 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__or4_4  _1017_
timestamp 1606120353
transform 1 0 24748 0 1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1606120353
transform 1 0 23552 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A
timestamp 1606120353
transform 1 0 24564 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__B
timestamp 1606120353
transform 1 0 24196 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_25_248
timestamp 1606120353
transform 1 0 23920 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_25_253
timestamp 1606120353
transform 1 0 24380 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _1021_
timestamp 1606120353
transform 1 0 26312 0 1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__B
timestamp 1606120353
transform 1 0 26128 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__A
timestamp 1606120353
transform 1 0 25760 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__A
timestamp 1606120353
transform 1 0 27324 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_266
timestamp 1606120353
transform 1 0 25576 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_270
timestamp 1606120353
transform 1 0 25944 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_283
timestamp 1606120353
transform 1 0 27140 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_297
timestamp 1606120353
transform 1 0 28428 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_25_291
timestamp 1606120353
transform 1 0 27876 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_25_287
timestamp 1606120353
transform 1 0 27508 0 1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__B
timestamp 1606120353
transform 1 0 27968 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0986_
timestamp 1606120353
transform 1 0 28152 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_25_306
timestamp 1606120353
transform 1 0 29256 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_301
timestamp 1606120353
transform 1 0 28796 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__A
timestamp 1606120353
transform 1 0 28980 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A
timestamp 1606120353
transform 1 0 28612 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1606120353
transform 1 0 29164 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__nor3_4  _1011_
timestamp 1606120353
transform 1 0 29440 0 1 15776
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A
timestamp 1606120353
transform 1 0 30820 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A
timestamp 1606120353
transform 1 0 31188 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_321
timestamp 1606120353
transform 1 0 30636 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_325
timestamp 1606120353
transform 1 0 31004 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_25_329
timestamp 1606120353
transform 1 0 31372 0 1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__o21a_4  _0989_
timestamp 1606120353
transform 1 0 32292 0 1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A2
timestamp 1606120353
transform 1 0 32108 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__B1
timestamp 1606120353
transform 1 0 31740 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_335
timestamp 1606120353
transform 1 0 31924 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_351
timestamp 1606120353
transform 1 0 33396 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_25_359
timestamp 1606120353
transform 1 0 34132 0 1 15776
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_25_355
timestamp 1606120353
transform 1 0 33764 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__B1
timestamp 1606120353
transform 1 0 33948 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A1
timestamp 1606120353
transform 1 0 33580 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_370
timestamp 1606120353
transform 1 0 35144 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_25_365
timestamp 1606120353
transform 1 0 34684 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A
timestamp 1606120353
transform 1 0 35328 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1606120353
transform 1 0 34776 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0985_
timestamp 1606120353
transform 1 0 34868 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_25_374
timestamp 1606120353
transform 1 0 35512 0 1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_25_386
timestamp 1606120353
transform 1 0 36616 0 1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606120353
transform -1 0 38548 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_25_398
timestamp 1606120353
transform 1 0 37720 0 1 15776
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606120353
transform 1 0 1104 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606120353
transform 1 0 1104 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1606120353
transform 1 0 1380 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1606120353
transform 1 0 1380 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__B2
timestamp 1606120353
transform 1 0 1564 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__CLK
timestamp 1606120353
transform 1 0 1564 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A1
timestamp 1606120353
transform 1 0 1932 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A2
timestamp 1606120353
transform 1 0 1932 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_7
timestamp 1606120353
transform 1 0 1748 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1606120353
transform 1 0 1748 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_11
timestamp 1606120353
transform 1 0 2116 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_19
timestamp 1606120353
transform 1 0 2852 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_15
timestamp 1606120353
transform 1 0 2484 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__B1
timestamp 1606120353
transform 1 0 2668 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__D
timestamp 1606120353
transform 1 0 2300 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__D
timestamp 1606120353
transform 1 0 3036 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1106_
timestamp 1606120353
transform 1 0 2116 0 1 16864
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_4  FILLER_27_30
timestamp 1606120353
transform 1 0 3864 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_26_32
timestamp 1606120353
transform 1 0 4048 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1606120353
transform 1 0 3588 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_23
timestamp 1606120353
transform 1 0 3220 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__D
timestamp 1606120353
transform 1 0 3404 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__B1
timestamp 1606120353
transform 1 0 3772 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1606120353
transform 1 0 3956 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_27_41
timestamp 1606120353
transform 1 0 4876 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_37
timestamp 1606120353
transform 1 0 4508 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_27_34
timestamp 1606120353
transform 1 0 4232 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__B
timestamp 1606120353
transform 1 0 4324 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__B
timestamp 1606120353
transform 1 0 4692 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__A
timestamp 1606120353
transform 1 0 5060 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__o41a_4  _0649_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 4324 0 -1 16864
box 0 -48 1564 592
use sky130_fd_sc_hd__fill_2  FILLER_27_53
timestamp 1606120353
transform 1 0 5980 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_27_45
timestamp 1606120353
transform 1 0 5244 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_26_52
timestamp 1606120353
transform 1 0 5888 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0591_
timestamp 1606120353
transform 1 0 5336 0 1 16864
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1606120353
transform 1 0 6808 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1606120353
transform 1 0 6348 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_56
timestamp 1606120353
transform 1 0 6256 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__B
timestamp 1606120353
transform 1 0 6072 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__C
timestamp 1606120353
transform 1 0 6440 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__A
timestamp 1606120353
transform 1 0 6164 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0535__A
timestamp 1606120353
transform 1 0 6532 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1606120353
transform 1 0 6716 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0541_
timestamp 1606120353
transform 1 0 6624 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_26_63
timestamp 1606120353
transform 1 0 6900 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A
timestamp 1606120353
transform 1 0 7084 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0690_
timestamp 1606120353
transform 1 0 6992 0 1 16864
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_27_73
timestamp 1606120353
transform 1 0 7820 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_26_71
timestamp 1606120353
transform 1 0 7636 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_26_67
timestamp 1606120353
transform 1 0 7268 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A
timestamp 1606120353
transform 1 0 8004 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__B
timestamp 1606120353
transform 1 0 7452 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0700_
timestamp 1606120353
transform 1 0 7728 0 -1 16864
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_27_84
timestamp 1606120353
transform 1 0 8832 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_77
timestamp 1606120353
transform 1 0 8188 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_26_81
timestamp 1606120353
transform 1 0 8556 0 -1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__C
timestamp 1606120353
transform 1 0 8372 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0539_
timestamp 1606120353
transform 1 0 8556 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_27_88
timestamp 1606120353
transform 1 0 9200 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_26_88
timestamp 1606120353
transform 1 0 9200 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_26_85
timestamp 1606120353
transform 1 0 8924 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__A
timestamp 1606120353
transform 1 0 9016 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0539__A
timestamp 1606120353
transform 1 0 9016 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp 1606120353
transform 1 0 10028 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_26_93
timestamp 1606120353
transform 1 0 9660 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__B
timestamp 1606120353
transform 1 0 9384 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__B
timestamp 1606120353
transform 1 0 10212 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__A
timestamp 1606120353
transform 1 0 9476 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1606120353
transform 1 0 9568 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0513_
timestamp 1606120353
transform 1 0 9752 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_27_106
timestamp 1606120353
transform 1 0 10856 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_26_101
timestamp 1606120353
transform 1 0 10396 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__B
timestamp 1606120353
transform 1 0 10580 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__B
timestamp 1606120353
transform 1 0 11224 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0694_
timestamp 1606120353
transform 1 0 10764 0 -1 16864
box 0 -48 828 592
use sky130_fd_sc_hd__nor3_4  _0611_
timestamp 1606120353
transform 1 0 9660 0 1 16864
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_4  FILLER_27_116
timestamp 1606120353
transform 1 0 11776 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_27_112
timestamp 1606120353
transform 1 0 11408 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_118
timestamp 1606120353
transform 1 0 11960 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_114
timestamp 1606120353
transform 1 0 11592 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__A
timestamp 1606120353
transform 1 0 11776 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__D
timestamp 1606120353
transform 1 0 11592 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__B
timestamp 1606120353
transform 1 0 12144 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__C
timestamp 1606120353
transform 1 0 12144 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1606120353
transform 1 0 12328 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _0633_
timestamp 1606120353
transform 1 0 12420 0 1 16864
box 0 -48 644 592
use sky130_fd_sc_hd__and3_4  _0619_
timestamp 1606120353
transform 1 0 12328 0 -1 16864
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_27_130
timestamp 1606120353
transform 1 0 13064 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_131
timestamp 1606120353
transform 1 0 13156 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__B
timestamp 1606120353
transform 1 0 13248 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_138
timestamp 1606120353
transform 1 0 13800 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_134
timestamp 1606120353
transform 1 0 13432 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_135
timestamp 1606120353
transform 1 0 13524 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__D
timestamp 1606120353
transform 1 0 13616 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__C
timestamp 1606120353
transform 1 0 13708 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__B
timestamp 1606120353
transform 1 0 13340 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0531_
timestamp 1606120353
transform 1 0 13892 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_27_143
timestamp 1606120353
transform 1 0 14260 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_146
timestamp 1606120353
transform 1 0 14536 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_142
timestamp 1606120353
transform 1 0 14168 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__B
timestamp 1606120353
transform 1 0 14352 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0530__A
timestamp 1606120353
transform 1 0 14444 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0530_
timestamp 1606120353
transform 1 0 13984 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_27_147
timestamp 1606120353
transform 1 0 14628 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_26_150
timestamp 1606120353
transform 1 0 14904 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__D
timestamp 1606120353
transform 1 0 14812 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__D
timestamp 1606120353
transform 1 0 14720 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1606120353
transform 1 0 15180 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _0525_
timestamp 1606120353
transform 1 0 14996 0 1 16864
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  FILLER_26_154
timestamp 1606120353
transform 1 0 15272 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_27_158
timestamp 1606120353
transform 1 0 15640 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_160
timestamp 1606120353
transform 1 0 15824 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0525__B
timestamp 1606120353
transform 1 0 15824 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0533_
timestamp 1606120353
transform 1 0 15548 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_27_162
timestamp 1606120353
transform 1 0 16008 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_164
timestamp 1606120353
transform 1 0 16192 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__C1
timestamp 1606120353
transform 1 0 16376 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__B1
timestamp 1606120353
transform 1 0 16008 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__A2
timestamp 1606120353
transform 1 0 16192 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0608_
timestamp 1606120353
transform 1 0 16376 0 1 16864
box 0 -48 644 592
use sky130_fd_sc_hd__and2_4  _0524_
timestamp 1606120353
transform 1 0 16560 0 -1 16864
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_27_173
timestamp 1606120353
transform 1 0 17020 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_175
timestamp 1606120353
transform 1 0 17204 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__B
timestamp 1606120353
transform 1 0 17204 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1606120353
transform 1 0 17756 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_177
timestamp 1606120353
transform 1 0 17388 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_26_183
timestamp 1606120353
transform 1 0 17940 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_26_179
timestamp 1606120353
transform 1 0 17572 0 -1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__A
timestamp 1606120353
transform 1 0 17388 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__D1
timestamp 1606120353
transform 1 0 17572 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1606120353
transform 1 0 17940 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_27_187
timestamp 1606120353
transform 1 0 18308 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_186
timestamp 1606120353
transform 1 0 18216 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__C
timestamp 1606120353
transform 1 0 18400 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0582__A
timestamp 1606120353
transform 1 0 18492 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__C
timestamp 1606120353
transform 1 0 18032 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0582_
timestamp 1606120353
transform 1 0 18032 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__or2_4  _0527_
timestamp 1606120353
transform 1 0 18584 0 -1 16864
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_27_191
timestamp 1606120353
transform 1 0 18676 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1606120353
transform 1 0 19228 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__A1
timestamp 1606120353
transform 1 0 18860 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0490_
timestamp 1606120353
transform 1 0 19044 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_27_198
timestamp 1606120353
transform 1 0 19320 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0490__A
timestamp 1606120353
transform 1 0 19504 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__A1
timestamp 1606120353
transform 1 0 19412 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_201
timestamp 1606120353
transform 1 0 19596 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__D
timestamp 1606120353
transform 1 0 19780 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__B1
timestamp 1606120353
transform 1 0 19872 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_202
timestamp 1606120353
transform 1 0 19688 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0528_
timestamp 1606120353
transform 1 0 20056 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_26_205
timestamp 1606120353
transform 1 0 19964 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A2
timestamp 1606120353
transform 1 0 20240 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1606120353
transform 1 0 20332 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_217
timestamp 1606120353
transform 1 0 21068 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_213
timestamp 1606120353
transform 1 0 20700 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1606120353
transform 1 0 20424 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__B1
timestamp 1606120353
transform 1 0 20884 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__B1
timestamp 1606120353
transform 1 0 20608 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__A1
timestamp 1606120353
transform 1 0 21252 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0528__A
timestamp 1606120353
transform 1 0 20516 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1606120353
transform 1 0 20792 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _0805_
timestamp 1606120353
transform 1 0 20884 0 -1 16864
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_26_229
timestamp 1606120353
transform 1 0 22172 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A1
timestamp 1606120353
transform 1 0 22356 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_242
timestamp 1606120353
transform 1 0 23368 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_238
timestamp 1606120353
transform 1 0 23000 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_234
timestamp 1606120353
transform 1 0 22632 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_233
timestamp 1606120353
transform 1 0 22540 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A2
timestamp 1606120353
transform 1 0 22724 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__A2
timestamp 1606120353
transform 1 0 23184 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__A1
timestamp 1606120353
transform 1 0 22816 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1080_
timestamp 1606120353
transform 1 0 21436 0 1 16864
box 0 -48 1196 592
use sky130_fd_sc_hd__o21a_4  _1079_
timestamp 1606120353
transform 1 0 22908 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_27_245
timestamp 1606120353
transform 1 0 23644 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_26_249
timestamp 1606120353
transform 1 0 24012 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__D
timestamp 1606120353
transform 1 0 24012 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__D
timestamp 1606120353
transform 1 0 24196 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1606120353
transform 1 0 23552 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0970_
timestamp 1606120353
transform 1 0 24196 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_27_259
timestamp 1606120353
transform 1 0 24932 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_27_254
timestamp 1606120353
transform 1 0 24472 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1606120353
transform 1 0 24380 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__A
timestamp 1606120353
transform 1 0 24748 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__C
timestamp 1606120353
transform 1 0 24564 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _1005_
timestamp 1606120353
transform 1 0 24748 0 -1 16864
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A
timestamp 1606120353
transform 1 0 25300 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_265
timestamp 1606120353
transform 1 0 25484 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_271
timestamp 1606120353
transform 1 0 26036 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_26_266
timestamp 1606120353
transform 1 0 25576 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__C
timestamp 1606120353
transform 1 0 26220 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__B
timestamp 1606120353
transform 1 0 25852 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__C
timestamp 1606120353
transform 1 0 25668 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0982_
timestamp 1606120353
transform 1 0 25852 0 1 16864
box 0 -48 828 592
use sky130_fd_sc_hd__decap_4  FILLER_27_282
timestamp 1606120353
transform 1 0 27048 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1606120353
transform 1 0 26680 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__C
timestamp 1606120353
transform 1 0 26864 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1606120353
transform 1 0 26404 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__or4_4  _0973_
timestamp 1606120353
transform 1 0 26496 0 -1 16864
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILLER_26_285
timestamp 1606120353
transform 1 0 27324 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__B
timestamp 1606120353
transform 1 0 27416 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_26_294
timestamp 1606120353
transform 1 0 28152 0 -1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_26_290
timestamp 1606120353
transform 1 0 27784 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__C
timestamp 1606120353
transform 1 0 27600 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__B
timestamp 1606120353
transform 1 0 27968 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _1074_
timestamp 1606120353
transform 1 0 27600 0 1 16864
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_27_301
timestamp 1606120353
transform 1 0 28796 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_297
timestamp 1606120353
transform 1 0 28428 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_26_298
timestamp 1606120353
transform 1 0 28520 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__D
timestamp 1606120353
transform 1 0 28612 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A
timestamp 1606120353
transform 1 0 28980 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__C
timestamp 1606120353
transform 1 0 28612 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _1055_
timestamp 1606120353
transform 1 0 28796 0 -1 16864
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1606120353
transform 1 0 29164 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _1045_
timestamp 1606120353
transform 1 0 29256 0 1 16864
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_27_319
timestamp 1606120353
transform 1 0 30452 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_315
timestamp 1606120353
transform 1 0 30084 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_318
timestamp 1606120353
transform 1 0 30360 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_314
timestamp 1606120353
transform 1 0 29992 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_310
timestamp 1606120353
transform 1 0 29624 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__B
timestamp 1606120353
transform 1 0 30176 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A
timestamp 1606120353
transform 1 0 30268 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__C
timestamp 1606120353
transform 1 0 29808 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_27_323
timestamp 1606120353
transform 1 0 30820 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_26_329
timestamp 1606120353
transform 1 0 31372 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_325
timestamp 1606120353
transform 1 0 31004 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__B
timestamp 1606120353
transform 1 0 30544 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A2
timestamp 1606120353
transform 1 0 31188 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A
timestamp 1606120353
transform 1 0 30636 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0974_
timestamp 1606120353
transform 1 0 30728 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__o21a_4  _1019_
timestamp 1606120353
transform 1 0 31096 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_27_338
timestamp 1606120353
transform 1 0 32200 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_26_341
timestamp 1606120353
transform 1 0 32476 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_26_337
timestamp 1606120353
transform 1 0 32108 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_26_333
timestamp 1606120353
transform 1 0 31740 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__A
timestamp 1606120353
transform 1 0 31556 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A1
timestamp 1606120353
transform 1 0 32292 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A1
timestamp 1606120353
transform 1 0 32476 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1606120353
transform 1 0 32016 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_27_343
timestamp 1606120353
transform 1 0 32660 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__B1
timestamp 1606120353
transform 1 0 32752 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _1012_
timestamp 1606120353
transform 1 0 32936 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__o21ai_4  _0990_
timestamp 1606120353
transform 1 0 32936 0 -1 16864
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_27_362
timestamp 1606120353
transform 1 0 34408 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_358
timestamp 1606120353
transform 1 0 34040 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_26_359
timestamp 1606120353
transform 1 0 34132 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A2
timestamp 1606120353
transform 1 0 34408 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A2
timestamp 1606120353
transform 1 0 34224 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_367
timestamp 1606120353
transform 1 0 34868 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_364
timestamp 1606120353
transform 1 0 34592 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__B1
timestamp 1606120353
transform 1 0 34776 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A1
timestamp 1606120353
transform 1 0 35052 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A1
timestamp 1606120353
transform 1 0 34592 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1606120353
transform 1 0 34776 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_27_371
timestamp 1606120353
transform 1 0 35236 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_26_368
timestamp 1606120353
transform 1 0 34960 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_26_380
timestamp 1606120353
transform 1 0 36064 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_26_392
timestamp 1606120353
transform 1 0 37168 0 -1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_26_396
timestamp 1606120353
transform 1 0 37536 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_27_383
timestamp 1606120353
transform 1 0 36340 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_27_395
timestamp 1606120353
transform 1 0 37444 0 1 16864
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606120353
transform -1 0 38548 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606120353
transform -1 0 38548 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1606120353
transform 1 0 37628 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_26_398
timestamp 1606120353
transform 1 0 37720 0 -1 16864
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_27_403
timestamp 1606120353
transform 1 0 38180 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _0811_
timestamp 1606120353
transform 1 0 1932 0 -1 17952
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606120353
transform 1 0 1104 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__CLK
timestamp 1606120353
transform 1 0 1748 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1606120353
transform 1 0 1380 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__nor3_4  _0636_
timestamp 1606120353
transform 1 0 5060 0 -1 17952
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1606120353
transform 1 0 3956 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__C
timestamp 1606120353
transform 1 0 4876 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__B
timestamp 1606120353
transform 1 0 4508 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__A
timestamp 1606120353
transform 1 0 3772 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_28_23
timestamp 1606120353
transform 1 0 3220 0 -1 17952
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILLER_28_32
timestamp 1606120353
transform 1 0 4048 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_28_36
timestamp 1606120353
transform 1 0 4416 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_28_39
timestamp 1606120353
transform 1 0 4692 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0535_
timestamp 1606120353
transform 1 0 6992 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__B
timestamp 1606120353
transform 1 0 6808 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__C
timestamp 1606120353
transform 1 0 6440 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_56
timestamp 1606120353
transform 1 0 6256 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_60
timestamp 1606120353
transform 1 0 6624 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0705_
timestamp 1606120353
transform 1 0 8004 0 -1 17952
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__A
timestamp 1606120353
transform 1 0 7636 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__C
timestamp 1606120353
transform 1 0 9016 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_28_67
timestamp 1606120353
transform 1 0 7268 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_28_73
timestamp 1606120353
transform 1 0 7820 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_84
timestamp 1606120353
transform 1 0 8832 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_88
timestamp 1606120353
transform 1 0 9200 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__or3_4  _0597_
timestamp 1606120353
transform 1 0 9660 0 -1 17952
box 0 -48 828 592
use sky130_fd_sc_hd__and4_4  _0616_
timestamp 1606120353
transform 1 0 11224 0 -1 17952
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1606120353
transform 1 0 9568 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__C
timestamp 1606120353
transform 1 0 10672 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__A
timestamp 1606120353
transform 1 0 11040 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__C
timestamp 1606120353
transform 1 0 9384 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_102
timestamp 1606120353
transform 1 0 10488 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_106
timestamp 1606120353
transform 1 0 10856 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0595_
timestamp 1606120353
transform 1 0 13064 0 -1 17952
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__B
timestamp 1606120353
transform 1 0 12236 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__C
timestamp 1606120353
transform 1 0 12604 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_119
timestamp 1606120353
transform 1 0 12052 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_123
timestamp 1606120353
transform 1 0 12420 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_28_127
timestamp 1606120353
transform 1 0 12788 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1606120353
transform 1 0 15180 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0526__A
timestamp 1606120353
transform 1 0 14168 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0525__A
timestamp 1606120353
transform 1 0 14996 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__A
timestamp 1606120353
transform 1 0 14536 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_28_137
timestamp 1606120353
transform 1 0 13708 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_28_141
timestamp 1606120353
transform 1 0 14076 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_28_144
timestamp 1606120353
transform 1 0 14352 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_28_148
timestamp 1606120353
transform 1 0 14720 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_28_154
timestamp 1606120353
transform 1 0 15272 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__a2111oi_4  _0610_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 15824 0 -1 17952
box 0 -48 2024 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__A
timestamp 1606120353
transform 1 0 15456 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_158
timestamp 1606120353
transform 1 0 15640 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0489_
timestamp 1606120353
transform 1 0 18768 0 -1 17952
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__A1
timestamp 1606120353
transform 1 0 18032 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__A
timestamp 1606120353
transform 1 0 18400 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_182
timestamp 1606120353
transform 1 0 17848 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_186
timestamp 1606120353
transform 1 0 18216 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_190
timestamp 1606120353
transform 1 0 18584 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1606120353
transform 1 0 20792 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0581__B
timestamp 1606120353
transform 1 0 19780 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0489__A
timestamp 1606120353
transform 1 0 20148 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0555__A
timestamp 1606120353
transform 1 0 20516 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_201
timestamp 1606120353
transform 1 0 19596 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_205
timestamp 1606120353
transform 1 0 19964 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_209
timestamp 1606120353
transform 1 0 20332 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1606120353
transform 1 0 20700 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_28_215
timestamp 1606120353
transform 1 0 20884 0 -1 17952
box 0 -48 552 592
use sky130_fd_sc_hd__o21a_4  _1076_
timestamp 1606120353
transform 1 0 22540 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__B1
timestamp 1606120353
transform 1 0 22356 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__A2
timestamp 1606120353
transform 1 0 21436 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__B1
timestamp 1606120353
transform 1 0 21988 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_28_223
timestamp 1606120353
transform 1 0 21620 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_28_229
timestamp 1606120353
transform 1 0 22172 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _1067_
timestamp 1606120353
transform 1 0 24380 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A2
timestamp 1606120353
transform 1 0 24196 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A1
timestamp 1606120353
transform 1 0 23828 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_245
timestamp 1606120353
transform 1 0 23644 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_249
timestamp 1606120353
transform 1 0 24012 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_28_265
timestamp 1606120353
transform 1 0 25484 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_28_271
timestamp 1606120353
transform 1 0 26036 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__D
timestamp 1606120353
transform 1 0 25852 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__B
timestamp 1606120353
transform 1 0 26220 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1606120353
transform 1 0 26404 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0971_
timestamp 1606120353
transform 1 0 26496 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_28_279
timestamp 1606120353
transform 1 0 26772 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_283
timestamp 1606120353
transform 1 0 27140 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1606120353
transform 1 0 26956 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__C
timestamp 1606120353
transform 1 0 27324 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _1065_
timestamp 1606120353
transform 1 0 27968 0 -1 17952
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__C
timestamp 1606120353
transform 1 0 29256 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__D
timestamp 1606120353
transform 1 0 27692 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_287
timestamp 1606120353
transform 1 0 27508 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_28_291
timestamp 1606120353
transform 1 0 27876 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_28_301
timestamp 1606120353
transform 1 0 28796 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_28_305
timestamp 1606120353
transform 1 0 29164 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_28_308
timestamp 1606120353
transform 1 0 29440 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0983_
timestamp 1606120353
transform 1 0 29532 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_28_312
timestamp 1606120353
transform 1 0 29808 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__D
timestamp 1606120353
transform 1 0 29992 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_316
timestamp 1606120353
transform 1 0 30176 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_28_320
timestamp 1606120353
transform 1 0 30544 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__B
timestamp 1606120353
transform 1 0 30360 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0968_
timestamp 1606120353
transform 1 0 30636 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_28_324
timestamp 1606120353
transform 1 0 30912 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A1
timestamp 1606120353
transform 1 0 31096 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_328
timestamp 1606120353
transform 1 0 31280 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__B1
timestamp 1606120353
transform 1 0 31464 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1054_
timestamp 1606120353
transform 1 0 32476 0 -1 17952
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1606120353
transform 1 0 32016 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A2
timestamp 1606120353
transform 1 0 32292 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_28_332
timestamp 1606120353
transform 1 0 31648 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_28_337
timestamp 1606120353
transform 1 0 32108 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1013_
timestamp 1606120353
transform 1 0 34408 0 -1 17952
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_8  FILLER_28_354
timestamp 1606120353
transform 1 0 33672 0 -1 17952
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_28_375
timestamp 1606120353
transform 1 0 35604 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_28_387
timestamp 1606120353
transform 1 0 36708 0 -1 17952
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_28_395
timestamp 1606120353
transform 1 0 37444 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606120353
transform -1 0 38548 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1606120353
transform 1 0 37628 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_28_398
timestamp 1606120353
transform 1 0 37720 0 -1 17952
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606120353
transform 1 0 1104 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__D
timestamp 1606120353
transform 1 0 1564 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__CLK
timestamp 1606120353
transform 1 0 1932 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1606120353
transform 1 0 1380 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_7
timestamp 1606120353
transform 1 0 1748 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_29_11
timestamp 1606120353
transform 1 0 2116 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__D
timestamp 1606120353
transform 1 0 5152 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__C
timestamp 1606120353
transform 1 0 4784 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__D
timestamp 1606120353
transform 1 0 4416 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__D
timestamp 1606120353
transform 1 0 4048 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_29_23
timestamp 1606120353
transform 1 0 3220 0 1 17952
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_29_31
timestamp 1606120353
transform 1 0 3956 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_29_34
timestamp 1606120353
transform 1 0 4232 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_38
timestamp 1606120353
transform 1 0 4600 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_42
timestamp 1606120353
transform 1 0 4968 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1606120353
transform 1 0 5980 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_46
timestamp 1606120353
transform 1 0 5336 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0536__A
timestamp 1606120353
transform 1 0 5520 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0520_
timestamp 1606120353
transform 1 0 5704 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1606120353
transform 1 0 6808 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1606120353
transform 1 0 6348 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__A
timestamp 1606120353
transform 1 0 6532 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0520__A
timestamp 1606120353
transform 1 0 6164 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1606120353
transform 1 0 6716 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0514__A
timestamp 1606120353
transform 1 0 6992 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0686_
timestamp 1606120353
transform 1 0 7176 0 1 17952
box 0 -48 828 592
use sky130_fd_sc_hd__and4_4  _0724_
timestamp 1606120353
transform 1 0 8832 0 1 17952
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__A
timestamp 1606120353
transform 1 0 8648 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__B
timestamp 1606120353
transform 1 0 8280 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_29_75
timestamp 1606120353
transform 1 0 8004 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_29_80
timestamp 1606120353
transform 1 0 8464 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0617_
timestamp 1606120353
transform 1 0 10396 0 1 17952
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__B
timestamp 1606120353
transform 1 0 10028 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__A
timestamp 1606120353
transform 1 0 11224 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_29_93
timestamp 1606120353
transform 1 0 9660 0 1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_29_99
timestamp 1606120353
transform 1 0 10212 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_108
timestamp 1606120353
transform 1 0 11040 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1606120353
transform 1 0 12144 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_116
timestamp 1606120353
transform 1 0 11776 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_112
timestamp 1606120353
transform 1 0 11408 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__B
timestamp 1606120353
transform 1 0 11592 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__A
timestamp 1606120353
transform 1 0 11960 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_128
timestamp 1606120353
transform 1 0 12880 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_29_123
timestamp 1606120353
transform 1 0 12420 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__A2
timestamp 1606120353
transform 1 0 12696 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__C1
timestamp 1606120353
transform 1 0 13064 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1606120353
transform 1 0 12328 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__a2111oi_4  _0596_
timestamp 1606120353
transform 1 0 13248 0 1 17952
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_3  FILLER_29_154
timestamp 1606120353
transform 1 0 15272 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__and2_4  _0607_
timestamp 1606120353
transform 1 0 16560 0 1 17952
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__B
timestamp 1606120353
transform 1 0 16376 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A
timestamp 1606120353
transform 1 0 15916 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__B
timestamp 1606120353
transform 1 0 15548 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_159
timestamp 1606120353
transform 1 0 15732 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_29_163
timestamp 1606120353
transform 1 0 16100 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_29_175
timestamp 1606120353
transform 1 0 17204 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0529_
timestamp 1606120353
transform 1 0 18032 0 1 17952
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1606120353
transform 1 0 17940 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0529__A
timestamp 1606120353
transform 1 0 17756 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__B
timestamp 1606120353
transform 1 0 17388 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0630__A
timestamp 1606120353
transform 1 0 19044 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_179
timestamp 1606120353
transform 1 0 17572 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_193
timestamp 1606120353
transform 1 0 18860 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_29_197
timestamp 1606120353
transform 1 0 19228 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1102_
timestamp 1606120353
transform 1 0 19688 0 1 17952
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__D
timestamp 1606120353
transform 1 0 19504 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1070_
timestamp 1606120353
transform 1 0 22356 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A1
timestamp 1606120353
transform 1 0 23092 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A
timestamp 1606120353
transform 1 0 22172 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_29_221
timestamp 1606120353
transform 1 0 21436 0 1 17952
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_29_234
timestamp 1606120353
transform 1 0 22632 0 1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_29_238
timestamp 1606120353
transform 1 0 23000 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_29_241
timestamp 1606120353
transform 1 0 23276 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_29_253
timestamp 1606120353
transform 1 0 24380 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_29_249
timestamp 1606120353
transform 1 0 24012 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_29_245
timestamp 1606120353
transform 1 0 23644 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A2
timestamp 1606120353
transform 1 0 23828 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1606120353
transform 1 0 23552 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _1006_
timestamp 1606120353
transform 1 0 24104 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_29_257
timestamp 1606120353
transform 1 0 24748 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A
timestamp 1606120353
transform 1 0 24564 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__A1
timestamp 1606120353
transform 1 0 24932 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1063_
timestamp 1606120353
transform 1 0 25116 0 1 17952
box 0 -48 1196 592
use sky130_fd_sc_hd__and4_4  _1064_
timestamp 1606120353
transform 1 0 27324 0 1 17952
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__D
timestamp 1606120353
transform 1 0 27140 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A
timestamp 1606120353
transform 1 0 26772 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_29_274
timestamp 1606120353
transform 1 0 26312 0 1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_29_278
timestamp 1606120353
transform 1 0 26680 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1606120353
transform 1 0 26956 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0944_
timestamp 1606120353
transform 1 0 29256 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1606120353
transform 1 0 29164 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A
timestamp 1606120353
transform 1 0 28336 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__C
timestamp 1606120353
transform 1 0 28704 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_294
timestamp 1606120353
transform 1 0 28152 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_298
timestamp 1606120353
transform 1 0 28520 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_29_302
timestamp 1606120353
transform 1 0 28888 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _0993_
timestamp 1606120353
transform 1 0 31188 0 1 17952
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__A
timestamp 1606120353
transform 1 0 29716 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A1
timestamp 1606120353
transform 1 0 31004 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__B1
timestamp 1606120353
transform 1 0 30636 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__A
timestamp 1606120353
transform 1 0 30084 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_309
timestamp 1606120353
transform 1 0 29532 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_313
timestamp 1606120353
transform 1 0 29900 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_29_317
timestamp 1606120353
transform 1 0 30268 0 1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_29_323
timestamp 1606120353
transform 1 0 30820 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A1
timestamp 1606120353
transform 1 0 32936 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__B1
timestamp 1606120353
transform 1 0 33304 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__B1
timestamp 1606120353
transform 1 0 32568 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_340
timestamp 1606120353
transform 1 0 32384 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_344
timestamp 1606120353
transform 1 0 32752 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_348
timestamp 1606120353
transform 1 0 33120 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_352
timestamp 1606120353
transform 1 0 33488 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1606120353
transform 1 0 34776 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A2
timestamp 1606120353
transform 1 0 33672 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_29_356
timestamp 1606120353
transform 1 0 33856 0 1 17952
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_29_364
timestamp 1606120353
transform 1 0 34592 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_29_367
timestamp 1606120353
transform 1 0 34868 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_29_379
timestamp 1606120353
transform 1 0 35972 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_29_391
timestamp 1606120353
transform 1 0 37076 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606120353
transform -1 0 38548 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_29_403
timestamp 1606120353
transform 1 0 38180 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1216_
timestamp 1606120353
transform 1 0 1380 0 -1 19040
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606120353
transform 1 0 1104 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_30_22
timestamp 1606120353
transform 1 0 3128 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__D
timestamp 1606120353
transform 1 0 3404 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1606120353
transform 1 0 3588 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__D
timestamp 1606120353
transform 1 0 3772 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_30_32
timestamp 1606120353
transform 1 0 4048 0 -1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1606120353
transform 1 0 3956 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_30_38
timestamp 1606120353
transform 1 0 4600 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__D
timestamp 1606120353
transform 1 0 4416 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_42
timestamp 1606120353
transform 1 0 4968 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__C
timestamp 1606120353
transform 1 0 4784 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__A
timestamp 1606120353
transform 1 0 5152 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0514_
timestamp 1606120353
transform 1 0 6624 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0536_
timestamp 1606120353
transform 1 0 5612 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__A
timestamp 1606120353
transform 1 0 6072 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__B
timestamp 1606120353
transform 1 0 6440 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_30_46
timestamp 1606120353
transform 1 0 5336 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_30_52
timestamp 1606120353
transform 1 0 5888 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_56
timestamp 1606120353
transform 1 0 6256 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_30_63
timestamp 1606120353
transform 1 0 6900 0 -1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__and3_4  _0689_
timestamp 1606120353
transform 1 0 7636 0 -1 19040
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__B
timestamp 1606120353
transform 1 0 9108 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__C
timestamp 1606120353
transform 1 0 7268 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__B
timestamp 1606120353
transform 1 0 8648 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_69
timestamp 1606120353
transform 1 0 7452 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_80
timestamp 1606120353
transform 1 0 8464 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_30_84
timestamp 1606120353
transform 1 0 8832 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__and4_4  _0742_
timestamp 1606120353
transform 1 0 10028 0 -1 19040
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1606120353
transform 1 0 9568 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__A
timestamp 1606120353
transform 1 0 11040 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__C
timestamp 1606120353
transform 1 0 9844 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_30_89
timestamp 1606120353
transform 1 0 9292 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1606120353
transform 1 0 9660 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_106
timestamp 1606120353
transform 1 0 10856 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_30_110
timestamp 1606120353
transform 1 0 11224 0 -1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__nor3_4  _0635_
timestamp 1606120353
transform 1 0 11960 0 -1 19040
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__B1
timestamp 1606120353
transform 1 0 11592 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_116
timestamp 1606120353
transform 1 0 11776 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_131
timestamp 1606120353
transform 1 0 13156 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_135
timestamp 1606120353
transform 1 0 13524 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__B1
timestamp 1606120353
transform 1 0 13340 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__D1
timestamp 1606120353
transform 1 0 13708 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_30_139
timestamp 1606120353
transform 1 0 13892 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0526_
timestamp 1606120353
transform 1 0 14168 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_30_145
timestamp 1606120353
transform 1 0 14444 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__C
timestamp 1606120353
transform 1 0 14628 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_149
timestamp 1606120353
transform 1 0 14812 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A2
timestamp 1606120353
transform 1 0 14996 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1606120353
transform 1 0 15180 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_30_154
timestamp 1606120353
transform 1 0 15272 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0609_
timestamp 1606120353
transform 1 0 17296 0 -1 19040
box 0 -48 644 592
use sky130_fd_sc_hd__or2_4  _0688_
timestamp 1606120353
transform 1 0 15916 0 -1 19040
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__A1_N
timestamp 1606120353
transform 1 0 16744 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__B1
timestamp 1606120353
transform 1 0 17112 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__D
timestamp 1606120353
transform 1 0 15456 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_30_158
timestamp 1606120353
transform 1 0 15640 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_30_168
timestamp 1606120353
transform 1 0 16560 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_172
timestamp 1606120353
transform 1 0 16928 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0630_
timestamp 1606120353
transform 1 0 18676 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__A
timestamp 1606120353
transform 1 0 18124 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__A
timestamp 1606120353
transform 1 0 18492 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_183
timestamp 1606120353
transform 1 0 17940 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_187
timestamp 1606120353
transform 1 0 18308 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_30_194
timestamp 1606120353
transform 1 0 18952 0 -1 19040
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1606120353
transform 1 0 20792 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__CLK
timestamp 1606120353
transform 1 0 19688 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_30_204
timestamp 1606120353
transform 1 0 19872 0 -1 19040
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1606120353
transform 1 0 20608 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1606120353
transform 1 0 20884 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__o21ai_4  _1068_
timestamp 1606120353
transform 1 0 23092 0 -1 19040
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__B1
timestamp 1606120353
transform 1 0 22908 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A
timestamp 1606120353
transform 1 0 22540 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_30_227
timestamp 1606120353
transform 1 0 21988 0 -1 19040
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_30_235
timestamp 1606120353
transform 1 0 22724 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1022_
timestamp 1606120353
transform 1 0 25116 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__A
timestamp 1606120353
transform 1 0 24472 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__B1
timestamp 1606120353
transform 1 0 24932 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_252
timestamp 1606120353
transform 1 0 24288 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_30_256
timestamp 1606120353
transform 1 0 24656 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_30_264
timestamp 1606120353
transform 1 0 25392 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0992_
timestamp 1606120353
transform 1 0 26772 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1606120353
transform 1 0 26404 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__A
timestamp 1606120353
transform 1 0 27324 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A
timestamp 1606120353
transform 1 0 25576 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__A2
timestamp 1606120353
transform 1 0 25944 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_268
timestamp 1606120353
transform 1 0 25760 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_30_272
timestamp 1606120353
transform 1 0 26128 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_30_276
timestamp 1606120353
transform 1 0 26496 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_30_282
timestamp 1606120353
transform 1 0 27048 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__nor3_4  _1075_
timestamp 1606120353
transform 1 0 28152 0 -1 19040
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__B
timestamp 1606120353
transform 1 0 27692 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_287
timestamp 1606120353
transform 1 0 27508 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_30_291
timestamp 1606120353
transform 1 0 27876 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_30_307
timestamp 1606120353
transform 1 0 29348 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__B
timestamp 1606120353
transform 1 0 29532 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_311
timestamp 1606120353
transform 1 0 29716 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__B
timestamp 1606120353
transform 1 0 29900 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_315
timestamp 1606120353
transform 1 0 30084 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__C
timestamp 1606120353
transform 1 0 30268 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_319
timestamp 1606120353
transform 1 0 30452 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A
timestamp 1606120353
transform 1 0 30636 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_323
timestamp 1606120353
transform 1 0 30820 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A2
timestamp 1606120353
transform 1 0 31004 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_327
timestamp 1606120353
transform 1 0 31188 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A2
timestamp 1606120353
transform 1 0 31372 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0980_
timestamp 1606120353
transform 1 0 32936 0 -1 19040
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1606120353
transform 1 0 32016 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__B1
timestamp 1606120353
transform 1 0 32752 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_30_331
timestamp 1606120353
transform 1 0 31556 0 -1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_30_335
timestamp 1606120353
transform 1 0 31924 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_30_337
timestamp 1606120353
transform 1 0 32108 0 -1 19040
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_30_343
timestamp 1606120353
transform 1 0 32660 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_30_359
timestamp 1606120353
transform 1 0 34132 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_30_371
timestamp 1606120353
transform 1 0 35236 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_30_383
timestamp 1606120353
transform 1 0 36340 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_30_395
timestamp 1606120353
transform 1 0 37444 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606120353
transform -1 0 38548 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1606120353
transform 1 0 37628 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_30_398
timestamp 1606120353
transform 1 0 37720 0 -1 19040
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1105_
timestamp 1606120353
transform 1 0 2300 0 1 19040
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606120353
transform 1 0 1104 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__D
timestamp 1606120353
transform 1 0 2116 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__CLK
timestamp 1606120353
transform 1 0 1748 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1606120353
transform 1 0 1380 0 1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_31_9
timestamp 1606120353
transform 1 0 1932 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0544_
timestamp 1606120353
transform 1 0 5152 0 1 19040
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__B
timestamp 1606120353
transform 1 0 4968 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__A
timestamp 1606120353
transform 1 0 4600 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__D
timestamp 1606120353
transform 1 0 4232 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_32
timestamp 1606120353
transform 1 0 4048 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_36
timestamp 1606120353
transform 1 0 4416 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_40
timestamp 1606120353
transform 1 0 4784 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0542_
timestamp 1606120353
transform 1 0 6808 0 1 19040
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1606120353
transform 1 0 6716 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__B
timestamp 1606120353
transform 1 0 6532 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__A
timestamp 1606120353
transform 1 0 6164 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_53
timestamp 1606120353
transform 1 0 5980 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1606120353
transform 1 0 6348 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0741_
timestamp 1606120353
transform 1 0 9108 0 1 19040
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A
timestamp 1606120353
transform 1 0 8924 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__B
timestamp 1606120353
transform 1 0 7820 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__A
timestamp 1606120353
transform 1 0 8188 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__C
timestamp 1606120353
transform 1 0 8556 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_71
timestamp 1606120353
transform 1 0 7636 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_75
timestamp 1606120353
transform 1 0 8004 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_79
timestamp 1606120353
transform 1 0 8372 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_83
timestamp 1606120353
transform 1 0 8740 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0725_
timestamp 1606120353
transform 1 0 10764 0 1 19040
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__B
timestamp 1606120353
transform 1 0 10580 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__B
timestamp 1606120353
transform 1 0 10120 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_96
timestamp 1606120353
transform 1 0 9936 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_31_100
timestamp 1606120353
transform 1 0 10304 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__and2_4  _0634_
timestamp 1606120353
transform 1 0 12788 0 1 19040
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1606120353
transform 1 0 12328 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__A1
timestamp 1606120353
transform 1 0 11776 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__A2
timestamp 1606120353
transform 1 0 12144 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__B
timestamp 1606120353
transform 1 0 12604 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_114
timestamp 1606120353
transform 1 0 11592 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1606120353
transform 1 0 11960 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_123
timestamp 1606120353
transform 1 0 12420 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0532_
timestamp 1606120353
transform 1 0 14168 0 1 19040
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0532__B
timestamp 1606120353
transform 1 0 14996 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__B
timestamp 1606120353
transform 1 0 13800 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_31_134
timestamp 1606120353
transform 1 0 13432 0 1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_31_140
timestamp 1606120353
transform 1 0 13984 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_149
timestamp 1606120353
transform 1 0 14812 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_153
timestamp 1606120353
transform 1 0 15180 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0766_
timestamp 1606120353
transform 1 0 16100 0 1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__A1
timestamp 1606120353
transform 1 0 15916 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__B
timestamp 1606120353
transform 1 0 15364 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_31_157
timestamp 1606120353
transform 1 0 15548 0 1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_31_175
timestamp 1606120353
transform 1 0 17204 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1606120353
transform 1 0 17940 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__A2_N
timestamp 1606120353
transform 1 0 17388 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__B2
timestamp 1606120353
transform 1 0 17756 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__A
timestamp 1606120353
transform 1 0 18216 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__A
timestamp 1606120353
transform 1 0 18584 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_179
timestamp 1606120353
transform 1 0 17572 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_184
timestamp 1606120353
transform 1 0 18032 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_188
timestamp 1606120353
transform 1 0 18400 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_31_192
timestamp 1606120353
transform 1 0 18768 0 1 19040
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1207_
timestamp 1606120353
transform 1 0 19688 0 1 19040
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__D
timestamp 1606120353
transform 1 0 19504 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1606120353
transform 1 0 21436 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A1
timestamp 1606120353
transform 1 0 21620 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1606120353
transform 1 0 21804 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A2
timestamp 1606120353
transform 1 0 21988 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_229
timestamp 1606120353
transform 1 0 22172 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__B1
timestamp 1606120353
transform 1 0 22356 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_31_233
timestamp 1606120353
transform 1 0 22540 0 1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_31_240
timestamp 1606120353
transform 1 0 23184 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_31_237
timestamp 1606120353
transform 1 0 22908 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__B1
timestamp 1606120353
transform 1 0 23000 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A2
timestamp 1606120353
transform 1 0 23368 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_31_249
timestamp 1606120353
transform 1 0 24012 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_31_245
timestamp 1606120353
transform 1 0 23644 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A1
timestamp 1606120353
transform 1 0 23828 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1606120353
transform 1 0 23552 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _1059_
timestamp 1606120353
transform 1 0 24288 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_31_259
timestamp 1606120353
transform 1 0 24932 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_255
timestamp 1606120353
transform 1 0 24564 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__A
timestamp 1606120353
transform 1 0 24748 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A1
timestamp 1606120353
transform 1 0 25116 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1062_
timestamp 1606120353
transform 1 0 25300 0 1 19040
box 0 -48 1196 592
use sky130_fd_sc_hd__nor3_4  _1066_
timestamp 1606120353
transform 1 0 27232 0 1 19040
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A
timestamp 1606120353
transform 1 0 27048 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__C
timestamp 1606120353
transform 1 0 26680 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_276
timestamp 1606120353
transform 1 0 26496 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_280
timestamp 1606120353
transform 1 0 26864 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _1046_
timestamp 1606120353
transform 1 0 29256 0 1 19040
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1606120353
transform 1 0 29164 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__C
timestamp 1606120353
transform 1 0 28980 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__A
timestamp 1606120353
transform 1 0 28612 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_297
timestamp 1606120353
transform 1 0 28428 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_301
timestamp 1606120353
transform 1 0 28796 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0976_
timestamp 1606120353
transform 1 0 31004 0 1 19040
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A1
timestamp 1606120353
transform 1 0 30820 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__A
timestamp 1606120353
transform 1 0 30268 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_315
timestamp 1606120353
transform 1 0 30084 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_31_319
timestamp 1606120353
transform 1 0 30452 0 1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__o21a_4  _1052_
timestamp 1606120353
transform 1 0 32936 0 1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A1
timestamp 1606120353
transform 1 0 32752 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A2
timestamp 1606120353
transform 1 0 32384 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_338
timestamp 1606120353
transform 1 0 32200 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_342
timestamp 1606120353
transform 1 0 32568 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1606120353
transform 1 0 34776 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__A2
timestamp 1606120353
transform 1 0 35052 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A1
timestamp 1606120353
transform 1 0 34224 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__A1
timestamp 1606120353
transform 1 0 35420 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__B1
timestamp 1606120353
transform 1 0 34592 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_358
timestamp 1606120353
transform 1 0 34040 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_362
timestamp 1606120353
transform 1 0 34408 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_367
timestamp 1606120353
transform 1 0 34868 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_371
timestamp 1606120353
transform 1 0 35236 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__B1
timestamp 1606120353
transform 1 0 35788 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_375
timestamp 1606120353
transform 1 0 35604 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_31_379
timestamp 1606120353
transform 1 0 35972 0 1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_31_391
timestamp 1606120353
transform 1 0 37076 0 1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606120353
transform -1 0 38548 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_31_403
timestamp 1606120353
transform 1 0 38180 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1606120353
transform 1 0 1380 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606120353
transform 1 0 1104 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_32_7
timestamp 1606120353
transform 1 0 1748 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__D
timestamp 1606120353
transform 1 0 1564 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_32_11
timestamp 1606120353
transform 1 0 2116 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__CLK
timestamp 1606120353
transform 1 0 1932 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_16
timestamp 1606120353
transform 1 0 2576 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__B2
timestamp 1606120353
transform 1 0 2392 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_32_20
timestamp 1606120353
transform 1 0 2944 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__B1
timestamp 1606120353
transform 1 0 2760 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_32_24
timestamp 1606120353
transform 1 0 3312 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__D
timestamp 1606120353
transform 1 0 3404 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1606120353
transform 1 0 3588 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__D
timestamp 1606120353
transform 1 0 3772 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_32_32
timestamp 1606120353
transform 1 0 4048 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1606120353
transform 1 0 3956 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_32_36
timestamp 1606120353
transform 1 0 4416 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__D
timestamp 1606120353
transform 1 0 4508 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_42
timestamp 1606120353
transform 1 0 4968 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0680_
timestamp 1606120353
transform 1 0 4692 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__C
timestamp 1606120353
transform 1 0 5152 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__or3_4  _0545_
timestamp 1606120353
transform 1 0 5704 0 -1 20128
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__B
timestamp 1606120353
transform 1 0 7084 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__C
timestamp 1606120353
transform 1 0 6716 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__C
timestamp 1606120353
transform 1 0 5520 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_46
timestamp 1606120353
transform 1 0 5336 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_59
timestamp 1606120353
transform 1 0 6532 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_63
timestamp 1606120353
transform 1 0 6900 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0540_
timestamp 1606120353
transform 1 0 7268 0 -1 20128
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__B
timestamp 1606120353
transform 1 0 8740 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__C
timestamp 1606120353
transform 1 0 8280 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_76
timestamp 1606120353
transform 1 0 8096 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_32_80
timestamp 1606120353
transform 1 0 8464 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_32_85
timestamp 1606120353
transform 1 0 8924 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__or4_4  _0743_
timestamp 1606120353
transform 1 0 9936 0 -1 20128
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1606120353
transform 1 0 9568 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__A
timestamp 1606120353
transform 1 0 9384 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__C
timestamp 1606120353
transform 1 0 10948 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_32_89
timestamp 1606120353
transform 1 0 9292 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_32_93
timestamp 1606120353
transform 1 0 9660 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_32_105
timestamp 1606120353
transform 1 0 10764 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_109
timestamp 1606120353
transform 1 0 11132 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0537_
timestamp 1606120353
transform 1 0 11592 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__A
timestamp 1606120353
transform 1 0 11316 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__B1
timestamp 1606120353
transform 1 0 13156 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_32_113
timestamp 1606120353
transform 1 0 11500 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_32_126
timestamp 1606120353
transform 1 0 12696 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_32_130
timestamp 1606120353
transform 1 0 13064 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_32_137
timestamp 1606120353
transform 1 0 13708 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_32_133
timestamp 1606120353
transform 1 0 13340 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__B1
timestamp 1606120353
transform 1 0 13524 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0594_
timestamp 1606120353
transform 1 0 13800 0 -1 20128
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_32_145
timestamp 1606120353
transform 1 0 14444 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_149
timestamp 1606120353
transform 1 0 14812 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__A
timestamp 1606120353
transform 1 0 14996 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__D
timestamp 1606120353
transform 1 0 14628 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1606120353
transform 1 0 15180 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _0687_
timestamp 1606120353
transform 1 0 15272 0 -1 20128
box 0 -48 644 592
use sky130_fd_sc_hd__a2bb2o_4  _0765_
timestamp 1606120353
transform 1 0 16744 0 -1 20128
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__B1
timestamp 1606120353
transform 1 0 16100 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__A2
timestamp 1606120353
transform 1 0 16468 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_161
timestamp 1606120353
transform 1 0 15916 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_165
timestamp 1606120353
transform 1 0 16284 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_32_169
timestamp 1606120353
transform 1 0 16652 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0532__A
timestamp 1606120353
transform 1 0 18400 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__CLK
timestamp 1606120353
transform 1 0 19136 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_186
timestamp 1606120353
transform 1 0 18216 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_32_190
timestamp 1606120353
transform 1 0 18584 0 -1 20128
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILLER_32_198
timestamp 1606120353
transform 1 0 19320 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1606120353
transform 1 0 20792 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__CLK
timestamp 1606120353
transform 1 0 19688 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_32_204
timestamp 1606120353
transform 1 0 19872 0 -1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_32_212
timestamp 1606120353
transform 1 0 20608 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_32_215
timestamp 1606120353
transform 1 0 20884 0 -1 20128
box 0 -48 552 592
use sky130_fd_sc_hd__o21ai_4  _1077_
timestamp 1606120353
transform 1 0 21528 0 -1 20128
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_1  FILLER_32_221
timestamp 1606120353
transform 1 0 21436 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_32_235
timestamp 1606120353
transform 1 0 22724 0 -1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _1018_
timestamp 1606120353
transform 1 0 25392 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _1069_
timestamp 1606120353
transform 1 0 23460 0 -1 20128
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__B1
timestamp 1606120353
transform 1 0 25116 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_32_256
timestamp 1606120353
transform 1 0 24656 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_32_260
timestamp 1606120353
transform 1 0 25024 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_32_263
timestamp 1606120353
transform 1 0 25300 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_32_267
timestamp 1606120353
transform 1 0 25668 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A2
timestamp 1606120353
transform 1 0 25852 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_271
timestamp 1606120353
transform 1 0 26036 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__B1
timestamp 1606120353
transform 1 0 26220 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_276
timestamp 1606120353
transform 1 0 26496 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1606120353
transform 1 0 26404 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__C
timestamp 1606120353
transform 1 0 26680 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_280
timestamp 1606120353
transform 1 0 26864 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A1
timestamp 1606120353
transform 1 0 27048 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_32_284
timestamp 1606120353
transform 1 0 27232 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__nor3_4  _1048_
timestamp 1606120353
transform 1 0 29440 0 -1 20128
box 0 -48 1196 592
use sky130_fd_sc_hd__nor3_4  _1056_
timestamp 1606120353
transform 1 0 27508 0 -1 20128
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A1
timestamp 1606120353
transform 1 0 29256 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__B1
timestamp 1606120353
transform 1 0 28888 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_300
timestamp 1606120353
transform 1 0 28704 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_304
timestamp 1606120353
transform 1 0 29072 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__B1
timestamp 1606120353
transform 1 0 31004 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A2
timestamp 1606120353
transform 1 0 31372 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_32_321
timestamp 1606120353
transform 1 0 30636 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_32_327
timestamp 1606120353
transform 1 0 31188 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1053_
timestamp 1606120353
transform 1 0 33120 0 -1 20128
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1606120353
transform 1 0 32016 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A2
timestamp 1606120353
transform 1 0 32936 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__B1
timestamp 1606120353
transform 1 0 32292 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_32_331
timestamp 1606120353
transform 1 0 31556 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_32_335
timestamp 1606120353
transform 1 0 31924 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_32_337
timestamp 1606120353
transform 1 0 32108 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_32_341
timestamp 1606120353
transform 1 0 32476 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_32_345
timestamp 1606120353
transform 1 0 32844 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__o21a_4  _1049_
timestamp 1606120353
transform 1 0 35052 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_32_361
timestamp 1606120353
transform 1 0 34316 0 -1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_32_381
timestamp 1606120353
transform 1 0 36156 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_32_393
timestamp 1606120353
transform 1 0 37260 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606120353
transform -1 0 38548 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1606120353
transform 1 0 37628 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_32_398
timestamp 1606120353
transform 1 0 37720 0 -1 20128
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_34_3
timestamp 1606120353
transform 1 0 1380 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_33_10
timestamp 1606120353
transform 1 0 2024 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_33_7
timestamp 1606120353
transform 1 0 1748 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1606120353
transform 1 0 1380 0 1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A2
timestamp 1606120353
transform 1 0 1840 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1606120353
transform 1 0 1104 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1606120353
transform 1 0 1104 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A1
timestamp 1606120353
transform 1 0 2208 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1104_
timestamp 1606120353
transform 1 0 1472 0 -1 21216
box 0 -48 1748 592
use sky130_fd_sc_hd__o22a_4  _0810_
timestamp 1606120353
transform 1 0 2392 0 1 20128
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_34_32
timestamp 1606120353
transform 1 0 4048 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_34_23
timestamp 1606120353
transform 1 0 3220 0 -1 21216
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_33_32
timestamp 1606120353
transform 1 0 4048 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_28
timestamp 1606120353
transform 1 0 3680 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__C
timestamp 1606120353
transform 1 0 3772 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__D
timestamp 1606120353
transform 1 0 3864 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1606120353
transform 1 0 3956 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_34_36
timestamp 1606120353
transform 1 0 4416 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_43
timestamp 1606120353
transform 1 0 5060 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_39
timestamp 1606120353
transform 1 0 4692 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__D
timestamp 1606120353
transform 1 0 4232 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__D
timestamp 1606120353
transform 1 0 4600 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__B
timestamp 1606120353
transform 1 0 4232 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0491__A
timestamp 1606120353
transform 1 0 4876 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0491_
timestamp 1606120353
transform 1 0 4416 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__nor4_4  _0546_
timestamp 1606120353
transform 1 0 4784 0 -1 21216
box 0 -48 1564 592
use sky130_fd_sc_hd__fill_2  FILLER_33_50
timestamp 1606120353
transform 1 0 5704 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0511__A
timestamp 1606120353
transform 1 0 5888 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__A
timestamp 1606120353
transform 1 0 5244 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0511_
timestamp 1606120353
transform 1 0 5428 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_34_61
timestamp 1606120353
transform 1 0 6716 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_34_57
timestamp 1606120353
transform 1 0 6348 0 -1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_33_62
timestamp 1606120353
transform 1 0 6808 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_33_58
timestamp 1606120353
transform 1 0 6440 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_33_54
timestamp 1606120353
transform 1 0 6072 0 1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__B
timestamp 1606120353
transform 1 0 6808 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__B
timestamp 1606120353
transform 1 0 6532 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1606120353
transform 1 0 6716 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_34_64
timestamp 1606120353
transform 1 0 6992 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__A
timestamp 1606120353
transform 1 0 6992 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0738_
timestamp 1606120353
transform 1 0 7176 0 1 20128
box 0 -48 828 592
use sky130_fd_sc_hd__and4_4  _0682_
timestamp 1606120353
transform 1 0 7084 0 -1 21216
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_34_74
timestamp 1606120353
transform 1 0 7912 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_75
timestamp 1606120353
transform 1 0 8004 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_34_82
timestamp 1606120353
transform 1 0 8648 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_34_78
timestamp 1606120353
transform 1 0 8280 0 -1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_33_79
timestamp 1606120353
transform 1 0 8372 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A
timestamp 1606120353
transform 1 0 8096 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__D
timestamp 1606120353
transform 1 0 8740 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__C
timestamp 1606120353
transform 1 0 8188 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A
timestamp 1606120353
transform 1 0 8556 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0726_
timestamp 1606120353
transform 1 0 8740 0 1 20128
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1606120353
transform 1 0 8924 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__B
timestamp 1606120353
transform 1 0 9108 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_34_89
timestamp 1606120353
transform 1 0 9292 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_33_96
timestamp 1606120353
transform 1 0 9936 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_92
timestamp 1606120353
transform 1 0 9568 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__B
timestamp 1606120353
transform 1 0 9752 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1606120353
transform 1 0 9568 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0739_
timestamp 1606120353
transform 1 0 9660 0 -1 21216
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_34_106
timestamp 1606120353
transform 1 0 10856 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_102
timestamp 1606120353
transform 1 0 10488 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__C
timestamp 1606120353
transform 1 0 10672 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A
timestamp 1606120353
transform 1 0 10120 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0727_
timestamp 1606120353
transform 1 0 10304 0 1 20128
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_33_109
timestamp 1606120353
transform 1 0 11132 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__D
timestamp 1606120353
transform 1 0 11040 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0507_
timestamp 1606120353
transform 1 0 11224 0 -1 21216
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_34_119
timestamp 1606120353
transform 1 0 12052 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1606120353
transform 1 0 12236 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_33_117
timestamp 1606120353
transform 1 0 11868 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1606120353
transform 1 0 11500 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__D
timestamp 1606120353
transform 1 0 12236 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__B
timestamp 1606120353
transform 1 0 12052 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__D
timestamp 1606120353
transform 1 0 11684 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0507__A
timestamp 1606120353
transform 1 0 11316 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_34_127
timestamp 1606120353
transform 1 0 12788 0 -1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_34_123
timestamp 1606120353
transform 1 0 12420 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_127
timestamp 1606120353
transform 1 0 12788 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_123
timestamp 1606120353
transform 1 0 12420 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__A
timestamp 1606120353
transform 1 0 12604 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__C
timestamp 1606120353
transform 1 0 12604 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A1
timestamp 1606120353
transform 1 0 13156 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A1
timestamp 1606120353
transform 1 0 12972 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1606120353
transform 1 0 12328 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__a21o_4  _0751_
timestamp 1606120353
transform 1 0 13156 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_33_143
timestamp 1606120353
transform 1 0 14260 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A2
timestamp 1606120353
transform 1 0 14444 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_145
timestamp 1606120353
transform 1 0 14444 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A1
timestamp 1606120353
transform 1 0 14812 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__B
timestamp 1606120353
transform 1 0 14628 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_147
timestamp 1606120353
transform 1 0 14628 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_149
timestamp 1606120353
transform 1 0 14812 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__D
timestamp 1606120353
transform 1 0 14996 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_151
timestamp 1606120353
transform 1 0 14996 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0654_
timestamp 1606120353
transform 1 0 15272 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1606120353
transform 1 0 15180 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0654__A
timestamp 1606120353
transform 1 0 15180 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0752_
timestamp 1606120353
transform 1 0 13340 0 -1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_34_165
timestamp 1606120353
transform 1 0 16284 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_34_161
timestamp 1606120353
transform 1 0 15916 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_157
timestamp 1606120353
transform 1 0 15548 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__B2
timestamp 1606120353
transform 1 0 16100 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__B1
timestamp 1606120353
transform 1 0 15732 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_175
timestamp 1606120353
transform 1 0 17204 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_171
timestamp 1606120353
transform 1 0 16836 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_167
timestamp 1606120353
transform 1 0 16468 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__B1
timestamp 1606120353
transform 1 0 17020 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A2
timestamp 1606120353
transform 1 0 16652 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0758_
timestamp 1606120353
transform 1 0 15364 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__o22a_4  _0754_
timestamp 1606120353
transform 1 0 16560 0 -1 21216
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  FILLER_34_187
timestamp 1606120353
transform 1 0 18308 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_34_182
timestamp 1606120353
transform 1 0 17848 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_33_184
timestamp 1606120353
transform 1 0 18032 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_179
timestamp 1606120353
transform 1 0 17572 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A1
timestamp 1606120353
transform 1 0 18124 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A1
timestamp 1606120353
transform 1 0 18216 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A2
timestamp 1606120353
transform 1 0 17756 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__B2
timestamp 1606120353
transform 1 0 17388 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1606120353
transform 1 0 17940 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_33_192
timestamp 1606120353
transform 1 0 18768 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_188
timestamp 1606120353
transform 1 0 18400 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1606120353
transform 1 0 18584 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__D
timestamp 1606120353
transform 1 0 18952 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 18584 0 -1 21216
box 0 -48 1840 592
use sky130_fd_sc_hd__dfxtp_4  _1209_
timestamp 1606120353
transform 1 0 19136 0 1 20128
box 0 -48 1748 592
use sky130_fd_sc_hd__buf_1  _0695_
timestamp 1606120353
transform 1 0 20424 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1606120353
transform 1 0 20792 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A1
timestamp 1606120353
transform 1 0 21160 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__A
timestamp 1606120353
transform 1 0 21068 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1606120353
transform 1 0 20884 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_33_219
timestamp 1606120353
transform 1 0 21252 0 1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_34_213
timestamp 1606120353
transform 1 0 20700 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_34_215
timestamp 1606120353
transform 1 0 20884 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_34_220
timestamp 1606120353
transform 1 0 21344 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_34_224
timestamp 1606120353
transform 1 0 21712 0 -1 21216
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILLER_33_227
timestamp 1606120353
transform 1 0 21988 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0552__A
timestamp 1606120353
transform 1 0 21528 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A1
timestamp 1606120353
transform 1 0 22264 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_33_240
timestamp 1606120353
transform 1 0 23184 0 1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_33_236
timestamp 1606120353
transform 1 0 22816 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_232
timestamp 1606120353
transform 1 0 22448 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__B1
timestamp 1606120353
transform 1 0 23000 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A2
timestamp 1606120353
transform 1 0 22632 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1078_
timestamp 1606120353
transform 1 0 22264 0 -1 21216
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1606120353
transform 1 0 23552 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_34_243
timestamp 1606120353
transform 1 0 23460 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A2
timestamp 1606120353
transform 1 0 23644 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_245
timestamp 1606120353
transform 1 0 23644 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__B1
timestamp 1606120353
transform 1 0 23828 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_247
timestamp 1606120353
transform 1 0 23828 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__B1
timestamp 1606120353
transform 1 0 24012 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_249
timestamp 1606120353
transform 1 0 24012 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A1
timestamp 1606120353
transform 1 0 24196 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_253
timestamp 1606120353
transform 1 0 24380 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_34_263
timestamp 1606120353
transform 1 0 25300 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_33_257
timestamp 1606120353
transform 1 0 24748 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A2
timestamp 1606120353
transform 1 0 24564 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A1
timestamp 1606120353
transform 1 0 24932 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _1071_
timestamp 1606120353
transform 1 0 24196 0 -1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__o21ai_4  _1060_
timestamp 1606120353
transform 1 0 25116 0 1 20128
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_3  FILLER_34_272
timestamp 1606120353
transform 1 0 26128 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_34_268
timestamp 1606120353
transform 1 0 25760 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_274
timestamp 1606120353
transform 1 0 26312 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A2
timestamp 1606120353
transform 1 0 25944 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A2
timestamp 1606120353
transform 1 0 25576 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1606120353
transform 1 0 26404 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_34_284
timestamp 1606120353
transform 1 0 27232 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_34_279
timestamp 1606120353
transform 1 0 26772 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1606120353
transform 1 0 26680 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__B1
timestamp 1606120353
transform 1 0 27048 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__A
timestamp 1606120353
transform 1 0 26496 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A2
timestamp 1606120353
transform 1 0 26864 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1043_
timestamp 1606120353
transform 1 0 26496 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__o21a_4  _1061_
timestamp 1606120353
transform 1 0 27048 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_34_289
timestamp 1606120353
transform 1 0 27692 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_294
timestamp 1606120353
transform 1 0 28152 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__B
timestamp 1606120353
transform 1 0 27508 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A1
timestamp 1606120353
transform 1 0 27876 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A2
timestamp 1606120353
transform 1 0 28336 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 1606120353
transform 1 0 29256 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_33_302
timestamp 1606120353
transform 1 0 28888 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_33_298
timestamp 1606120353
transform 1 0 28520 0 1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__B1
timestamp 1606120353
transform 1 0 29440 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A2
timestamp 1606120353
transform 1 0 28980 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1606120353
transform 1 0 29164 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__o21ai_4  _1047_
timestamp 1606120353
transform 1 0 28060 0 -1 21216
box 0 -48 1196 592
use sky130_fd_sc_hd__o21ai_4  _0959_
timestamp 1606120353
transform 1 0 29256 0 1 20128
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_1  FILLER_34_314
timestamp 1606120353
transform 1 0 29992 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_34_310
timestamp 1606120353
transform 1 0 29624 0 -1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_33_319
timestamp 1606120353
transform 1 0 30452 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A2
timestamp 1606120353
transform 1 0 30084 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1044_
timestamp 1606120353
transform 1 0 30268 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_34_330
timestamp 1606120353
transform 1 0 31464 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_34_324
timestamp 1606120353
transform 1 0 30912 0 -1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_34_320
timestamp 1606120353
transform 1 0 30544 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_323
timestamp 1606120353
transform 1 0 30820 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__B1
timestamp 1606120353
transform 1 0 30728 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__B1
timestamp 1606120353
transform 1 0 31280 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A1
timestamp 1606120353
transform 1 0 31004 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__A
timestamp 1606120353
transform 1 0 30636 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1050_
timestamp 1606120353
transform 1 0 31188 0 1 20128
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_1  FILLER_34_337
timestamp 1606120353
transform 1 0 32108 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_34_334
timestamp 1606120353
transform 1 0 31832 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_340
timestamp 1606120353
transform 1 0 32384 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__B1
timestamp 1606120353
transform 1 0 31648 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1606120353
transform 1 0 32016 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_33_344
timestamp 1606120353
transform 1 0 32752 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A2
timestamp 1606120353
transform 1 0 32936 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A1
timestamp 1606120353
transform 1 0 32568 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_34_351
timestamp 1606120353
transform 1 0 33396 0 -1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_33_348
timestamp 1606120353
transform 1 0 33120 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__o21ai_4  _1051_
timestamp 1606120353
transform 1 0 32200 0 -1 21216
box 0 -48 1196 592
use sky130_fd_sc_hd__dfxtp_4  _1194_
timestamp 1606120353
transform 1 0 34868 0 -1 21216
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1606120353
transform 1 0 34776 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__D
timestamp 1606120353
transform 1 0 35052 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__CLK
timestamp 1606120353
transform 1 0 35420 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_33_360
timestamp 1606120353
transform 1 0 34224 0 1 20128
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_33_367
timestamp 1606120353
transform 1 0 34868 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_371
timestamp 1606120353
transform 1 0 35236 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_34_363
timestamp 1606120353
transform 1 0 34500 0 -1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_33_375
timestamp 1606120353
transform 1 0 35604 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_33_387
timestamp 1606120353
transform 1 0 36708 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_34_386
timestamp 1606120353
transform 1 0 36616 0 -1 21216
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_34_394
timestamp 1606120353
transform 1 0 37352 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1606120353
transform -1 0 38548 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1606120353
transform -1 0 38548 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1606120353
transform 1 0 37628 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_33_399
timestamp 1606120353
transform 1 0 37812 0 1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_33_403
timestamp 1606120353
transform 1 0 38180 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_34_398
timestamp 1606120353
transform 1 0 37720 0 -1 21216
box 0 -48 552 592
use sky130_fd_sc_hd__o22a_4  _0809_
timestamp 1606120353
transform 1 0 1932 0 1 21216
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1606120353
transform 1 0 1104 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A1
timestamp 1606120353
transform 1 0 1748 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1606120353
transform 1 0 1380 0 1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_35_23
timestamp 1606120353
transform 1 0 3220 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A2
timestamp 1606120353
transform 1 0 3404 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1606120353
transform 1 0 3588 0 1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_35_31
timestamp 1606120353
transform 1 0 3956 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A
timestamp 1606120353
transform 1 0 4048 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0808_
timestamp 1606120353
transform 1 0 4232 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_35_37
timestamp 1606120353
transform 1 0 4508 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_41
timestamp 1606120353
transform 1 0 4876 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0512__A
timestamp 1606120353
transform 1 0 4692 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__B
timestamp 1606120353
transform 1 0 5060 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_53
timestamp 1606120353
transform 1 0 5980 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_35_49
timestamp 1606120353
transform 1 0 5612 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_35_45
timestamp 1606120353
transform 1 0 5244 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__A
timestamp 1606120353
transform 1 0 5428 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0515_
timestamp 1606120353
transform 1 0 5704 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1606120353
transform 1 0 6348 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0515__A
timestamp 1606120353
transform 1 0 6164 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A
timestamp 1606120353
transform 1 0 6532 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1606120353
transform 1 0 6716 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0679_
timestamp 1606120353
transform 1 0 6808 0 1 21216
box 0 -48 828 592
use sky130_fd_sc_hd__buf_1  _0508_
timestamp 1606120353
transform 1 0 8556 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0508__A
timestamp 1606120353
transform 1 0 9016 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A
timestamp 1606120353
transform 1 0 7820 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__A
timestamp 1606120353
transform 1 0 8372 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_71
timestamp 1606120353
transform 1 0 7636 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_35_75
timestamp 1606120353
transform 1 0 8004 0 1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_35_84
timestamp 1606120353
transform 1 0 8832 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_88
timestamp 1606120353
transform 1 0 9200 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0510_
timestamp 1606120353
transform 1 0 11132 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__or4_4  _0744_
timestamp 1606120353
transform 1 0 9568 0 1 21216
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__B
timestamp 1606120353
transform 1 0 9384 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__A
timestamp 1606120353
transform 1 0 10580 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__D
timestamp 1606120353
transform 1 0 10948 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_101
timestamp 1606120353
transform 1 0 10396 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_105
timestamp 1606120353
transform 1 0 10764 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_112
timestamp 1606120353
transform 1 0 11408 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_116
timestamp 1606120353
transform 1 0 11776 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__B
timestamp 1606120353
transform 1 0 11592 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__C
timestamp 1606120353
transform 1 0 11960 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_120
timestamp 1606120353
transform 1 0 12144 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1606120353
transform 1 0 12328 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_35_123
timestamp 1606120353
transform 1 0 12420 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0506_
timestamp 1606120353
transform 1 0 12512 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_35_127
timestamp 1606120353
transform 1 0 12788 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_131
timestamp 1606120353
transform 1 0 13156 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0506__A
timestamp 1606120353
transform 1 0 12972 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0757_
timestamp 1606120353
transform 1 0 13524 0 1 21216
box 0 -48 644 592
use sky130_fd_sc_hd__o21a_4  _0759_
timestamp 1606120353
transform 1 0 14904 0 1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__B
timestamp 1606120353
transform 1 0 13340 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__B
timestamp 1606120353
transform 1 0 14352 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B1
timestamp 1606120353
transform 1 0 14720 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_142
timestamp 1606120353
transform 1 0 14168 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_146
timestamp 1606120353
transform 1 0 14536 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__A2
timestamp 1606120353
transform 1 0 16192 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A2
timestamp 1606120353
transform 1 0 16560 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__B1
timestamp 1606120353
transform 1 0 16928 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__A
timestamp 1606120353
transform 1 0 17296 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_162
timestamp 1606120353
transform 1 0 16008 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1606120353
transform 1 0 16376 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_170
timestamp 1606120353
transform 1 0 16744 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_174
timestamp 1606120353
transform 1 0 17112 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1121_
timestamp 1606120353
transform 1 0 18768 0 1 21216
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1606120353
transform 1 0 17940 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__D
timestamp 1606120353
transform 1 0 18584 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A2
timestamp 1606120353
transform 1 0 18216 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__B1
timestamp 1606120353
transform 1 0 17756 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_35_178
timestamp 1606120353
transform 1 0 17480 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_35_184
timestamp 1606120353
transform 1 0 18032 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_188
timestamp 1606120353
transform 1 0 18400 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0552_
timestamp 1606120353
transform 1 0 21252 0 1 21216
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__B1_N
timestamp 1606120353
transform 1 0 21068 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A2
timestamp 1606120353
transform 1 0 20700 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_211
timestamp 1606120353
transform 1 0 20516 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_215
timestamp 1606120353
transform 1 0 20884 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A1
timestamp 1606120353
transform 1 0 23368 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__A1
timestamp 1606120353
transform 1 0 23000 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__A2
timestamp 1606120353
transform 1 0 22632 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__B1
timestamp 1606120353
transform 1 0 22264 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_228
timestamp 1606120353
transform 1 0 22080 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_232
timestamp 1606120353
transform 1 0 22448 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1606120353
transform 1 0 22816 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1606120353
transform 1 0 23184 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1072_
timestamp 1606120353
transform 1 0 23644 0 1 21216
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1606120353
transform 1 0 23552 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A1
timestamp 1606120353
transform 1 0 25392 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_35_258
timestamp 1606120353
transform 1 0 24840 0 1 21216
box 0 -48 552 592
use sky130_fd_sc_hd__o21ai_4  _1058_
timestamp 1606120353
transform 1 0 25576 0 1 21216
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A2
timestamp 1606120353
transform 1 0 26956 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A1
timestamp 1606120353
transform 1 0 27324 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_279
timestamp 1606120353
transform 1 0 26772 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_283
timestamp 1606120353
transform 1 0 27140 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_287
timestamp 1606120353
transform 1 0 27508 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__B1
timestamp 1606120353
transform 1 0 27692 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_35_291
timestamp 1606120353
transform 1 0 27876 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0879_
timestamp 1606120353
transform 1 0 27968 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_35_295
timestamp 1606120353
transform 1 0 28244 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A
timestamp 1606120353
transform 1 0 28428 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_299
timestamp 1606120353
transform 1 0 28612 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A
timestamp 1606120353
transform 1 0 28796 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_303
timestamp 1606120353
transform 1 0 28980 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1606120353
transform 1 0 29164 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0984_
timestamp 1606120353
transform 1 0 29256 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_35_313
timestamp 1606120353
transform 1 0 29900 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_309
timestamp 1606120353
transform 1 0 29532 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A1
timestamp 1606120353
transform 1 0 30084 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A
timestamp 1606120353
transform 1 0 29716 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0998_
timestamp 1606120353
transform 1 0 30268 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_35_324
timestamp 1606120353
transform 1 0 30912 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_320
timestamp 1606120353
transform 1 0 30544 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A1
timestamp 1606120353
transform 1 0 31096 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A
timestamp 1606120353
transform 1 0 30728 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1023_
timestamp 1606120353
transform 1 0 31280 0 1 21216
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__D
timestamp 1606120353
transform 1 0 32660 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__CLK
timestamp 1606120353
transform 1 0 33028 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_341
timestamp 1606120353
transform 1 0 32476 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_345
timestamp 1606120353
transform 1 0 32844 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1606120353
transform 1 0 33212 0 1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1606120353
transform 1 0 34776 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__CLK
timestamp 1606120353
transform 1 0 35236 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_35_361
timestamp 1606120353
transform 1 0 34316 0 1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_35_365
timestamp 1606120353
transform 1 0 34684 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_35_367
timestamp 1606120353
transform 1 0 34868 0 1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_35_373
timestamp 1606120353
transform 1 0 35420 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1228_
timestamp 1606120353
transform 1 0 35788 0 1 21216
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__D
timestamp 1606120353
transform 1 0 35604 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_35_396
timestamp 1606120353
transform 1 0 37536 0 1 21216
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1606120353
transform -1 0 38548 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1606120353
transform 1 0 1380 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1606120353
transform 1 0 1104 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_36_7
timestamp 1606120353
transform 1 0 1748 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__B1
timestamp 1606120353
transform 1 0 1564 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_36_11
timestamp 1606120353
transform 1 0 2116 0 -1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__B2
timestamp 1606120353
transform 1 0 1932 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_36_15
timestamp 1606120353
transform 1 0 2484 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A1
timestamp 1606120353
transform 1 0 2576 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_18
timestamp 1606120353
transform 1 0 2760 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A2
timestamp 1606120353
transform 1 0 2944 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_36_22
timestamp 1606120353
transform 1 0 3128 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__D
timestamp 1606120353
transform 1 0 3404 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1606120353
transform 1 0 3588 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__D
timestamp 1606120353
transform 1 0 3772 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1606120353
transform 1 0 3956 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_36_32
timestamp 1606120353
transform 1 0 4048 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A1_N
timestamp 1606120353
transform 1 0 4232 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0512_
timestamp 1606120353
transform 1 0 4416 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_36_39
timestamp 1606120353
transform 1 0 4692 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_43
timestamp 1606120353
transform 1 0 5060 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__B1
timestamp 1606120353
transform 1 0 4876 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0521_
timestamp 1606120353
transform 1 0 5428 0 -1 22304
box 0 -48 828 592
use sky130_fd_sc_hd__or4_4  _0683_
timestamp 1606120353
transform 1 0 6992 0 -1 22304
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__C
timestamp 1606120353
transform 1 0 5244 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__C
timestamp 1606120353
transform 1 0 6808 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__A
timestamp 1606120353
transform 1 0 6440 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_56
timestamp 1606120353
transform 1 0 6256 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_60
timestamp 1606120353
transform 1 0 6624 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0652_
timestamp 1606120353
transform 1 0 8556 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A
timestamp 1606120353
transform 1 0 9016 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__A
timestamp 1606120353
transform 1 0 8004 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__D
timestamp 1606120353
transform 1 0 8372 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_73
timestamp 1606120353
transform 1 0 7820 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_77
timestamp 1606120353
transform 1 0 8188 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_84
timestamp 1606120353
transform 1 0 8832 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_88
timestamp 1606120353
transform 1 0 9200 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0722_
timestamp 1606120353
transform 1 0 9660 0 -1 22304
box 0 -48 828 592
use sky130_fd_sc_hd__or2_4  _0737_
timestamp 1606120353
transform 1 0 11224 0 -1 22304
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1606120353
transform 1 0 9568 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__C
timestamp 1606120353
transform 1 0 9384 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__C
timestamp 1606120353
transform 1 0 10672 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__A
timestamp 1606120353
transform 1 0 11040 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_102
timestamp 1606120353
transform 1 0 10488 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_106
timestamp 1606120353
transform 1 0 10856 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _0720_
timestamp 1606120353
transform 1 0 12604 0 -1 22304
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A2
timestamp 1606120353
transform 1 0 12420 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__B
timestamp 1606120353
transform 1 0 12052 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_117
timestamp 1606120353
transform 1 0 11868 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_121
timestamp 1606120353
transform 1 0 12236 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_36_132
timestamp 1606120353
transform 1 0 13248 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A
timestamp 1606120353
transform 1 0 13524 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_137
timestamp 1606120353
transform 1 0 13708 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__B
timestamp 1606120353
transform 1 0 13892 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1606120353
transform 1 0 14076 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A3
timestamp 1606120353
transform 1 0 14260 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_145
timestamp 1606120353
transform 1 0 14444 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__C
timestamp 1606120353
transform 1 0 14628 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_149
timestamp 1606120353
transform 1 0 14812 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A1
timestamp 1606120353
transform 1 0 14996 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_154
timestamp 1606120353
transform 1 0 15272 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1606120353
transform 1 0 15180 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _0768_
timestamp 1606120353
transform 1 0 16100 0 -1 22304
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A2
timestamp 1606120353
transform 1 0 15456 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__B1
timestamp 1606120353
transform 1 0 15824 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_158
timestamp 1606120353
transform 1 0 15640 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_36_162
timestamp 1606120353
transform 1 0 16008 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__o21a_4  _0753_
timestamp 1606120353
transform 1 0 18124 0 -1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__A1
timestamp 1606120353
transform 1 0 17572 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0510__A
timestamp 1606120353
transform 1 0 17940 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_177
timestamp 1606120353
transform 1 0 17388 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_181
timestamp 1606120353
transform 1 0 17756 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1606120353
transform 1 0 19228 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0929_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 21160 0 -1 22304
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1606120353
transform 1 0 20792 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__CLK
timestamp 1606120353
transform 1 0 20148 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__CLK
timestamp 1606120353
transform 1 0 19412 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_36_201
timestamp 1606120353
transform 1 0 19596 0 -1 22304
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILLER_36_209
timestamp 1606120353
transform 1 0 20332 0 -1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_36_213
timestamp 1606120353
transform 1 0 20700 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_36_215
timestamp 1606120353
transform 1 0 20884 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _1073_
timestamp 1606120353
transform 1 0 23092 0 -1 22304
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_8  FILLER_36_231
timestamp 1606120353
transform 1 0 22356 0 -1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_36_252
timestamp 1606120353
transform 1 0 24288 0 -1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1606120353
transform 1 0 25392 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _1057_
timestamp 1606120353
transform 1 0 26496 0 -1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1606120353
transform 1 0 26404 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__C
timestamp 1606120353
transform 1 0 26220 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__B1
timestamp 1606120353
transform 1 0 25576 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_36_268
timestamp 1606120353
transform 1 0 25760 0 -1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_36_272
timestamp 1606120353
transform 1 0 26128 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _0878_
timestamp 1606120353
transform 1 0 28336 0 -1 22304
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILLER_36_288
timestamp 1606120353
transform 1 0 27600 0 -1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_36_305
timestamp 1606120353
transform 1 0 29164 0 -1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__o21ai_4  _1020_
timestamp 1606120353
transform 1 0 30084 0 -1 22304
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A2
timestamp 1606120353
transform 1 0 31464 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_313
timestamp 1606120353
transform 1 0 29900 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_328
timestamp 1606120353
transform 1 0 31280 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1134_
timestamp 1606120353
transform 1 0 32660 0 -1 22304
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1606120353
transform 1 0 32016 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_36_332
timestamp 1606120353
transform 1 0 31648 0 -1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_36_337
timestamp 1606120353
transform 1 0 32108 0 -1 22304
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_36_362
timestamp 1606120353
transform 1 0 34408 0 -1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_36_374
timestamp 1606120353
transform 1 0 35512 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__CLK
timestamp 1606120353
transform 1 0 35788 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_36_379
timestamp 1606120353
transform 1 0 35972 0 -1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_36_391
timestamp 1606120353
transform 1 0 37076 0 -1 22304
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1606120353
transform -1 0 38548 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1606120353
transform 1 0 37628 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_36_398
timestamp 1606120353
transform 1 0 37720 0 -1 22304
box 0 -48 552 592
use sky130_fd_sc_hd__o22a_4  _0780_
timestamp 1606120353
transform 1 0 2576 0 1 22304
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1606120353
transform 1 0 1104 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__B1
timestamp 1606120353
transform 1 0 2392 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__B2
timestamp 1606120353
transform 1 0 2024 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__D
timestamp 1606120353
transform 1 0 1564 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1606120353
transform 1 0 1380 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_37_7
timestamp 1606120353
transform 1 0 1748 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_37_12
timestamp 1606120353
transform 1 0 2208 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0656_
timestamp 1606120353
transform 1 0 4876 0 1 22304
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__B2
timestamp 1606120353
transform 1 0 4048 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A2_N
timestamp 1606120353
transform 1 0 4416 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_30
timestamp 1606120353
transform 1 0 3864 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_34
timestamp 1606120353
transform 1 0 4232 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_37_38
timestamp 1606120353
transform 1 0 4600 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1606120353
transform 1 0 6716 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__D
timestamp 1606120353
transform 1 0 7084 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__B
timestamp 1606120353
transform 1 0 5704 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__C
timestamp 1606120353
transform 1 0 6256 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_48
timestamp 1606120353
transform 1 0 5520 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1606120353
transform 1 0 5888 0 1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_37_58
timestamp 1606120353
transform 1 0 6440 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_37_62
timestamp 1606120353
transform 1 0 6808 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__and4_4  _0681_
timestamp 1606120353
transform 1 0 7268 0 1 22304
box 0 -48 828 592
use sky130_fd_sc_hd__and4_4  _0740_
timestamp 1606120353
transform 1 0 8832 0 1 22304
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B
timestamp 1606120353
transform 1 0 8648 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__B
timestamp 1606120353
transform 1 0 8280 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_76
timestamp 1606120353
transform 1 0 8096 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_80
timestamp 1606120353
transform 1 0 8464 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0728_
timestamp 1606120353
transform 1 0 10396 0 1 22304
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__A
timestamp 1606120353
transform 1 0 9844 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__C
timestamp 1606120353
transform 1 0 10212 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_93
timestamp 1606120353
transform 1 0 9660 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_97
timestamp 1606120353
transform 1 0 10028 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1606120353
transform 1 0 11224 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_118
timestamp 1606120353
transform 1 0 11960 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_114
timestamp 1606120353
transform 1 0 11592 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__B
timestamp 1606120353
transform 1 0 11776 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A
timestamp 1606120353
transform 1 0 11408 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_127
timestamp 1606120353
transform 1 0 12788 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_123
timestamp 1606120353
transform 1 0 12420 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A1
timestamp 1606120353
transform 1 0 12144 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__A
timestamp 1606120353
transform 1 0 12604 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1606120353
transform 1 0 12328 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__C
timestamp 1606120353
transform 1 0 12972 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0718_
timestamp 1606120353
transform 1 0 13156 0 1 22304
box 0 -48 828 592
use sky130_fd_sc_hd__and2_4  _0717_
timestamp 1606120353
transform 1 0 14720 0 1 22304
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__A
timestamp 1606120353
transform 1 0 14536 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__B2
timestamp 1606120353
transform 1 0 14168 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_140
timestamp 1606120353
transform 1 0 13984 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_144
timestamp 1606120353
transform 1 0 14352 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0767_
timestamp 1606120353
transform 1 0 16100 0 1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A2
timestamp 1606120353
transform 1 0 15916 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__B
timestamp 1606120353
transform 1 0 15548 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_155
timestamp 1606120353
transform 1 0 15364 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_159
timestamp 1606120353
transform 1 0 15732 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_175
timestamp 1606120353
transform 1 0 17204 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_179
timestamp 1606120353
transform 1 0 17572 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__B1
timestamp 1606120353
transform 1 0 17388 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A1
timestamp 1606120353
transform 1 0 17756 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1606120353
transform 1 0 17940 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0801_
timestamp 1606120353
transform 1 0 18032 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_37_187
timestamp 1606120353
transform 1 0 18308 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_191
timestamp 1606120353
transform 1 0 18676 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__A
timestamp 1606120353
transform 1 0 18492 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A1
timestamp 1606120353
transform 1 0 18860 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_195
timestamp 1606120353
transform 1 0 19044 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__B1
timestamp 1606120353
transform 1 0 19228 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1099_
timestamp 1606120353
transform 1 0 20148 0 1 22304
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__D
timestamp 1606120353
transform 1 0 19964 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A2
timestamp 1606120353
transform 1 0 19596 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_199
timestamp 1606120353
transform 1 0 19412 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_203
timestamp 1606120353
transform 1 0 19780 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__D
timestamp 1606120353
transform 1 0 22448 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__CLK
timestamp 1606120353
transform 1 0 22816 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_37_226
timestamp 1606120353
transform 1 0 21896 0 1 22304
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_37_234
timestamp 1606120353
transform 1 0 22632 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_37_238
timestamp 1606120353
transform 1 0 23000 0 1 22304
box 0 -48 552 592
use sky130_fd_sc_hd__inv_8  _0840_
timestamp 1606120353
transform 1 0 24748 0 1 22304
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1606120353
transform 1 0 23552 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A
timestamp 1606120353
transform 1 0 24564 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_37_245
timestamp 1606120353
transform 1 0 23644 0 1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_37_253
timestamp 1606120353
transform 1 0 24380 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__or3_4  _0837_
timestamp 1606120353
transform 1 0 27048 0 1 22304
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__B
timestamp 1606120353
transform 1 0 26496 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__B
timestamp 1606120353
transform 1 0 26864 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__C
timestamp 1606120353
transform 1 0 26128 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__A
timestamp 1606120353
transform 1 0 25760 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_266
timestamp 1606120353
transform 1 0 25576 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_270
timestamp 1606120353
transform 1 0 25944 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_274
timestamp 1606120353
transform 1 0 26312 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1606120353
transform 1 0 26680 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0842_
timestamp 1606120353
transform 1 0 29256 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1606120353
transform 1 0 29164 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__B1
timestamp 1606120353
transform 1 0 28520 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A1
timestamp 1606120353
transform 1 0 28888 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A
timestamp 1606120353
transform 1 0 28060 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_291
timestamp 1606120353
transform 1 0 27876 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_37_295
timestamp 1606120353
transform 1 0 28244 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_37_300
timestamp 1606120353
transform 1 0 28704 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_37_304
timestamp 1606120353
transform 1 0 29072 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _0843_
timestamp 1606120353
transform 1 0 30268 0 1 22304
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A2
timestamp 1606120353
transform 1 0 29716 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__A
timestamp 1606120353
transform 1 0 30084 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_309
timestamp 1606120353
transform 1 0 29532 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_313
timestamp 1606120353
transform 1 0 29900 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_37_326
timestamp 1606120353
transform 1 0 31096 0 1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__B1_N
timestamp 1606120353
transform 1 0 32108 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A2
timestamp 1606120353
transform 1 0 32476 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A1
timestamp 1606120353
transform 1 0 32844 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_37_334
timestamp 1606120353
transform 1 0 31832 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_37_339
timestamp 1606120353
transform 1 0 32292 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_343
timestamp 1606120353
transform 1 0 32660 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_37_347
timestamp 1606120353
transform 1 0 33028 0 1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1606120353
transform 1 0 34776 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_37_359
timestamp 1606120353
transform 1 0 34132 0 1 22304
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_37_365
timestamp 1606120353
transform 1 0 34684 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_37_367
timestamp 1606120353
transform 1 0 34868 0 1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1189_
timestamp 1606120353
transform 1 0 35788 0 1 22304
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__D
timestamp 1606120353
transform 1 0 35604 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_37_396
timestamp 1606120353
transform 1 0 37536 0 1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1606120353
transform -1 0 38548 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1091_
timestamp 1606120353
transform 1 0 1472 0 -1 23392
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1606120353
transform 1 0 1104 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_38_3
timestamp 1606120353
transform 1 0 1380 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__a2bb2o_4  _0778_
timestamp 1606120353
transform 1 0 4048 0 -1 23392
box 0 -48 1472 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1606120353
transform 1 0 3956 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__D
timestamp 1606120353
transform 1 0 3772 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__D
timestamp 1606120353
transform 1 0 3404 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_23
timestamp 1606120353
transform 1 0 3220 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_27
timestamp 1606120353
transform 1 0 3588 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0675_
timestamp 1606120353
transform 1 0 6256 0 -1 23392
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__A
timestamp 1606120353
transform 1 0 5704 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__B
timestamp 1606120353
transform 1 0 6072 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_48
timestamp 1606120353
transform 1 0 5520 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_52
timestamp 1606120353
transform 1 0 5888 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_65
timestamp 1606120353
transform 1 0 7084 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0723_
timestamp 1606120353
transform 1 0 8004 0 -1 23392
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__B
timestamp 1606120353
transform 1 0 7268 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A
timestamp 1606120353
transform 1 0 7636 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__B
timestamp 1606120353
transform 1 0 9016 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_69
timestamp 1606120353
transform 1 0 7452 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_73
timestamp 1606120353
transform 1 0 7820 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_84
timestamp 1606120353
transform 1 0 8832 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_88
timestamp 1606120353
transform 1 0 9200 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__C
timestamp 1606120353
transform 1 0 9384 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1606120353
transform 1 0 9568 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0669_
timestamp 1606120353
transform 1 0 9660 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_38_96
timestamp 1606120353
transform 1 0 9936 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_100
timestamp 1606120353
transform 1 0 10304 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A2
timestamp 1606120353
transform 1 0 10120 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A3
timestamp 1606120353
transform 1 0 10488 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_104
timestamp 1606120353
transform 1 0 10672 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__B1
timestamp 1606120353
transform 1 0 10856 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_38_108
timestamp 1606120353
transform 1 0 11040 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__and3_4  _0729_
timestamp 1606120353
transform 1 0 11316 0 -1 23392
box 0 -48 828 592
use sky130_fd_sc_hd__a32o_4  _0731_
timestamp 1606120353
transform 1 0 12880 0 -1 23392
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__D
timestamp 1606120353
transform 1 0 12696 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__D
timestamp 1606120353
transform 1 0 12328 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_120
timestamp 1606120353
transform 1 0 12144 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_124
timestamp 1606120353
transform 1 0 12512 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1606120353
transform 1 0 15180 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__B2
timestamp 1606120353
transform 1 0 14996 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A2
timestamp 1606120353
transform 1 0 14628 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_145
timestamp 1606120353
transform 1 0 14444 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_149
timestamp 1606120353
transform 1 0 14812 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_38_154
timestamp 1606120353
transform 1 0 15272 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _0761_
timestamp 1606120353
transform 1 0 15364 0 -1 23392
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__B1
timestamp 1606120353
transform 1 0 16836 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A1
timestamp 1606120353
transform 1 0 17204 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_169
timestamp 1606120353
transform 1 0 16652 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_173
timestamp 1606120353
transform 1 0 17020 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0777_
timestamp 1606120353
transform 1 0 18400 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__D
timestamp 1606120353
transform 1 0 17572 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__CLK
timestamp 1606120353
transform 1 0 17940 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_177
timestamp 1606120353
transform 1 0 17388 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_181
timestamp 1606120353
transform 1 0 17756 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_38_185
timestamp 1606120353
transform 1 0 18124 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0487_
timestamp 1606120353
transform 1 0 20884 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1606120353
transform 1 0 20792 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__B2
timestamp 1606120353
transform 1 0 20516 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0487__A
timestamp 1606120353
transform 1 0 21344 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_38_200
timestamp 1606120353
transform 1 0 19504 0 -1 23392
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_38_208
timestamp 1606120353
transform 1 0 20240 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_38_213
timestamp 1606120353
transform 1 0 20700 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_38_218
timestamp 1606120353
transform 1 0 21160 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1157_
timestamp 1606120353
transform 1 0 22448 0 -1 23392
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_8  FILLER_38_222
timestamp 1606120353
transform 1 0 21528 0 -1 23392
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_38_230
timestamp 1606120353
transform 1 0 22264 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0825_
timestamp 1606120353
transform 1 0 25392 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_38_251
timestamp 1606120353
transform 1 0 24196 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_38_263
timestamp 1606120353
transform 1 0 25300 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__or4_4  _0943_
timestamp 1606120353
transform 1 0 26496 0 -1 23392
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1606120353
transform 1 0 26404 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__D
timestamp 1606120353
transform 1 0 26220 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A
timestamp 1606120353
transform 1 0 25852 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_267
timestamp 1606120353
transform 1 0 25668 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_271
timestamp 1606120353
transform 1 0 26036 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_38_285
timestamp 1606120353
transform 1 0 27324 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__o21a_4  _0958_
timestamp 1606120353
transform 1 0 28520 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__C
timestamp 1606120353
transform 1 0 27600 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__B
timestamp 1606120353
transform 1 0 27968 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__A
timestamp 1606120353
transform 1 0 28336 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_290
timestamp 1606120353
transform 1 0 27784 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_294
timestamp 1606120353
transform 1 0 28152 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__A
timestamp 1606120353
transform 1 0 31004 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A
timestamp 1606120353
transform 1 0 30268 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A1
timestamp 1606120353
transform 1 0 31372 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__B
timestamp 1606120353
transform 1 0 29808 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_310
timestamp 1606120353
transform 1 0 29624 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_38_314
timestamp 1606120353
transform 1 0 29992 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_38_319
timestamp 1606120353
transform 1 0 30452 0 -1 23392
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_38_327
timestamp 1606120353
transform 1 0 31188 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0930_
timestamp 1606120353
transform 1 0 32108 0 -1 23392
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1606120353
transform 1 0 32016 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__B1
timestamp 1606120353
transform 1 0 31740 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_331
timestamp 1606120353
transform 1 0 31556 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_38_335
timestamp 1606120353
transform 1 0 31924 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_38_350
timestamp 1606120353
transform 1 0 33304 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_38_362
timestamp 1606120353
transform 1 0 34408 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_38_374
timestamp 1606120353
transform 1 0 35512 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__CLK
timestamp 1606120353
transform 1 0 35788 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_38_379
timestamp 1606120353
transform 1 0 35972 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_38_391
timestamp 1606120353
transform 1 0 37076 0 -1 23392
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1606120353
transform -1 0 38548 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1606120353
transform 1 0 37628 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_38_398
timestamp 1606120353
transform 1 0 37720 0 -1 23392
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_39_11
timestamp 1606120353
transform 1 0 2116 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_7
timestamp 1606120353
transform 1 0 1748 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1606120353
transform 1 0 1380 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__CLK
timestamp 1606120353
transform 1 0 1932 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__D
timestamp 1606120353
transform 1 0 1564 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1606120353
transform 1 0 1104 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1606120353
transform 1 0 1104 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_40_22
timestamp 1606120353
transform 1 0 3128 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_39_22
timestamp 1606120353
transform 1 0 3128 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_39_19
timestamp 1606120353
transform 1 0 2852 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_39_15
timestamp 1606120353
transform 1 0 2484 0 1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__CLK
timestamp 1606120353
transform 1 0 2300 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__D
timestamp 1606120353
transform 1 0 2944 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1123_
timestamp 1606120353
transform 1 0 1380 0 -1 24480
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__C
timestamp 1606120353
transform 1 0 3312 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__A2
timestamp 1606120353
transform 1 0 3404 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__A
timestamp 1606120353
transform 1 0 3680 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_26
timestamp 1606120353
transform 1 0 3496 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_27
timestamp 1606120353
transform 1 0 3588 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1606120353
transform 1 0 3956 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__D
timestamp 1606120353
transform 1 0 3772 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_30
timestamp 1606120353
transform 1 0 3864 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__C1
timestamp 1606120353
transform 1 0 4048 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_40_32
timestamp 1606120353
transform 1 0 4048 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_39_42
timestamp 1606120353
transform 1 0 4968 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_38
timestamp 1606120353
transform 1 0 4600 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_34
timestamp 1606120353
transform 1 0 4232 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__B1
timestamp 1606120353
transform 1 0 5152 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__A1
timestamp 1606120353
transform 1 0 4784 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__A2
timestamp 1606120353
transform 1 0 4416 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__a211o_4  _0657_
timestamp 1606120353
transform 1 0 4324 0 -1 24480
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_40_53
timestamp 1606120353
transform 1 0 5980 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_49
timestamp 1606120353
transform 1 0 5612 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_53
timestamp 1606120353
transform 1 0 5980 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_46
timestamp 1606120353
transform 1 0 5336 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__D
timestamp 1606120353
transform 1 0 5796 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__B
timestamp 1606120353
transform 1 0 5520 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__A
timestamp 1606120353
transform 1 0 6164 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__A
timestamp 1606120353
transform 1 0 6164 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0653_
timestamp 1606120353
transform 1 0 5704 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1606120353
transform 1 0 6348 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__C
timestamp 1606120353
transform 1 0 6532 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1606120353
transform 1 0 6716 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0677_
timestamp 1606120353
transform 1 0 6808 0 1 23392
box 0 -48 828 592
use sky130_fd_sc_hd__nor4_4  _0684_
timestamp 1606120353
transform 1 0 6348 0 -1 24480
box 0 -48 1564 592
use sky130_fd_sc_hd__fill_2  FILLER_40_74
timestamp 1606120353
transform 1 0 7912 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_39_71
timestamp 1606120353
transform 1 0 7636 0 1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A
timestamp 1606120353
transform 1 0 8004 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_83
timestamp 1606120353
transform 1 0 8740 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_40_78
timestamp 1606120353
transform 1 0 8280 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_39_77
timestamp 1606120353
transform 1 0 8188 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__B2
timestamp 1606120353
transform 1 0 8096 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__C
timestamp 1606120353
transform 1 0 8556 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__B
timestamp 1606120353
transform 1 0 8372 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0721_
timestamp 1606120353
transform 1 0 8556 0 1 23392
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_40_87
timestamp 1606120353
transform 1 0 9108 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__B1
timestamp 1606120353
transform 1 0 8924 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_40_91
timestamp 1606120353
transform 1 0 9476 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_39_99
timestamp 1606120353
transform 1 0 10212 0 1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_39_95
timestamp 1606120353
transform 1 0 9844 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_39_90
timestamp 1606120353
transform 1 0 9384 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A3
timestamp 1606120353
transform 1 0 9292 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__B2
timestamp 1606120353
transform 1 0 10028 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A1
timestamp 1606120353
transform 1 0 9660 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1606120353
transform 1 0 9568 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1606120353
transform 1 0 11224 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__A
timestamp 1606120353
transform 1 0 10580 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _0745_
timestamp 1606120353
transform 1 0 10764 0 1 23392
box 0 -48 828 592
use sky130_fd_sc_hd__a32o_4  _0735_
timestamp 1606120353
transform 1 0 9660 0 -1 24480
box 0 -48 1564 592
use sky130_fd_sc_hd__decap_3  FILLER_40_118
timestamp 1606120353
transform 1 0 11960 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_40_114
timestamp 1606120353
transform 1 0 11592 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1606120353
transform 1 0 11960 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_114
timestamp 1606120353
transform 1 0 11592 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__C1
timestamp 1606120353
transform 1 0 11776 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__C1
timestamp 1606120353
transform 1 0 12236 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__C
timestamp 1606120353
transform 1 0 11776 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A1
timestamp 1606120353
transform 1 0 11408 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A
timestamp 1606120353
transform 1 0 12144 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_130
timestamp 1606120353
transform 1 0 13064 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_39_123
timestamp 1606120353
transform 1 0 12420 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__A1
timestamp 1606120353
transform 1 0 13248 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A2
timestamp 1606120353
transform 1 0 12696 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1606120353
transform 1 0 12328 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _0716_
timestamp 1606120353
transform 1 0 12420 0 -1 24480
box 0 -48 644 592
use sky130_fd_sc_hd__a211o_4  _0730_
timestamp 1606120353
transform 1 0 12880 0 1 23392
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_40_134
timestamp 1606120353
transform 1 0 13432 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_142
timestamp 1606120353
transform 1 0 14168 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__B1
timestamp 1606120353
transform 1 0 13616 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0771_
timestamp 1606120353
transform 1 0 13800 0 -1 24480
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_40_149
timestamp 1606120353
transform 1 0 14812 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_145
timestamp 1606120353
transform 1 0 14444 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_39_146
timestamp 1606120353
transform 1 0 14536 0 1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__B
timestamp 1606120353
transform 1 0 14628 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A1
timestamp 1606120353
transform 1 0 14996 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__B1
timestamp 1606120353
transform 1 0 14904 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__B
timestamp 1606120353
transform 1 0 14352 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1606120353
transform 1 0 15180 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0750_
timestamp 1606120353
transform 1 0 15088 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__o21a_4  _0773_
timestamp 1606120353
transform 1 0 15272 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_39_159
timestamp 1606120353
transform 1 0 15732 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_155
timestamp 1606120353
transform 1 0 15364 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__A
timestamp 1606120353
transform 1 0 15548 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A2
timestamp 1606120353
transform 1 0 15916 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_174
timestamp 1606120353
transform 1 0 17112 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_170
timestamp 1606120353
transform 1 0 16744 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1606120353
transform 1 0 16376 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_175
timestamp 1606120353
transform 1 0 17204 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__A1
timestamp 1606120353
transform 1 0 17296 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A1
timestamp 1606120353
transform 1 0 16928 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__B1
timestamp 1606120353
transform 1 0 16560 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0760_
timestamp 1606120353
transform 1 0 16100 0 1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_40_178
timestamp 1606120353
transform 1 0 17480 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_39_184
timestamp 1606120353
transform 1 0 18032 0 1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_39_179
timestamp 1606120353
transform 1 0 17572 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A1
timestamp 1606120353
transform 1 0 17756 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__A
timestamp 1606120353
transform 1 0 17388 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1606120353
transform 1 0 17940 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_40_198
timestamp 1606120353
transform 1 0 19320 0 -1 24480
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_39_197
timestamp 1606120353
transform 1 0 19228 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__B
timestamp 1606120353
transform 1 0 18400 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0776_
timestamp 1606120353
transform 1 0 18584 0 1 23392
box 0 -48 644 592
use sky130_fd_sc_hd__dfxtp_4  _1090_
timestamp 1606120353
transform 1 0 17572 0 -1 24480
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_4  FILLER_40_206
timestamp 1606120353
transform 1 0 20056 0 -1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_39_207
timestamp 1606120353
transform 1 0 20148 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_39_201
timestamp 1606120353
transform 1 0 19596 0 1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__CLK
timestamp 1606120353
transform 1 0 19872 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__B1
timestamp 1606120353
transform 1 0 19964 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A1
timestamp 1606120353
transform 1 0 20332 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__A
timestamp 1606120353
transform 1 0 19412 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_219
timestamp 1606120353
transform 1 0 21252 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_215
timestamp 1606120353
transform 1 0 20884 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_40_213
timestamp 1606120353
transform 1 0 20700 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_40_210
timestamp 1606120353
transform 1 0 20424 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A2
timestamp 1606120353
transform 1 0 20516 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__B1
timestamp 1606120353
transform 1 0 21068 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1606120353
transform 1 0 20792 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _0802_
timestamp 1606120353
transform 1 0 20516 0 1 23392
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  FILLER_40_231
timestamp 1606120353
transform 1 0 22356 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_40_223
timestamp 1606120353
transform 1 0 21620 0 -1 24480
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_39_225
timestamp 1606120353
transform 1 0 21804 0 1 23392
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__B2
timestamp 1606120353
transform 1 0 21436 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_39_240
timestamp 1606120353
transform 1 0 23184 0 1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_39_236
timestamp 1606120353
transform 1 0 22816 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_39_233
timestamp 1606120353
transform 1 0 22540 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__CLK
timestamp 1606120353
transform 1 0 23000 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__D
timestamp 1606120353
transform 1 0 22632 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1149_
timestamp 1606120353
transform 1 0 22632 0 -1 24480
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_6  FILLER_40_253
timestamp 1606120353
transform 1 0 24380 0 -1 24480
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1606120353
transform 1 0 23552 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_40_261
timestamp 1606120353
transform 1 0 25116 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_39_263
timestamp 1606120353
transform 1 0 25300 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_39_257
timestamp 1606120353
transform 1 0 24748 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A
timestamp 1606120353
transform 1 0 24840 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__A
timestamp 1606120353
transform 1 0 24932 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0885_
timestamp 1606120353
transform 1 0 25392 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0824_
timestamp 1606120353
transform 1 0 25024 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_39_245
timestamp 1606120353
transform 1 0 23644 0 1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 1606120353
transform 1 0 26036 0 -1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_40_267
timestamp 1606120353
transform 1 0 25668 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_267
timestamp 1606120353
transform 1 0 25668 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A
timestamp 1606120353
transform 1 0 25852 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__A
timestamp 1606120353
transform 1 0 25484 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A
timestamp 1606120353
transform 1 0 25852 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0836_
timestamp 1606120353
transform 1 0 26036 0 1 23392
box 0 -48 828 592
use sky130_fd_sc_hd__decap_4  FILLER_40_276
timestamp 1606120353
transform 1 0 26496 0 -1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_39_280
timestamp 1606120353
transform 1 0 26864 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A
timestamp 1606120353
transform 1 0 27048 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1606120353
transform 1 0 26404 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _0834_
timestamp 1606120353
transform 1 0 26864 0 -1 24480
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_39_284
timestamp 1606120353
transform 1 0 27232 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__A
timestamp 1606120353
transform 1 0 27416 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_293
timestamp 1606120353
transform 1 0 28060 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_289
timestamp 1606120353
transform 1 0 27692 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__A
timestamp 1606120353
transform 1 0 28244 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__C
timestamp 1606120353
transform 1 0 27876 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__or3_4  _0835_
timestamp 1606120353
transform 1 0 27600 0 1 23392
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_39_301
timestamp 1606120353
transform 1 0 28796 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_297
timestamp 1606120353
transform 1 0 28428 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__C
timestamp 1606120353
transform 1 0 28612 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__B
timestamp 1606120353
transform 1 0 28980 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__or3_4  _0841_
timestamp 1606120353
transform 1 0 28428 0 -1 24480
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILLER_40_306
timestamp 1606120353
transform 1 0 29256 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_39_306
timestamp 1606120353
transform 1 0 29256 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1606120353
transform 1 0 29164 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_40_317
timestamp 1606120353
transform 1 0 30268 0 -1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_40_311
timestamp 1606120353
transform 1 0 29716 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_39_316
timestamp 1606120353
transform 1 0 30176 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A
timestamp 1606120353
transform 1 0 29532 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__A
timestamp 1606120353
transform 1 0 30360 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0838_
timestamp 1606120353
transform 1 0 29532 0 1 23392
box 0 -48 644 592
use sky130_fd_sc_hd__buf_1  _0832_
timestamp 1606120353
transform 1 0 29992 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_40_328
timestamp 1606120353
transform 1 0 31280 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_323
timestamp 1606120353
transform 1 0 30820 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_320
timestamp 1606120353
transform 1 0 30544 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__B1
timestamp 1606120353
transform 1 0 31464 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__B
timestamp 1606120353
transform 1 0 30636 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A2
timestamp 1606120353
transform 1 0 30728 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0839_
timestamp 1606120353
transform 1 0 31004 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _0874_
timestamp 1606120353
transform 1 0 30912 0 1 23392
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_40_340
timestamp 1606120353
transform 1 0 32384 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_40_332
timestamp 1606120353
transform 1 0 31648 0 -1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1606120353
transform 1 0 32108 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__A
timestamp 1606120353
transform 1 0 32292 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1606120353
transform 1 0 32016 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0822_
timestamp 1606120353
transform 1 0 32108 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_40_344
timestamp 1606120353
transform 1 0 32752 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A
timestamp 1606120353
transform 1 0 32936 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__B
timestamp 1606120353
transform 1 0 32568 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_40_348
timestamp 1606120353
transform 1 0 33120 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_39_341
timestamp 1606120353
transform 1 0 32476 0 1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1606120353
transform 1 0 34776 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_39_353
timestamp 1606120353
transform 1 0 33580 0 1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_39_365
timestamp 1606120353
transform 1 0 34684 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_39_367
timestamp 1606120353
transform 1 0 34868 0 1 23392
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_40_360
timestamp 1606120353
transform 1 0 34224 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_40_372
timestamp 1606120353
transform 1 0 35328 0 -1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1154_
timestamp 1606120353
transform 1 0 35788 0 1 23392
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__D
timestamp 1606120353
transform 1 0 35604 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__CLK
timestamp 1606120353
transform 1 0 35788 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_39_396
timestamp 1606120353
transform 1 0 37536 0 1 23392
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_40_376
timestamp 1606120353
transform 1 0 35696 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_40_379
timestamp 1606120353
transform 1 0 35972 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_40_391
timestamp 1606120353
transform 1 0 37076 0 -1 24480
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1606120353
transform -1 0 38548 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1606120353
transform -1 0 38548 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1606120353
transform 1 0 37628 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_40_398
timestamp 1606120353
transform 1 0 37720 0 -1 24480
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1606120353
transform 1 0 1104 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1606120353
transform 1 0 1380 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_41_15
timestamp 1606120353
transform 1 0 2484 0 1 24480
box 0 -48 736 592
use sky130_fd_sc_hd__inv_8  _0502_
timestamp 1606120353
transform 1 0 3496 0 1 24480
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__A1
timestamp 1606120353
transform 1 0 4508 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0509__B
timestamp 1606120353
transform 1 0 5060 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0502__A
timestamp 1606120353
transform 1 0 3312 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_41_23
timestamp 1606120353
transform 1 0 3220 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_41_35
timestamp 1606120353
transform 1 0 4324 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_41_39
timestamp 1606120353
transform 1 0 4692 0 1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _0509_
timestamp 1606120353
transform 1 0 5244 0 1 24480
box 0 -48 644 592
use sky130_fd_sc_hd__and4_4  _0676_
timestamp 1606120353
transform 1 0 6808 0 1 24480
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1606120353
transform 1 0 6716 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__B
timestamp 1606120353
transform 1 0 6532 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0509__A
timestamp 1606120353
transform 1 0 6072 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_52
timestamp 1606120353
transform 1 0 5888 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_41_56
timestamp 1606120353
transform 1 0 6256 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__a32o_4  _0772_
timestamp 1606120353
transform 1 0 8924 0 1 24480
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__B1
timestamp 1606120353
transform 1 0 7820 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A1
timestamp 1606120353
transform 1 0 8740 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A1
timestamp 1606120353
transform 1 0 8188 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_71
timestamp 1606120353
transform 1 0 7636 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_75
timestamp 1606120353
transform 1 0 8004 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_41_79
timestamp 1606120353
transform 1 0 8372 0 1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__B1
timestamp 1606120353
transform 1 0 10672 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A
timestamp 1606120353
transform 1 0 11132 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_102
timestamp 1606120353
transform 1 0 10488 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_41_106
timestamp 1606120353
transform 1 0 10856 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0668_
timestamp 1606120353
transform 1 0 11316 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__a211o_4  _0746_
timestamp 1606120353
transform 1 0 12420 0 1 24480
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1606120353
transform 1 0 12328 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__B2
timestamp 1606120353
transform 1 0 12144 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__B1
timestamp 1606120353
transform 1 0 11776 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_114
timestamp 1606120353
transform 1 0 11592 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1606120353
transform 1 0 11960 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0719_
timestamp 1606120353
transform 1 0 14444 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__A
timestamp 1606120353
transform 1 0 14904 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__B1
timestamp 1606120353
transform 1 0 13892 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__A2
timestamp 1606120353
transform 1 0 14260 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__A3
timestamp 1606120353
transform 1 0 15272 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_137
timestamp 1606120353
transform 1 0 13708 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_141
timestamp 1606120353
transform 1 0 14076 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_148
timestamp 1606120353
transform 1 0 14720 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_152
timestamp 1606120353
transform 1 0 15088 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _0775_
timestamp 1606120353
transform 1 0 15640 0 1 24480
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A2
timestamp 1606120353
transform 1 0 17112 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_156
timestamp 1606120353
transform 1 0 15456 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_172
timestamp 1606120353
transform 1 0 16928 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_176
timestamp 1606120353
transform 1 0 17296 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1606120353
transform 1 0 17940 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__B1
timestamp 1606120353
transform 1 0 17480 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_41_180
timestamp 1606120353
transform 1 0 17664 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1606120353
transform 1 0 18032 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_41_196
timestamp 1606120353
transform 1 0 19136 0 1 24480
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1100_
timestamp 1606120353
transform 1 0 19872 0 1 24480
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__D
timestamp 1606120353
transform 1 0 19688 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A1
timestamp 1606120353
transform 1 0 21804 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A2
timestamp 1606120353
transform 1 0 22172 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_223
timestamp 1606120353
transform 1 0 21620 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_227
timestamp 1606120353
transform 1 0 21988 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_41_231
timestamp 1606120353
transform 1 0 22356 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__nand4_4  _1042_
timestamp 1606120353
transform 1 0 24932 0 1 24480
box 0 -48 1564 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1606120353
transform 1 0 23552 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__C
timestamp 1606120353
transform 1 0 24748 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__D
timestamp 1606120353
transform 1 0 24380 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_41_243
timestamp 1606120353
transform 1 0 23460 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_41_245
timestamp 1606120353
transform 1 0 23644 0 1 24480
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_41_255
timestamp 1606120353
transform 1 0 24564 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__A1
timestamp 1606120353
transform 1 0 27232 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__A2
timestamp 1606120353
transform 1 0 26864 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1606120353
transform 1 0 26496 0 1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_41_282
timestamp 1606120353
transform 1 0 27048 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_286
timestamp 1606120353
transform 1 0 27416 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__or3_4  _0831_
timestamp 1606120353
transform 1 0 27600 0 1 24480
box 0 -48 828 592
use sky130_fd_sc_hd__buf_1  _0858_
timestamp 1606120353
transform 1 0 29256 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1606120353
transform 1 0 29164 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__B
timestamp 1606120353
transform 1 0 28980 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__B1
timestamp 1606120353
transform 1 0 28612 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_297
timestamp 1606120353
transform 1 0 28428 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_301
timestamp 1606120353
transform 1 0 28796 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0873_
timestamp 1606120353
transform 1 0 30636 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A
timestamp 1606120353
transform 1 0 29716 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A2
timestamp 1606120353
transform 1 0 30452 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__C
timestamp 1606120353
transform 1 0 30084 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_309
timestamp 1606120353
transform 1 0 29532 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_313
timestamp 1606120353
transform 1 0 29900 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_317
timestamp 1606120353
transform 1 0 30268 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0872_
timestamp 1606120353
transform 1 0 32476 0 1 24480
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__A
timestamp 1606120353
transform 1 0 32108 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__A
timestamp 1606120353
transform 1 0 33488 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_41_333
timestamp 1606120353
transform 1 0 31740 0 1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_41_339
timestamp 1606120353
transform 1 0 32292 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_350
timestamp 1606120353
transform 1 0 33304 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1606120353
transform 1 0 34776 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_41_354
timestamp 1606120353
transform 1 0 33672 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_41_367
timestamp 1606120353
transform 1 0 34868 0 1 24480
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1162_
timestamp 1606120353
transform 1 0 35788 0 1 24480
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__D
timestamp 1606120353
transform 1 0 35604 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_41_396
timestamp 1606120353
transform 1 0 37536 0 1 24480
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1606120353
transform -1 0 38548 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1606120353
transform 1 0 1104 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__D
timestamp 1606120353
transform 1 0 1564 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1606120353
transform 1 0 1380 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_42_7
timestamp 1606120353
transform 1 0 1748 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_42_19
timestamp 1606120353
transform 1 0 2852 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__a21oi_4  _0648_
timestamp 1606120353
transform 1 0 4416 0 -1 25568
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1606120353
transform 1 0 3956 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__B1
timestamp 1606120353
transform 1 0 4232 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_32
timestamp 1606120353
transform 1 0 4048 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__a32o_4  _0671_
timestamp 1606120353
transform 1 0 7176 0 -1 25568
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A
timestamp 1606120353
transform 1 0 6808 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__C
timestamp 1606120353
transform 1 0 6440 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A2
timestamp 1606120353
transform 1 0 6072 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_42_49
timestamp 1606120353
transform 1 0 5612 0 -1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_42_53
timestamp 1606120353
transform 1 0 5980 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_42_56
timestamp 1606120353
transform 1 0 6256 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_60
timestamp 1606120353
transform 1 0 6624 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_64
timestamp 1606120353
transform 1 0 6992 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A2
timestamp 1606120353
transform 1 0 8924 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_83
timestamp 1606120353
transform 1 0 8740 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_42_87
timestamp 1606120353
transform 1 0 9108 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__a211o_4  _0736_
timestamp 1606120353
transform 1 0 10580 0 -1 25568
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1606120353
transform 1 0 9568 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__A2
timestamp 1606120353
transform 1 0 9844 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A1
timestamp 1606120353
transform 1 0 10304 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__B
timestamp 1606120353
transform 1 0 9384 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_93
timestamp 1606120353
transform 1 0 9660 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_42_97
timestamp 1606120353
transform 1 0 10028 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_42_102
timestamp 1606120353
transform 1 0 10488 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__a32o_4  _0747_
timestamp 1606120353
transform 1 0 12604 0 -1 25568
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A2
timestamp 1606120353
transform 1 0 12420 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A3
timestamp 1606120353
transform 1 0 12052 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_117
timestamp 1606120353
transform 1 0 11868 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_121
timestamp 1606120353
transform 1 0 12236 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1606120353
transform 1 0 15180 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__A
timestamp 1606120353
transform 1 0 14352 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__B2
timestamp 1606120353
transform 1 0 14996 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_142
timestamp 1606120353
transform 1 0 14168 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_42_146
timestamp 1606120353
transform 1 0 14536 0 -1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_42_150
timestamp 1606120353
transform 1 0 14904 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_42_154
timestamp 1606120353
transform 1 0 15272 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0798_
timestamp 1606120353
transform 1 0 16652 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__B1
timestamp 1606120353
transform 1 0 15456 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__A2
timestamp 1606120353
transform 1 0 15824 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__B1
timestamp 1606120353
transform 1 0 16192 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_158
timestamp 1606120353
transform 1 0 15640 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_162
timestamp 1606120353
transform 1 0 16008 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_42_166
timestamp 1606120353
transform 1 0 16376 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__D
timestamp 1606120353
transform 1 0 18216 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_42_181
timestamp 1606120353
transform 1 0 17756 0 -1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_42_185
timestamp 1606120353
transform 1 0 18124 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_42_188
timestamp 1606120353
transform 1 0 18400 0 -1 25568
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_42_196
timestamp 1606120353
transform 1 0 19136 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__o22a_4  _0803_
timestamp 1606120353
transform 1 0 20884 0 -1 25568
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1606120353
transform 1 0 20792 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__B
timestamp 1606120353
transform 1 0 19412 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_42_201
timestamp 1606120353
transform 1 0 19596 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_42_213
timestamp 1606120353
transform 1 0 20700 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_42_229
timestamp 1606120353
transform 1 0 22172 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_42_241
timestamp 1606120353
transform 1 0 23276 0 -1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _0823_
timestamp 1606120353
transform 1 0 25392 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__B
timestamp 1606120353
transform 1 0 24932 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__CLK
timestamp 1606120353
transform 1 0 23644 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_42_247
timestamp 1606120353
transform 1 0 23828 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_42_261
timestamp 1606120353
transform 1 0 25116 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__o21a_4  _0826_
timestamp 1606120353
transform 1 0 27232 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1606120353
transform 1 0 26404 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__B
timestamp 1606120353
transform 1 0 27048 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A1
timestamp 1606120353
transform 1 0 26680 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_42_267
timestamp 1606120353
transform 1 0 25668 0 -1 25568
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_42_276
timestamp 1606120353
transform 1 0 26496 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_280
timestamp 1606120353
transform 1 0 26864 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _0845_
timestamp 1606120353
transform 1 0 29072 0 -1 25568
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__C1
timestamp 1606120353
transform 1 0 28888 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_42_296
timestamp 1606120353
transform 1 0 28336 0 -1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _0859_
timestamp 1606120353
transform 1 0 30636 0 -1 25568
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__A
timestamp 1606120353
transform 1 0 30084 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__A
timestamp 1606120353
transform 1 0 31464 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A1
timestamp 1606120353
transform 1 0 30452 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_313
timestamp 1606120353
transform 1 0 29900 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_317
timestamp 1606120353
transform 1 0 30268 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_328
timestamp 1606120353
transform 1 0 31280 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0833_
timestamp 1606120353
transform 1 0 33488 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__and2_4  _0844_
timestamp 1606120353
transform 1 0 32108 0 -1 25568
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1606120353
transform 1 0 32016 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A
timestamp 1606120353
transform 1 0 31832 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_332
timestamp 1606120353
transform 1 0 31648 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_42_344
timestamp 1606120353
transform 1 0 32752 0 -1 25568
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_42_355
timestamp 1606120353
transform 1 0 33764 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_42_367
timestamp 1606120353
transform 1 0 34868 0 -1 25568
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__CLK
timestamp 1606120353
transform 1 0 35788 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_375
timestamp 1606120353
transform 1 0 35604 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_42_379
timestamp 1606120353
transform 1 0 35972 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_42_391
timestamp 1606120353
transform 1 0 37076 0 -1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1606120353
transform -1 0 38548 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1606120353
transform 1 0 37628 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_42_398
timestamp 1606120353
transform 1 0 37720 0 -1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1205_
timestamp 1606120353
transform 1 0 1380 0 1 25568
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1606120353
transform 1 0 1104 0 1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_43_22
timestamp 1606120353
transform 1 0 3128 0 1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__inv_8  _0673_
timestamp 1606120353
transform 1 0 3864 0 1 25568
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__B1
timestamp 1606120353
transform 1 0 4876 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A
timestamp 1606120353
transform 1 0 3680 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_39
timestamp 1606120353
transform 1 0 4692 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_43
timestamp 1606120353
transform 1 0 5060 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0685_
timestamp 1606120353
transform 1 0 6808 0 1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1606120353
transform 1 0 6716 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__A1
timestamp 1606120353
transform 1 0 6532 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__A2
timestamp 1606120353
transform 1 0 6164 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__B1
timestamp 1606120353
transform 1 0 5796 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A2
timestamp 1606120353
transform 1 0 5244 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_43_47
timestamp 1606120353
transform 1 0 5428 0 1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_43_53
timestamp 1606120353
transform 1 0 5980 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1606120353
transform 1 0 6348 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0655_
timestamp 1606120353
transform 1 0 8648 0 1 25568
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__B1
timestamp 1606120353
transform 1 0 8096 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__B
timestamp 1606120353
transform 1 0 8464 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_74
timestamp 1606120353
transform 1 0 7912 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_78
timestamp 1606120353
transform 1 0 8280 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__a211o_4  _0672_
timestamp 1606120353
transform 1 0 10304 0 1 25568
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__B1
timestamp 1606120353
transform 1 0 10120 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__B1
timestamp 1606120353
transform 1 0 9660 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_43_89
timestamp 1606120353
transform 1 0 9292 0 1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_43_95
timestamp 1606120353
transform 1 0 9844 0 1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_43_114
timestamp 1606120353
transform 1 0 11592 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__B1
timestamp 1606120353
transform 1 0 11776 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_118
timestamp 1606120353
transform 1 0 11960 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A1
timestamp 1606120353
transform 1 0 12144 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_123
timestamp 1606120353
transform 1 0 12420 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1606120353
transform 1 0 12328 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A2
timestamp 1606120353
transform 1 0 12604 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_127
timestamp 1606120353
transform 1 0 12788 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__B2
timestamp 1606120353
transform 1 0 12972 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_131
timestamp 1606120353
transform 1 0 13156 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_135
timestamp 1606120353
transform 1 0 13524 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__C1
timestamp 1606120353
transform 1 0 13340 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A1
timestamp 1606120353
transform 1 0 13708 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_139
timestamp 1606120353
transform 1 0 13892 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0496__A
timestamp 1606120353
transform 1 0 14076 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_43_143
timestamp 1606120353
transform 1 0 14260 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0711_
timestamp 1606120353
transform 1 0 14352 0 1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_43_147
timestamp 1606120353
transform 1 0 14628 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A2
timestamp 1606120353
transform 1 0 14812 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_151
timestamp 1606120353
transform 1 0 14996 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0495__A
timestamp 1606120353
transform 1 0 15180 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0774_
timestamp 1606120353
transform 1 0 15364 0 1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A1
timestamp 1606120353
transform 1 0 16928 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__B1
timestamp 1606120353
transform 1 0 17296 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_43_167
timestamp 1606120353
transform 1 0 16468 0 1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_43_171
timestamp 1606120353
transform 1 0 16836 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_43_174
timestamp 1606120353
transform 1 0 17112 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1084_
timestamp 1606120353
transform 1 0 18216 0 1 25568
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1606120353
transform 1 0 17940 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__B2
timestamp 1606120353
transform 1 0 17664 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_178
timestamp 1606120353
transform 1 0 17480 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_43_182
timestamp 1606120353
transform 1 0 17848 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_43_184
timestamp 1606120353
transform 1 0 18032 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A
timestamp 1606120353
transform 1 0 20148 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A1
timestamp 1606120353
transform 1 0 20884 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A2
timestamp 1606120353
transform 1 0 21252 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_205
timestamp 1606120353
transform 1 0 19964 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_43_209
timestamp 1606120353
transform 1 0 20332 0 1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_43_217
timestamp 1606120353
transform 1 0 21068 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0830_
timestamp 1606120353
transform 1 0 21988 0 1 25568
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__D
timestamp 1606120353
transform 1 0 23368 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__B1
timestamp 1606120353
transform 1 0 21620 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_221
timestamp 1606120353
transform 1 0 21436 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1606120353
transform 1 0 21804 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_43_236
timestamp 1606120353
transform 1 0 22816 0 1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1116_
timestamp 1606120353
transform 1 0 23644 0 1 25568
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1606120353
transform 1 0 23552 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_43_264
timestamp 1606120353
transform 1 0 25392 0 1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__buf_1  _0883_
timestamp 1606120353
transform 1 0 26588 0 1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__A
timestamp 1606120353
transform 1 0 27048 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A2
timestamp 1606120353
transform 1 0 26404 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__B1_N
timestamp 1606120353
transform 1 0 26036 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_43_270
timestamp 1606120353
transform 1 0 25944 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_43_273
timestamp 1606120353
transform 1 0 26220 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_280
timestamp 1606120353
transform 1 0 26864 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_43_284
timestamp 1606120353
transform 1 0 27232 0 1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _0846_
timestamp 1606120353
transform 1 0 29256 0 1 25568
box 0 -48 644 592
use sky130_fd_sc_hd__buf_1  _0881_
timestamp 1606120353
transform 1 0 27600 0 1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1606120353
transform 1 0 29164 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A1
timestamp 1606120353
transform 1 0 28980 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__A
timestamp 1606120353
transform 1 0 28060 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A2
timestamp 1606120353
transform 1 0 28612 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_291
timestamp 1606120353
transform 1 0 27876 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_43_295
timestamp 1606120353
transform 1 0 28244 0 1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_43_301
timestamp 1606120353
transform 1 0 28796 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0852_
timestamp 1606120353
transform 1 0 30636 0 1 25568
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__B1
timestamp 1606120353
transform 1 0 30084 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__B
timestamp 1606120353
transform 1 0 31464 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__B
timestamp 1606120353
transform 1 0 30452 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_313
timestamp 1606120353
transform 1 0 29900 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_317
timestamp 1606120353
transform 1 0 30268 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_328
timestamp 1606120353
transform 1 0 31280 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0921_
timestamp 1606120353
transform 1 0 32384 0 1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A1
timestamp 1606120353
transform 1 0 32200 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__B1
timestamp 1606120353
transform 1 0 31832 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_332
timestamp 1606120353
transform 1 0 31648 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_336
timestamp 1606120353
transform 1 0 32016 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_352
timestamp 1606120353
transform 1 0 33488 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1606120353
transform 1 0 34776 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__A
timestamp 1606120353
transform 1 0 33672 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__A
timestamp 1606120353
transform 1 0 34500 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_43_356
timestamp 1606120353
transform 1 0 33856 0 1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_43_362
timestamp 1606120353
transform 1 0 34408 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_43_365
timestamp 1606120353
transform 1 0 34684 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_43_367
timestamp 1606120353
transform 1 0 34868 0 1 25568
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1195_
timestamp 1606120353
transform 1 0 35788 0 1 25568
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__D
timestamp 1606120353
transform 1 0 35604 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_43_396
timestamp 1606120353
transform 1 0 37536 0 1 25568
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1606120353
transform -1 0 38548 0 1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1606120353
transform 1 0 1104 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__CLK
timestamp 1606120353
transform 1 0 1564 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1606120353
transform 1 0 1380 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_44_7
timestamp 1606120353
transform 1 0 1748 0 -1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_44_19
timestamp 1606120353
transform 1 0 2852 0 -1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__a21oi_4  _0706_
timestamp 1606120353
transform 1 0 4692 0 -1 26656
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1606120353
transform 1 0 3956 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A2_N
timestamp 1606120353
transform 1 0 3312 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A1
timestamp 1606120353
transform 1 0 4508 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_44_23
timestamp 1606120353
transform 1 0 3220 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_44_26
timestamp 1606120353
transform 1 0 3496 0 -1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_44_30
timestamp 1606120353
transform 1 0 3864 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_44_32
timestamp 1606120353
transform 1 0 4048 0 -1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_44_36
timestamp 1606120353
transform 1 0 4416 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__o21ai_4  _0551_
timestamp 1606120353
transform 1 0 6624 0 -1 26656
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A
timestamp 1606120353
transform 1 0 6440 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A1
timestamp 1606120353
transform 1 0 6072 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_52
timestamp 1606120353
transform 1 0 5888 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_56
timestamp 1606120353
transform 1 0 6256 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__B
timestamp 1606120353
transform 1 0 8004 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A2
timestamp 1606120353
transform 1 0 8372 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A1
timestamp 1606120353
transform 1 0 8740 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A2
timestamp 1606120353
transform 1 0 9108 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_73
timestamp 1606120353
transform 1 0 7820 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_77
timestamp 1606120353
transform 1 0 8188 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_81
timestamp 1606120353
transform 1 0 8556 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1606120353
transform 1 0 8924 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0707_
timestamp 1606120353
transform 1 0 9660 0 -1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1606120353
transform 1 0 9568 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__C1
timestamp 1606120353
transform 1 0 10948 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_44_89
timestamp 1606120353
transform 1 0 9292 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_44_105
timestamp 1606120353
transform 1 0 10764 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_109
timestamp 1606120353
transform 1 0 11132 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__a32o_4  _0712_
timestamp 1606120353
transform 1 0 11776 0 -1 26656
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__C
timestamp 1606120353
transform 1 0 11316 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_44_113
timestamp 1606120353
transform 1 0 11500 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0495_
timestamp 1606120353
transform 1 0 15272 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0496_
timestamp 1606120353
transform 1 0 14076 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1606120353
transform 1 0 15180 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A1
timestamp 1606120353
transform 1 0 13524 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_133
timestamp 1606120353
transform 1 0 13340 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_44_137
timestamp 1606120353
transform 1 0 13708 0 -1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_44_144
timestamp 1606120353
transform 1 0 14352 0 -1 26656
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_44_152
timestamp 1606120353
transform 1 0 15088 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _0800_
timestamp 1606120353
transform 1 0 16928 0 -1 26656
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A1
timestamp 1606120353
transform 1 0 15732 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__D
timestamp 1606120353
transform 1 0 16284 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A2
timestamp 1606120353
transform 1 0 16744 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_157
timestamp 1606120353
transform 1 0 15548 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_44_161
timestamp 1606120353
transform 1 0 15916 0 -1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_44_167
timestamp 1606120353
transform 1 0 16468 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A1
timestamp 1606120353
transform 1 0 19044 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__CLK
timestamp 1606120353
transform 1 0 18400 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_186
timestamp 1606120353
transform 1 0 18216 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_44_190
timestamp 1606120353
transform 1 0 18584 0 -1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_44_194
timestamp 1606120353
transform 1 0 18952 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1606120353
transform 1 0 19228 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0714_
timestamp 1606120353
transform 1 0 19412 0 -1 26656
box 0 -48 644 592
use sky130_fd_sc_hd__o21ai_4  _0850_
timestamp 1606120353
transform 1 0 20884 0 -1 26656
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1606120353
transform 1 0 20792 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_44_206
timestamp 1606120353
transform 1 0 20056 0 -1 26656
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A
timestamp 1606120353
transform 1 0 22264 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_228
timestamp 1606120353
transform 1 0 22080 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_44_232
timestamp 1606120353
transform 1 0 22448 0 -1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A2
timestamp 1606120353
transform 1 0 23644 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__B1_N
timestamp 1606120353
transform 1 0 24012 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__B1_N
timestamp 1606120353
transform 1 0 24380 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_44_244
timestamp 1606120353
transform 1 0 23552 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_44_247
timestamp 1606120353
transform 1 0 23828 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_251
timestamp 1606120353
transform 1 0 24196 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_44_255
timestamp 1606120353
transform 1 0 24564 0 -1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__a21bo_4  _0898_
timestamp 1606120353
transform 1 0 26496 0 -1 26656
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1606120353
transform 1 0 26404 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A1
timestamp 1606120353
transform 1 0 26220 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_clk_A
timestamp 1606120353
transform 1 0 25852 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_267
timestamp 1606120353
transform 1 0 25668 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_271
timestamp 1606120353
transform 1 0 26036 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__a211o_4  _0847_
timestamp 1606120353
transform 1 0 29072 0 -1 26656
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__B1_N
timestamp 1606120353
transform 1 0 27876 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__A
timestamp 1606120353
transform 1 0 28888 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A1
timestamp 1606120353
transform 1 0 28244 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_289
timestamp 1606120353
transform 1 0 27692 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_293
timestamp 1606120353
transform 1 0 28060 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_44_297
timestamp 1606120353
transform 1 0 28428 0 -1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_44_301
timestamp 1606120353
transform 1 0 28796 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_clk
timestamp 1606120353
transform 1 0 31096 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A1
timestamp 1606120353
transform 1 0 30544 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__A
timestamp 1606120353
transform 1 0 30912 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_318
timestamp 1606120353
transform 1 0 30360 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_322
timestamp 1606120353
transform 1 0 30728 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_44_329
timestamp 1606120353
transform 1 0 31372 0 -1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _0875_
timestamp 1606120353
transform 1 0 32936 0 -1 26656
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1606120353
transform 1 0 32016 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A2
timestamp 1606120353
transform 1 0 32384 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__B
timestamp 1606120353
transform 1 0 32752 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A
timestamp 1606120353
transform 1 0 31832 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_44_333
timestamp 1606120353
transform 1 0 31740 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_44_337
timestamp 1606120353
transform 1 0 32108 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_44_342
timestamp 1606120353
transform 1 0 32568 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0907_
timestamp 1606120353
transform 1 0 34500 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A
timestamp 1606120353
transform 1 0 34960 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_44_355
timestamp 1606120353
transform 1 0 33764 0 -1 26656
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_44_366
timestamp 1606120353
transform 1 0 34776 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_44_370
timestamp 1606120353
transform 1 0 35144 0 -1 26656
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__B1_N
timestamp 1606120353
transform 1 0 35696 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A2
timestamp 1606120353
transform 1 0 36064 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_378
timestamp 1606120353
transform 1 0 35880 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_44_382
timestamp 1606120353
transform 1 0 36248 0 -1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_44_394
timestamp 1606120353
transform 1 0 37352 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1606120353
transform -1 0 38548 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1606120353
transform 1 0 37628 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_44_398
timestamp 1606120353
transform 1 0 37720 0 -1 26656
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1606120353
transform 1 0 1380 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__D
timestamp 1606120353
transform 1 0 1564 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1606120353
transform 1 0 1104 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_45_11
timestamp 1606120353
transform 1 0 2116 0 1 26656
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_45_7
timestamp 1606120353
transform 1 0 1748 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__CLK
timestamp 1606120353
transform 1 0 1932 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_45_17
timestamp 1606120353
transform 1 0 2668 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A1_N
timestamp 1606120353
transform 1 0 2760 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_20
timestamp 1606120353
transform 1 0 2944 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__B2
timestamp 1606120353
transform 1 0 3128 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__a2bb2o_4  _0781_
timestamp 1606120353
transform 1 0 3312 0 1 26656
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__A1
timestamp 1606120353
transform 1 0 5152 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_45_40
timestamp 1606120353
transform 1 0 4784 0 1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _0674_
timestamp 1606120353
transform 1 0 6808 0 1 26656
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1606120353
transform 1 0 6716 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__A2
timestamp 1606120353
transform 1 0 5520 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__A3
timestamp 1606120353
transform 1 0 5888 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__B1
timestamp 1606120353
transform 1 0 6256 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_46
timestamp 1606120353
transform 1 0 5336 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_50
timestamp 1606120353
transform 1 0 5704 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1606120353
transform 1 0 6072 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_45_58
timestamp 1606120353
transform 1 0 6440 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__a21oi_4  _0708_
timestamp 1606120353
transform 1 0 8280 0 1 26656
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__A
timestamp 1606120353
transform 1 0 8004 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__B
timestamp 1606120353
transform 1 0 7636 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_69
timestamp 1606120353
transform 1 0 7452 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_73
timestamp 1606120353
transform 1 0 7820 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_45_77
timestamp 1606120353
transform 1 0 8188 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__o21ai_4  _0710_
timestamp 1606120353
transform 1 0 10304 0 1 26656
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__A1
timestamp 1606120353
transform 1 0 10120 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__B1
timestamp 1606120353
transform 1 0 9660 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_91
timestamp 1606120353
transform 1 0 9476 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_45_95
timestamp 1606120353
transform 1 0 9844 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0709_
timestamp 1606120353
transform 1 0 12420 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1606120353
transform 1 0 12328 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0492__B
timestamp 1606120353
transform 1 0 11776 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0492__C
timestamp 1606120353
transform 1 0 12144 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A
timestamp 1606120353
transform 1 0 12880 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_45_113
timestamp 1606120353
transform 1 0 11500 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_45_118
timestamp 1606120353
transform 1 0 11960 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_126
timestamp 1606120353
transform 1 0 12696 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_45_130
timestamp 1606120353
transform 1 0 13064 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _0494_
timestamp 1606120353
transform 1 0 14076 0 1 26656
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0494__A
timestamp 1606120353
transform 1 0 13892 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0497__A
timestamp 1606120353
transform 1 0 15272 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0501__A
timestamp 1606120353
transform 1 0 13340 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_45_135
timestamp 1606120353
transform 1 0 13524 0 1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_45_150
timestamp 1606120353
transform 1 0 14904 0 1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _0797_
timestamp 1606120353
transform 1 0 16008 0 1 26656
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__B
timestamp 1606120353
transform 1 0 16836 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__A
timestamp 1606120353
transform 1 0 15824 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__CLK
timestamp 1606120353
transform 1 0 17204 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_45_156
timestamp 1606120353
transform 1 0 15456 0 1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1606120353
transform 1 0 16652 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_173
timestamp 1606120353
transform 1 0 17020 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0715_
timestamp 1606120353
transform 1 0 19044 0 1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1606120353
transform 1 0 17940 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__A
timestamp 1606120353
transform 1 0 18768 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__B1
timestamp 1606120353
transform 1 0 18400 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_45_177
timestamp 1606120353
transform 1 0 17388 0 1 26656
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILLER_45_184
timestamp 1606120353
transform 1 0 18032 0 1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_45_190
timestamp 1606120353
transform 1 0 18584 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_45_194
timestamp 1606120353
transform 1 0 18952 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A1
timestamp 1606120353
transform 1 0 21252 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__B1
timestamp 1606120353
transform 1 0 20884 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_45_207
timestamp 1606120353
transform 1 0 20148 0 1 26656
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_45_217
timestamp 1606120353
transform 1 0 21068 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0849_
timestamp 1606120353
transform 1 0 21436 0 1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__A
timestamp 1606120353
transform 1 0 22724 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A2
timestamp 1606120353
transform 1 0 23368 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_233
timestamp 1606120353
transform 1 0 22540 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_45_237
timestamp 1606120353
transform 1 0 22908 0 1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_45_241
timestamp 1606120353
transform 1 0 23276 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__a21bo_4  _0915_
timestamp 1606120353
transform 1 0 23644 0 1 26656
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1606120353
transform 1 0 23552 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A1
timestamp 1606120353
transform 1 0 25024 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_258
timestamp 1606120353
transform 1 0 24840 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_45_262
timestamp 1606120353
transform 1 0 25208 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__a21o_4  _0896_
timestamp 1606120353
transform 1 0 26312 0 1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_clk
timestamp 1606120353
transform 1 0 26036 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A2
timestamp 1606120353
transform 1 0 25852 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__B1
timestamp 1606120353
transform 1 0 25484 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_267
timestamp 1606120353
transform 1 0 25668 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_45_286
timestamp 1606120353
transform 1 0 27416 0 1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _0877_
timestamp 1606120353
transform 1 0 28152 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1606120353
transform 1 0 29164 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A
timestamp 1606120353
transform 1 0 28612 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A2
timestamp 1606120353
transform 1 0 27876 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_45_290
timestamp 1606120353
transform 1 0 27784 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_45_293
timestamp 1606120353
transform 1 0 28060 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_45_297
timestamp 1606120353
transform 1 0 28428 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_45_301
timestamp 1606120353
transform 1 0 28796 0 1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_45_306
timestamp 1606120353
transform 1 0 29256 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__a211o_4  _0853_
timestamp 1606120353
transform 1 0 30084 0 1 26656
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A2
timestamp 1606120353
transform 1 0 29900 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__C1
timestamp 1606120353
transform 1 0 29532 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_311
timestamp 1606120353
transform 1 0 29716 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_45_329
timestamp 1606120353
transform 1 0 31372 0 1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _0920_
timestamp 1606120353
transform 1 0 32384 0 1 26656
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__B
timestamp 1606120353
transform 1 0 32108 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A
timestamp 1606120353
transform 1 0 31740 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__A
timestamp 1606120353
transform 1 0 33488 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_335
timestamp 1606120353
transform 1 0 31924 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_45_339
timestamp 1606120353
transform 1 0 32292 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_45_347
timestamp 1606120353
transform 1 0 33028 0 1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_45_351
timestamp 1606120353
transform 1 0 33396 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0926_
timestamp 1606120353
transform 1 0 33764 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1196_
timestamp 1606120353
transform 1 0 34868 0 1 26656
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1606120353
transform 1 0 34776 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__D
timestamp 1606120353
transform 1 0 34592 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A
timestamp 1606120353
transform 1 0 34224 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_45_354
timestamp 1606120353
transform 1 0 33672 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_45_358
timestamp 1606120353
transform 1 0 34040 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_362
timestamp 1606120353
transform 1 0 34408 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A1
timestamp 1606120353
transform 1 0 36800 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_386
timestamp 1606120353
transform 1 0 36616 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_45_390
timestamp 1606120353
transform 1 0 36984 0 1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1606120353
transform -1 0 38548 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_45_402
timestamp 1606120353
transform 1 0 38088 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1180_
timestamp 1606120353
transform 1 0 1380 0 -1 27744
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1606120353
transform 1 0 1104 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1606120353
transform 1 0 1104 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__D
timestamp 1606120353
transform 1 0 1564 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__CLK
timestamp 1606120353
transform 1 0 1932 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_22
timestamp 1606120353
transform 1 0 3128 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1606120353
transform 1 0 1380 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_7
timestamp 1606120353
transform 1 0 1748 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_47_11
timestamp 1606120353
transform 1 0 2116 0 1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_46_32
timestamp 1606120353
transform 1 0 4048 0 -1 27744
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_46_30
timestamp 1606120353
transform 1 0 3864 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_46_26
timestamp 1606120353
transform 1 0 3496 0 -1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__B1
timestamp 1606120353
transform 1 0 3312 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1606120353
transform 1 0 3956 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_47_41
timestamp 1606120353
transform 1 0 4876 0 1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_47_35
timestamp 1606120353
transform 1 0 4324 0 1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_46_40
timestamp 1606120353
transform 1 0 4784 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A
timestamp 1606120353
transform 1 0 4692 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__B2
timestamp 1606120353
transform 1 0 4968 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_47_23
timestamp 1606120353
transform 1 0 3220 0 1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__a32oi_4  _0658_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 5152 0 -1 27744
box 0 -48 2024 592
use sky130_fd_sc_hd__fill_2  FILLER_47_47
timestamp 1606120353
transform 1 0 5428 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__C1
timestamp 1606120353
transform 1 0 5244 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_51
timestamp 1606120353
transform 1 0 5796 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__A2
timestamp 1606120353
transform 1 0 5612 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_55
timestamp 1606120353
transform 1 0 6164 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__B1
timestamp 1606120353
transform 1 0 5980 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_59
timestamp 1606120353
transform 1 0 6532 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__A1
timestamp 1606120353
transform 1 0 6348 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_47_62
timestamp 1606120353
transform 1 0 6808 0 1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1606120353
transform 1 0 6716 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_47_66
timestamp 1606120353
transform 1 0 7176 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_46_66
timestamp 1606120353
transform 1 0 7176 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_47_76
timestamp 1606120353
transform 1 0 8096 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_47_72
timestamp 1606120353
transform 1 0 7728 0 1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_46_71
timestamp 1606120353
transform 1 0 7636 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__A
timestamp 1606120353
transform 1 0 7820 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0550__A
timestamp 1606120353
transform 1 0 7452 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0549__A
timestamp 1606120353
transform 1 0 7268 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__A2
timestamp 1606120353
transform 1 0 8188 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _0659_
timestamp 1606120353
transform 1 0 8004 0 -1 27744
box 0 -48 644 592
use sky130_fd_sc_hd__buf_1  _0550_
timestamp 1606120353
transform 1 0 7452 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_47_79
timestamp 1606120353
transform 1 0 8372 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_86
timestamp 1606120353
transform 1 0 9016 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1606120353
transform 1 0 8648 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__B2
timestamp 1606120353
transform 1 0 9200 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__B1_N
timestamp 1606120353
transform 1 0 8832 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__A1
timestamp 1606120353
transform 1 0 8556 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0660_
timestamp 1606120353
transform 1 0 8740 0 1 27744
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_46_90
timestamp 1606120353
transform 1 0 9384 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1606120353
transform 1 0 9568 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_47_96
timestamp 1606120353
transform 1 0 9936 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_93
timestamp 1606120353
transform 1 0 9660 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__A1
timestamp 1606120353
transform 1 0 9844 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_100
timestamp 1606120353
transform 1 0 10304 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_46_97
timestamp 1606120353
transform 1 0 10028 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__A2
timestamp 1606120353
transform 1 0 10304 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__A1
timestamp 1606120353
transform 1 0 10120 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_104
timestamp 1606120353
transform 1 0 10672 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_102
timestamp 1606120353
transform 1 0 10488 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__B1
timestamp 1606120353
transform 1 0 10672 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__B1
timestamp 1606120353
transform 1 0 10488 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_108
timestamp 1606120353
transform 1 0 11040 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_106
timestamp 1606120353
transform 1 0 10856 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A2
timestamp 1606120353
transform 1 0 10856 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A2
timestamp 1606120353
transform 1 0 11040 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_46_110
timestamp 1606120353
transform 1 0 11224 0 -1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__A2
timestamp 1606120353
transform 1 0 11224 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_47_118
timestamp 1606120353
transform 1 0 11960 0 1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_47_112
timestamp 1606120353
transform 1 0 11408 0 1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0492__A
timestamp 1606120353
transform 1 0 11776 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0492__D
timestamp 1606120353
transform 1 0 11592 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0492_
timestamp 1606120353
transform 1 0 11776 0 -1 27744
box 0 -48 828 592
use sky130_fd_sc_hd__decap_4  FILLER_47_127
timestamp 1606120353
transform 1 0 12788 0 1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_47_123
timestamp 1606120353
transform 1 0 12420 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_46_125
timestamp 1606120353
transform 1 0 12604 0 -1 27744
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__A
timestamp 1606120353
transform 1 0 12604 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1606120353
transform 1 0 12328 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__B1_N
timestamp 1606120353
transform 1 0 13156 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_140
timestamp 1606120353
transform 1 0 13984 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_136
timestamp 1606120353
transform 1 0 13616 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A1
timestamp 1606120353
transform 1 0 14168 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0493__A
timestamp 1606120353
transform 1 0 13800 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0501_
timestamp 1606120353
transform 1 0 13340 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_47_146
timestamp 1606120353
transform 1 0 14536 0 1 27744
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_46_152
timestamp 1606120353
transform 1 0 15088 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_46_144
timestamp 1606120353
transform 1 0 14352 0 -1 27744
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__D
timestamp 1606120353
transform 1 0 15272 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1606120353
transform 1 0 15180 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0497_
timestamp 1606120353
transform 1 0 15272 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__a21bo_4  _0934_
timestamp 1606120353
transform 1 0 13340 0 1 27744
box 0 -48 1196 592
use sky130_fd_sc_hd__dfxtp_4  _1098_
timestamp 1606120353
transform 1 0 16284 0 -1 27744
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__CLK
timestamp 1606120353
transform 1 0 15640 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_46_157
timestamp 1606120353
transform 1 0 15548 0 -1 27744
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_47_156
timestamp 1606120353
transform 1 0 15456 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_47_160
timestamp 1606120353
transform 1 0 15824 0 1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_47_172
timestamp 1606120353
transform 1 0 16928 0 1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_47_176
timestamp 1606120353
transform 1 0 17296 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_47_184
timestamp 1606120353
transform 1 0 18032 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_179
timestamp 1606120353
transform 1 0 17572 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_46_184
timestamp 1606120353
transform 1 0 18032 0 -1 27744
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__CLK
timestamp 1606120353
transform 1 0 17388 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__D
timestamp 1606120353
transform 1 0 17756 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__B1
timestamp 1606120353
transform 1 0 18216 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1606120353
transform 1 0 17940 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_47_188
timestamp 1606120353
transform 1 0 18400 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_195
timestamp 1606120353
transform 1 0 19044 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A2
timestamp 1606120353
transform 1 0 19228 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__A1
timestamp 1606120353
transform 1 0 18584 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0664_
timestamp 1606120353
transform 1 0 18768 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__a21o_4  _0756_
timestamp 1606120353
transform 1 0 18768 0 1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_47_208
timestamp 1606120353
transform 1 0 20240 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_204
timestamp 1606120353
transform 1 0 19872 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__A2
timestamp 1606120353
transform 1 0 20056 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_212
timestamp 1606120353
transform 1 0 20608 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_219
timestamp 1606120353
transform 1 0 21252 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_215
timestamp 1606120353
transform 1 0 20884 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_46_211
timestamp 1606120353
transform 1 0 20516 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A1
timestamp 1606120353
transform 1 0 21068 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__B1
timestamp 1606120353
transform 1 0 20424 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A2
timestamp 1606120353
transform 1 0 20792 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1606120353
transform 1 0 20792 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_46_199
timestamp 1606120353
transform 1 0 19412 0 -1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__o21a_4  _0870_
timestamp 1606120353
transform 1 0 20976 0 1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_47_228
timestamp 1606120353
transform 1 0 22080 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_46_223
timestamp 1606120353
transform 1 0 21620 0 -1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A1
timestamp 1606120353
transform 1 0 21988 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A2
timestamp 1606120353
transform 1 0 21436 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0848_
timestamp 1606120353
transform 1 0 22172 0 -1 27744
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_47_236
timestamp 1606120353
transform 1 0 22816 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_232
timestamp 1606120353
transform 1 0 22448 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_46_238
timestamp 1606120353
transform 1 0 23000 0 -1 27744
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A1
timestamp 1606120353
transform 1 0 23000 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A2
timestamp 1606120353
transform 1 0 22632 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__B1_N
timestamp 1606120353
transform 1 0 22264 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_240
timestamp 1606120353
transform 1 0 23184 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__A
timestamp 1606120353
transform 1 0 23368 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A1
timestamp 1606120353
transform 1 0 23552 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1606120353
transform 1 0 23552 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__nor2_4  _0914_
timestamp 1606120353
transform 1 0 23644 0 1 27744
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILLER_47_258
timestamp 1606120353
transform 1 0 24840 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_47_254
timestamp 1606120353
transform 1 0 24472 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_46_259
timestamp 1606120353
transform 1 0 24932 0 -1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__B
timestamp 1606120353
transform 1 0 25300 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A2
timestamp 1606120353
transform 1 0 24656 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A
timestamp 1606120353
transform 1 0 25116 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0897_
timestamp 1606120353
transform 1 0 25300 0 1 27744
box 0 -48 828 592
use sky130_fd_sc_hd__a21bo_4  _0938_
timestamp 1606120353
transform 1 0 23736 0 -1 27744
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_4  FILLER_47_272
timestamp 1606120353
transform 1 0 26128 0 1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_46_271
timestamp 1606120353
transform 1 0 26036 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_46_265
timestamp 1606120353
transform 1 0 25484 0 -1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__D
timestamp 1606120353
transform 1 0 25852 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__D
timestamp 1606120353
transform 1 0 26220 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_47_278
timestamp 1606120353
transform 1 0 26680 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_46_276
timestamp 1606120353
transform 1 0 26496 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__B
timestamp 1606120353
transform 1 0 26680 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__A
timestamp 1606120353
transform 1 0 26956 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__A
timestamp 1606120353
transform 1 0 26496 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1606120353
transform 1 0 26404 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0890_
timestamp 1606120353
transform 1 0 26864 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_46_283
timestamp 1606120353
transform 1 0 27140 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__A
timestamp 1606120353
transform 1 0 27324 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0891_
timestamp 1606120353
transform 1 0 27140 0 1 27744
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_47_296
timestamp 1606120353
transform 1 0 28336 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_292
timestamp 1606120353
transform 1 0 27968 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_287
timestamp 1606120353
transform 1 0 27508 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__C
timestamp 1606120353
transform 1 0 27692 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__C
timestamp 1606120353
transform 1 0 28152 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_306
timestamp 1606120353
transform 1 0 29256 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_300
timestamp 1606120353
transform 1 0 28704 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_308
timestamp 1606120353
transform 1 0 29440 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_304
timestamp 1606120353
transform 1 0 29072 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__B1
timestamp 1606120353
transform 1 0 29256 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__A2
timestamp 1606120353
transform 1 0 28520 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A2
timestamp 1606120353
transform 1 0 29440 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_clk
timestamp 1606120353
transform 1 0 28888 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1606120353
transform 1 0 29164 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__a21bo_4  _0894_
timestamp 1606120353
transform 1 0 27876 0 -1 27744
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_47_310
timestamp 1606120353
transform 1 0 29624 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_317
timestamp 1606120353
transform 1 0 30268 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_46_312
timestamp 1606120353
transform 1 0 29808 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_clk_A
timestamp 1606120353
transform 1 0 29624 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__B1
timestamp 1606120353
transform 1 0 30084 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__B1
timestamp 1606120353
transform 1 0 29808 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0827_
timestamp 1606120353
transform 1 0 30452 0 -1 27744
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_47_330
timestamp 1606120353
transform 1 0 31464 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_326
timestamp 1606120353
transform 1 0 31096 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_328
timestamp 1606120353
transform 1 0 31280 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_clk_A
timestamp 1606120353
transform 1 0 31464 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A
timestamp 1606120353
transform 1 0 31280 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0865_
timestamp 1606120353
transform 1 0 29992 0 1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_47_334
timestamp 1606120353
transform 1 0 31832 0 1 27744
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILLER_46_332
timestamp 1606120353
transform 1 0 31648 0 -1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__B
timestamp 1606120353
transform 1 0 31648 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1606120353
transform 1 0 32016 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _0828_
timestamp 1606120353
transform 1 0 32108 0 -1 27744
box 0 -48 644 592
use sky130_fd_sc_hd__fill_1  FILLER_47_340
timestamp 1606120353
transform 1 0 32384 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_46_344
timestamp 1606120353
transform 1 0 32752 0 -1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A2
timestamp 1606120353
transform 1 0 33120 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A
timestamp 1606120353
transform 1 0 32476 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0922_
timestamp 1606120353
transform 1 0 32660 0 1 27744
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_47_352
timestamp 1606120353
transform 1 0 33488 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_350
timestamp 1606120353
transform 1 0 33304 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0932_
timestamp 1606120353
transform 1 0 33488 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_47_360
timestamp 1606120353
transform 1 0 34224 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_356
timestamp 1606120353
transform 1 0 33856 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_46_355
timestamp 1606120353
transform 1 0 33764 0 -1 27744
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__C1
timestamp 1606120353
transform 1 0 34040 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__B1
timestamp 1606120353
transform 1 0 33672 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_47_367
timestamp 1606120353
transform 1 0 34868 0 1 27744
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_47_364
timestamp 1606120353
transform 1 0 34592 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_366
timestamp 1606120353
transform 1 0 34776 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__CLK
timestamp 1606120353
transform 1 0 34960 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A1
timestamp 1606120353
transform 1 0 34408 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1606120353
transform 1 0 34776 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0876_
timestamp 1606120353
transform 1 0 34500 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_46_370
timestamp 1606120353
transform 1 0 35144 0 -1 27744
box 0 -48 552 592
use sky130_fd_sc_hd__a21bo_4  _0937_
timestamp 1606120353
transform 1 0 35696 0 -1 27744
box 0 -48 1196 592
use sky130_fd_sc_hd__dfxtp_4  _1225_
timestamp 1606120353
transform 1 0 35788 0 1 27744
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__D
timestamp 1606120353
transform 1 0 35604 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_46_389
timestamp 1606120353
transform 1 0 36892 0 -1 27744
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_47_396
timestamp 1606120353
transform 1 0 37536 0 1 27744
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1606120353
transform -1 0 38548 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1606120353
transform -1 0 38548 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1606120353
transform 1 0 37628 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_46_398
timestamp 1606120353
transform 1 0 37720 0 -1 27744
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1126_
timestamp 1606120353
transform 1 0 1472 0 -1 28832
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1606120353
transform 1 0 1104 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_48_3
timestamp 1606120353
transform 1 0 1380 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0779_
timestamp 1606120353
transform 1 0 4692 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1606120353
transform 1 0 3956 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_48_23
timestamp 1606120353
transform 1 0 3220 0 -1 28832
box 0 -48 736 592
use sky130_fd_sc_hd__decap_6  FILLER_48_32
timestamp 1606120353
transform 1 0 4048 0 -1 28832
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_48_38
timestamp 1606120353
transform 1 0 4600 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_48_42
timestamp 1606120353
transform 1 0 4968 0 -1 28832
box 0 -48 736 592
use sky130_fd_sc_hd__a211o_4  _0650_
timestamp 1606120353
transform 1 0 5980 0 -1 28832
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  FILLER_48_50
timestamp 1606120353
transform 1 0 5704 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _0549_
timestamp 1606120353
transform 1 0 8004 0 -1 28832
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A3
timestamp 1606120353
transform 1 0 9016 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_48_67
timestamp 1606120353
transform 1 0 7268 0 -1 28832
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_48_84
timestamp 1606120353
transform 1 0 8832 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_48_88
timestamp 1606120353
transform 1 0 9200 0 -1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__a21o_4  _0666_
timestamp 1606120353
transform 1 0 10120 0 -1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1606120353
transform 1 0 9568 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_48_93
timestamp 1606120353
transform 1 0 9660 0 -1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_48_97
timestamp 1606120353
transform 1 0 10028 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_48_110
timestamp 1606120353
transform 1 0 11224 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0651_
timestamp 1606120353
transform 1 0 12236 0 -1 28832
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__A
timestamp 1606120353
transform 1 0 11408 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_48_114
timestamp 1606120353
transform 1 0 11592 0 -1 28832
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_48_120
timestamp 1606120353
transform 1 0 12144 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_48_130
timestamp 1606120353
transform 1 0 13064 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0493_
timestamp 1606120353
transform 1 0 13800 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1156_
timestamp 1606120353
transform 1 0 15272 0 -1 28832
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1606120353
transform 1 0 15180 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A2
timestamp 1606120353
transform 1 0 13340 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__CLK
timestamp 1606120353
transform 1 0 14260 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_48_135
timestamp 1606120353
transform 1 0 13524 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1606120353
transform 1 0 14076 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_48_145
timestamp 1606120353
transform 1 0 14444 0 -1 28832
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_48_173
timestamp 1606120353
transform 1 0 17020 0 -1 28832
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1087_
timestamp 1606120353
transform 1 0 17756 0 -1 28832
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1606120353
transform 1 0 20792 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A1
timestamp 1606120353
transform 1 0 20332 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A
timestamp 1606120353
transform 1 0 19688 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_200
timestamp 1606120353
transform 1 0 19504 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_48_204
timestamp 1606120353
transform 1 0 19872 0 -1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_48_208
timestamp 1606120353
transform 1 0 20240 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_48_211
timestamp 1606120353
transform 1 0 20516 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_48_215
timestamp 1606120353
transform 1 0 20884 0 -1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__a21bo_4  _0924_
timestamp 1606120353
transform 1 0 21988 0 -1 28832
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_4  FILLER_48_240
timestamp 1606120353
transform 1 0 23184 0 -1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__a21o_4  _0913_
timestamp 1606120353
transform 1 0 24472 0 -1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__B1
timestamp 1606120353
transform 1 0 24288 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__B
timestamp 1606120353
transform 1 0 23644 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_48_244
timestamp 1606120353
transform 1 0 23552 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_48_247
timestamp 1606120353
transform 1 0 23828 0 -1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1606120353
transform 1 0 24196 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0895_
timestamp 1606120353
transform 1 0 26496 0 -1 28832
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1606120353
transform 1 0 26404 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A1
timestamp 1606120353
transform 1 0 26220 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_48_266
timestamp 1606120353
transform 1 0 25576 0 -1 28832
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_48_272
timestamp 1606120353
transform 1 0 26128 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_48_285
timestamp 1606120353
transform 1 0 27324 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0892_
timestamp 1606120353
transform 1 0 28152 0 -1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__A
timestamp 1606120353
transform 1 0 27968 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__B
timestamp 1606120353
transform 1 0 27508 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__A1
timestamp 1606120353
transform 1 0 29440 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_48_289
timestamp 1606120353
transform 1 0 27692 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_48_306
timestamp 1606120353
transform 1 0 29256 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0893_
timestamp 1606120353
transform 1 0 29992 0 -1 28832
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__A2
timestamp 1606120353
transform 1 0 31096 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A1
timestamp 1606120353
transform 1 0 29808 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_310
timestamp 1606120353
transform 1 0 29624 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_48_323
timestamp 1606120353
transform 1 0 30820 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_48_328
timestamp 1606120353
transform 1 0 31280 0 -1 28832
box 0 -48 736 592
use sky130_fd_sc_hd__a211o_4  _0923_
timestamp 1606120353
transform 1 0 33120 0 -1 28832
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1606120353
transform 1 0 32016 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__B
timestamp 1606120353
transform 1 0 32660 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_48_337
timestamp 1606120353
transform 1 0 32108 0 -1 28832
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILLER_48_345
timestamp 1606120353
transform 1 0 32844 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__D
timestamp 1606120353
transform 1 0 35144 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_48_362
timestamp 1606120353
transform 1 0 34408 0 -1 28832
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_48_372
timestamp 1606120353
transform 1 0 35328 0 -1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__CLK
timestamp 1606120353
transform 1 0 35788 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_48_376
timestamp 1606120353
transform 1 0 35696 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_48_379
timestamp 1606120353
transform 1 0 35972 0 -1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_48_391
timestamp 1606120353
transform 1 0 37076 0 -1 28832
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1606120353
transform -1 0 38548 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1606120353
transform 1 0 37628 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_48_398
timestamp 1606120353
transform 1 0 37720 0 -1 28832
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1606120353
transform 1 0 1104 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__D
timestamp 1606120353
transform 1 0 3128 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__D
timestamp 1606120353
transform 1 0 1564 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__CLK
timestamp 1606120353
transform 1 0 1932 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1606120353
transform 1 0 1380 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_7
timestamp 1606120353
transform 1 0 1748 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_49_11
timestamp 1606120353
transform 1 0 2116 0 1 28832
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_49_19
timestamp 1606120353
transform 1 0 2852 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1115_
timestamp 1606120353
transform 1 0 3312 0 1 28832
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_12  FILLER_49_43
timestamp 1606120353
transform 1 0 5060 0 1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1606120353
transform 1 0 6716 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__A1
timestamp 1606120353
transform 1 0 6992 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_49_55
timestamp 1606120353
transform 1 0 6164 0 1 28832
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_49_62
timestamp 1606120353
transform 1 0 6808 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_66
timestamp 1606120353
transform 1 0 7176 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1083_
timestamp 1606120353
transform 1 0 8556 0 1 28832
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__A2
timestamp 1606120353
transform 1 0 7360 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__B1
timestamp 1606120353
transform 1 0 7728 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__D
timestamp 1606120353
transform 1 0 8372 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_70
timestamp 1606120353
transform 1 0 7544 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_49_74
timestamp 1606120353
transform 1 0 7912 0 1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_49_78
timestamp 1606120353
transform 1 0 8280 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0548__A
timestamp 1606120353
transform 1 0 11132 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__B
timestamp 1606120353
transform 1 0 10488 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_100
timestamp 1606120353
transform 1 0 10304 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_49_104
timestamp 1606120353
transform 1 0 10672 0 1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_49_108
timestamp 1606120353
transform 1 0 11040 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0548_
timestamp 1606120353
transform 1 0 11316 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_49_114
timestamp 1606120353
transform 1 0 11592 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__B
timestamp 1606120353
transform 1 0 11776 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_118
timestamp 1606120353
transform 1 0 11960 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__C
timestamp 1606120353
transform 1 0 12144 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1606120353
transform 1 0 12328 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_49_123
timestamp 1606120353
transform 1 0 12420 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0498__A
timestamp 1606120353
transform 1 0 12604 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0500_
timestamp 1606120353
transform 1 0 12788 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_49_130
timestamp 1606120353
transform 1 0 13064 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0500__A
timestamp 1606120353
transform 1 0 13248 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1148_
timestamp 1606120353
transform 1 0 13800 0 1 28832
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__D
timestamp 1606120353
transform 1 0 13616 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_134
timestamp 1606120353
transform 1 0 13432 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__D
timestamp 1606120353
transform 1 0 16192 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__CLK
timestamp 1606120353
transform 1 0 16560 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_49_157
timestamp 1606120353
transform 1 0 15548 0 1 28832
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_49_163
timestamp 1606120353
transform 1 0 16100 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1606120353
transform 1 0 16376 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_49_170
timestamp 1606120353
transform 1 0 16744 0 1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__and2_4  _0755_
timestamp 1606120353
transform 1 0 18768 0 1 28832
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1606120353
transform 1 0 17940 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__B
timestamp 1606120353
transform 1 0 18584 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_49_182
timestamp 1606120353
transform 1 0 17848 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_49_184
timestamp 1606120353
transform 1 0 18032 0 1 28832
box 0 -48 552 592
use sky130_fd_sc_hd__o21ai_4  _0871_
timestamp 1606120353
transform 1 0 20332 0 1 28832
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A
timestamp 1606120353
transform 1 0 19596 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A2
timestamp 1606120353
transform 1 0 20148 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_199
timestamp 1606120353
transform 1 0 19412 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_49_203
timestamp 1606120353
transform 1 0 19780 0 1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_49_222
timestamp 1606120353
transform 1 0 21528 0 1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_49_226
timestamp 1606120353
transform 1 0 21896 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A1
timestamp 1606120353
transform 1 0 21988 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_229
timestamp 1606120353
transform 1 0 22172 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A2
timestamp 1606120353
transform 1 0 22356 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_233
timestamp 1606120353
transform 1 0 22540 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__B1_N
timestamp 1606120353
transform 1 0 22724 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_49_237
timestamp 1606120353
transform 1 0 22908 0 1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_49_241
timestamp 1606120353
transform 1 0 23276 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__B1_N
timestamp 1606120353
transform 1 0 23368 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0912_
timestamp 1606120353
transform 1 0 24840 0 1 28832
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1606120353
transform 1 0 23552 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A2
timestamp 1606120353
transform 1 0 24288 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__A
timestamp 1606120353
transform 1 0 24656 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__B
timestamp 1606120353
transform 1 0 23920 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_49_245
timestamp 1606120353
transform 1 0 23644 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_49_250
timestamp 1606120353
transform 1 0 24104 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_254
timestamp 1606120353
transform 1 0 24472 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_267
timestamp 1606120353
transform 1 0 25668 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__C
timestamp 1606120353
transform 1 0 25852 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_271
timestamp 1606120353
transform 1 0 26036 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__D
timestamp 1606120353
transform 1 0 26220 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0884_
timestamp 1606120353
transform 1 0 26404 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1606120353
transform 1 0 26680 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_282
timestamp 1606120353
transform 1 0 27048 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A
timestamp 1606120353
transform 1 0 26864 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__A
timestamp 1606120353
transform 1 0 27232 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0886_
timestamp 1606120353
transform 1 0 27416 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__o21a_4  _0860_
timestamp 1606120353
transform 1 0 29256 0 1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1606120353
transform 1 0 29164 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__B1
timestamp 1606120353
transform 1 0 28980 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A2
timestamp 1606120353
transform 1 0 28612 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__C
timestamp 1606120353
transform 1 0 27968 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_49_289
timestamp 1606120353
transform 1 0 27692 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_49_294
timestamp 1606120353
transform 1 0 28152 0 1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_49_298
timestamp 1606120353
transform 1 0 28520 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_49_301
timestamp 1606120353
transform 1 0 28796 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0829_
timestamp 1606120353
transform 1 0 31096 0 1 28832
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__A
timestamp 1606120353
transform 1 0 30544 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__A1
timestamp 1606120353
transform 1 0 30912 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_318
timestamp 1606120353
transform 1 0 30360 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_322
timestamp 1606120353
transform 1 0 30728 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_49_339
timestamp 1606120353
transform 1 0 32292 0 1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_49_351
timestamp 1606120353
transform 1 0 33396 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1187_
timestamp 1606120353
transform 1 0 35144 0 1 28832
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1606120353
transform 1 0 34776 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__B1_N
timestamp 1606120353
transform 1 0 33948 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A2
timestamp 1606120353
transform 1 0 34316 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A1
timestamp 1606120353
transform 1 0 33580 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_355
timestamp 1606120353
transform 1 0 33764 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_359
timestamp 1606120353
transform 1 0 34132 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_49_363
timestamp 1606120353
transform 1 0 34500 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_49_367
timestamp 1606120353
transform 1 0 34868 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_49_389
timestamp 1606120353
transform 1 0 36892 0 1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1606120353
transform -1 0 38548 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_49_401
timestamp 1606120353
transform 1 0 37996 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1164_
timestamp 1606120353
transform 1 0 1380 0 -1 29920
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1606120353
transform 1 0 1104 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_50_22
timestamp 1606120353
transform 1 0 3128 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1606120353
transform 1 0 3956 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__CLK
timestamp 1606120353
transform 1 0 3312 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_50_26
timestamp 1606120353
transform 1 0 3496 0 -1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_50_30
timestamp 1606120353
transform 1 0 3864 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_50_32
timestamp 1606120353
transform 1 0 4048 0 -1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_50_44
timestamp 1606120353
transform 1 0 5152 0 -1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__o21ai_4  _0621_
timestamp 1606120353
transform 1 0 6992 0 -1 29920
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__B1
timestamp 1606120353
transform 1 0 6808 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_50_56
timestamp 1606120353
transform 1 0 6256 0 -1 29920
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__CLK
timestamp 1606120353
transform 1 0 8556 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_50_77
timestamp 1606120353
transform 1 0 8188 0 -1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_50_83
timestamp 1606120353
transform 1 0 8740 0 -1 29920
box 0 -48 736 592
use sky130_fd_sc_hd__and2_4  _0665_
timestamp 1606120353
transform 1 0 10028 0 -1 29920
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1606120353
transform 1 0 9568 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__A
timestamp 1606120353
transform 1 0 10856 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_50_91
timestamp 1606120353
transform 1 0 9476 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_50_93
timestamp 1606120353
transform 1 0 9660 0 -1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_50_104
timestamp 1606120353
transform 1 0 10672 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_50_108
timestamp 1606120353
transform 1 0 11040 0 -1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _0498_
timestamp 1606120353
transform 1 0 12972 0 -1 29920
box 0 -48 828 592
use sky130_fd_sc_hd__or3_4  _0547_
timestamp 1606120353
transform 1 0 11408 0 -1 29920
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0499__B
timestamp 1606120353
transform 1 0 12420 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__A
timestamp 1606120353
transform 1 0 12788 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_121
timestamp 1606120353
transform 1 0 12236 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_125
timestamp 1606120353
transform 1 0 12604 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1606120353
transform 1 0 15180 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_clk_A
timestamp 1606120353
transform 1 0 13984 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1606120353
transform 1 0 13800 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_50_142
timestamp 1606120353
transform 1 0 14168 0 -1 29920
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_50_150
timestamp 1606120353
transform 1 0 14904 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_50_154
timestamp 1606120353
transform 1 0 15272 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1089_
timestamp 1606120353
transform 1 0 16192 0 -1 29920
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__CLK
timestamp 1606120353
transform 1 0 15456 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_50_158
timestamp 1606120353
transform 1 0 15640 0 -1 29920
box 0 -48 552 592
use sky130_fd_sc_hd__inv_8  _0869_
timestamp 1606120353
transform 1 0 19228 0 -1 29920
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__B1
timestamp 1606120353
transform 1 0 18124 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__A2
timestamp 1606120353
transform 1 0 18492 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__CLK
timestamp 1606120353
transform 1 0 19044 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_183
timestamp 1606120353
transform 1 0 17940 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_187
timestamp 1606120353
transform 1 0 18308 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_50_191
timestamp 1606120353
transform 1 0 18676 0 -1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1606120353
transform 1 0 20792 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__B1
timestamp 1606120353
transform 1 0 20332 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__CLK
timestamp 1606120353
transform 1 0 21344 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_50_206
timestamp 1606120353
transform 1 0 20056 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_50_211
timestamp 1606120353
transform 1 0 20516 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_50_215
timestamp 1606120353
transform 1 0 20884 0 -1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_50_219
timestamp 1606120353
transform 1 0 21252 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__a21bo_4  _0919_
timestamp 1606120353
transform 1 0 22356 0 -1 29920
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__B
timestamp 1606120353
transform 1 0 21988 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_50_222
timestamp 1606120353
transform 1 0 21528 0 -1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_50_226
timestamp 1606120353
transform 1 0 21896 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_50_229
timestamp 1606120353
transform 1 0 22172 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0939_
timestamp 1606120353
transform 1 0 24288 0 -1 29920
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__B1
timestamp 1606120353
transform 1 0 24104 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A1
timestamp 1606120353
transform 1 0 23736 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_244
timestamp 1606120353
transform 1 0 23552 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_248
timestamp 1606120353
transform 1 0 23920 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_265
timestamp 1606120353
transform 1 0 25484 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__C
timestamp 1606120353
transform 1 0 25668 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_269
timestamp 1606120353
transform 1 0 25852 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_273
timestamp 1606120353
transform 1 0 26220 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A1
timestamp 1606120353
transform 1 0 26036 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1606120353
transform 1 0 26404 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0882_
timestamp 1606120353
transform 1 0 26496 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_50_279
timestamp 1606120353
transform 1 0 26772 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__A
timestamp 1606120353
transform 1 0 27048 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_284
timestamp 1606120353
transform 1 0 27232 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A
timestamp 1606120353
transform 1 0 27416 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__nor3_4  _0888_
timestamp 1606120353
transform 1 0 27968 0 -1 29920
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A1
timestamp 1606120353
transform 1 0 29348 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__B
timestamp 1606120353
transform 1 0 27784 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_288
timestamp 1606120353
transform 1 0 27600 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_305
timestamp 1606120353
transform 1 0 29164 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0880_
timestamp 1606120353
transform 1 0 29900 0 -1 29920
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__B1_N
timestamp 1606120353
transform 1 0 31096 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__B
timestamp 1606120353
transform 1 0 30728 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A2
timestamp 1606120353
transform 1 0 29716 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1606120353
transform 1 0 29532 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_320
timestamp 1606120353
transform 1 0 30544 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_324
timestamp 1606120353
transform 1 0 30912 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_50_328
timestamp 1606120353
transform 1 0 31280 0 -1 29920
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1606120353
transform 1 0 32016 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__B1
timestamp 1606120353
transform 1 0 32292 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_337
timestamp 1606120353
transform 1 0 32108 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_50_341
timestamp 1606120353
transform 1 0 32476 0 -1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__a21bo_4  _0928_
timestamp 1606120353
transform 1 0 33948 0 -1 29920
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__CLK
timestamp 1606120353
transform 1 0 35328 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_50_353
timestamp 1606120353
transform 1 0 33580 0 -1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_50_370
timestamp 1606120353
transform 1 0 35144 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_50_374
timestamp 1606120353
transform 1 0 35512 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__CLK
timestamp 1606120353
transform 1 0 35788 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_50_379
timestamp 1606120353
transform 1 0 35972 0 -1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_50_391
timestamp 1606120353
transform 1 0 37076 0 -1 29920
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1606120353
transform -1 0 38548 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1606120353
transform 1 0 37628 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_50_398
timestamp 1606120353
transform 1 0 37720 0 -1 29920
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1092_
timestamp 1606120353
transform 1 0 3128 0 1 29920
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1606120353
transform 1 0 1104 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__D
timestamp 1606120353
transform 1 0 2944 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__CLK
timestamp 1606120353
transform 1 0 2576 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1606120353
transform 1 0 1380 0 1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_51_15
timestamp 1606120353
transform 1 0 2484 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_51_18
timestamp 1606120353
transform 1 0 2760 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_51_41
timestamp 1606120353
transform 1 0 4876 0 1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__o21a_4  _0623_
timestamp 1606120353
transform 1 0 6808 0 1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1606120353
transform 1 0 6716 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__A2
timestamp 1606120353
transform 1 0 6532 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_51_53
timestamp 1606120353
transform 1 0 5980 0 1 29920
box 0 -48 552 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_clk
timestamp 1606120353
transform 1 0 8648 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_clk_A
timestamp 1606120353
transform 1 0 9108 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_51_74
timestamp 1606120353
transform 1 0 7912 0 1 29920
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_51_85
timestamp 1606120353
transform 1 0 8924 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__nand3_4  _0622_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 10304 0 1 29920
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__B
timestamp 1606120353
transform 1 0 10120 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__A
timestamp 1606120353
transform 1 0 9752 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_51_89
timestamp 1606120353
transform 1 0 9292 0 1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_51_93
timestamp 1606120353
transform 1 0 9660 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_51_96
timestamp 1606120353
transform 1 0 9936 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__or3_4  _0499_
timestamp 1606120353
transform 1 0 12420 0 1 29920
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1606120353
transform 1 0 12328 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0499__C
timestamp 1606120353
transform 1 0 12144 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0488__A
timestamp 1606120353
transform 1 0 11776 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_114
timestamp 1606120353
transform 1 0 11592 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_118
timestamp 1606120353
transform 1 0 11960 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_132
timestamp 1606120353
transform 1 0 13248 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0748_
timestamp 1606120353
transform 1 0 14720 0 1 29920
box 0 -48 644 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_clk
timestamp 1606120353
transform 1 0 13984 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__C
timestamp 1606120353
transform 1 0 13432 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__B
timestamp 1606120353
transform 1 0 14536 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__B
timestamp 1606120353
transform 1 0 13800 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_136
timestamp 1606120353
transform 1 0 13616 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_51_143
timestamp 1606120353
transform 1 0 14260 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__A
timestamp 1606120353
transform 1 0 15548 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__D
timestamp 1606120353
transform 1 0 15916 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_155
timestamp 1606120353
transform 1 0 15364 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_159
timestamp 1606120353
transform 1 0 15732 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_51_163
timestamp 1606120353
transform 1 0 16100 0 1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_51_175
timestamp 1606120353
transform 1 0 17204 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0769_
timestamp 1606120353
transform 1 0 18032 0 1 29920
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1606120353
transform 1 0 17940 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__D
timestamp 1606120353
transform 1 0 19228 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A
timestamp 1606120353
transform 1 0 18860 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__A1
timestamp 1606120353
transform 1 0 17756 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__B
timestamp 1606120353
transform 1 0 17388 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_179
timestamp 1606120353
transform 1 0 17572 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_191
timestamp 1606120353
transform 1 0 18676 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_195
timestamp 1606120353
transform 1 0 19044 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1179_
timestamp 1606120353
transform 1 0 19412 0 1 29920
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__D
timestamp 1606120353
transform 1 0 21344 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_218
timestamp 1606120353
transform 1 0 21160 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0918_
timestamp 1606120353
transform 1 0 21988 0 1 29920
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__A
timestamp 1606120353
transform 1 0 21804 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__D
timestamp 1606120353
transform 1 0 23368 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_51_222
timestamp 1606120353
transform 1 0 21528 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_51_236
timestamp 1606120353
transform 1 0 22816 0 1 29920
box 0 -48 552 592
use sky130_fd_sc_hd__a21o_4  _0917_
timestamp 1606120353
transform 1 0 25024 0 1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1606120353
transform 1 0 23552 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A2
timestamp 1606120353
transform 1 0 24840 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A
timestamp 1606120353
transform 1 0 24472 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__B
timestamp 1606120353
transform 1 0 24104 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_51_245
timestamp 1606120353
transform 1 0 23644 0 1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_51_249
timestamp 1606120353
transform 1 0 24012 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_51_252
timestamp 1606120353
transform 1 0 24288 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_256
timestamp 1606120353
transform 1 0 24656 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0889_
timestamp 1606120353
transform 1 0 26864 0 1 29920
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A2
timestamp 1606120353
transform 1 0 26680 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__B
timestamp 1606120353
transform 1 0 26312 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_272
timestamp 1606120353
transform 1 0 26128 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_276
timestamp 1606120353
transform 1 0 26496 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0931_
timestamp 1606120353
transform 1 0 29256 0 1 29920
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1606120353
transform 1 0 29164 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_clk
timestamp 1606120353
transform 1 0 28796 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__C
timestamp 1606120353
transform 1 0 28244 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__B1_N
timestamp 1606120353
transform 1 0 28612 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_293
timestamp 1606120353
transform 1 0 28060 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_297
timestamp 1606120353
transform 1 0 28428 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_51_304
timestamp 1606120353
transform 1 0 29072 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A
timestamp 1606120353
transform 1 0 30636 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_clk_A
timestamp 1606120353
transform 1 0 31004 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_319
timestamp 1606120353
transform 1 0 30452 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_323
timestamp 1606120353
transform 1 0 30820 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_51_327
timestamp 1606120353
transform 1 0 31188 0 1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__o21ai_4  _0868_
timestamp 1606120353
transform 1 0 32200 0 1 29920
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A2
timestamp 1606120353
transform 1 0 32016 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A1
timestamp 1606120353
transform 1 0 31648 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_51_331
timestamp 1606120353
transform 1 0 31556 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1606120353
transform 1 0 31832 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_51_351
timestamp 1606120353
transform 1 0 33396 0 1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1606120353
transform 1 0 34776 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_51_363
timestamp 1606120353
transform 1 0 34500 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_51_367
timestamp 1606120353
transform 1 0 34868 0 1 29920
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1184_
timestamp 1606120353
transform 1 0 35788 0 1 29920
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__D
timestamp 1606120353
transform 1 0 35604 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_51_396
timestamp 1606120353
transform 1 0 37536 0 1 29920
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1606120353
transform -1 0 38548 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1606120353
transform 1 0 1104 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1606120353
transform 1 0 1104 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_53_18
timestamp 1606120353
transform 1 0 2760 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_53_15
timestamp 1606120353
transform 1 0 2484 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_52_21
timestamp 1606120353
transform 1 0 3036 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_52_15
timestamp 1606120353
transform 1 0 2484 0 -1 31008
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A2
timestamp 1606120353
transform 1 0 2576 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A1
timestamp 1606120353
transform 1 0 3128 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__B1
timestamp 1606120353
transform 1 0 2944 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1606120353
transform 1 0 1380 0 1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1606120353
transform 1 0 1380 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__o22a_4  _0782_
timestamp 1606120353
transform 1 0 3128 0 1 31008
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1606120353
transform 1 0 3956 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_52_24
timestamp 1606120353
transform 1 0 3312 0 -1 31008
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_52_30
timestamp 1606120353
transform 1 0 3864 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_52_32
timestamp 1606120353
transform 1 0 4048 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_52_44
timestamp 1606120353
transform 1 0 5152 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_53_36
timestamp 1606120353
transform 1 0 4416 0 1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1606120353
transform 1 0 6716 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__A1
timestamp 1606120353
transform 1 0 6808 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_52_56
timestamp 1606120353
transform 1 0 6256 0 -1 31008
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_52_64
timestamp 1606120353
transform 1 0 6992 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_53_48
timestamp 1606120353
transform 1 0 5520 0 1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_53_60
timestamp 1606120353
transform 1 0 6624 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_53_62
timestamp 1606120353
transform 1 0 6808 0 1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_52_76
timestamp 1606120353
transform 1 0 8096 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_52_88
timestamp 1606120353
transform 1 0 9200 0 -1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_53_74
timestamp 1606120353
transform 1 0 7912 0 1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_53_86
timestamp 1606120353
transform 1 0 9016 0 1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_53_98
timestamp 1606120353
transform 1 0 10120 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_52_99
timestamp 1606120353
transform 1 0 10212 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_52_93
timestamp 1606120353
transform 1 0 9660 0 -1 31008
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1606120353
transform 1 0 9568 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_53_103
timestamp 1606120353
transform 1 0 10580 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_52_110
timestamp 1606120353
transform 1 0 11224 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_52_102
timestamp 1606120353
transform 1 0 10488 0 -1 31008
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_clk_A
timestamp 1606120353
transform 1 0 10764 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__C
timestamp 1606120353
transform 1 0 10304 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_clk
timestamp 1606120353
transform 1 0 10304 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_53_107
timestamp 1606120353
transform 1 0 10948 0 1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_53_119
timestamp 1606120353
transform 1 0 12052 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_52_120
timestamp 1606120353
transform 1 0 12144 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _0488_
timestamp 1606120353
transform 1 0 11316 0 -1 31008
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILLER_53_123
timestamp 1606120353
transform 1 0 12420 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_52_125
timestamp 1606120353
transform 1 0 12604 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__D
timestamp 1606120353
transform 1 0 12696 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0499__A
timestamp 1606120353
transform 1 0 12420 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1606120353
transform 1 0 12328 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__and3_4  _0620_
timestamp 1606120353
transform 1 0 12880 0 -1 31008
box 0 -48 828 592
use sky130_fd_sc_hd__dfxtp_4  _1086_
timestamp 1606120353
transform 1 0 12880 0 1 31008
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1088_
timestamp 1606120353
transform 1 0 15272 0 -1 31008
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1606120353
transform 1 0 15180 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A
timestamp 1606120353
transform 1 0 13892 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__B
timestamp 1606120353
transform 1 0 14260 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_137
timestamp 1606120353
transform 1 0 13708 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1606120353
transform 1 0 14076 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_52_145
timestamp 1606120353
transform 1 0 14444 0 -1 31008
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_53_147
timestamp 1606120353
transform 1 0 14628 0 1 31008
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_53_160
timestamp 1606120353
transform 1 0 15824 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_53_155
timestamp 1606120353
transform 1 0 15364 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__B
timestamp 1606120353
transform 1 0 15640 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_164
timestamp 1606120353
transform 1 0 16192 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__B1
timestamp 1606120353
transform 1 0 16008 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__A1
timestamp 1606120353
transform 1 0 16376 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0763_
timestamp 1606120353
transform 1 0 16560 0 1 31008
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_53_175
timestamp 1606120353
transform 1 0 17204 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_173
timestamp 1606120353
transform 1 0 17020 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__A2
timestamp 1606120353
transform 1 0 17204 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_187
timestamp 1606120353
transform 1 0 18308 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_53_179
timestamp 1606120353
transform 1 0 17572 0 1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_52_183
timestamp 1606120353
transform 1 0 17940 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_52_177
timestamp 1606120353
transform 1 0 17388 0 -1 31008
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A
timestamp 1606120353
transform 1 0 17388 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1606120353
transform 1 0 17940 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0762_
timestamp 1606120353
transform 1 0 18032 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_53_198
timestamp 1606120353
transform 1 0 19320 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_53_191
timestamp 1606120353
transform 1 0 18676 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_52_196
timestamp 1606120353
transform 1 0 19136 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__A
timestamp 1606120353
transform 1 0 18860 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A
timestamp 1606120353
transform 1 0 18492 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk
timestamp 1606120353
transform 1 0 19044 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__a21o_4  _0770_
timestamp 1606120353
transform 1 0 18032 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_52_209
timestamp 1606120353
transform 1 0 20332 0 -1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_52_205
timestamp 1606120353
transform 1 0 19964 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_201
timestamp 1606120353
transform 1 0 19596 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__CLK
timestamp 1606120353
transform 1 0 20148 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__D
timestamp 1606120353
transform 1 0 19780 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0663__A
timestamp 1606120353
transform 1 0 19412 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_52_219
timestamp 1606120353
transform 1 0 21252 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_52_215
timestamp 1606120353
transform 1 0 20884 0 -1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_52_213
timestamp 1606120353
transform 1 0 20700 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1606120353
transform 1 0 20792 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_53_220
timestamp 1606120353
transform 1 0 21344 0 1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1190_
timestamp 1606120353
transform 1 0 21344 0 -1 31008
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1147_
timestamp 1606120353
transform 1 0 19596 0 1 31008
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A2
timestamp 1606120353
transform 1 0 23368 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A1
timestamp 1606120353
transform 1 0 23000 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_52_239
timestamp 1606120353
transform 1 0 23092 0 -1 31008
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILLER_53_232
timestamp 1606120353
transform 1 0 22448 0 1 31008
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_53_240
timestamp 1606120353
transform 1 0 23184 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_252
timestamp 1606120353
transform 1 0 24288 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_52_247
timestamp 1606120353
transform 1 0 23828 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__D
timestamp 1606120353
transform 1 0 24104 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__B1_N
timestamp 1606120353
transform 1 0 23644 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1606120353
transform 1 0 23552 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_53_262
timestamp 1606120353
transform 1 0 25208 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_258
timestamp 1606120353
transform 1 0 24840 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_256
timestamp 1606120353
transform 1 0 24656 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__B1_N
timestamp 1606120353
transform 1 0 24472 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__B
timestamp 1606120353
transform 1 0 25024 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__A
timestamp 1606120353
transform 1 0 25392 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0916_
timestamp 1606120353
transform 1 0 24840 0 -1 31008
box 0 -48 828 592
use sky130_fd_sc_hd__a21bo_4  _0911_
timestamp 1606120353
transform 1 0 23644 0 1 31008
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_52_271
timestamp 1606120353
transform 1 0 26036 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_267
timestamp 1606120353
transform 1 0 25668 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__D
timestamp 1606120353
transform 1 0 26220 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__C
timestamp 1606120353
transform 1 0 25852 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0908_
timestamp 1606120353
transform 1 0 25576 0 1 31008
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_53_279
timestamp 1606120353
transform 1 0 26772 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_275
timestamp 1606120353
transform 1 0 26404 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_280
timestamp 1606120353
transform 1 0 26864 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_276
timestamp 1606120353
transform 1 0 26496 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__B
timestamp 1606120353
transform 1 0 26680 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A
timestamp 1606120353
transform 1 0 26956 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A
timestamp 1606120353
transform 1 0 26588 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1606120353
transform 1 0 26404 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0887_
timestamp 1606120353
transform 1 0 27048 0 -1 31008
box 0 -48 828 592
use sky130_fd_sc_hd__and4_4  _0899_
timestamp 1606120353
transform 1 0 27140 0 1 31008
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_53_292
timestamp 1606120353
transform 1 0 27968 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_52_295
timestamp 1606120353
transform 1 0 28244 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_52_291
timestamp 1606120353
transform 1 0 27876 0 -1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__C
timestamp 1606120353
transform 1 0 28152 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_53_300
timestamp 1606120353
transform 1 0 28704 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_53_296
timestamp 1606120353
transform 1 0 28336 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_52_302
timestamp 1606120353
transform 1 0 28888 0 -1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_52_298
timestamp 1606120353
transform 1 0 28520 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A1
timestamp 1606120353
transform 1 0 28704 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__B1
timestamp 1606120353
transform 1 0 28336 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A2
timestamp 1606120353
transform 1 0 28520 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__A
timestamp 1606120353
transform 1 0 28980 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_308
timestamp 1606120353
transform 1 0 29440 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__B1_N
timestamp 1606120353
transform 1 0 29256 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1606120353
transform 1 0 29164 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__nor2_4  _0910_
timestamp 1606120353
transform 1 0 29256 0 1 31008
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILLER_53_319
timestamp 1606120353
transform 1 0 30452 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_53_315
timestamp 1606120353
transform 1 0 30084 0 1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_52_316
timestamp 1606120353
transform 1 0 30176 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_52_312
timestamp 1606120353
transform 1 0 29808 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A1
timestamp 1606120353
transform 1 0 29992 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__B
timestamp 1606120353
transform 1 0 29624 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0866_
timestamp 1606120353
transform 1 0 30452 0 -1 31008
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_53_322
timestamp 1606120353
transform 1 0 30728 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_328
timestamp 1606120353
transform 1 0 31280 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__B1
timestamp 1606120353
transform 1 0 31464 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A1
timestamp 1606120353
transform 1 0 30544 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A2
timestamp 1606120353
transform 1 0 30912 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0867_
timestamp 1606120353
transform 1 0 31096 0 1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1606120353
transform 1 0 32016 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_52_332
timestamp 1606120353
transform 1 0 31648 0 -1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_52_337
timestamp 1606120353
transform 1 0 32108 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_52_349
timestamp 1606120353
transform 1 0 33212 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_53_338
timestamp 1606120353
transform 1 0 32200 0 1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_53_350
timestamp 1606120353
transform 1 0 33304 0 1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1606120353
transform 1 0 34776 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_52_361
timestamp 1606120353
transform 1 0 34316 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_52_373
timestamp 1606120353
transform 1 0 35420 0 -1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_53_362
timestamp 1606120353
transform 1 0 34408 0 1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_53_367
timestamp 1606120353
transform 1 0 34868 0 1 31008
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1173_
timestamp 1606120353
transform 1 0 35788 0 1 31008
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__D
timestamp 1606120353
transform 1 0 35604 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__CLK
timestamp 1606120353
transform 1 0 35788 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_52_379
timestamp 1606120353
transform 1 0 35972 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_52_391
timestamp 1606120353
transform 1 0 37076 0 -1 31008
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_53_396
timestamp 1606120353
transform 1 0 37536 0 1 31008
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1606120353
transform -1 0 38548 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1606120353
transform -1 0 38548 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1606120353
transform 1 0 37628 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_52_398
timestamp 1606120353
transform 1 0 37720 0 -1 31008
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1606120353
transform 1 0 1104 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__B2
timestamp 1606120353
transform 1 0 3128 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1606120353
transform 1 0 1380 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_54_15
timestamp 1606120353
transform 1 0 2484 0 -1 32096
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_54_21
timestamp 1606120353
transform 1 0 3036 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1606120353
transform 1 0 3956 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_54_24
timestamp 1606120353
transform 1 0 3312 0 -1 32096
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_54_30
timestamp 1606120353
transform 1 0 3864 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_54_32
timestamp 1606120353
transform 1 0 4048 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_54_44
timestamp 1606120353
transform 1 0 5152 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_54_56
timestamp 1606120353
transform 1 0 6256 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_54_68
timestamp 1606120353
transform 1 0 7360 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_54_80
timestamp 1606120353
transform 1 0 8464 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1606120353
transform 1 0 9568 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_54_93
timestamp 1606120353
transform 1 0 9660 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_54_105
timestamp 1606120353
transform 1 0 10764 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__CLK
timestamp 1606120353
transform 1 0 12880 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_54_117
timestamp 1606120353
transform 1 0 11868 0 -1 32096
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_54_125
timestamp 1606120353
transform 1 0 12604 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_54_130
timestamp 1606120353
transform 1 0 13064 0 -1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _0733_
timestamp 1606120353
transform 1 0 13800 0 -1 32096
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1606120353
transform 1 0 15180 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__B1
timestamp 1606120353
transform 1 0 13524 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_54_134
timestamp 1606120353
transform 1 0 13432 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_54_137
timestamp 1606120353
transform 1 0 13708 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_54_145
timestamp 1606120353
transform 1 0 14444 0 -1 32096
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_54_154
timestamp 1606120353
transform 1 0 15272 0 -1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__a21o_4  _0764_
timestamp 1606120353
transform 1 0 16560 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__D
timestamp 1606120353
transform 1 0 15732 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A2
timestamp 1606120353
transform 1 0 16100 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_54_158
timestamp 1606120353
transform 1 0 15640 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_54_161
timestamp 1606120353
transform 1 0 15916 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_54_165
timestamp 1606120353
transform 1 0 16284 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0732_
timestamp 1606120353
transform 1 0 18400 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__D
timestamp 1606120353
transform 1 0 19044 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_54_180
timestamp 1606120353
transform 1 0 17664 0 -1 32096
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_54_191
timestamp 1606120353
transform 1 0 18676 0 -1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1606120353
transform 1 0 19228 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0663_
timestamp 1606120353
transform 1 0 19412 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1606120353
transform 1 0 20792 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_clk_A
timestamp 1606120353
transform 1 0 19872 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_202
timestamp 1606120353
transform 1 0 19688 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_54_206
timestamp 1606120353
transform 1 0 20056 0 -1 32096
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_54_215
timestamp 1606120353
transform 1 0 20884 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_54_227
timestamp 1606120353
transform 1 0 21988 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_54_239
timestamp 1606120353
transform 1 0 23092 0 -1 32096
box 0 -48 552 592
use sky130_fd_sc_hd__a21bo_4  _0936_
timestamp 1606120353
transform 1 0 24472 0 -1 32096
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A2
timestamp 1606120353
transform 1 0 24288 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A1
timestamp 1606120353
transform 1 0 23644 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_54_247
timestamp 1606120353
transform 1 0 23828 0 -1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1606120353
transform 1 0 24196 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0903_
timestamp 1606120353
transform 1 0 26496 0 -1 32096
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1606120353
transform 1 0 26404 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__D
timestamp 1606120353
transform 1 0 26220 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__D
timestamp 1606120353
transform 1 0 25852 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_267
timestamp 1606120353
transform 1 0 25668 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_271
timestamp 1606120353
transform 1 0 26036 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_285
timestamp 1606120353
transform 1 0 27324 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0909_
timestamp 1606120353
transform 1 0 28336 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_clk
timestamp 1606120353
transform 1 0 28060 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__B
timestamp 1606120353
transform 1 0 27508 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__C
timestamp 1606120353
transform 1 0 27876 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_289
timestamp 1606120353
transform 1 0 27692 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_54_308
timestamp 1606120353
transform 1 0 29440 0 -1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _0864_
timestamp 1606120353
transform 1 0 30452 0 -1 32096
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A1
timestamp 1606120353
transform 1 0 30176 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A
timestamp 1606120353
transform 1 0 29808 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_314
timestamp 1606120353
transform 1 0 29992 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_54_318
timestamp 1606120353
transform 1 0 30360 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_54_328
timestamp 1606120353
transform 1 0 31280 0 -1 32096
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1606120353
transform 1 0 32016 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_54_337
timestamp 1606120353
transform 1 0 32108 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_54_349
timestamp 1606120353
transform 1 0 33212 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_54_361
timestamp 1606120353
transform 1 0 34316 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_54_373
timestamp 1606120353
transform 1 0 35420 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_54_385
timestamp 1606120353
transform 1 0 36524 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1606120353
transform -1 0 38548 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1606120353
transform 1 0 37628 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_54_398
timestamp 1606120353
transform 1 0 37720 0 -1 32096
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1606120353
transform 1 0 1104 0 1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1606120353
transform 1 0 1380 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1606120353
transform 1 0 2484 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1606120353
transform 1 0 3588 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1606120353
transform 1 0 4692 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1606120353
transform 1 0 6716 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__D
timestamp 1606120353
transform 1 0 5980 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__CLK
timestamp 1606120353
transform 1 0 6348 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_51
timestamp 1606120353
transform 1 0 5796 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_55
timestamp 1606120353
transform 1 0 6164 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_59
timestamp 1606120353
transform 1 0 6532 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_55_62
timestamp 1606120353
transform 1 0 6808 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_55_74
timestamp 1606120353
transform 1 0 7912 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_55_86
timestamp 1606120353
transform 1 0 9016 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_clk_A
timestamp 1606120353
transform 1 0 10856 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_55_98
timestamp 1606120353
transform 1 0 10120 0 1 32096
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_55_108
timestamp 1606120353
transform 1 0 11040 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1606120353
transform 1 0 12328 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__D
timestamp 1606120353
transform 1 0 12604 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A2
timestamp 1606120353
transform 1 0 12972 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__CLK
timestamp 1606120353
transform 1 0 12144 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_123
timestamp 1606120353
transform 1 0 12420 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_127
timestamp 1606120353
transform 1 0 12788 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_131
timestamp 1606120353
transform 1 0 13156 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0734_
timestamp 1606120353
transform 1 0 13524 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A1
timestamp 1606120353
transform 1 0 15180 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A1
timestamp 1606120353
transform 1 0 13340 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__B1
timestamp 1606120353
transform 1 0 14812 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_147
timestamp 1606120353
transform 1 0 14628 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_151
timestamp 1606120353
transform 1 0 14996 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0749_
timestamp 1606120353
transform 1 0 15364 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__CLK
timestamp 1606120353
transform 1 0 16652 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_167
timestamp 1606120353
transform 1 0 16468 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_55_171
timestamp 1606120353
transform 1 0 16836 0 1 32096
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _0815_
timestamp 1606120353
transform 1 0 18032 0 1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1155_
timestamp 1606120353
transform 1 0 19044 0 1 32096
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1606120353
transform 1 0 17940 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__D
timestamp 1606120353
transform 1 0 18492 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A
timestamp 1606120353
transform 1 0 18860 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__CLK
timestamp 1606120353
transform 1 0 17756 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_179
timestamp 1606120353
transform 1 0 17572 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_187
timestamp 1606120353
transform 1 0 18308 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_191
timestamp 1606120353
transform 1 0 18676 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_55_214
timestamp 1606120353
transform 1 0 20792 0 1 32096
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__D
timestamp 1606120353
transform 1 0 21620 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A
timestamp 1606120353
transform 1 0 23368 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__CLK
timestamp 1606120353
transform 1 0 21988 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_55_222
timestamp 1606120353
transform 1 0 21528 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1606120353
transform 1 0 21804 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_55_229
timestamp 1606120353
transform 1 0 22172 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_55_241
timestamp 1606120353
transform 1 0 23276 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _0861_
timestamp 1606120353
transform 1 0 23736 0 1 32096
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1606120353
transform 1 0 23552 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__A
timestamp 1606120353
transform 1 0 24840 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__B
timestamp 1606120353
transform 1 0 25208 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_55_245
timestamp 1606120353
transform 1 0 23644 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_55_255
timestamp 1606120353
transform 1 0 24564 0 1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_55_260
timestamp 1606120353
transform 1 0 25024 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_55_264
timestamp 1606120353
transform 1 0 25392 0 1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__a21o_4  _0900_
timestamp 1606120353
transform 1 0 27324 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A2
timestamp 1606120353
transform 1 0 26496 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A2
timestamp 1606120353
transform 1 0 27140 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__B1
timestamp 1606120353
transform 1 0 26128 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A1
timestamp 1606120353
transform 1 0 25760 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_270
timestamp 1606120353
transform 1 0 25944 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_274
timestamp 1606120353
transform 1 0 26312 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_55_278
timestamp 1606120353
transform 1 0 26680 0 1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_55_282
timestamp 1606120353
transform 1 0 27048 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1606120353
transform 1 0 29164 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__A
timestamp 1606120353
transform 1 0 28612 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__B
timestamp 1606120353
transform 1 0 28980 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_297
timestamp 1606120353
transform 1 0 28428 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_301
timestamp 1606120353
transform 1 0 28796 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_55_306
timestamp 1606120353
transform 1 0 29256 0 1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _0854_
timestamp 1606120353
transform 1 0 30176 0 1 32096
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A2
timestamp 1606120353
transform 1 0 29992 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A
timestamp 1606120353
transform 1 0 29624 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__B1
timestamp 1606120353
transform 1 0 31188 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_312
timestamp 1606120353
transform 1 0 29808 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_325
timestamp 1606120353
transform 1 0 31004 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_329
timestamp 1606120353
transform 1 0 31372 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_clk_A
timestamp 1606120353
transform 1 0 31556 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_55_333
timestamp 1606120353
transform 1 0 31740 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_55_345
timestamp 1606120353
transform 1 0 32844 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1606120353
transform 1 0 34776 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_55_357
timestamp 1606120353
transform 1 0 33948 0 1 32096
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_55_365
timestamp 1606120353
transform 1 0 34684 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_55_367
timestamp 1606120353
transform 1 0 34868 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_55_379
timestamp 1606120353
transform 1 0 35972 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_55_391
timestamp 1606120353
transform 1 0 37076 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1606120353
transform -1 0 38548 0 1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_55_403
timestamp 1606120353
transform 1 0 38180 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1606120353
transform 1 0 1104 0 -1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1606120353
transform 1 0 1380 0 -1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1606120353
transform 1 0 2484 0 -1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1606120353
transform 1 0 3956 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_56_27
timestamp 1606120353
transform 1 0 3588 0 -1 33184
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_56_32
timestamp 1606120353
transform 1 0 4048 0 -1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_56_44
timestamp 1606120353
transform 1 0 5152 0 -1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1145_
timestamp 1606120353
transform 1 0 5980 0 -1 33184
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_1  FILLER_56_52
timestamp 1606120353
transform 1 0 5888 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_56_72
timestamp 1606120353
transform 1 0 7728 0 -1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_56_84
timestamp 1606120353
transform 1 0 8832 0 -1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1606120353
transform 1 0 9568 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_clk
timestamp 1606120353
transform 1 0 10856 0 -1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_56_93
timestamp 1606120353
transform 1 0 9660 0 -1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_56_105
timestamp 1606120353
transform 1 0 10764 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1606120353
transform 1 0 11132 0 -1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1085_
timestamp 1606120353
transform 1 0 12604 0 -1 33184
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_4  FILLER_56_121
timestamp 1606120353
transform 1 0 12236 0 -1 33184
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1606120353
transform 1 0 15180 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__A2
timestamp 1606120353
transform 1 0 14996 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_56_144
timestamp 1606120353
transform 1 0 14352 0 -1 33184
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_56_150
timestamp 1606120353
transform 1 0 14904 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_56_154
timestamp 1606120353
transform 1 0 15272 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1113_
timestamp 1606120353
transform 1 0 15732 0 -1 33184
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__B2
timestamp 1606120353
transform 1 0 15456 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_56_158
timestamp 1606120353
transform 1 0 15640 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1186_
timestamp 1606120353
transform 1 0 18308 0 -1 33184
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_8  FILLER_56_178
timestamp 1606120353
transform 1 0 17480 0 -1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_56_186
timestamp 1606120353
transform 1 0 18216 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1606120353
transform 1 0 20792 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A2
timestamp 1606120353
transform 1 0 20332 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_56_206
timestamp 1606120353
transform 1 0 20056 0 -1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_56_211
timestamp 1606120353
transform 1 0 20516 0 -1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_56_215
timestamp 1606120353
transform 1 0 20884 0 -1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1197_
timestamp 1606120353
transform 1 0 21620 0 -1 33184
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_12  FILLER_56_242
timestamp 1606120353
transform 1 0 23368 0 -1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__nor2_4  _0905_
timestamp 1606120353
transform 1 0 24840 0 -1 33184
box 0 -48 828 592
use sky130_fd_sc_hd__decap_4  FILLER_56_254
timestamp 1606120353
transform 1 0 24472 0 -1 33184
box 0 -48 368 592
use sky130_fd_sc_hd__a21o_4  _0904_
timestamp 1606120353
transform 1 0 26496 0 -1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1606120353
transform 1 0 26404 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_56_267
timestamp 1606120353
transform 1 0 25668 0 -1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__nor2_4  _0901_
timestamp 1606120353
transform 1 0 28336 0 -1 33184
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__B1
timestamp 1606120353
transform 1 0 29440 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__B1
timestamp 1606120353
transform 1 0 27784 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A1
timestamp 1606120353
transform 1 0 28152 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_288
timestamp 1606120353
transform 1 0 27600 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_292
timestamp 1606120353
transform 1 0 27968 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_56_305
timestamp 1606120353
transform 1 0 29164 0 -1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__o21a_4  _0855_
timestamp 1606120353
transform 1 0 30176 0 -1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_clk
timestamp 1606120353
transform 1 0 29900 0 -1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_56_310
timestamp 1606120353
transform 1 0 29624 0 -1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_56_328
timestamp 1606120353
transform 1 0 31280 0 -1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1606120353
transform 1 0 32016 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_56_337
timestamp 1606120353
transform 1 0 32108 0 -1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_56_349
timestamp 1606120353
transform 1 0 33212 0 -1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_56_361
timestamp 1606120353
transform 1 0 34316 0 -1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_56_373
timestamp 1606120353
transform 1 0 35420 0 -1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_56_385
timestamp 1606120353
transform 1 0 36524 0 -1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1606120353
transform -1 0 38548 0 -1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1606120353
transform 1 0 37628 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_56_398
timestamp 1606120353
transform 1 0 37720 0 -1 33184
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1606120353
transform 1 0 1104 0 1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1606120353
transform 1 0 1380 0 1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1606120353
transform 1 0 2484 0 1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1606120353
transform 1 0 3588 0 1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1606120353
transform 1 0 4692 0 1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1606120353
transform 1 0 6716 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_57_51
timestamp 1606120353
transform 1 0 5796 0 1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_57_59
timestamp 1606120353
transform 1 0 6532 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_57_62
timestamp 1606120353
transform 1 0 6808 0 1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_57_74
timestamp 1606120353
transform 1 0 7912 0 1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_57_86
timestamp 1606120353
transform 1 0 9016 0 1 33184
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__D
timestamp 1606120353
transform 1 0 9660 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__CLK
timestamp 1606120353
transform 1 0 10028 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_57_92
timestamp 1606120353
transform 1 0 9568 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_57_95
timestamp 1606120353
transform 1 0 9844 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_57_99
timestamp 1606120353
transform 1 0 10212 0 1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1606120353
transform 1 0 12328 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_57_111
timestamp 1606120353
transform 1 0 11316 0 1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_57_119
timestamp 1606120353
transform 1 0 12052 0 1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_57_123
timestamp 1606120353
transform 1 0 12420 0 1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__A1
timestamp 1606120353
transform 1 0 15088 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__B2
timestamp 1606120353
transform 1 0 14720 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__B1
timestamp 1606120353
transform 1 0 14352 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_57_135
timestamp 1606120353
transform 1 0 13524 0 1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_57_143
timestamp 1606120353
transform 1 0 14260 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_57_146
timestamp 1606120353
transform 1 0 14536 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_150
timestamp 1606120353
transform 1 0 14904 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_154
timestamp 1606120353
transform 1 0 15272 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _0820_
timestamp 1606120353
transform 1 0 15916 0 1 33184
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A1
timestamp 1606120353
transform 1 0 15456 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_57_158
timestamp 1606120353
transform 1 0 15640 0 1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_57_175
timestamp 1606120353
transform 1 0 17204 0 1 33184
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_57_184
timestamp 1606120353
transform 1 0 18032 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_57_182
timestamp 1606120353
transform 1 0 17848 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_57_179
timestamp 1606120353
transform 1 0 17572 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__D
timestamp 1606120353
transform 1 0 17664 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1606120353
transform 1 0 17940 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_57_188
timestamp 1606120353
transform 1 0 18400 0 1 33184
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__CLK
timestamp 1606120353
transform 1 0 18216 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_57_197
timestamp 1606120353
transform 1 0 19228 0 1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_57_194
timestamp 1606120353
transform 1 0 18952 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__CLK
timestamp 1606120353
transform 1 0 19044 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0927_
timestamp 1606120353
transform 1 0 20332 0 1 33184
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__B1_N
timestamp 1606120353
transform 1 0 20148 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_205
timestamp 1606120353
transform 1 0 19964 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A2
timestamp 1606120353
transform 1 0 21712 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A1
timestamp 1606120353
transform 1 0 22080 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__B1
timestamp 1606120353
transform 1 0 23368 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__B1
timestamp 1606120353
transform 1 0 22448 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 1606120353
transform 1 0 21528 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_226
timestamp 1606120353
transform 1 0 21896 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_230
timestamp 1606120353
transform 1 0 22264 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_57_234
timestamp 1606120353
transform 1 0 22632 0 1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_57_253
timestamp 1606120353
transform 1 0 24380 0 1 33184
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_57_249
timestamp 1606120353
transform 1 0 24012 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_245
timestamp 1606120353
transform 1 0 23644 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__A1
timestamp 1606120353
transform 1 0 24196 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__A2
timestamp 1606120353
transform 1 0 23828 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1606120353
transform 1 0 23552 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_57_259
timestamp 1606120353
transform 1 0 24932 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A1
timestamp 1606120353
transform 1 0 24748 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A2
timestamp 1606120353
transform 1 0 25116 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0906_
timestamp 1606120353
transform 1 0 25300 0 1 33184
box 0 -48 1196 592
use sky130_fd_sc_hd__a21bo_4  _0902_
timestamp 1606120353
transform 1 0 27232 0 1 33184
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A2
timestamp 1606120353
transform 1 0 27048 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__B1_N
timestamp 1606120353
transform 1 0 26680 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_276
timestamp 1606120353
transform 1 0 26496 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_280
timestamp 1606120353
transform 1 0 26864 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0851_
timestamp 1606120353
transform 1 0 29256 0 1 33184
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1606120353
transform 1 0 29164 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A1
timestamp 1606120353
transform 1 0 28980 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_clk_A
timestamp 1606120353
transform 1 0 28612 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_297
timestamp 1606120353
transform 1 0 28428 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_301
timestamp 1606120353
transform 1 0 28796 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A2
timestamp 1606120353
transform 1 0 30268 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_315
timestamp 1606120353
transform 1 0 30084 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_57_319
timestamp 1606120353
transform 1 0 30452 0 1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_57_331
timestamp 1606120353
transform 1 0 31556 0 1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_57_343
timestamp 1606120353
transform 1 0 32660 0 1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1606120353
transform 1 0 34776 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_57_355
timestamp 1606120353
transform 1 0 33764 0 1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_57_363
timestamp 1606120353
transform 1 0 34500 0 1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_57_367
timestamp 1606120353
transform 1 0 34868 0 1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_57_379
timestamp 1606120353
transform 1 0 35972 0 1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_57_391
timestamp 1606120353
transform 1 0 37076 0 1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1606120353
transform -1 0 38548 0 1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_57_403
timestamp 1606120353
transform 1 0 38180 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1606120353
transform 1 0 1104 0 -1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1606120353
transform 1 0 1380 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1606120353
transform 1 0 2484 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1606120353
transform 1 0 3956 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_58_27
timestamp 1606120353
transform 1 0 3588 0 -1 34272
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_58_32
timestamp 1606120353
transform 1 0 4048 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_58_44
timestamp 1606120353
transform 1 0 5152 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_58_56
timestamp 1606120353
transform 1 0 6256 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_58_68
timestamp 1606120353
transform 1 0 7360 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_58_80
timestamp 1606120353
transform 1 0 8464 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1150_
timestamp 1606120353
transform 1 0 9660 0 -1 34272
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1606120353
transform 1 0 9568 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_58_112
timestamp 1606120353
transform 1 0 11408 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_58_124
timestamp 1606120353
transform 1 0 12512 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1606120353
transform 1 0 15180 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A2
timestamp 1606120353
transform 1 0 14996 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_58_136
timestamp 1606120353
transform 1 0 13616 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_58_148
timestamp 1606120353
transform 1 0 14720 0 -1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_58_154
timestamp 1606120353
transform 1 0 15272 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _0821_
timestamp 1606120353
transform 1 0 15456 0 -1 34272
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__B1
timestamp 1606120353
transform 1 0 16928 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_170
timestamp 1606120353
transform 1 0 16744 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_58_174
timestamp 1606120353
transform 1 0 17112 0 -1 34272
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1117_
timestamp 1606120353
transform 1 0 17664 0 -1 34272
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1606120353
transform 1 0 20792 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A1
timestamp 1606120353
transform 1 0 20332 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__CLK
timestamp 1606120353
transform 1 0 19780 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_58_199
timestamp 1606120353
transform 1 0 19412 0 -1 34272
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_58_205
timestamp 1606120353
transform 1 0 19964 0 -1 34272
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_58_211
timestamp 1606120353
transform 1 0 20516 0 -1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_58_215
timestamp 1606120353
transform 1 0 20884 0 -1 34272
box 0 -48 552 592
use sky130_fd_sc_hd__o21ai_4  _0863_
timestamp 1606120353
transform 1 0 21528 0 -1 34272
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_1  FILLER_58_221
timestamp 1606120353
transform 1 0 21436 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_58_235
timestamp 1606120353
transform 1 0 22724 0 -1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__o21a_4  _0862_
timestamp 1606120353
transform 1 0 23460 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__B1_N
timestamp 1606120353
transform 1 0 25300 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_58_255
timestamp 1606120353
transform 1 0 24564 0 -1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1606120353
transform 1 0 26404 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_clk
timestamp 1606120353
transform 1 0 27232 0 -1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_58_265
timestamp 1606120353
transform 1 0 25484 0 -1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_58_273
timestamp 1606120353
transform 1 0 26220 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_58_276
timestamp 1606120353
transform 1 0 26496 0 -1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__o21ai_4  _0856_
timestamp 1606120353
transform 1 0 29440 0 -1 34272
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A1
timestamp 1606120353
transform 1 0 27692 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A
timestamp 1606120353
transform 1 0 29256 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_clk_A
timestamp 1606120353
transform 1 0 28060 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_287
timestamp 1606120353
transform 1 0 27508 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_291
timestamp 1606120353
transform 1 0 27876 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_58_295
timestamp 1606120353
transform 1 0 28244 0 -1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_58_303
timestamp 1606120353
transform 1 0 28980 0 -1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1606120353
transform 1 0 30636 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1606120353
transform 1 0 32016 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_58_333
timestamp 1606120353
transform 1 0 31740 0 -1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_58_337
timestamp 1606120353
transform 1 0 32108 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_58_349
timestamp 1606120353
transform 1 0 33212 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_58_361
timestamp 1606120353
transform 1 0 34316 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_58_373
timestamp 1606120353
transform 1 0 35420 0 -1 34272
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__CLK
timestamp 1606120353
transform 1 0 35788 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_58_379
timestamp 1606120353
transform 1 0 35972 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_58_391
timestamp 1606120353
transform 1 0 37076 0 -1 34272
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1606120353
transform -1 0 38548 0 -1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1606120353
transform 1 0 37628 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_58_398
timestamp 1606120353
transform 1 0 37720 0 -1 34272
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1606120353
transform 1 0 1104 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1606120353
transform 1 0 1104 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1606120353
transform 1 0 1380 0 1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1606120353
transform 1 0 2484 0 1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1606120353
transform 1 0 1380 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1606120353
transform 1 0 2484 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1606120353
transform 1 0 3956 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1606120353
transform 1 0 3588 0 1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1606120353
transform 1 0 4692 0 1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_60_27
timestamp 1606120353
transform 1 0 3588 0 -1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_60_32
timestamp 1606120353
transform 1 0 4048 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_60_44
timestamp 1606120353
transform 1 0 5152 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1158_
timestamp 1606120353
transform 1 0 6992 0 -1 35360
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1606120353
transform 1 0 6716 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__D
timestamp 1606120353
transform 1 0 6992 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_59_51
timestamp 1606120353
transform 1 0 5796 0 1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_59_59
timestamp 1606120353
transform 1 0 6532 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_62
timestamp 1606120353
transform 1 0 6808 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_66
timestamp 1606120353
transform 1 0 7176 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_60_56
timestamp 1606120353
transform 1 0 6256 0 -1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__CLK
timestamp 1606120353
transform 1 0 7360 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_59_70
timestamp 1606120353
transform 1 0 7544 0 1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_59_82
timestamp 1606120353
transform 1 0 8648 0 1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_60_83
timestamp 1606120353
transform 1 0 8740 0 -1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1606120353
transform 1 0 9568 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_59_94
timestamp 1606120353
transform 1 0 9752 0 1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_59_106
timestamp 1606120353
transform 1 0 10856 0 1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_60_91
timestamp 1606120353
transform 1 0 9476 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_60_93
timestamp 1606120353
transform 1 0 9660 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_60_105
timestamp 1606120353
transform 1 0 10764 0 -1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_60_113
timestamp 1606120353
transform 1 0 11500 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_59_121
timestamp 1606120353
transform 1 0 12236 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_59_117
timestamp 1606120353
transform 1 0 11868 0 1 34272
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_59_114
timestamp 1606120353
transform 1 0 11592 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_clk_A
timestamp 1606120353
transform 1 0 11684 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_clk
timestamp 1606120353
transform 1 0 11684 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_60_130
timestamp 1606120353
transform 1 0 13064 0 -1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1606120353
transform 1 0 12328 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_60_118
timestamp 1606120353
transform 1 0 11960 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_59_123
timestamp 1606120353
transform 1 0 12420 0 1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_60_143
timestamp 1606120353
transform 1 0 14260 0 -1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1606120353
transform 1 0 13800 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_59_142
timestamp 1606120353
transform 1 0 14168 0 1 34272
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_59_139
timestamp 1606120353
transform 1 0 13892 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_59_135
timestamp 1606120353
transform 1 0 13524 0 1 34272
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_clk_A
timestamp 1606120353
transform 1 0 13984 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_clk
timestamp 1606120353
transform 1 0 13984 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_60_150
timestamp 1606120353
transform 1 0 14904 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_60_147
timestamp 1606120353
transform 1 0 14628 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__CLK
timestamp 1606120353
transform 1 0 14720 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__D
timestamp 1606120353
transform 1 0 14536 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1606120353
transform 1 0 15180 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_60_154
timestamp 1606120353
transform 1 0 15272 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1114_
timestamp 1606120353
transform 1 0 14720 0 1 34272
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_12  FILLER_59_167
timestamp 1606120353
transform 1 0 16468 0 1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_60_166
timestamp 1606120353
transform 1 0 16376 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1606120353
transform 1 0 17940 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__CLK
timestamp 1606120353
transform 1 0 18032 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_59_179
timestamp 1606120353
transform 1 0 17572 0 1 34272
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_59_184
timestamp 1606120353
transform 1 0 18032 0 1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_59_196
timestamp 1606120353
transform 1 0 19136 0 1 34272
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_60_178
timestamp 1606120353
transform 1 0 17480 0 -1 35360
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_60_186
timestamp 1606120353
transform 1 0 18216 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_60_198
timestamp 1606120353
transform 1 0 19320 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1151_
timestamp 1606120353
transform 1 0 19780 0 1 34272
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1606120353
transform 1 0 20792 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__D
timestamp 1606120353
transform 1 0 19596 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_59_200
timestamp 1606120353
transform 1 0 19504 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_60_210
timestamp 1606120353
transform 1 0 20424 0 -1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_60_215
timestamp 1606120353
transform 1 0 20884 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_59_222
timestamp 1606120353
transform 1 0 21528 0 1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_59_234
timestamp 1606120353
transform 1 0 22632 0 1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_59_242
timestamp 1606120353
transform 1 0 23368 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_60_227
timestamp 1606120353
transform 1 0 21988 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_60_239
timestamp 1606120353
transform 1 0 23092 0 -1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_60_250
timestamp 1606120353
transform 1 0 24104 0 -1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_60_247
timestamp 1606120353
transform 1 0 23828 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_59_245
timestamp 1606120353
transform 1 0 23644 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__A
timestamp 1606120353
transform 1 0 23920 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1606120353
transform 1 0 23552 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _0857_
timestamp 1606120353
transform 1 0 23920 0 1 34272
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILLER_60_258
timestamp 1606120353
transform 1 0 24840 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__CLK
timestamp 1606120353
transform 1 0 25116 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_60_263
timestamp 1606120353
transform 1 0 25300 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_59_257
timestamp 1606120353
transform 1 0 24748 0 1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1178_
timestamp 1606120353
transform 1 0 26404 0 1 34272
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1606120353
transform 1 0 26404 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__D
timestamp 1606120353
transform 1 0 26220 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__CLK
timestamp 1606120353
transform 1 0 25852 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_271
timestamp 1606120353
transform 1 0 26036 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_60_276
timestamp 1606120353
transform 1 0 26496 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1170_
timestamp 1606120353
transform 1 0 29256 0 1 34272
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1606120353
transform 1 0 29164 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__D
timestamp 1606120353
transform 1 0 28980 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__CLK
timestamp 1606120353
transform 1 0 29256 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_59_294
timestamp 1606120353
transform 1 0 28152 0 1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_59_302
timestamp 1606120353
transform 1 0 28888 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_60_288
timestamp 1606120353
transform 1 0 27600 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_60_300
timestamp 1606120353
transform 1 0 28704 0 -1 35360
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_60_308
timestamp 1606120353
transform 1 0 29440 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_59_325
timestamp 1606120353
transform 1 0 31004 0 1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_60_320
timestamp 1606120353
transform 1 0 30544 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1606120353
transform 1 0 32016 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1606120353
transform 1 0 32108 0 1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1606120353
transform 1 0 33212 0 1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_60_332
timestamp 1606120353
transform 1 0 31648 0 -1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_60_337
timestamp 1606120353
transform 1 0 32108 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_60_349
timestamp 1606120353
transform 1 0 33212 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1606120353
transform 1 0 34776 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_59_361
timestamp 1606120353
transform 1 0 34316 0 1 34272
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_59_365
timestamp 1606120353
transform 1 0 34684 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_59_367
timestamp 1606120353
transform 1 0 34868 0 1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_60_361
timestamp 1606120353
transform 1 0 34316 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_60_373
timestamp 1606120353
transform 1 0 35420 0 -1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1159_
timestamp 1606120353
transform 1 0 35788 0 1 34272
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__D
timestamp 1606120353
transform 1 0 35604 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__CLK
timestamp 1606120353
transform 1 0 35788 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_59_396
timestamp 1606120353
transform 1 0 37536 0 1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_60_379
timestamp 1606120353
transform 1 0 35972 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_60_391
timestamp 1606120353
transform 1 0 37076 0 -1 35360
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1606120353
transform -1 0 38548 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1606120353
transform -1 0 38548 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1606120353
transform 1 0 37628 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_60_398
timestamp 1606120353
transform 1 0 37720 0 -1 35360
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1606120353
transform 1 0 1104 0 1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1606120353
transform 1 0 1380 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1606120353
transform 1 0 2484 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__D
timestamp 1606120353
transform 1 0 4876 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1606120353
transform 1 0 3588 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_61_39
timestamp 1606120353
transform 1 0 4692 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_43
timestamp 1606120353
transform 1 0 5060 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1606120353
transform 1 0 6716 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__CLK
timestamp 1606120353
transform 1 0 5244 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_61_47
timestamp 1606120353
transform 1 0 5428 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_61_59
timestamp 1606120353
transform 1 0 6532 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_61_62
timestamp 1606120353
transform 1 0 6808 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_61_74
timestamp 1606120353
transform 1 0 7912 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_61_86
timestamp 1606120353
transform 1 0 9016 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_clk_A
timestamp 1606120353
transform 1 0 10396 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_61_98
timestamp 1606120353
transform 1 0 10120 0 1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_61_103
timestamp 1606120353
transform 1 0 10580 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1606120353
transform 1 0 12328 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_61_115
timestamp 1606120353
transform 1 0 11684 0 1 35360
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_61_121
timestamp 1606120353
transform 1 0 12236 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_61_123
timestamp 1606120353
transform 1 0 12420 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_61_135
timestamp 1606120353
transform 1 0 13524 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_61_147
timestamp 1606120353
transform 1 0 14628 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__D
timestamp 1606120353
transform 1 0 16376 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__CLK
timestamp 1606120353
transform 1 0 16744 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_61_159
timestamp 1606120353
transform 1 0 15732 0 1 35360
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_61_165
timestamp 1606120353
transform 1 0 16284 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_61_168
timestamp 1606120353
transform 1 0 16560 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_61_172
timestamp 1606120353
transform 1 0 16928 0 1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1172_
timestamp 1606120353
transform 1 0 18032 0 1 35360
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1606120353
transform 1 0 17940 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__D
timestamp 1606120353
transform 1 0 17756 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_61_180
timestamp 1606120353
transform 1 0 17664 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_61_203
timestamp 1606120353
transform 1 0 19780 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_61_215
timestamp 1606120353
transform 1 0 20884 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_61_227
timestamp 1606120353
transform 1 0 21988 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_61_239
timestamp 1606120353
transform 1 0 23092 0 1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1174_
timestamp 1606120353
transform 1 0 25116 0 1 35360
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1606120353
transform 1 0 23552 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__D
timestamp 1606120353
transform 1 0 24932 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_61_243
timestamp 1606120353
transform 1 0 23460 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_61_245
timestamp 1606120353
transform 1 0 23644 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_61_257
timestamp 1606120353
transform 1 0 24748 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_61_280
timestamp 1606120353
transform 1 0 26864 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1606120353
transform 1 0 29164 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_61_292
timestamp 1606120353
transform 1 0 27968 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_61_304
timestamp 1606120353
transform 1 0 29072 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_61_306
timestamp 1606120353
transform 1 0 29256 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_61_318
timestamp 1606120353
transform 1 0 30360 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_61_330
timestamp 1606120353
transform 1 0 31464 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_61_342
timestamp 1606120353
transform 1 0 32568 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1606120353
transform 1 0 34776 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_61_354
timestamp 1606120353
transform 1 0 33672 0 1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_61_367
timestamp 1606120353
transform 1 0 34868 0 1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1222_
timestamp 1606120353
transform 1 0 35788 0 1 35360
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__D
timestamp 1606120353
transform 1 0 35604 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_61_396
timestamp 1606120353
transform 1 0 37536 0 1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1606120353
transform -1 0 38548 0 1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1606120353
transform 1 0 1104 0 -1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0486__A
timestamp 1606120353
transform 1 0 1564 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1606120353
transform 1 0 1380 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_62_7
timestamp 1606120353
transform 1 0 1748 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_62_19
timestamp 1606120353
transform 1 0 2852 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1221_
timestamp 1606120353
transform 1 0 4876 0 -1 36448
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1606120353
transform 1 0 3956 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_62_32
timestamp 1606120353
transform 1 0 4048 0 -1 36448
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_62_40
timestamp 1606120353
transform 1 0 4784 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_62_60
timestamp 1606120353
transform 1 0 6624 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_62_72
timestamp 1606120353
transform 1 0 7728 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_62_84
timestamp 1606120353
transform 1 0 8832 0 -1 36448
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1606120353
transform 1 0 9568 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_clk
timestamp 1606120353
transform 1 0 10396 0 -1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_62_93
timestamp 1606120353
transform 1 0 9660 0 -1 36448
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_62_104
timestamp 1606120353
transform 1 0 10672 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_62_116
timestamp 1606120353
transform 1 0 11776 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_62_128
timestamp 1606120353
transform 1 0 12880 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1606120353
transform 1 0 15180 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_62_140
timestamp 1606120353
transform 1 0 13984 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_62_152
timestamp 1606120353
transform 1 0 15088 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_62_154
timestamp 1606120353
transform 1 0 15272 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1199_
timestamp 1606120353
transform 1 0 16376 0 -1 36448
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__CLK
timestamp 1606120353
transform 1 0 19136 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__CLK
timestamp 1606120353
transform 1 0 18308 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_185
timestamp 1606120353
transform 1 0 18124 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1606120353
transform 1 0 18492 0 -1 36448
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1606120353
transform 1 0 19044 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_62_198
timestamp 1606120353
transform 1 0 19320 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1606120353
transform 1 0 20792 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_62_210
timestamp 1606120353
transform 1 0 20424 0 -1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_62_215
timestamp 1606120353
transform 1 0 20884 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_62_227
timestamp 1606120353
transform 1 0 21988 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_62_239
timestamp 1606120353
transform 1 0 23092 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__CLK
timestamp 1606120353
transform 1 0 25300 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_62_251
timestamp 1606120353
transform 1 0 24196 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1606120353
transform 1 0 26404 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_62_265
timestamp 1606120353
transform 1 0 25484 0 -1 36448
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_62_273
timestamp 1606120353
transform 1 0 26220 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_62_276
timestamp 1606120353
transform 1 0 26496 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_62_288
timestamp 1606120353
transform 1 0 27600 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_62_300
timestamp 1606120353
transform 1 0 28704 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_62_312
timestamp 1606120353
transform 1 0 29808 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_62_324
timestamp 1606120353
transform 1 0 30912 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1606120353
transform 1 0 32016 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_62_337
timestamp 1606120353
transform 1 0 32108 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_62_349
timestamp 1606120353
transform 1 0 33212 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_62_361
timestamp 1606120353
transform 1 0 34316 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_62_373
timestamp 1606120353
transform 1 0 35420 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A2
timestamp 1606120353
transform 1 0 35604 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1606120353
transform 1 0 35788 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_62_389
timestamp 1606120353
transform 1 0 36892 0 -1 36448
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1606120353
transform -1 0 38548 0 -1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1606120353
transform 1 0 37628 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_62_398
timestamp 1606120353
transform 1 0 37720 0 -1 36448
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _0486_
timestamp 1606120353
transform 1 0 1380 0 1 36448
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1606120353
transform 1 0 1104 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0486__B
timestamp 1606120353
transform 1 0 2208 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_10
timestamp 1606120353
transform 1 0 2024 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_63_14
timestamp 1606120353
transform 1 0 2392 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_63_26
timestamp 1606120353
transform 1 0 3496 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_63_38
timestamp 1606120353
transform 1 0 4600 0 1 36448
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1606120353
transform 1 0 6716 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__D
timestamp 1606120353
transform 1 0 5612 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__CLK
timestamp 1606120353
transform 1 0 5980 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_63_46
timestamp 1606120353
transform 1 0 5336 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_63_51
timestamp 1606120353
transform 1 0 5796 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_63_55
timestamp 1606120353
transform 1 0 6164 0 1 36448
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_63_62
timestamp 1606120353
transform 1 0 6808 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_63_74
timestamp 1606120353
transform 1 0 7912 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_63_86
timestamp 1606120353
transform 1 0 9016 0 1 36448
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__D
timestamp 1606120353
transform 1 0 9660 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__CLK
timestamp 1606120353
transform 1 0 10028 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_63_92
timestamp 1606120353
transform 1 0 9568 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_63_95
timestamp 1606120353
transform 1 0 9844 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_63_99
timestamp 1606120353
transform 1 0 10212 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1606120353
transform 1 0 12328 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__D
timestamp 1606120353
transform 1 0 12144 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__CLK
timestamp 1606120353
transform 1 0 12604 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_63_111
timestamp 1606120353
transform 1 0 11316 0 1 36448
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_63_119
timestamp 1606120353
transform 1 0 12052 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_63_123
timestamp 1606120353
transform 1 0 12420 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_63_127
timestamp 1606120353
transform 1 0 12788 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__D
timestamp 1606120353
transform 1 0 15272 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_63_139
timestamp 1606120353
transform 1 0 13892 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_63_151
timestamp 1606120353
transform 1 0 14996 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__CLK
timestamp 1606120353
transform 1 0 15640 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_156
timestamp 1606120353
transform 1 0 15456 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_63_160
timestamp 1606120353
transform 1 0 15824 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_63_172
timestamp 1606120353
transform 1 0 16928 0 1 36448
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1153_
timestamp 1606120353
transform 1 0 19136 0 1 36448
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1606120353
transform 1 0 17940 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__D
timestamp 1606120353
transform 1 0 18308 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__D
timestamp 1606120353
transform 1 0 18952 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_63_180
timestamp 1606120353
transform 1 0 17664 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_63_184
timestamp 1606120353
transform 1 0 18032 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_63_189
timestamp 1606120353
transform 1 0 18492 0 1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_63_193
timestamp 1606120353
transform 1 0 18860 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_63_215
timestamp 1606120353
transform 1 0 20884 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_63_227
timestamp 1606120353
transform 1 0 21988 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_63_239
timestamp 1606120353
transform 1 0 23092 0 1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1213_
timestamp 1606120353
transform 1 0 25300 0 1 36448
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1606120353
transform 1 0 23552 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__D
timestamp 1606120353
transform 1 0 25116 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_63_243
timestamp 1606120353
transform 1 0 23460 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_63_245
timestamp 1606120353
transform 1 0 23644 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_63_257
timestamp 1606120353
transform 1 0 24748 0 1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_63_282
timestamp 1606120353
transform 1 0 27048 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1606120353
transform 1 0 29164 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_63_294
timestamp 1606120353
transform 1 0 28152 0 1 36448
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_63_302
timestamp 1606120353
transform 1 0 28888 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_63_306
timestamp 1606120353
transform 1 0 29256 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_63_318
timestamp 1606120353
transform 1 0 30360 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_63_330
timestamp 1606120353
transform 1 0 31464 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_63_342
timestamp 1606120353
transform 1 0 32568 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_63_354
timestamp 1606120353
transform 1 0 33672 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__D
timestamp 1606120353
transform 1 0 33764 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_357
timestamp 1606120353
transform 1 0 33948 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__CLK
timestamp 1606120353
transform 1 0 34132 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_63_361
timestamp 1606120353
transform 1 0 34316 0 1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_63_367
timestamp 1606120353
transform 1 0 34868 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_63_365
timestamp 1606120353
transform 1 0 34684 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1606120353
transform 1 0 34776 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_63_371
timestamp 1606120353
transform 1 0 35236 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A1
timestamp 1606120353
transform 1 0 35052 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__B1_N
timestamp 1606120353
transform 1 0 35420 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0925_
timestamp 1606120353
transform 1 0 35604 0 1 36448
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILLER_63_388
timestamp 1606120353
transform 1 0 36800 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1606120353
transform -1 0 38548 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_63_400
timestamp 1606120353
transform 1 0 37904 0 1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1606120353
transform 1 0 1104 0 -1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1606120353
transform 1 0 1380 0 -1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1606120353
transform 1 0 2484 0 -1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1606120353
transform 1 0 3956 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1606120353
transform 1 0 3588 0 -1 37536
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_64_32
timestamp 1606120353
transform 1 0 4048 0 -1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_64_44
timestamp 1606120353
transform 1 0 5152 0 -1 37536
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1127_
timestamp 1606120353
transform 1 0 5612 0 -1 37536
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_1  FILLER_64_48
timestamp 1606120353
transform 1 0 5520 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_64_68
timestamp 1606120353
transform 1 0 7360 0 -1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_64_80
timestamp 1606120353
transform 1 0 8464 0 -1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1141_
timestamp 1606120353
transform 1 0 9660 0 -1 37536
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1606120353
transform 1 0 9568 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1192_
timestamp 1606120353
transform 1 0 12144 0 -1 37536
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_8  FILLER_64_112
timestamp 1606120353
transform 1 0 11408 0 -1 37536
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1128_
timestamp 1606120353
transform 1 0 15272 0 -1 37536
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1606120353
transform 1 0 15180 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_64_139
timestamp 1606120353
transform 1 0 13892 0 -1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_64_151
timestamp 1606120353
transform 1 0 14996 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_64_173
timestamp 1606120353
transform 1 0 17020 0 -1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1161_
timestamp 1606120353
transform 1 0 18308 0 -1 37536
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_2  FILLER_64_185
timestamp 1606120353
transform 1 0 18124 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1606120353
transform 1 0 20792 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_64_206
timestamp 1606120353
transform 1 0 20056 0 -1 37536
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_64_215
timestamp 1606120353
transform 1 0 20884 0 -1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_64_227
timestamp 1606120353
transform 1 0 21988 0 -1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_64_239
timestamp 1606120353
transform 1 0 23092 0 -1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_64_251
timestamp 1606120353
transform 1 0 24196 0 -1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_64_263
timestamp 1606120353
transform 1 0 25300 0 -1 37536
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1606120353
transform 1 0 26404 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__D
timestamp 1606120353
transform 1 0 26680 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__CLK
timestamp 1606120353
transform 1 0 26220 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_271
timestamp 1606120353
transform 1 0 26036 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_276
timestamp 1606120353
transform 1 0 26496 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_64_280
timestamp 1606120353
transform 1 0 26864 0 -1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_64_292
timestamp 1606120353
transform 1 0 27968 0 -1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_64_304
timestamp 1606120353
transform 1 0 29072 0 -1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_64_316
timestamp 1606120353
transform 1 0 30176 0 -1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_64_328
timestamp 1606120353
transform 1 0 31280 0 -1 37536
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1606120353
transform 1 0 32016 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A2
timestamp 1606120353
transform 1 0 32292 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__CLK
timestamp 1606120353
transform 1 0 32660 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1606120353
transform 1 0 32108 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_341
timestamp 1606120353
transform 1 0 32476 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_64_345
timestamp 1606120353
transform 1 0 32844 0 -1 37536
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1183_
timestamp 1606120353
transform 1 0 33764 0 -1 37536
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_2  FILLER_64_353
timestamp 1606120353
transform 1 0 33580 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_64_374
timestamp 1606120353
transform 1 0 35512 0 -1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__CLK
timestamp 1606120353
transform 1 0 35788 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_64_379
timestamp 1606120353
transform 1 0 35972 0 -1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_64_391
timestamp 1606120353
transform 1 0 37076 0 -1 37536
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1606120353
transform -1 0 38548 0 -1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1606120353
transform 1 0 37628 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_64_398
timestamp 1606120353
transform 1 0 37720 0 -1 37536
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1606120353
transform 1 0 1104 0 1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__D
timestamp 1606120353
transform 1 0 1564 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__CLK
timestamp 1606120353
transform 1 0 1932 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_3
timestamp 1606120353
transform 1 0 1380 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_7
timestamp 1606120353
transform 1 0 1748 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_65_11
timestamp 1606120353
transform 1 0 2116 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_65_23
timestamp 1606120353
transform 1 0 3220 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_65_35
timestamp 1606120353
transform 1 0 4324 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1606120353
transform 1 0 6716 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__D
timestamp 1606120353
transform 1 0 7176 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__D
timestamp 1606120353
transform 1 0 5428 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__CLK
timestamp 1606120353
transform 1 0 5796 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_49
timestamp 1606120353
transform 1 0 5612 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_65_53
timestamp 1606120353
transform 1 0 5980 0 1 37536
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_65_62
timestamp 1606120353
transform 1 0 6808 0 1 37536
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1146_
timestamp 1606120353
transform 1 0 7360 0 1 37536
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_12  FILLER_65_87
timestamp 1606120353
transform 1 0 9108 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__or2_4  _1082_
timestamp 1606120353
transform 1 0 10580 0 1 37536
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__B
timestamp 1606120353
transform 1 0 10396 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_99
timestamp 1606120353
transform 1 0 10212 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_110
timestamp 1606120353
transform 1 0 11224 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1606120353
transform 1 0 12328 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A
timestamp 1606120353
transform 1 0 11408 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__D
timestamp 1606120353
transform 1 0 11776 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__CLK
timestamp 1606120353
transform 1 0 12144 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_114
timestamp 1606120353
transform 1 0 11592 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_118
timestamp 1606120353
transform 1 0 11960 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_65_123
timestamp 1606120353
transform 1 0 12420 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_65_135
timestamp 1606120353
transform 1 0 13524 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_65_147
timestamp 1606120353
transform 1 0 14628 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__D
timestamp 1606120353
transform 1 0 17204 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_65_159
timestamp 1606120353
transform 1 0 15732 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_65_171
timestamp 1606120353
transform 1 0 16836 0 1 37536
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1132_
timestamp 1606120353
transform 1 0 19320 0 1 37536
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1606120353
transform 1 0 17940 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__D
timestamp 1606120353
transform 1 0 19136 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__CLK
timestamp 1606120353
transform 1 0 17572 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_177
timestamp 1606120353
transform 1 0 17388 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_181
timestamp 1606120353
transform 1 0 17756 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_65_184
timestamp 1606120353
transform 1 0 18032 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_65_217
timestamp 1606120353
transform 1 0 21068 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__D
timestamp 1606120353
transform 1 0 22908 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__CLK
timestamp 1606120353
transform 1 0 23276 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_65_229
timestamp 1606120353
transform 1 0 22172 0 1 37536
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_65_239
timestamp 1606120353
transform 1 0 23092 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1606120353
transform 1 0 23552 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_65_243
timestamp 1606120353
transform 1 0 23460 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_65_245
timestamp 1606120353
transform 1 0 23644 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_65_257
timestamp 1606120353
transform 1 0 24748 0 1 37536
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1226_
timestamp 1606120353
transform 1 0 26220 0 1 37536
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__D
timestamp 1606120353
transform 1 0 26036 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__CLK
timestamp 1606120353
transform 1 0 25668 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_265
timestamp 1606120353
transform 1 0 25484 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_269
timestamp 1606120353
transform 1 0 25852 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1606120353
transform 1 0 29164 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_65_292
timestamp 1606120353
transform 1 0 27968 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_65_304
timestamp 1606120353
transform 1 0 29072 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_65_306
timestamp 1606120353
transform 1 0 29256 0 1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__D
timestamp 1606120353
transform 1 0 29532 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A1
timestamp 1606120353
transform 1 0 31280 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__CLK
timestamp 1606120353
transform 1 0 29900 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_311
timestamp 1606120353
transform 1 0 29716 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_65_315
timestamp 1606120353
transform 1 0 30084 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_65_327
timestamp 1606120353
transform 1 0 31188 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_65_330
timestamp 1606120353
transform 1 0 31464 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0933_
timestamp 1606120353
transform 1 0 32200 0 1 37536
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__D
timestamp 1606120353
transform 1 0 32016 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__B1_N
timestamp 1606120353
transform 1 0 31648 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_334
timestamp 1606120353
transform 1 0 31832 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_65_351
timestamp 1606120353
transform 1 0 33396 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1606120353
transform 1 0 34776 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_65_363
timestamp 1606120353
transform 1 0 34500 0 1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_65_367
timestamp 1606120353
transform 1 0 34868 0 1 37536
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1185_
timestamp 1606120353
transform 1 0 35788 0 1 37536
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__D
timestamp 1606120353
transform 1 0 35604 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_65_396
timestamp 1606120353
transform 1 0 37536 0 1 37536
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1606120353
transform -1 0 38548 0 1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1165_
timestamp 1606120353
transform 1 0 1472 0 -1 38624
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1606120353
transform 1 0 1104 0 -1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1606120353
transform 1 0 1104 0 1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_66_3
timestamp 1606120353
transform 1 0 1380 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1606120353
transform 1 0 1380 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_67_15
timestamp 1606120353
transform 1 0 2484 0 1 38624
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_67_27
timestamp 1606120353
transform 1 0 3588 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_23
timestamp 1606120353
transform 1 0 3220 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_66_23
timestamp 1606120353
transform 1 0 3220 0 -1 38624
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__CLK
timestamp 1606120353
transform 1 0 3404 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__D
timestamp 1606120353
transform 1 0 3772 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1606120353
transform 1 0 3956 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1606120353
transform 1 0 3956 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_66_44
timestamp 1606120353
transform 1 0 5152 0 -1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_66_32
timestamp 1606120353
transform 1 0 4048 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1193_
timestamp 1606120353
transform 1 0 4048 0 1 38624
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1606120353
transform 1 0 6164 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1606120353
transform 1 0 5796 0 1 38624
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_67_63
timestamp 1606120353
transform 1 0 6900 0 1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_67_58
timestamp 1606120353
transform 1 0 6440 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_66
timestamp 1606120353
transform 1 0 7176 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__CLK
timestamp 1606120353
transform 1 0 6256 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__D
timestamp 1606120353
transform 1 0 6624 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1606120353
transform 1 0 6808 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1181_
timestamp 1606120353
transform 1 0 7176 0 1 38624
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1122_
timestamp 1606120353
transform 1 0 5428 0 -1 38624
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__CLK
timestamp 1606120353
transform 1 0 7360 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_66_70
timestamp 1606120353
transform 1 0 7544 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_66_82
timestamp 1606120353
transform 1 0 8648 0 -1 38624
box 0 -48 736 592
use sky130_fd_sc_hd__decap_6  FILLER_67_85
timestamp 1606120353
transform 1 0 8924 0 1 38624
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_67_94
timestamp 1606120353
transform 1 0 9752 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_66_93
timestamp 1606120353
transform 1 0 9660 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_90
timestamp 1606120353
transform 1 0 9384 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__CLK
timestamp 1606120353
transform 1 0 9844 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__D
timestamp 1606120353
transform 1 0 9476 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1606120353
transform 1 0 9660 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1606120353
transform 1 0 9568 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_66_109
timestamp 1606120353
transform 1 0 11132 0 -1 38624
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1606120353
transform 1 0 10028 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1203_
timestamp 1606120353
transform 1 0 9844 0 1 38624
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1163_
timestamp 1606120353
transform 1 0 11684 0 -1 38624
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1606120353
transform 1 0 12512 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__B1_N
timestamp 1606120353
transform 1 0 13156 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__A2
timestamp 1606120353
transform 1 0 12788 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_67_114
timestamp 1606120353
transform 1 0 11592 0 1 38624
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_67_122
timestamp 1606120353
transform 1 0 12328 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_125
timestamp 1606120353
transform 1 0 12604 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_129
timestamp 1606120353
transform 1 0 12972 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_134
timestamp 1606120353
transform 1 0 13432 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__A1
timestamp 1606120353
transform 1 0 13616 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_67_152
timestamp 1606120353
transform 1 0 15088 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_67_146
timestamp 1606120353
transform 1 0 14536 0 1 38624
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_66_154
timestamp 1606120353
transform 1 0 15272 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_66_150
timestamp 1606120353
transform 1 0 14904 0 -1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__D
timestamp 1606120353
transform 1 0 15180 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1606120353
transform 1 0 15180 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_66_138
timestamp 1606120353
transform 1 0 13800 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__a21bo_4  _0935_
timestamp 1606120353
transform 1 0 13340 0 1 38624
box 0 -48 1196 592
use sky130_fd_sc_hd__dfxtp_4  _1130_
timestamp 1606120353
transform 1 0 17204 0 -1 38624
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1138_
timestamp 1606120353
transform 1 0 15456 0 1 38624
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1606120353
transform 1 0 15364 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__CLK
timestamp 1606120353
transform 1 0 15456 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_66_158
timestamp 1606120353
transform 1 0 15640 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_66_170
timestamp 1606120353
transform 1 0 16744 0 -1 38624
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_66_174
timestamp 1606120353
transform 1 0 17112 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_67_175
timestamp 1606120353
transform 1 0 17204 0 1 38624
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1606120353
transform 1 0 18216 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__CLK
timestamp 1606120353
transform 1 0 19320 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_66_194
timestamp 1606120353
transform 1 0 18952 0 -1 38624
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_67_183
timestamp 1606120353
transform 1 0 17940 0 1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_67_187
timestamp 1606120353
transform 1 0 18308 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1606120353
transform 1 0 20792 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1606120353
transform 1 0 21068 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_66_200
timestamp 1606120353
transform 1 0 19504 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_66_212
timestamp 1606120353
transform 1 0 20608 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_66_215
timestamp 1606120353
transform 1 0 20884 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_67_199
timestamp 1606120353
transform 1 0 19412 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_67_211
timestamp 1606120353
transform 1 0 20516 0 1 38624
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_67_218
timestamp 1606120353
transform 1 0 21160 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1224_
timestamp 1606120353
transform 1 0 22908 0 -1 38624
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_8  FILLER_66_227
timestamp 1606120353
transform 1 0 21988 0 -1 38624
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_66_235
timestamp 1606120353
transform 1 0 22724 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_67_230
timestamp 1606120353
transform 1 0 22264 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_67_242
timestamp 1606120353
transform 1 0 23368 0 1 38624
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1606120353
transform 1 0 23920 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_66_256
timestamp 1606120353
transform 1 0 24656 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_67_249
timestamp 1606120353
transform 1 0 24012 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_67_261
timestamp 1606120353
transform 1 0 25116 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_67_275
timestamp 1606120353
transform 1 0 26404 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_66_274
timestamp 1606120353
transform 1 0 26312 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_66_268
timestamp 1606120353
transform 1 0 25760 0 -1 38624
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__CLK
timestamp 1606120353
transform 1 0 26220 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1606120353
transform 1 0 26404 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_67_280
timestamp 1606120353
transform 1 0 26864 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__D
timestamp 1606120353
transform 1 0 26588 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1606120353
transform 1 0 26772 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1177_
timestamp 1606120353
transform 1 0 26496 0 -1 38624
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1171_
timestamp 1606120353
transform 1 0 27048 0 1 38624
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_12  FILLER_66_295
timestamp 1606120353
transform 1 0 28244 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_66_307
timestamp 1606120353
transform 1 0 29348 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_67_301
timestamp 1606120353
transform 1 0 28796 0 1 38624
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1182_
timestamp 1606120353
transform 1 0 29532 0 -1 38624
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1606120353
transform 1 0 29624 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_66_328
timestamp 1606120353
transform 1 0 31280 0 -1 38624
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_67_309
timestamp 1606120353
transform 1 0 29532 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_67_311
timestamp 1606120353
transform 1 0 29716 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_67_323
timestamp 1606120353
transform 1 0 30820 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1191_
timestamp 1606120353
transform 1 0 32108 0 -1 38624
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1606120353
transform 1 0 32016 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1606120353
transform 1 0 32476 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_67_335
timestamp 1606120353
transform 1 0 31924 0 1 38624
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_67_342
timestamp 1606120353
transform 1 0 32568 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1606120353
transform 1 0 35328 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_66_356
timestamp 1606120353
transform 1 0 33856 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_66_368
timestamp 1606120353
transform 1 0 34960 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_67_354
timestamp 1606120353
transform 1 0 33672 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_67_366
timestamp 1606120353
transform 1 0 34776 0 1 38624
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1606120353
transform 1 0 35420 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_66_380
timestamp 1606120353
transform 1 0 36064 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_66_392
timestamp 1606120353
transform 1 0 37168 0 -1 38624
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_66_396
timestamp 1606120353
transform 1 0 37536 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_67_385
timestamp 1606120353
transform 1 0 36524 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1606120353
transform -1 0 38548 0 -1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1606120353
transform -1 0 38548 0 1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1606120353
transform 1 0 37628 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1606120353
transform 1 0 38180 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_66_398
timestamp 1606120353
transform 1 0 37720 0 -1 38624
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILLER_67_397
timestamp 1606120353
transform 1 0 37628 0 1 38624
box 0 -48 552 592
<< labels >>
rlabel metal2 s 30838 0 30894 800 6 addr_r[0]
port 0 nsew default input
rlabel metal3 s 38852 36048 39652 36168 6 addr_r[10]
port 1 nsew default input
rlabel metal3 s 38852 9528 39652 9648 6 addr_r[11]
port 2 nsew default input
rlabel metal2 s 24398 40996 24454 41796 6 addr_r[12]
port 3 nsew default input
rlabel metal3 s 38852 28568 39652 28688 6 addr_r[13]
port 4 nsew default input
rlabel metal3 s 0 35368 800 35488 6 addr_r[1]
port 5 nsew default input
rlabel metal2 s 23018 40996 23074 41796 6 addr_r[2]
port 6 nsew default input
rlabel metal2 s 22558 0 22614 800 6 addr_r[3]
port 7 nsew default input
rlabel metal3 s 0 21088 800 21208 6 addr_r[4]
port 8 nsew default input
rlabel metal2 s 7838 40996 7894 41796 6 addr_r[5]
port 9 nsew default input
rlabel metal3 s 0 6128 800 6248 6 addr_r[6]
port 10 nsew default input
rlabel metal3 s 0 10888 800 11008 6 addr_r[7]
port 11 nsew default input
rlabel metal2 s 7378 0 7434 800 6 addr_r[8]
port 12 nsew default input
rlabel metal2 s 4158 40996 4214 41796 6 addr_r[9]
port 13 nsew default input
rlabel metal2 s 20718 0 20774 800 6 addr_w[0]
port 14 nsew default input
rlabel metal3 s 0 8168 800 8288 6 addr_w[10]
port 15 nsew default input
rlabel metal3 s 0 40808 800 40928 6 addr_w[11]
port 16 nsew default input
rlabel metal2 s 29458 0 29514 800 6 addr_w[12]
port 17 nsew default input
rlabel metal2 s 11978 0 12034 800 6 addr_w[13]
port 18 nsew default input
rlabel metal2 s 15658 0 15714 800 6 addr_w[1]
port 19 nsew default input
rlabel metal3 s 38852 4768 39652 4888 6 addr_w[2]
port 20 nsew default input
rlabel metal2 s 24398 0 24454 800 6 addr_w[3]
port 21 nsew default input
rlabel metal2 s 33138 0 33194 800 6 addr_w[4]
port 22 nsew default input
rlabel metal2 s 9678 40996 9734 41796 6 addr_w[5]
port 23 nsew default input
rlabel metal3 s 0 1368 800 1488 6 addr_w[6]
port 24 nsew default input
rlabel metal2 s 2778 0 2834 800 6 addr_w[7]
port 25 nsew default input
rlabel metal2 s 938 40996 994 41796 6 addr_w[8]
port 26 nsew default input
rlabel metal3 s 0 41488 800 41608 6 addr_w[9]
port 27 nsew default input
rlabel metal3 s 38852 17008 39652 17128 6 baseaddr_r_sync[0]
port 28 nsew default tristate
rlabel metal2 s 27618 40996 27674 41796 6 baseaddr_r_sync[1]
port 29 nsew default tristate
rlabel metal2 s 36358 0 36414 800 6 baseaddr_r_sync[2]
port 30 nsew default tristate
rlabel metal2 s 14278 0 14334 800 6 baseaddr_r_sync[3]
port 31 nsew default tristate
rlabel metal3 s 38852 2048 39652 2168 6 baseaddr_r_sync[4]
port 32 nsew default tristate
rlabel metal2 s 16118 0 16174 800 6 baseaddr_r_sync[5]
port 33 nsew default tristate
rlabel metal2 s 39118 0 39174 800 6 baseaddr_r_sync[6]
port 34 nsew default tristate
rlabel metal2 s 5538 40996 5594 41796 6 baseaddr_r_sync[7]
port 35 nsew default tristate
rlabel metal2 s 28538 40996 28594 41796 6 baseaddr_r_sync[8]
port 36 nsew default tristate
rlabel metal2 s 13818 40996 13874 41796 6 baseaddr_w_sync[0]
port 37 nsew default tristate
rlabel metal3 s 38852 36728 39652 36848 6 baseaddr_w_sync[1]
port 38 nsew default tristate
rlabel metal2 s 4618 0 4674 800 6 baseaddr_w_sync[2]
port 39 nsew default tristate
rlabel metal2 s 10598 40996 10654 41796 6 baseaddr_w_sync[3]
port 40 nsew default tristate
rlabel metal2 s 16118 40996 16174 41796 6 baseaddr_w_sync[4]
port 41 nsew default tristate
rlabel metal2 s 34518 40996 34574 41796 6 baseaddr_w_sync[5]
port 42 nsew default tristate
rlabel metal2 s 19798 0 19854 800 6 baseaddr_w_sync[6]
port 43 nsew default tristate
rlabel metal3 s 0 26528 800 26648 6 baseaddr_w_sync[7]
port 44 nsew default tristate
rlabel metal2 s 31298 0 31354 800 6 baseaddr_w_sync[8]
port 45 nsew default tristate
rlabel metal3 s 0 18368 800 18488 6 clk
port 46 nsew default input
rlabel metal2 s 26698 40996 26754 41796 6 conf[0]
port 47 nsew default input
rlabel metal2 s 14738 0 14794 800 6 conf[1]
port 48 nsew default input
rlabel metal3 s 38852 14288 39652 14408 6 conf[2]
port 49 nsew default input
rlabel metal2 s 34978 0 35034 800 6 csb
port 50 nsew default input
rlabel metal2 s 37738 40996 37794 41796 6 csb0_sync
port 51 nsew default tristate
rlabel metal2 s 3698 40996 3754 41796 6 csb1_sync
port 52 nsew default tristate
rlabel metal2 s 32218 0 32274 800 6 d_fabric_in[0]
port 53 nsew default input
rlabel metal2 s 25778 0 25834 800 6 d_fabric_in[10]
port 54 nsew default input
rlabel metal2 s 23478 40996 23534 41796 6 d_fabric_in[11]
port 55 nsew default input
rlabel metal3 s 38852 40128 39652 40248 6 d_fabric_in[12]
port 56 nsew default input
rlabel metal3 s 0 25168 800 25288 6 d_fabric_in[13]
port 57 nsew default input
rlabel metal3 s 0 688 800 808 6 d_fabric_in[14]
port 58 nsew default input
rlabel metal2 s 6458 40996 6514 41796 6 d_fabric_in[15]
port 59 nsew default input
rlabel metal2 s 29458 40996 29514 41796 6 d_fabric_in[16]
port 60 nsew default input
rlabel metal3 s 38852 39448 39652 39568 6 d_fabric_in[17]
port 61 nsew default input
rlabel metal3 s 38852 31288 39652 31408 6 d_fabric_in[18]
port 62 nsew default input
rlabel metal2 s 38198 40996 38254 41796 6 d_fabric_in[19]
port 63 nsew default input
rlabel metal3 s 0 5448 800 5568 6 d_fabric_in[1]
port 64 nsew default input
rlabel metal2 s 17038 0 17094 800 6 d_fabric_in[20]
port 65 nsew default input
rlabel metal3 s 38852 29248 39652 29368 6 d_fabric_in[21]
port 66 nsew default input
rlabel metal2 s 32678 0 32734 800 6 d_fabric_in[22]
port 67 nsew default input
rlabel metal3 s 38852 22448 39652 22568 6 d_fabric_in[23]
port 68 nsew default input
rlabel metal3 s 0 30608 800 30728 6 d_fabric_in[24]
port 69 nsew default input
rlabel metal2 s 31758 40996 31814 41796 6 d_fabric_in[25]
port 70 nsew default input
rlabel metal2 s 11058 40996 11114 41796 6 d_fabric_in[26]
port 71 nsew default input
rlabel metal2 s 2778 40996 2834 41796 6 d_fabric_in[27]
port 72 nsew default input
rlabel metal3 s 38852 19728 39652 19848 6 d_fabric_in[28]
port 73 nsew default input
rlabel metal3 s 38852 25168 39652 25288 6 d_fabric_in[29]
port 74 nsew default input
rlabel metal2 s 22098 0 22154 800 6 d_fabric_in[2]
port 75 nsew default input
rlabel metal2 s 35898 0 35954 800 6 d_fabric_in[30]
port 76 nsew default input
rlabel metal3 s 0 33328 800 33448 6 d_fabric_in[31]
port 77 nsew default input
rlabel metal2 s 27618 0 27674 800 6 d_fabric_in[3]
port 78 nsew default input
rlabel metal2 s 29918 40996 29974 41796 6 d_fabric_in[4]
port 79 nsew default input
rlabel metal2 s 26238 40996 26294 41796 6 d_fabric_in[5]
port 80 nsew default input
rlabel metal3 s 0 36048 800 36168 6 d_fabric_in[6]
port 81 nsew default input
rlabel metal3 s 38852 41488 39652 41608 6 d_fabric_in[7]
port 82 nsew default input
rlabel metal3 s 0 36728 800 36848 6 d_fabric_in[8]
port 83 nsew default input
rlabel metal2 s 938 0 994 800 6 d_fabric_in[9]
port 84 nsew default input
rlabel metal2 s 10598 0 10654 800 6 d_fabric_out[0]
port 85 nsew default tristate
rlabel metal3 s 0 2728 800 2848 6 d_fabric_out[10]
port 86 nsew default tristate
rlabel metal2 s 24858 0 24914 800 6 d_fabric_out[11]
port 87 nsew default tristate
rlabel metal3 s 38852 34008 39652 34128 6 d_fabric_out[12]
port 88 nsew default tristate
rlabel metal2 s 12438 0 12494 800 6 d_fabric_out[13]
port 89 nsew default tristate
rlabel metal2 s 26238 0 26294 800 6 d_fabric_out[14]
port 90 nsew default tristate
rlabel metal2 s 16578 40996 16634 41796 6 d_fabric_out[15]
port 91 nsew default tristate
rlabel metal3 s 38852 24488 39652 24608 6 d_fabric_out[16]
port 92 nsew default tristate
rlabel metal2 s 25778 40996 25834 41796 6 d_fabric_out[17]
port 93 nsew default tristate
rlabel metal2 s 21178 0 21234 800 6 d_fabric_out[18]
port 94 nsew default tristate
rlabel metal3 s 38852 3408 39652 3528 6 d_fabric_out[19]
port 95 nsew default tristate
rlabel metal2 s 23938 0 23994 800 6 d_fabric_out[1]
port 96 nsew default tristate
rlabel metal2 s 11058 0 11114 800 6 d_fabric_out[20]
port 97 nsew default tristate
rlabel metal3 s 0 23128 800 23248 6 d_fabric_out[21]
port 98 nsew default tristate
rlabel metal3 s 0 21768 800 21888 6 d_fabric_out[22]
port 99 nsew default tristate
rlabel metal3 s 0 17688 800 17808 6 d_fabric_out[23]
port 100 nsew default tristate
rlabel metal3 s 38852 14968 39652 15088 6 d_fabric_out[24]
port 101 nsew default tristate
rlabel metal3 s 0 3408 800 3528 6 d_fabric_out[25]
port 102 nsew default tristate
rlabel metal3 s 0 6808 800 6928 6 d_fabric_out[26]
port 103 nsew default tristate
rlabel metal3 s 0 11568 800 11688 6 d_fabric_out[27]
port 104 nsew default tristate
rlabel metal2 s 17498 40996 17554 41796 6 d_fabric_out[28]
port 105 nsew default tristate
rlabel metal3 s 0 38768 800 38888 6 d_fabric_out[29]
port 106 nsew default tristate
rlabel metal2 s 14278 40996 14334 41796 6 d_fabric_out[2]
port 107 nsew default tristate
rlabel metal2 s 19798 40996 19854 41796 6 d_fabric_out[30]
port 108 nsew default tristate
rlabel metal2 s 39578 40996 39634 41796 6 d_fabric_out[31]
port 109 nsew default tristate
rlabel metal2 s 32678 40996 32734 41796 6 d_fabric_out[3]
port 110 nsew default tristate
rlabel metal2 s 28078 0 28134 800 6 d_fabric_out[4]
port 111 nsew default tristate
rlabel metal3 s 38852 32648 39652 32768 6 d_fabric_out[5]
port 112 nsew default tristate
rlabel metal3 s 38852 29928 39652 30048 6 d_fabric_out[6]
port 113 nsew default tristate
rlabel metal3 s 38852 21088 39652 21208 6 d_fabric_out[7]
port 114 nsew default tristate
rlabel metal3 s 0 20408 800 20528 6 d_fabric_out[8]
port 115 nsew default tristate
rlabel metal3 s 0 38088 800 38208 6 d_fabric_out[9]
port 116 nsew default tristate
rlabel metal2 s 478 0 534 800 6 d_sram_in[0]
port 117 nsew default tristate
rlabel metal3 s 38852 12248 39652 12368 6 d_sram_in[10]
port 118 nsew default tristate
rlabel metal3 s 38852 11568 39652 11688 6 d_sram_in[11]
port 119 nsew default tristate
rlabel metal2 s 20718 40996 20774 41796 6 d_sram_in[12]
port 120 nsew default tristate
rlabel metal2 s 1398 40996 1454 41796 6 d_sram_in[13]
port 121 nsew default tristate
rlabel metal3 s 0 4088 800 4208 6 d_sram_in[14]
port 122 nsew default tristate
rlabel metal3 s 0 25848 800 25968 6 d_sram_in[15]
port 123 nsew default tristate
rlabel metal3 s 38852 7488 39652 7608 6 d_sram_in[16]
port 124 nsew default tristate
rlabel metal3 s 38852 8 39652 128 6 d_sram_in[17]
port 125 nsew default tristate
rlabel metal2 s 1858 0 1914 800 6 d_sram_in[18]
port 126 nsew default tristate
rlabel metal3 s 38852 37408 39652 37528 6 d_sram_in[19]
port 127 nsew default tristate
rlabel metal2 s 14738 40996 14794 41796 6 d_sram_in[1]
port 128 nsew default tristate
rlabel metal2 s 8758 40996 8814 41796 6 d_sram_in[20]
port 129 nsew default tristate
rlabel metal3 s 38852 27208 39652 27328 6 d_sram_in[21]
port 130 nsew default tristate
rlabel metal2 s 13818 0 13874 800 6 d_sram_in[22]
port 131 nsew default tristate
rlabel metal2 s 17498 0 17554 800 6 d_sram_in[23]
port 132 nsew default tristate
rlabel metal2 s 37278 0 37334 800 6 d_sram_in[24]
port 133 nsew default tristate
rlabel metal2 s 36358 40996 36414 41796 6 d_sram_in[25]
port 134 nsew default tristate
rlabel metal2 s 6918 0 6974 800 6 d_sram_in[26]
port 135 nsew default tristate
rlabel metal2 s 12898 40996 12954 41796 6 d_sram_in[27]
port 136 nsew default tristate
rlabel metal3 s 0 31288 800 31408 6 d_sram_in[28]
port 137 nsew default tristate
rlabel metal2 s 37738 0 37794 800 6 d_sram_in[29]
port 138 nsew default tristate
rlabel metal2 s 5538 0 5594 800 6 d_sram_in[2]
port 139 nsew default tristate
rlabel metal2 s 21178 40996 21234 41796 6 d_sram_in[30]
port 140 nsew default tristate
rlabel metal3 s 38852 6128 39652 6248 6 d_sram_in[31]
port 141 nsew default tristate
rlabel metal2 s 478 40996 534 41796 6 d_sram_in[3]
port 142 nsew default tristate
rlabel metal2 s 17958 40996 18014 41796 6 d_sram_in[4]
port 143 nsew default tristate
rlabel metal3 s 38852 10208 39652 10328 6 d_sram_in[5]
port 144 nsew default tristate
rlabel metal2 s 7378 40996 7434 41796 6 d_sram_in[6]
port 145 nsew default tristate
rlabel metal2 s 28998 0 29054 800 6 d_sram_in[7]
port 146 nsew default tristate
rlabel metal2 s 27158 0 27214 800 6 d_sram_in[8]
port 147 nsew default tristate
rlabel metal3 s 38852 13608 39652 13728 6 d_sram_in[9]
port 148 nsew default tristate
rlabel metal3 s 0 28568 800 28688 6 d_sram_out[0]
port 149 nsew default input
rlabel metal2 s 7838 0 7894 800 6 d_sram_out[10]
port 150 nsew default input
rlabel metal3 s 0 29248 800 29368 6 d_sram_out[11]
port 151 nsew default input
rlabel metal2 s 5998 40996 6054 41796 6 d_sram_out[12]
port 152 nsew default input
rlabel metal2 s 22558 40996 22614 41796 6 d_sram_out[13]
port 153 nsew default input
rlabel metal3 s 0 12928 800 13048 6 d_sram_out[14]
port 154 nsew default input
rlabel metal2 s 34978 40996 35034 41796 6 d_sram_out[15]
port 155 nsew default input
rlabel metal2 s 9218 0 9274 800 6 d_sram_out[16]
port 156 nsew default input
rlabel metal3 s 38852 38768 39652 38888 6 d_sram_out[17]
port 157 nsew default input
rlabel metal2 s 19338 0 19394 800 6 d_sram_out[18]
port 158 nsew default input
rlabel metal2 s 33138 40996 33194 41796 6 d_sram_out[19]
port 159 nsew default input
rlabel metal3 s 38852 26528 39652 26648 6 d_sram_out[1]
port 160 nsew default input
rlabel metal2 s 39578 0 39634 800 6 d_sram_out[20]
port 161 nsew default input
rlabel metal3 s 0 13608 800 13728 6 d_sram_out[21]
port 162 nsew default input
rlabel metal2 s 2318 0 2374 800 6 d_sram_out[22]
port 163 nsew default input
rlabel metal2 s 33598 40996 33654 41796 6 d_sram_out[23]
port 164 nsew default input
rlabel metal2 s 34058 0 34114 800 6 d_sram_out[24]
port 165 nsew default input
rlabel metal3 s 0 10208 800 10328 6 d_sram_out[25]
port 166 nsew default input
rlabel metal2 s 35898 40996 35954 41796 6 d_sram_out[26]
port 167 nsew default input
rlabel metal2 s 38198 0 38254 800 6 d_sram_out[27]
port 168 nsew default input
rlabel metal2 s 9678 0 9734 800 6 d_sram_out[28]
port 169 nsew default input
rlabel metal2 s 23018 0 23074 800 6 d_sram_out[29]
port 170 nsew default input
rlabel metal3 s 38852 34688 39652 34808 6 d_sram_out[2]
port 171 nsew default input
rlabel metal3 s 0 32648 800 32768 6 d_sram_out[30]
port 172 nsew default input
rlabel metal3 s 0 40128 800 40248 6 d_sram_out[31]
port 173 nsew default input
rlabel metal3 s 38852 8848 39652 8968 6 d_sram_out[3]
port 174 nsew default input
rlabel metal2 s 8758 0 8814 800 6 d_sram_out[4]
port 175 nsew default input
rlabel metal2 s 3698 0 3754 800 6 d_sram_out[5]
port 176 nsew default input
rlabel metal3 s 38852 21768 39652 21888 6 d_sram_out[6]
port 177 nsew default input
rlabel metal2 s 4618 40996 4674 41796 6 d_sram_out[7]
port 178 nsew default input
rlabel metal3 s 0 23808 800 23928 6 d_sram_out[8]
port 179 nsew default input
rlabel metal3 s 0 16328 800 16448 6 d_sram_out[9]
port 180 nsew default input
rlabel metal2 s 30838 40996 30894 41796 6 out_reg
port 181 nsew default input
rlabel metal3 s 0 19048 800 19168 6 reb
port 182 nsew default input
rlabel metal2 s 34518 0 34574 800 6 w_mask[0]
port 183 nsew default tristate
rlabel metal2 s 19338 40996 19394 41796 6 w_mask[10]
port 184 nsew default tristate
rlabel metal3 s 38852 31968 39652 32088 6 w_mask[11]
port 185 nsew default tristate
rlabel metal2 s 18 0 74 800 6 w_mask[12]
port 186 nsew default tristate
rlabel metal3 s 0 15648 800 15768 6 w_mask[13]
port 187 nsew default tristate
rlabel metal2 s 12898 0 12954 800 6 w_mask[14]
port 188 nsew default tristate
rlabel metal2 s 5998 0 6054 800 6 w_mask[15]
port 189 nsew default tristate
rlabel metal2 s 31298 40996 31354 41796 6 w_mask[16]
port 190 nsew default tristate
rlabel metal2 s 38658 40996 38714 41796 6 w_mask[17]
port 191 nsew default tristate
rlabel metal3 s 38852 23808 39652 23928 6 w_mask[18]
port 192 nsew default tristate
rlabel metal2 s 18878 0 18934 800 6 w_mask[19]
port 193 nsew default tristate
rlabel metal2 s 29918 0 29974 800 6 w_mask[1]
port 194 nsew default tristate
rlabel metal2 s 12438 40996 12494 41796 6 w_mask[20]
port 195 nsew default tristate
rlabel metal2 s 2318 40996 2374 41796 6 w_mask[21]
port 196 nsew default tristate
rlabel metal2 s 28078 40996 28134 41796 6 w_mask[22]
port 197 nsew default tristate
rlabel metal3 s 0 8848 800 8968 6 w_mask[23]
port 198 nsew default tristate
rlabel metal2 s 4158 0 4214 800 6 w_mask[24]
port 199 nsew default tristate
rlabel metal3 s 0 34008 800 34128 6 w_mask[25]
port 200 nsew default tristate
rlabel metal2 s 24858 40996 24914 41796 6 w_mask[26]
port 201 nsew default tristate
rlabel metal2 s 11518 40996 11574 41796 6 w_mask[27]
port 202 nsew default tristate
rlabel metal2 s 21638 40996 21694 41796 6 w_mask[28]
port 203 nsew default tristate
rlabel metal2 s 36818 40996 36874 41796 6 w_mask[29]
port 204 nsew default tristate
rlabel metal2 s 15658 40996 15714 41796 6 w_mask[2]
port 205 nsew default tristate
rlabel metal2 s 17958 0 18014 800 6 w_mask[30]
port 206 nsew default tristate
rlabel metal3 s 0 14288 800 14408 6 w_mask[31]
port 207 nsew default tristate
rlabel metal3 s 38852 19048 39652 19168 6 w_mask[3]
port 208 nsew default tristate
rlabel metal3 s 38852 16328 39652 16448 6 w_mask[4]
port 209 nsew default tristate
rlabel metal2 s 18418 40996 18474 41796 6 w_mask[5]
port 210 nsew default tristate
rlabel metal3 s 38852 6808 39652 6928 6 w_mask[6]
port 211 nsew default tristate
rlabel metal3 s 38852 1368 39652 1488 6 w_mask[7]
port 212 nsew default tristate
rlabel metal3 s 38852 17688 39652 17808 6 w_mask[8]
port 213 nsew default tristate
rlabel metal3 s 38852 4088 39652 4208 6 w_mask[9]
port 214 nsew default tristate
rlabel metal2 s 9218 40996 9274 41796 6 web
port 215 nsew default input
rlabel metal3 s 0 27888 800 28008 6 web0_sync
port 216 nsew default tristate
rlabel metal5 s 1104 5298 38548 5618 6 VPWR
port 217 nsew default input
rlabel metal5 s 1104 20616 38548 20936 6 VGND
port 218 nsew default input
<< end >>
