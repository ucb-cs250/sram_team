magic
tech sky130A
magscale 1 2
timestamp 1607420259
<< checkpaint >>
rect -3932 -3652 23932 83593
<< locali >>
rect 9689 70295 9723 70533
rect 11345 64855 11379 65161
rect 11345 63767 11379 63869
rect 3157 61591 3191 61897
rect 9045 56695 9079 57001
rect 12817 55675 12851 55913
rect 5917 51255 5951 51561
rect 5457 50779 5491 51017
rect 6193 50711 6227 51017
rect 8769 50847 8803 51017
rect 13185 50711 13219 51017
rect 14473 50847 14507 51017
rect 9229 49623 9263 49929
rect 9505 49623 9539 49929
rect 14933 49623 14967 49929
rect 7205 47991 7239 48229
rect 10517 42619 10551 42857
rect 14289 42551 14323 42857
rect 10057 38267 10091 38437
rect 14473 36635 14507 36805
rect 15853 30583 15887 30821
rect 12449 25687 12483 25857
rect 13645 25143 13679 25449
rect 12909 21335 12943 21437
rect 6377 18071 6411 18173
rect 14473 14807 14507 14909
rect 12265 14263 12299 14569
rect 11345 13855 11379 14025
<< viali >>
rect 4353 75429 4387 75463
rect 5181 75361 5215 75395
rect 7113 75361 7147 75395
rect 4905 75293 4939 75327
rect 5365 75293 5399 75327
rect 2237 75157 2271 75191
rect 4169 75157 4203 75191
rect 7297 75157 7331 75191
rect 3525 74953 3559 74987
rect 5825 74953 5859 74987
rect 7021 74953 7055 74987
rect 2053 74885 2087 74919
rect 2145 74817 2179 74851
rect 3893 74817 3927 74851
rect 2697 74749 2731 74783
rect 2973 74749 3007 74783
rect 3157 74749 3191 74783
rect 4445 74749 4479 74783
rect 4721 74749 4755 74783
rect 6469 74749 6503 74783
rect 6929 74749 6963 74783
rect 7481 74749 7515 74783
rect 6837 74681 6871 74715
rect 4261 74613 4295 74647
rect 4261 74409 4295 74443
rect 6469 74409 6503 74443
rect 5181 74341 5215 74375
rect 7665 74341 7699 74375
rect 2973 74273 3007 74307
rect 5365 74273 5399 74307
rect 7757 74273 7791 74307
rect 2697 74205 2731 74239
rect 4997 74205 5031 74239
rect 4721 74137 4755 74171
rect 7021 74137 7055 74171
rect 2237 74069 2271 74103
rect 5457 74069 5491 74103
rect 6193 74069 6227 74103
rect 10149 74069 10183 74103
rect 2145 73865 2179 73899
rect 2881 73865 2915 73899
rect 3525 73797 3559 73831
rect 3893 73729 3927 73763
rect 6101 73729 6135 73763
rect 6377 73729 6411 73763
rect 10701 73729 10735 73763
rect 2513 73661 2547 73695
rect 2789 73661 2823 73695
rect 4813 73661 4847 73695
rect 5089 73661 5123 73695
rect 5273 73661 5307 73695
rect 5641 73661 5675 73695
rect 9505 73661 9539 73695
rect 10057 73661 10091 73695
rect 10609 73661 10643 73695
rect 10793 73661 10827 73695
rect 2605 73593 2639 73627
rect 4261 73593 4295 73627
rect 8033 73593 8067 73627
rect 9965 73593 9999 73627
rect 5917 73525 5951 73559
rect 7481 73525 7515 73559
rect 2697 73321 2731 73355
rect 9321 73321 9355 73355
rect 2973 73253 3007 73287
rect 4813 73253 4847 73287
rect 3801 73185 3835 73219
rect 4353 73185 4387 73219
rect 5365 73185 5399 73219
rect 5641 73185 5675 73219
rect 6929 73185 6963 73219
rect 7389 73185 7423 73219
rect 8953 73185 8987 73219
rect 9689 73185 9723 73219
rect 10057 73185 10091 73219
rect 3525 73117 3559 73151
rect 3985 73117 4019 73151
rect 5825 73117 5859 73151
rect 9045 73117 9079 73151
rect 10885 73117 10919 73151
rect 6929 73049 6963 73083
rect 4721 72981 4755 73015
rect 6469 72981 6503 73015
rect 8217 72981 8251 73015
rect 11161 72981 11195 73015
rect 2697 72777 2731 72811
rect 3065 72777 3099 72811
rect 3893 72777 3927 72811
rect 7757 72777 7791 72811
rect 8401 72777 8435 72811
rect 11161 72709 11195 72743
rect 4537 72641 4571 72675
rect 5089 72641 5123 72675
rect 6377 72641 6411 72675
rect 10333 72641 10367 72675
rect 5365 72573 5399 72607
rect 5549 72573 5583 72607
rect 6653 72573 6687 72607
rect 10885 72573 10919 72607
rect 11437 72573 11471 72607
rect 11805 72573 11839 72607
rect 11989 72573 12023 72607
rect 4445 72505 4479 72539
rect 8861 72505 8895 72539
rect 12725 72505 12759 72539
rect 3433 72437 3467 72471
rect 5825 72437 5859 72471
rect 6193 72437 6227 72471
rect 9229 72437 9263 72471
rect 9965 72437 9999 72471
rect 10701 72437 10735 72471
rect 4997 72233 5031 72267
rect 5549 72233 5583 72267
rect 6193 72233 6227 72267
rect 10885 72233 10919 72267
rect 3617 72097 3651 72131
rect 3893 72097 3927 72131
rect 7113 72097 7147 72131
rect 8677 72097 8711 72131
rect 9321 72097 9355 72131
rect 9689 72097 9723 72131
rect 8585 72029 8619 72063
rect 8861 72029 8895 72063
rect 6561 71961 6595 71995
rect 7297 71961 7331 71995
rect 7757 71893 7791 71927
rect 11253 71893 11287 71927
rect 3249 71689 3283 71723
rect 4629 71689 4663 71723
rect 6193 71689 6227 71723
rect 6837 71689 6871 71723
rect 9137 71689 9171 71723
rect 17509 71689 17543 71723
rect 4813 71553 4847 71587
rect 7205 71553 7239 71587
rect 10609 71553 10643 71587
rect 12909 71553 12943 71587
rect 5089 71485 5123 71519
rect 7665 71485 7699 71519
rect 8217 71485 8251 71519
rect 8585 71485 8619 71519
rect 11161 71485 11195 71519
rect 11253 71485 11287 71519
rect 11437 71485 11471 71519
rect 11713 71485 11747 71519
rect 11897 71485 11931 71519
rect 12817 71485 12851 71519
rect 13001 71485 13035 71519
rect 16129 71485 16163 71519
rect 16405 71485 16439 71519
rect 8769 71417 8803 71451
rect 10517 71417 10551 71451
rect 3709 71349 3743 71383
rect 7481 71349 7515 71383
rect 9413 71349 9447 71383
rect 10149 71349 10183 71383
rect 16037 71349 16071 71383
rect 5457 71145 5491 71179
rect 8217 71145 8251 71179
rect 11069 71145 11103 71179
rect 10701 71077 10735 71111
rect 4353 71009 4387 71043
rect 4721 71009 4755 71043
rect 5181 71009 5215 71043
rect 7481 71009 7515 71043
rect 8953 71009 8987 71043
rect 6837 70941 6871 70975
rect 9597 70941 9631 70975
rect 4169 70873 4203 70907
rect 8493 70805 8527 70839
rect 9965 70805 9999 70839
rect 10241 70805 10275 70839
rect 11897 70805 11931 70839
rect 16129 70805 16163 70839
rect 2053 70601 2087 70635
rect 4353 70601 4387 70635
rect 5917 70601 5951 70635
rect 7113 70601 7147 70635
rect 11897 70601 11931 70635
rect 9505 70533 9539 70567
rect 9689 70533 9723 70567
rect 5733 70465 5767 70499
rect 7849 70465 7883 70499
rect 8309 70465 8343 70499
rect 9045 70465 9079 70499
rect 5917 70397 5951 70431
rect 6561 70397 6595 70431
rect 8217 70397 8251 70431
rect 8585 70397 8619 70431
rect 8677 70397 8711 70431
rect 10793 70465 10827 70499
rect 9965 70397 9999 70431
rect 10149 70397 10183 70431
rect 10517 70397 10551 70431
rect 11989 70397 12023 70431
rect 12173 70397 12207 70431
rect 12541 70397 12575 70431
rect 1685 70261 1719 70295
rect 4629 70261 4663 70295
rect 7481 70261 7515 70295
rect 9689 70261 9723 70295
rect 11713 70261 11747 70295
rect 6653 70057 6687 70091
rect 8769 70057 8803 70091
rect 11069 69989 11103 70023
rect 1501 69921 1535 69955
rect 5089 69921 5123 69955
rect 7113 69921 7147 69955
rect 9505 69921 9539 69955
rect 9689 69921 9723 69955
rect 10057 69921 10091 69955
rect 10609 69921 10643 69955
rect 1777 69853 1811 69887
rect 6837 69853 6871 69887
rect 9781 69853 9815 69887
rect 12173 69785 12207 69819
rect 2881 69717 2915 69751
rect 4169 69717 4203 69751
rect 5273 69717 5307 69751
rect 5825 69717 5859 69751
rect 8401 69717 8435 69751
rect 9229 69717 9263 69751
rect 11897 69717 11931 69751
rect 5733 69513 5767 69547
rect 9873 69513 9907 69547
rect 4169 69445 4203 69479
rect 1777 69377 1811 69411
rect 5825 69377 5859 69411
rect 6837 69377 6871 69411
rect 7665 69377 7699 69411
rect 9137 69377 9171 69411
rect 12173 69377 12207 69411
rect 2329 69309 2363 69343
rect 4077 69309 4111 69343
rect 4629 69309 4663 69343
rect 6377 69309 6411 69343
rect 6653 69309 6687 69343
rect 7573 69309 7607 69343
rect 8217 69309 8251 69343
rect 9965 69309 9999 69343
rect 10149 69309 10183 69343
rect 10517 69309 10551 69343
rect 11253 69309 11287 69343
rect 12081 69309 12115 69343
rect 12449 69309 12483 69343
rect 12817 69309 12851 69343
rect 2145 69241 2179 69275
rect 8769 69241 8803 69275
rect 11621 69241 11655 69275
rect 2421 69173 2455 69207
rect 3065 69173 3099 69207
rect 3433 69173 3467 69207
rect 3801 69173 3835 69207
rect 5089 69173 5123 69207
rect 7205 69173 7239 69207
rect 9505 69173 9539 69207
rect 11897 69173 11931 69207
rect 5549 68969 5583 69003
rect 6285 68969 6319 69003
rect 3525 68901 3559 68935
rect 13829 68901 13863 68935
rect 2237 68833 2271 68867
rect 2513 68833 2547 68867
rect 4353 68833 4387 68867
rect 5365 68833 5399 68867
rect 8033 68833 8067 68867
rect 8401 68833 8435 68867
rect 9689 68833 9723 68867
rect 9781 68833 9815 68867
rect 10425 68833 10459 68867
rect 10701 68833 10735 68867
rect 12449 68833 12483 68867
rect 14013 68833 14047 68867
rect 1685 68765 1719 68799
rect 2697 68765 2731 68799
rect 4077 68765 4111 68799
rect 4537 68765 4571 68799
rect 7389 68765 7423 68799
rect 7941 68765 7975 68799
rect 8309 68765 8343 68799
rect 10057 68765 10091 68799
rect 14381 68765 14415 68799
rect 4905 68697 4939 68731
rect 5917 68697 5951 68731
rect 8953 68697 8987 68731
rect 2973 68629 3007 68663
rect 3433 68629 3467 68663
rect 6561 68629 6595 68663
rect 7297 68629 7331 68663
rect 9229 68629 9263 68663
rect 11253 68629 11287 68663
rect 11621 68629 11655 68663
rect 12081 68629 12115 68663
rect 12633 68629 12667 68663
rect 12909 68629 12943 68663
rect 13369 68629 13403 68663
rect 16129 68629 16163 68663
rect 6745 68425 6779 68459
rect 7481 68425 7515 68459
rect 17509 68425 17543 68459
rect 7113 68357 7147 68391
rect 1501 68289 1535 68323
rect 1777 68289 1811 68323
rect 3893 68289 3927 68323
rect 9137 68289 9171 68323
rect 11713 68289 11747 68323
rect 16037 68289 16071 68323
rect 4077 68221 4111 68255
rect 4353 68221 4387 68255
rect 6469 68221 6503 68255
rect 6561 68221 6595 68255
rect 7665 68221 7699 68255
rect 9781 68221 9815 68255
rect 11069 68221 11103 68255
rect 11161 68221 11195 68255
rect 11529 68221 11563 68255
rect 12817 68221 12851 68255
rect 13185 68221 13219 68255
rect 13369 68221 13403 68255
rect 16129 68221 16163 68255
rect 16405 68221 16439 68255
rect 3433 68153 3467 68187
rect 6009 68153 6043 68187
rect 10333 68153 10367 68187
rect 2881 68085 2915 68119
rect 5457 68085 5491 68119
rect 8033 68085 8067 68119
rect 8677 68085 8711 68119
rect 9505 68085 9539 68119
rect 9965 68085 9999 68119
rect 10701 68085 10735 68119
rect 12449 68085 12483 68119
rect 13921 68085 13955 68119
rect 14289 68085 14323 68119
rect 1685 67881 1719 67915
rect 3525 67881 3559 67915
rect 4077 67881 4111 67915
rect 4905 67881 4939 67915
rect 7941 67881 7975 67915
rect 9781 67881 9815 67915
rect 3065 67813 3099 67847
rect 7573 67813 7607 67847
rect 10241 67813 10275 67847
rect 2605 67745 2639 67779
rect 3617 67745 3651 67779
rect 4813 67745 4847 67779
rect 5457 67745 5491 67779
rect 7481 67745 7515 67779
rect 9321 67745 9355 67779
rect 10609 67745 10643 67779
rect 10977 67745 11011 67779
rect 11345 67745 11379 67779
rect 12449 67745 12483 67779
rect 13001 67745 13035 67779
rect 13185 67745 13219 67779
rect 15761 67745 15795 67779
rect 1777 67677 1811 67711
rect 2329 67677 2363 67711
rect 2789 67677 2823 67711
rect 5641 67677 5675 67711
rect 11529 67677 11563 67711
rect 12173 67677 12207 67711
rect 15485 67677 15519 67711
rect 17141 67677 17175 67711
rect 3801 67609 3835 67643
rect 4721 67609 4755 67643
rect 9505 67609 9539 67643
rect 6193 67541 6227 67575
rect 8217 67541 8251 67575
rect 12541 67541 12575 67575
rect 2881 67337 2915 67371
rect 4905 67337 4939 67371
rect 6745 67337 6779 67371
rect 7297 67337 7331 67371
rect 13645 67337 13679 67371
rect 14381 67269 14415 67303
rect 5365 67201 5399 67235
rect 6377 67201 6411 67235
rect 8217 67201 8251 67235
rect 10517 67201 10551 67235
rect 16037 67201 16071 67235
rect 1869 67133 1903 67167
rect 4261 67133 4295 67167
rect 5917 67133 5951 67167
rect 6193 67133 6227 67167
rect 7205 67133 7239 67167
rect 7941 67133 7975 67167
rect 9689 67133 9723 67167
rect 10057 67133 10091 67167
rect 10425 67133 10459 67167
rect 12173 67133 12207 67167
rect 12541 67133 12575 67167
rect 12909 67133 12943 67167
rect 14197 67133 14231 67167
rect 14657 67133 14691 67167
rect 15117 67133 15151 67167
rect 16129 67133 16163 67167
rect 16405 67133 16439 67167
rect 2237 67065 2271 67099
rect 7113 67065 7147 67099
rect 13277 67065 13311 67099
rect 2605 66997 2639 67031
rect 3617 66997 3651 67031
rect 4445 66997 4479 67031
rect 5181 66997 5215 67031
rect 8585 66997 8619 67031
rect 9045 66997 9079 67031
rect 9505 66997 9539 67031
rect 11253 66997 11287 67031
rect 11621 66997 11655 67031
rect 11989 66997 12023 67031
rect 14013 66997 14047 67031
rect 15485 66997 15519 67031
rect 17509 66997 17543 67031
rect 2053 66793 2087 66827
rect 2513 66793 2547 66827
rect 3801 66793 3835 66827
rect 4261 66793 4295 66827
rect 9321 66793 9355 66827
rect 16957 66793 16991 66827
rect 2237 66725 2271 66759
rect 2421 66657 2455 66691
rect 3617 66657 3651 66691
rect 5273 66657 5307 66691
rect 5825 66657 5859 66691
rect 7481 66657 7515 66691
rect 8493 66657 8527 66691
rect 9597 66657 9631 66691
rect 9873 66657 9907 66691
rect 10241 66657 10275 66691
rect 12449 66657 12483 66691
rect 12909 66657 12943 66691
rect 13185 66657 13219 66691
rect 15025 66657 15059 66691
rect 5549 66589 5583 66623
rect 6193 66589 6227 66623
rect 9689 66589 9723 66623
rect 11897 66589 11931 66623
rect 15301 66589 15335 66623
rect 16681 66589 16715 66623
rect 8677 66521 8711 66555
rect 1685 66453 1719 66487
rect 4997 66453 5031 66487
rect 6653 66453 6687 66487
rect 7113 66453 7147 66487
rect 7665 66453 7699 66487
rect 11069 66453 11103 66487
rect 12265 66453 12299 66487
rect 12541 66453 12575 66487
rect 1777 66249 1811 66283
rect 2513 66249 2547 66283
rect 2881 66249 2915 66283
rect 6837 66249 6871 66283
rect 14381 66249 14415 66283
rect 4997 66181 5031 66215
rect 11529 66181 11563 66215
rect 13645 66181 13679 66215
rect 4445 66113 4479 66147
rect 5733 66113 5767 66147
rect 6469 66113 6503 66147
rect 13001 66113 13035 66147
rect 15117 66113 15151 66147
rect 15577 66113 15611 66147
rect 1593 66045 1627 66079
rect 2973 66045 3007 66079
rect 5089 66045 5123 66079
rect 5549 66045 5583 66079
rect 7297 66045 7331 66079
rect 7573 66045 7607 66079
rect 8125 66045 8159 66079
rect 8585 66045 8619 66079
rect 10141 66045 10175 66079
rect 10609 66045 10643 66079
rect 11345 66045 11379 66079
rect 12081 66045 12115 66079
rect 12633 66045 12667 66079
rect 13277 66045 13311 66079
rect 15301 66045 15335 66079
rect 4813 65977 4847 66011
rect 2053 65909 2087 65943
rect 3157 65909 3191 65943
rect 3617 65909 3651 65943
rect 7849 65909 7883 65943
rect 9137 65909 9171 65943
rect 9413 65909 9447 65943
rect 9965 65909 9999 65943
rect 10333 65909 10367 65943
rect 11253 65909 11287 65943
rect 12541 65909 12575 65943
rect 14749 65909 14783 65943
rect 16681 65909 16715 65943
rect 2605 65705 2639 65739
rect 7113 65705 7147 65739
rect 11069 65705 11103 65739
rect 13001 65705 13035 65739
rect 14749 65705 14783 65739
rect 15393 65705 15427 65739
rect 16129 65705 16163 65739
rect 2973 65637 3007 65671
rect 10977 65637 11011 65671
rect 11161 65637 11195 65671
rect 12725 65637 12759 65671
rect 3157 65569 3191 65603
rect 4169 65569 4203 65603
rect 6653 65569 6687 65603
rect 7481 65569 7515 65603
rect 7941 65569 7975 65603
rect 8217 65569 8251 65603
rect 8677 65569 8711 65603
rect 9045 65569 9079 65603
rect 13369 65569 13403 65603
rect 4445 65501 4479 65535
rect 8033 65501 8067 65535
rect 10793 65501 10827 65535
rect 11529 65501 11563 65535
rect 13645 65501 13679 65535
rect 3341 65433 3375 65467
rect 9689 65433 9723 65467
rect 2237 65365 2271 65399
rect 3709 65365 3743 65399
rect 4077 65365 4111 65399
rect 5549 65365 5583 65399
rect 6101 65365 6135 65399
rect 10149 65365 10183 65399
rect 11897 65365 11931 65399
rect 3249 65161 3283 65195
rect 5273 65161 5307 65195
rect 7021 65161 7055 65195
rect 7941 65161 7975 65195
rect 9505 65161 9539 65195
rect 11345 65161 11379 65195
rect 13185 65161 13219 65195
rect 17509 65161 17543 65195
rect 2697 65025 2731 65059
rect 5641 65025 5675 65059
rect 5917 65025 5951 65059
rect 10609 65025 10643 65059
rect 2237 64957 2271 64991
rect 2421 64957 2455 64991
rect 4353 64957 4387 64991
rect 4629 64957 4663 64991
rect 4813 64957 4847 64991
rect 8585 64957 8619 64991
rect 10149 64957 10183 64991
rect 10701 64957 10735 64991
rect 2145 64889 2179 64923
rect 3893 64889 3927 64923
rect 9045 64889 9079 64923
rect 10057 64889 10091 64923
rect 16037 65025 16071 65059
rect 12357 64957 12391 64991
rect 12449 64957 12483 64991
rect 13277 64957 13311 64991
rect 14105 64957 14139 64991
rect 16129 64957 16163 64991
rect 16405 64957 16439 64991
rect 13829 64889 13863 64923
rect 1777 64821 1811 64855
rect 7573 64821 7607 64855
rect 8401 64821 8435 64855
rect 8769 64821 8803 64855
rect 11161 64821 11195 64855
rect 11345 64821 11379 64855
rect 11621 64821 11655 64855
rect 13461 64821 13495 64855
rect 6653 64617 6687 64651
rect 9965 64617 9999 64651
rect 7113 64549 7147 64583
rect 2789 64481 2823 64515
rect 5273 64481 5307 64515
rect 7573 64481 7607 64515
rect 8401 64481 8435 64515
rect 8861 64481 8895 64515
rect 10149 64481 10183 64515
rect 10333 64481 10367 64515
rect 10701 64481 10735 64515
rect 11253 64481 11287 64515
rect 13277 64481 13311 64515
rect 15485 64481 15519 64515
rect 3065 64413 3099 64447
rect 7849 64413 7883 64447
rect 11621 64413 11655 64447
rect 13001 64413 13035 64447
rect 14381 64413 14415 64447
rect 15761 64413 15795 64447
rect 16865 64413 16899 64447
rect 2237 64345 2271 64379
rect 6285 64345 6319 64379
rect 8125 64345 8159 64379
rect 1685 64277 1719 64311
rect 2605 64277 2639 64311
rect 4169 64277 4203 64311
rect 4997 64277 5031 64311
rect 5457 64277 5491 64311
rect 5825 64277 5859 64311
rect 9321 64277 9355 64311
rect 9781 64277 9815 64311
rect 6377 64073 6411 64107
rect 9505 64073 9539 64107
rect 15117 64073 15151 64107
rect 2053 64005 2087 64039
rect 3893 64005 3927 64039
rect 11069 63937 11103 63971
rect 16037 63937 16071 63971
rect 2697 63869 2731 63903
rect 2973 63869 3007 63903
rect 3157 63869 3191 63903
rect 4537 63869 4571 63903
rect 5273 63869 5307 63903
rect 5457 63869 5491 63903
rect 7113 63869 7147 63903
rect 7297 63869 7331 63903
rect 7941 63869 7975 63903
rect 8125 63869 8159 63903
rect 8493 63869 8527 63903
rect 9781 63869 9815 63903
rect 10333 63869 10367 63903
rect 10517 63869 10551 63903
rect 11345 63869 11379 63903
rect 11621 63869 11655 63903
rect 12081 63869 12115 63903
rect 12449 63869 12483 63903
rect 13093 63869 13127 63903
rect 13553 63869 13587 63903
rect 14013 63869 14047 63903
rect 14565 63869 14599 63903
rect 16129 63869 16163 63903
rect 16405 63869 16439 63903
rect 2145 63801 2179 63835
rect 3525 63801 3559 63835
rect 7205 63801 7239 63835
rect 9137 63801 9171 63835
rect 13369 63801 13403 63835
rect 1685 63733 1719 63767
rect 4813 63733 4847 63767
rect 5089 63733 5123 63767
rect 6745 63733 6779 63767
rect 9781 63733 9815 63767
rect 11345 63733 11379 63767
rect 11437 63733 11471 63767
rect 11713 63733 11747 63767
rect 13645 63733 13679 63767
rect 15577 63733 15611 63767
rect 17509 63733 17543 63767
rect 5641 63529 5675 63563
rect 6193 63529 6227 63563
rect 6653 63529 6687 63563
rect 11713 63529 11747 63563
rect 15577 63529 15611 63563
rect 16497 63529 16531 63563
rect 7941 63461 7975 63495
rect 11161 63461 11195 63495
rect 1501 63393 1535 63427
rect 4261 63393 4295 63427
rect 7481 63393 7515 63427
rect 7573 63393 7607 63427
rect 9229 63393 9263 63427
rect 9413 63393 9447 63427
rect 9781 63393 9815 63427
rect 10149 63393 10183 63427
rect 10701 63393 10735 63427
rect 12449 63393 12483 63427
rect 13553 63393 13587 63427
rect 16037 63393 16071 63427
rect 1777 63325 1811 63359
rect 4537 63325 4571 63359
rect 13829 63325 13863 63359
rect 3433 63257 3467 63291
rect 9229 63257 9263 63291
rect 2881 63189 2915 63223
rect 4077 63189 4111 63223
rect 8309 63189 8343 63223
rect 12633 63189 12667 63223
rect 13001 63189 13035 63223
rect 13369 63189 13403 63223
rect 14933 63189 14967 63223
rect 16221 63189 16255 63223
rect 3157 62985 3191 63019
rect 3893 62985 3927 63019
rect 4353 62985 4387 63019
rect 4997 62985 5031 63019
rect 8125 62985 8159 63019
rect 9965 62985 9999 63019
rect 11437 62985 11471 63019
rect 14749 62985 14783 63019
rect 15025 62985 15059 63019
rect 16957 62985 16991 63019
rect 8493 62917 8527 62951
rect 2053 62849 2087 62883
rect 9137 62849 9171 62883
rect 12633 62849 12667 62883
rect 15669 62849 15703 62883
rect 2329 62781 2363 62815
rect 2513 62781 2547 62815
rect 2789 62781 2823 62815
rect 4261 62781 4295 62815
rect 6193 62781 6227 62815
rect 6653 62781 6687 62815
rect 8585 62781 8619 62815
rect 10057 62781 10091 62815
rect 10241 62781 10275 62815
rect 10701 62781 10735 62815
rect 12725 62781 12759 62815
rect 13001 62781 13035 62815
rect 15393 62781 15427 62815
rect 1501 62713 1535 62747
rect 4077 62713 4111 62747
rect 7757 62713 7791 62747
rect 9413 62713 9447 62747
rect 5273 62645 5307 62679
rect 6561 62645 6595 62679
rect 7297 62645 7331 62679
rect 8769 62645 8803 62679
rect 12265 62645 12299 62679
rect 14105 62645 14139 62679
rect 2421 62441 2455 62475
rect 4629 62441 4663 62475
rect 8953 62441 8987 62475
rect 9689 62441 9723 62475
rect 10241 62441 10275 62475
rect 12633 62441 12667 62475
rect 2973 62373 3007 62407
rect 1593 62305 1627 62339
rect 1777 62305 1811 62339
rect 3801 62305 3835 62339
rect 8769 62305 8803 62339
rect 9781 62305 9815 62339
rect 11345 62305 11379 62339
rect 12449 62305 12483 62339
rect 12909 62305 12943 62339
rect 13737 62305 13771 62339
rect 2145 62237 2179 62271
rect 2789 62237 2823 62271
rect 3525 62237 3559 62271
rect 3985 62237 4019 62271
rect 11529 62237 11563 62271
rect 14013 62237 14047 62271
rect 15209 62237 15243 62271
rect 16037 62237 16071 62271
rect 4353 62169 4387 62203
rect 9321 62169 9355 62203
rect 9965 62101 9999 62135
rect 10701 62101 10735 62135
rect 13645 62101 13679 62135
rect 3065 61897 3099 61931
rect 3157 61897 3191 61931
rect 9413 61897 9447 61931
rect 11161 61897 11195 61931
rect 11805 61897 11839 61931
rect 14749 61897 14783 61931
rect 2053 61761 2087 61795
rect 2513 61761 2547 61795
rect 2329 61693 2363 61727
rect 1501 61625 1535 61659
rect 8861 61829 8895 61863
rect 12265 61829 12299 61863
rect 14289 61829 14323 61863
rect 4077 61761 4111 61795
rect 13553 61761 13587 61795
rect 15117 61761 15151 61795
rect 4353 61693 4387 61727
rect 9965 61693 9999 61727
rect 10149 61693 10183 61727
rect 10517 61693 10551 61727
rect 11529 61693 11563 61727
rect 12541 61693 12575 61727
rect 12725 61693 12759 61727
rect 13277 61693 13311 61727
rect 15301 61693 15335 61727
rect 15577 61693 15611 61727
rect 3709 61625 3743 61659
rect 3157 61557 3191 61591
rect 3433 61557 3467 61591
rect 5457 61557 5491 61591
rect 8493 61557 8527 61591
rect 9965 61557 9999 61591
rect 13921 61557 13955 61591
rect 16681 61557 16715 61591
rect 3065 61353 3099 61387
rect 4261 61353 4295 61387
rect 4813 61353 4847 61387
rect 9781 61353 9815 61387
rect 3525 61285 3559 61319
rect 1501 61217 1535 61251
rect 3985 61217 4019 61251
rect 4169 61217 4203 61251
rect 8309 61217 8343 61251
rect 8769 61217 8803 61251
rect 8953 61217 8987 61251
rect 10517 61217 10551 61251
rect 11069 61217 11103 61251
rect 13001 61217 13035 61251
rect 13185 61217 13219 61251
rect 14749 61217 14783 61251
rect 1777 61149 1811 61183
rect 3801 61149 3835 61183
rect 10885 61149 10919 61183
rect 13461 61149 13495 61183
rect 15025 61149 15059 61183
rect 8309 61013 8343 61047
rect 10149 61013 10183 61047
rect 11989 61013 12023 61047
rect 16129 61013 16163 61047
rect 3433 60809 3467 60843
rect 3801 60809 3835 60843
rect 9413 60809 9447 60843
rect 10149 60809 10183 60843
rect 11437 60809 11471 60843
rect 13737 60809 13771 60843
rect 10425 60741 10459 60775
rect 2145 60673 2179 60707
rect 12541 60673 12575 60707
rect 15485 60673 15519 60707
rect 16037 60673 16071 60707
rect 2697 60605 2731 60639
rect 2973 60605 3007 60639
rect 3157 60605 3191 60639
rect 4261 60605 4295 60639
rect 5273 60605 5307 60639
rect 8309 60605 8343 60639
rect 10609 60605 10643 60639
rect 10885 60605 10919 60639
rect 11897 60605 11931 60639
rect 12449 60605 12483 60639
rect 12725 60605 12759 60639
rect 16129 60605 16163 60639
rect 16405 60605 16439 60639
rect 2053 60537 2087 60571
rect 4077 60537 4111 60571
rect 4905 60537 4939 60571
rect 1685 60469 1719 60503
rect 4353 60469 4387 60503
rect 7849 60469 7883 60503
rect 8401 60469 8435 60503
rect 9045 60469 9079 60503
rect 11805 60469 11839 60503
rect 13461 60469 13495 60503
rect 14841 60469 14875 60503
rect 17509 60469 17543 60503
rect 2237 60265 2271 60299
rect 4629 60265 4663 60299
rect 7113 60265 7147 60299
rect 8033 60265 8067 60299
rect 10149 60265 10183 60299
rect 11989 60265 12023 60299
rect 14013 60265 14047 60299
rect 16129 60265 16163 60299
rect 3249 60129 3283 60163
rect 6101 60129 6135 60163
rect 6377 60129 6411 60163
rect 8769 60129 8803 60163
rect 10885 60129 10919 60163
rect 12725 60129 12759 60163
rect 12817 60129 12851 60163
rect 13185 60129 13219 60163
rect 2973 60061 3007 60095
rect 3525 60061 3559 60095
rect 9413 60061 9447 60095
rect 11529 60061 11563 60095
rect 13001 60061 13035 60095
rect 6193 59993 6227 60027
rect 1685 59925 1719 59959
rect 2605 59925 2639 59959
rect 8309 59925 8343 59959
rect 10609 59925 10643 59959
rect 3709 59721 3743 59755
rect 4905 59721 4939 59755
rect 5641 59721 5675 59755
rect 6285 59721 6319 59755
rect 6837 59721 6871 59755
rect 9413 59721 9447 59755
rect 12173 59721 12207 59755
rect 13461 59721 13495 59755
rect 14013 59721 14047 59755
rect 17509 59721 17543 59755
rect 1685 59653 1719 59687
rect 2329 59653 2363 59687
rect 11805 59653 11839 59687
rect 7113 59585 7147 59619
rect 10057 59585 10091 59619
rect 10793 59585 10827 59619
rect 14381 59585 14415 59619
rect 16037 59585 16071 59619
rect 2513 59517 2547 59551
rect 2881 59517 2915 59551
rect 4445 59517 4479 59551
rect 5089 59517 5123 59551
rect 5273 59517 5307 59551
rect 7297 59517 7331 59551
rect 7389 59517 7423 59551
rect 7757 59517 7791 59551
rect 10149 59517 10183 59551
rect 10701 59517 10735 59551
rect 10885 59517 10919 59551
rect 12541 59517 12575 59551
rect 12725 59517 12759 59551
rect 13001 59517 13035 59551
rect 13553 59517 13587 59551
rect 16129 59517 16163 59551
rect 16405 59517 16439 59551
rect 9045 59449 9079 59483
rect 2145 59381 2179 59415
rect 3341 59381 3375 59415
rect 4813 59381 4847 59415
rect 8677 59381 8711 59415
rect 3525 59177 3559 59211
rect 3893 59177 3927 59211
rect 10333 59177 10367 59211
rect 10885 59177 10919 59211
rect 11437 59177 11471 59211
rect 12265 59177 12299 59211
rect 13185 59177 13219 59211
rect 1593 59109 1627 59143
rect 11897 59109 11931 59143
rect 1501 59041 1535 59075
rect 2329 59041 2363 59075
rect 3341 59041 3375 59075
rect 5365 59041 5399 59075
rect 5733 59041 5767 59075
rect 5825 59041 5859 59075
rect 7481 59041 7515 59075
rect 7941 59041 7975 59075
rect 8493 59041 8527 59075
rect 9045 59041 9079 59075
rect 9229 59041 9263 59075
rect 9781 59041 9815 59075
rect 11253 59041 11287 59075
rect 13369 59041 13403 59075
rect 2421 58973 2455 59007
rect 4813 58973 4847 59007
rect 8677 58973 8711 59007
rect 13461 58973 13495 59007
rect 13737 58973 13771 59007
rect 14841 58973 14875 59007
rect 2881 58905 2915 58939
rect 3249 58905 3283 58939
rect 5181 58905 5215 58939
rect 6193 58905 6227 58939
rect 6653 58837 6687 58871
rect 7113 58837 7147 58871
rect 7665 58837 7699 58871
rect 8309 58837 8343 58871
rect 12817 58837 12851 58871
rect 16129 58837 16163 58871
rect 2881 58633 2915 58667
rect 4629 58633 4663 58667
rect 4997 58633 5031 58667
rect 7665 58633 7699 58667
rect 14657 58633 14691 58667
rect 5549 58565 5583 58599
rect 7297 58565 7331 58599
rect 10425 58565 10459 58599
rect 1501 58497 1535 58531
rect 1777 58497 1811 58531
rect 8677 58497 8711 58531
rect 11805 58497 11839 58531
rect 12725 58497 12759 58531
rect 3525 58429 3559 58463
rect 4077 58429 4111 58463
rect 5733 58429 5767 58463
rect 6009 58429 6043 58463
rect 6377 58429 6411 58463
rect 6653 58429 6687 58463
rect 8217 58429 8251 58463
rect 8585 58429 8619 58463
rect 9689 58429 9723 58463
rect 10149 58429 10183 58463
rect 10517 58429 10551 58463
rect 12449 58429 12483 58463
rect 13001 58429 13035 58463
rect 3893 58361 3927 58395
rect 7757 58361 7791 58395
rect 4261 58293 4295 58327
rect 5365 58293 5399 58327
rect 9137 58293 9171 58327
rect 9505 58293 9539 58327
rect 11345 58293 11379 58327
rect 12081 58293 12115 58327
rect 12265 58293 12299 58327
rect 14105 58293 14139 58327
rect 5549 58089 5583 58123
rect 6469 58089 6503 58123
rect 11161 58089 11195 58123
rect 15945 58089 15979 58123
rect 1593 58021 1627 58055
rect 3985 58021 4019 58055
rect 6837 58021 6871 58055
rect 8861 58021 8895 58055
rect 2329 57953 2363 57987
rect 4813 57953 4847 57987
rect 6653 57953 6687 57987
rect 7481 57953 7515 57987
rect 7849 57953 7883 57987
rect 9689 57953 9723 57987
rect 11069 57953 11103 57987
rect 12541 57953 12575 57987
rect 12817 57953 12851 57987
rect 13185 57953 13219 57987
rect 1501 57885 1535 57919
rect 2421 57885 2455 57919
rect 2881 57885 2915 57919
rect 3893 57885 3927 57919
rect 4537 57885 4571 57919
rect 4997 57885 5031 57919
rect 7297 57885 7331 57919
rect 7757 57885 7791 57919
rect 9413 57885 9447 57919
rect 9873 57885 9907 57919
rect 11713 57885 11747 57919
rect 13553 57885 13587 57919
rect 14289 57885 14323 57919
rect 5917 57817 5951 57851
rect 3157 57749 3191 57783
rect 6285 57749 6319 57783
rect 8585 57749 8619 57783
rect 10149 57749 10183 57783
rect 10609 57749 10643 57783
rect 14013 57749 14047 57783
rect 4997 57545 5031 57579
rect 8953 57545 8987 57579
rect 10609 57545 10643 57579
rect 12725 57545 12759 57579
rect 2145 57409 2179 57443
rect 3157 57409 3191 57443
rect 4261 57409 4295 57443
rect 5365 57409 5399 57443
rect 6469 57409 6503 57443
rect 11805 57409 11839 57443
rect 15853 57409 15887 57443
rect 2697 57341 2731 57375
rect 2973 57341 3007 57375
rect 6377 57341 6411 57375
rect 7205 57341 7239 57375
rect 7389 57341 7423 57375
rect 10149 57341 10183 57375
rect 11069 57341 11103 57375
rect 11437 57341 11471 57375
rect 11713 57341 11747 57375
rect 12173 57341 12207 57375
rect 15945 57341 15979 57375
rect 16221 57341 16255 57375
rect 5641 57273 5675 57307
rect 13001 57273 13035 57307
rect 1685 57205 1719 57239
rect 2053 57205 2087 57239
rect 3525 57205 3559 57239
rect 3893 57205 3927 57239
rect 6745 57205 6779 57239
rect 7941 57205 7975 57239
rect 8401 57205 8435 57239
rect 9229 57205 9263 57239
rect 9965 57205 9999 57239
rect 10333 57205 10367 57239
rect 13461 57205 13495 57239
rect 17325 57205 17359 57239
rect 4077 57001 4111 57035
rect 5641 57001 5675 57035
rect 6193 57001 6227 57035
rect 9045 57001 9079 57035
rect 11529 57001 11563 57035
rect 12173 57001 12207 57035
rect 8217 56933 8251 56967
rect 1869 56865 1903 56899
rect 4537 56865 4571 56899
rect 7205 56865 7239 56899
rect 7665 56865 7699 56899
rect 1593 56797 1627 56831
rect 4261 56797 4295 56831
rect 6929 56797 6963 56831
rect 7665 56729 7699 56763
rect 12449 56933 12483 56967
rect 9229 56865 9263 56899
rect 9597 56865 9631 56899
rect 10241 56865 10275 56899
rect 10701 56865 10735 56899
rect 11713 56865 11747 56899
rect 13001 56865 13035 56899
rect 9321 56797 9355 56831
rect 15301 56797 15335 56831
rect 15577 56797 15611 56831
rect 2973 56661 3007 56695
rect 3617 56661 3651 56695
rect 6653 56661 6687 56695
rect 8861 56661 8895 56695
rect 9045 56661 9079 56695
rect 11253 56661 11287 56695
rect 13461 56661 13495 56695
rect 13921 56661 13955 56695
rect 16681 56661 16715 56695
rect 1593 56457 1627 56491
rect 2329 56457 2363 56491
rect 3893 56457 3927 56491
rect 5641 56457 5675 56491
rect 7941 56457 7975 56491
rect 8493 56457 8527 56491
rect 11897 56457 11931 56491
rect 7389 56389 7423 56423
rect 9965 56389 9999 56423
rect 11621 56389 11655 56423
rect 10241 56321 10275 56355
rect 16037 56321 16071 56355
rect 2513 56253 2547 56287
rect 2881 56253 2915 56287
rect 4077 56253 4111 56287
rect 4353 56253 4387 56287
rect 6561 56253 6595 56287
rect 7021 56253 7055 56287
rect 7389 56253 7423 56287
rect 8585 56253 8619 56287
rect 11069 56253 11103 56287
rect 11161 56253 11195 56287
rect 12541 56253 12575 56287
rect 16129 56253 16163 56287
rect 16405 56253 16439 56287
rect 2145 56185 2179 56219
rect 10333 56185 10367 56219
rect 13553 56185 13587 56219
rect 13829 56185 13863 56219
rect 3525 56117 3559 56151
rect 6101 56117 6135 56151
rect 6469 56117 6503 56151
rect 8769 56117 8803 56151
rect 9321 56117 9355 56151
rect 12541 56117 12575 56151
rect 13093 56117 13127 56151
rect 14197 56117 14231 56151
rect 14657 56117 14691 56151
rect 15025 56117 15059 56151
rect 15577 56117 15611 56151
rect 17509 56117 17543 56151
rect 1685 55913 1719 55947
rect 2329 55913 2363 55947
rect 4537 55913 4571 55947
rect 6469 55913 6503 55947
rect 8309 55913 8343 55947
rect 8861 55913 8895 55947
rect 9413 55913 9447 55947
rect 11529 55913 11563 55947
rect 12081 55913 12115 55947
rect 12817 55913 12851 55947
rect 13001 55913 13035 55947
rect 3709 55845 3743 55879
rect 7941 55845 7975 55879
rect 9321 55845 9355 55879
rect 4813 55777 4847 55811
rect 4997 55777 5031 55811
rect 5181 55777 5215 55811
rect 6653 55777 6687 55811
rect 7205 55777 7239 55811
rect 7665 55777 7699 55811
rect 9597 55777 9631 55811
rect 9781 55777 9815 55811
rect 10057 55777 10091 55811
rect 10425 55777 10459 55811
rect 12265 55777 12299 55811
rect 12449 55777 12483 55811
rect 6929 55709 6963 55743
rect 10609 55709 10643 55743
rect 11253 55709 11287 55743
rect 13461 55845 13495 55879
rect 15577 55777 15611 55811
rect 16957 55777 16991 55811
rect 13645 55709 13679 55743
rect 13921 55709 13955 55743
rect 16129 55709 16163 55743
rect 16681 55709 16715 55743
rect 17141 55709 17175 55743
rect 12817 55641 12851 55675
rect 16037 55641 16071 55675
rect 4169 55573 4203 55607
rect 5733 55573 5767 55607
rect 6101 55573 6135 55607
rect 11897 55573 11931 55607
rect 12633 55573 12667 55607
rect 15209 55573 15243 55607
rect 1685 55369 1719 55403
rect 3433 55369 3467 55403
rect 3801 55369 3835 55403
rect 5365 55369 5399 55403
rect 9045 55369 9079 55403
rect 9413 55369 9447 55403
rect 10517 55369 10551 55403
rect 17233 55369 17267 55403
rect 6285 55301 6319 55335
rect 8769 55301 8803 55335
rect 13277 55301 13311 55335
rect 4813 55233 4847 55267
rect 5641 55233 5675 55267
rect 6929 55233 6963 55267
rect 7941 55233 7975 55267
rect 11529 55233 11563 55267
rect 13921 55233 13955 55267
rect 15117 55233 15151 55267
rect 17601 55233 17635 55267
rect 2973 55165 3007 55199
rect 4261 55165 4295 55199
rect 6009 55165 6043 55199
rect 6285 55165 6319 55199
rect 8217 55165 8251 55199
rect 8401 55165 8435 55199
rect 9689 55165 9723 55199
rect 10149 55165 10183 55199
rect 11069 55165 11103 55199
rect 11805 55165 11839 55199
rect 11897 55165 11931 55199
rect 12265 55165 12299 55199
rect 14197 55165 14231 55199
rect 14381 55165 14415 55199
rect 15301 55165 15335 55199
rect 15577 55165 15611 55199
rect 7389 55097 7423 55131
rect 10977 55097 11011 55131
rect 13369 55097 13403 55131
rect 3157 55029 3191 55063
rect 4445 55029 4479 55063
rect 7297 55029 7331 55063
rect 9873 55029 9907 55063
rect 12817 55029 12851 55063
rect 14749 55029 14783 55063
rect 16681 55029 16715 55063
rect 4721 54825 4755 54859
rect 11805 54825 11839 54859
rect 13185 54825 13219 54859
rect 2421 54689 2455 54723
rect 2881 54689 2915 54723
rect 5549 54689 5583 54723
rect 7205 54689 7239 54723
rect 7941 54689 7975 54723
rect 8861 54689 8895 54723
rect 9229 54689 9263 54723
rect 9873 54689 9907 54723
rect 10977 54689 11011 54723
rect 13277 54689 13311 54723
rect 16589 54689 16623 54723
rect 16865 54689 16899 54723
rect 7297 54621 7331 54655
rect 9505 54621 9539 54655
rect 10885 54621 10919 54655
rect 11437 54621 11471 54655
rect 13553 54621 13587 54655
rect 16129 54621 16163 54655
rect 1685 54553 1719 54587
rect 2329 54553 2363 54587
rect 5089 54553 5123 54587
rect 12173 54553 12207 54587
rect 15393 54553 15427 54587
rect 16957 54553 16991 54587
rect 1961 54485 1995 54519
rect 4261 54485 4295 54519
rect 5641 54485 5675 54519
rect 6285 54485 6319 54519
rect 6653 54485 6687 54519
rect 8309 54485 8343 54519
rect 8769 54485 8803 54519
rect 10517 54485 10551 54519
rect 12633 54485 12667 54519
rect 14657 54485 14691 54519
rect 15761 54485 15795 54519
rect 2881 54281 2915 54315
rect 5365 54281 5399 54315
rect 5733 54281 5767 54315
rect 9413 54281 9447 54315
rect 11437 54281 11471 54315
rect 17785 54281 17819 54315
rect 6837 54213 6871 54247
rect 10517 54213 10551 54247
rect 1593 54145 1627 54179
rect 2421 54145 2455 54179
rect 9873 54145 9907 54179
rect 12541 54145 12575 54179
rect 14013 54145 14047 54179
rect 15853 54145 15887 54179
rect 1501 54077 1535 54111
rect 2329 54077 2363 54111
rect 3893 54077 3927 54111
rect 4261 54077 4295 54111
rect 6101 54077 6135 54111
rect 6377 54077 6411 54111
rect 6653 54077 6687 54111
rect 7113 54077 7147 54111
rect 7941 54077 7975 54111
rect 8125 54077 8159 54111
rect 8493 54077 8527 54111
rect 9137 54077 9171 54111
rect 10057 54077 10091 54111
rect 10517 54077 10551 54111
rect 11805 54077 11839 54111
rect 12081 54077 12115 54111
rect 12633 54077 12667 54111
rect 12909 54077 12943 54111
rect 14105 54077 14139 54111
rect 14565 54077 14599 54111
rect 15301 54077 15335 54111
rect 15945 54077 15979 54111
rect 16313 54077 16347 54111
rect 16681 54077 16715 54111
rect 4077 54009 4111 54043
rect 4905 54009 4939 54043
rect 7573 54009 7607 54043
rect 4353 53941 4387 53975
rect 6193 53941 6227 53975
rect 8585 53941 8619 53975
rect 11161 53941 11195 53975
rect 11621 53941 11655 53975
rect 13645 53941 13679 53975
rect 14289 53941 14323 53975
rect 15117 53941 15151 53975
rect 17049 53941 17083 53975
rect 17417 53941 17451 53975
rect 1685 53737 1719 53771
rect 5641 53737 5675 53771
rect 9781 53737 9815 53771
rect 12081 53737 12115 53771
rect 14013 53737 14047 53771
rect 4721 53669 4755 53703
rect 6009 53669 6043 53703
rect 3433 53601 3467 53635
rect 3709 53601 3743 53635
rect 4905 53601 4939 53635
rect 6285 53601 6319 53635
rect 7021 53601 7055 53635
rect 8217 53601 8251 53635
rect 8677 53601 8711 53635
rect 8861 53601 8895 53635
rect 9505 53601 9539 53635
rect 10609 53601 10643 53635
rect 10793 53601 10827 53635
rect 11345 53601 11379 53635
rect 12541 53601 12575 53635
rect 12817 53601 12851 53635
rect 13185 53601 13219 53635
rect 15301 53601 15335 53635
rect 15945 53601 15979 53635
rect 16221 53601 16255 53635
rect 16589 53601 16623 53635
rect 2881 53533 2915 53567
rect 3893 53533 3927 53567
rect 9413 53533 9447 53567
rect 10149 53533 10183 53567
rect 11529 53533 11563 53567
rect 12909 53533 12943 53567
rect 4353 53465 4387 53499
rect 14749 53465 14783 53499
rect 15117 53465 15151 53499
rect 2329 53397 2363 53431
rect 2789 53397 2823 53431
rect 4997 53397 5031 53431
rect 6101 53397 6135 53431
rect 6653 53397 6687 53431
rect 7205 53397 7239 53431
rect 7757 53397 7791 53431
rect 14473 53397 14507 53431
rect 16497 53397 16531 53431
rect 17049 53397 17083 53431
rect 2881 53193 2915 53227
rect 3893 53193 3927 53227
rect 5641 53193 5675 53227
rect 6653 53193 6687 53227
rect 8585 53193 8619 53227
rect 8861 53193 8895 53227
rect 9965 53193 9999 53227
rect 6929 53125 6963 53159
rect 8217 53125 8251 53159
rect 11529 53125 11563 53159
rect 13921 53125 13955 53159
rect 1777 53057 1811 53091
rect 7573 53057 7607 53091
rect 9505 53057 9539 53091
rect 10241 53057 10275 53091
rect 13185 53057 13219 53091
rect 15485 53057 15519 53091
rect 17141 53057 17175 53091
rect 1501 52989 1535 53023
rect 4261 52989 4295 53023
rect 4537 52989 4571 53023
rect 6745 52989 6779 53023
rect 7297 52989 7331 53023
rect 10609 52989 10643 53023
rect 10885 52989 10919 53023
rect 11989 52989 12023 53023
rect 12633 52989 12667 53023
rect 12725 52989 12759 53023
rect 14013 52989 14047 53023
rect 14473 52989 14507 53023
rect 15577 52989 15611 53023
rect 15945 52989 15979 53023
rect 16129 52989 16163 53023
rect 16681 52989 16715 53023
rect 17969 52989 18003 53023
rect 11161 52921 11195 52955
rect 15117 52921 15151 52955
rect 3525 52853 3559 52887
rect 6193 52853 6227 52887
rect 11897 52853 11931 52887
rect 13461 52853 13495 52887
rect 14197 52853 14231 52887
rect 17509 52853 17543 52887
rect 2973 52649 3007 52683
rect 4721 52649 4755 52683
rect 5181 52649 5215 52683
rect 5825 52649 5859 52683
rect 7757 52649 7791 52683
rect 9137 52649 9171 52683
rect 9505 52649 9539 52683
rect 16221 52649 16255 52683
rect 1685 52581 1719 52615
rect 5457 52581 5491 52615
rect 3157 52513 3191 52547
rect 5641 52513 5675 52547
rect 7389 52513 7423 52547
rect 8125 52513 8159 52547
rect 8493 52513 8527 52547
rect 10333 52513 10367 52547
rect 10793 52513 10827 52547
rect 11069 52513 11103 52547
rect 13001 52513 13035 52547
rect 13369 52513 13403 52547
rect 14657 52513 14691 52547
rect 15025 52513 15059 52547
rect 15209 52513 15243 52547
rect 15669 52513 15703 52547
rect 16957 52513 16991 52547
rect 3433 52445 3467 52479
rect 6653 52445 6687 52479
rect 7481 52445 7515 52479
rect 10149 52445 10183 52479
rect 12633 52445 12667 52479
rect 10425 52377 10459 52411
rect 11989 52377 12023 52411
rect 13369 52377 13403 52411
rect 14197 52377 14231 52411
rect 17141 52377 17175 52411
rect 2053 52309 2087 52343
rect 6101 52309 6135 52343
rect 9873 52309 9907 52343
rect 13921 52309 13955 52343
rect 14473 52309 14507 52343
rect 16497 52309 16531 52343
rect 3893 52105 3927 52139
rect 5457 52105 5491 52139
rect 8401 52105 8435 52139
rect 10057 52105 10091 52139
rect 14749 52105 14783 52139
rect 17601 52105 17635 52139
rect 17969 52105 18003 52139
rect 3525 52037 3559 52071
rect 7021 52037 7055 52071
rect 7665 52037 7699 52071
rect 13277 52037 13311 52071
rect 4077 51969 4111 52003
rect 4629 51969 4663 52003
rect 5089 51969 5123 52003
rect 6009 51969 6043 52003
rect 9505 51969 9539 52003
rect 12909 51969 12943 52003
rect 14381 51969 14415 52003
rect 17233 51969 17267 52003
rect 4905 51901 4939 51935
rect 6101 51901 6135 51935
rect 6561 51901 6595 51935
rect 6653 51901 6687 51935
rect 8585 51901 8619 51935
rect 9045 51901 9079 51935
rect 10701 51901 10735 51935
rect 11069 51901 11103 51935
rect 11437 51901 11471 51935
rect 12081 51901 12115 51935
rect 12541 51901 12575 51935
rect 13921 51901 13955 51935
rect 14197 51901 14231 51935
rect 15485 51901 15519 51935
rect 15853 51901 15887 51935
rect 16221 51901 16255 51935
rect 16773 51901 16807 51935
rect 10609 51833 10643 51867
rect 13369 51833 13403 51867
rect 15117 51833 15151 51867
rect 16681 51833 16715 51867
rect 2789 51765 2823 51799
rect 3157 51765 3191 51799
rect 5825 51765 5859 51799
rect 8033 51765 8067 51799
rect 8769 51765 8803 51799
rect 10425 51765 10459 51799
rect 1685 51561 1719 51595
rect 3157 51561 3191 51595
rect 4629 51561 4663 51595
rect 5917 51561 5951 51595
rect 6193 51561 6227 51595
rect 7113 51561 7147 51595
rect 10701 51561 10735 51595
rect 11069 51561 11103 51595
rect 12817 51561 12851 51595
rect 14933 51561 14967 51595
rect 17141 51561 17175 51595
rect 17509 51561 17543 51595
rect 5181 51425 5215 51459
rect 5549 51425 5583 51459
rect 4813 51357 4847 51391
rect 5641 51289 5675 51323
rect 7297 51493 7331 51527
rect 7665 51493 7699 51527
rect 8401 51493 8435 51527
rect 10241 51493 10275 51527
rect 11161 51493 11195 51527
rect 12173 51493 12207 51527
rect 14565 51493 14599 51527
rect 7205 51425 7239 51459
rect 7941 51425 7975 51459
rect 8953 51425 8987 51459
rect 9229 51425 9263 51459
rect 9321 51425 9355 51459
rect 9965 51425 9999 51459
rect 10977 51425 11011 51459
rect 15577 51425 15611 51459
rect 16037 51425 16071 51459
rect 16221 51425 16255 51459
rect 16773 51425 16807 51459
rect 6929 51357 6963 51391
rect 8493 51357 8527 51391
rect 9597 51357 9631 51391
rect 10793 51357 10827 51391
rect 11529 51357 11563 51391
rect 11805 51357 11839 51391
rect 12909 51357 12943 51391
rect 13185 51357 13219 51391
rect 15301 51357 15335 51391
rect 4077 51221 4111 51255
rect 5917 51221 5951 51255
rect 6653 51221 6687 51255
rect 15485 51221 15519 51255
rect 3065 51017 3099 51051
rect 3893 51017 3927 51051
rect 4997 51017 5031 51051
rect 5457 51017 5491 51051
rect 3525 50881 3559 50915
rect 1501 50813 1535 50847
rect 1777 50813 1811 50847
rect 4077 50813 4111 50847
rect 4537 50813 4571 50847
rect 5365 50813 5399 50847
rect 5457 50745 5491 50779
rect 6193 51017 6227 51051
rect 6745 51017 6779 51051
rect 8769 51017 8803 51051
rect 9321 51017 9355 51051
rect 10057 51017 10091 51051
rect 12449 51017 12483 51051
rect 13185 51017 13219 51051
rect 7757 50813 7791 50847
rect 7849 50813 7883 50847
rect 8125 50813 8159 50847
rect 8309 50813 8343 50847
rect 8493 50813 8527 50847
rect 8769 50813 8803 50847
rect 10517 50813 10551 50847
rect 10977 50813 11011 50847
rect 11253 50813 11287 50847
rect 11529 50813 11563 50847
rect 12725 50813 12759 50847
rect 11989 50745 12023 50779
rect 14473 51017 14507 51051
rect 14749 51017 14783 51051
rect 14381 50881 14415 50915
rect 17509 50949 17543 50983
rect 15853 50881 15887 50915
rect 13921 50813 13955 50847
rect 14197 50813 14231 50847
rect 14473 50813 14507 50847
rect 15301 50813 15335 50847
rect 16129 50813 16163 50847
rect 16681 50813 16715 50847
rect 17141 50813 17175 50847
rect 17509 50813 17543 50847
rect 13369 50745 13403 50779
rect 4261 50677 4295 50711
rect 5181 50677 5215 50711
rect 5641 50677 5675 50711
rect 6193 50677 6227 50711
rect 6377 50677 6411 50711
rect 7021 50677 7055 50711
rect 7297 50677 7331 50711
rect 8953 50677 8987 50711
rect 10333 50677 10367 50711
rect 12541 50677 12575 50711
rect 13093 50677 13127 50711
rect 13185 50677 13219 50711
rect 15025 50677 15059 50711
rect 15485 50677 15519 50711
rect 16589 50677 16623 50711
rect 18061 50677 18095 50711
rect 4721 50473 4755 50507
rect 5089 50473 5123 50507
rect 5549 50473 5583 50507
rect 6653 50473 6687 50507
rect 7481 50473 7515 50507
rect 8401 50473 8435 50507
rect 10793 50473 10827 50507
rect 11805 50473 11839 50507
rect 13001 50473 13035 50507
rect 15485 50473 15519 50507
rect 17325 50473 17359 50507
rect 3341 50405 3375 50439
rect 5917 50405 5951 50439
rect 7849 50405 7883 50439
rect 11161 50405 11195 50439
rect 4077 50337 4111 50371
rect 4169 50337 4203 50371
rect 8309 50337 8343 50371
rect 8585 50337 8619 50371
rect 9045 50337 9079 50371
rect 9229 50337 9263 50371
rect 9413 50337 9447 50371
rect 9689 50337 9723 50371
rect 11345 50337 11379 50371
rect 12265 50337 12299 50371
rect 13369 50337 13403 50371
rect 15117 50337 15151 50371
rect 15577 50337 15611 50371
rect 15945 50337 15979 50371
rect 16313 50337 16347 50371
rect 16865 50337 16899 50371
rect 3249 50269 3283 50303
rect 8677 50269 8711 50303
rect 13093 50269 13127 50303
rect 15853 50269 15887 50303
rect 7113 50201 7147 50235
rect 11529 50201 11563 50235
rect 1685 50133 1719 50167
rect 6285 50133 6319 50167
rect 10057 50133 10091 50167
rect 10517 50133 10551 50167
rect 14473 50133 14507 50167
rect 2237 49929 2271 49963
rect 3525 49929 3559 49963
rect 4905 49929 4939 49963
rect 9229 49929 9263 49963
rect 6101 49861 6135 49895
rect 7113 49861 7147 49895
rect 2789 49793 2823 49827
rect 3801 49793 3835 49827
rect 2513 49725 2547 49759
rect 2973 49725 3007 49759
rect 4537 49725 4571 49759
rect 4997 49725 5031 49759
rect 5181 49725 5215 49759
rect 5641 49725 5675 49759
rect 5733 49725 5767 49759
rect 7205 49725 7239 49759
rect 7757 49725 7791 49759
rect 7849 49725 7883 49759
rect 8033 49725 8067 49759
rect 8217 49725 8251 49759
rect 8493 49725 8527 49759
rect 9045 49725 9079 49759
rect 9505 49929 9539 49963
rect 11897 49929 11931 49963
rect 12449 49929 12483 49963
rect 13185 49929 13219 49963
rect 13553 49929 13587 49963
rect 13645 49929 13679 49963
rect 14933 49929 14967 49963
rect 14657 49861 14691 49895
rect 10149 49793 10183 49827
rect 9689 49725 9723 49759
rect 10333 49725 10367 49759
rect 10609 49725 10643 49759
rect 10977 49725 11011 49759
rect 11529 49725 11563 49759
rect 12081 49725 12115 49759
rect 12173 49725 12207 49759
rect 12265 49725 12299 49759
rect 13829 49725 13863 49759
rect 13921 49725 13955 49759
rect 14381 49657 14415 49691
rect 6745 49589 6779 49623
rect 9229 49589 9263 49623
rect 9321 49589 9355 49623
rect 9505 49589 9539 49623
rect 16221 49861 16255 49895
rect 17601 49793 17635 49827
rect 15301 49725 15335 49759
rect 15761 49725 15795 49759
rect 16681 49725 16715 49759
rect 17233 49725 17267 49759
rect 17509 49725 17543 49759
rect 14933 49589 14967 49623
rect 15025 49589 15059 49623
rect 15485 49589 15519 49623
rect 16589 49589 16623 49623
rect 2513 49385 2547 49419
rect 4537 49385 4571 49419
rect 6285 49385 6319 49419
rect 6653 49385 6687 49419
rect 8769 49385 8803 49419
rect 9505 49385 9539 49419
rect 10425 49385 10459 49419
rect 11161 49385 11195 49419
rect 12081 49385 12115 49419
rect 14105 49385 14139 49419
rect 15945 49385 15979 49419
rect 17509 49385 17543 49419
rect 5917 49317 5951 49351
rect 8401 49317 8435 49351
rect 10517 49317 10551 49351
rect 10885 49317 10919 49351
rect 12633 49317 12667 49351
rect 14381 49317 14415 49351
rect 14749 49317 14783 49351
rect 15301 49317 15335 49351
rect 15669 49317 15703 49351
rect 3065 49249 3099 49283
rect 3433 49249 3467 49283
rect 6837 49249 6871 49283
rect 7481 49249 7515 49283
rect 7849 49249 7883 49283
rect 8861 49249 8895 49283
rect 10333 49249 10367 49283
rect 12449 49249 12483 49283
rect 12725 49249 12759 49283
rect 14841 49249 14875 49283
rect 16957 49249 16991 49283
rect 17141 49249 17175 49283
rect 3157 49181 3191 49215
rect 7573 49181 7607 49215
rect 7941 49181 7975 49215
rect 10149 49181 10183 49215
rect 16129 49181 16163 49215
rect 16681 49181 16715 49215
rect 5549 49113 5583 49147
rect 1593 49045 1627 49079
rect 5181 49045 5215 49079
rect 9045 49045 9079 49079
rect 9873 49045 9907 49079
rect 11621 49045 11655 49079
rect 12909 49045 12943 49079
rect 13645 49045 13679 49079
rect 14565 49045 14599 49079
rect 3065 48841 3099 48875
rect 3525 48841 3559 48875
rect 4905 48841 4939 48875
rect 8217 48841 8251 48875
rect 11529 48841 11563 48875
rect 12265 48841 12299 48875
rect 14289 48841 14323 48875
rect 15025 48841 15059 48875
rect 15485 48841 15519 48875
rect 13277 48773 13311 48807
rect 1501 48705 1535 48739
rect 6745 48705 6779 48739
rect 7481 48705 7515 48739
rect 10609 48705 10643 48739
rect 17325 48705 17359 48739
rect 17785 48705 17819 48739
rect 1777 48637 1811 48671
rect 4905 48637 4939 48671
rect 5365 48637 5399 48671
rect 6285 48637 6319 48671
rect 6653 48637 6687 48671
rect 7389 48637 7423 48671
rect 7757 48637 7791 48671
rect 7849 48637 7883 48671
rect 9505 48637 9539 48671
rect 9873 48637 9907 48671
rect 10149 48637 10183 48671
rect 10793 48637 10827 48671
rect 11253 48637 11287 48671
rect 11897 48637 11931 48671
rect 12081 48637 12115 48671
rect 12909 48637 12943 48671
rect 15301 48637 15335 48671
rect 15761 48637 15795 48671
rect 17601 48637 17635 48671
rect 4721 48569 4755 48603
rect 12541 48569 12575 48603
rect 16221 48569 16255 48603
rect 16773 48569 16807 48603
rect 3801 48501 3835 48535
rect 5917 48501 5951 48535
rect 8953 48501 8987 48535
rect 13829 48501 13863 48535
rect 14657 48501 14691 48535
rect 16589 48501 16623 48535
rect 6285 48297 6319 48331
rect 9137 48297 9171 48331
rect 12725 48297 12759 48331
rect 17417 48297 17451 48331
rect 6653 48229 6687 48263
rect 7205 48229 7239 48263
rect 9781 48229 9815 48263
rect 11713 48229 11747 48263
rect 12081 48229 12115 48263
rect 15853 48229 15887 48263
rect 16405 48229 16439 48263
rect 16773 48229 16807 48263
rect 17141 48229 17175 48263
rect 5825 48161 5859 48195
rect 5917 48093 5951 48127
rect 7021 48093 7055 48127
rect 7389 48161 7423 48195
rect 8033 48161 8067 48195
rect 9229 48161 9263 48195
rect 10425 48161 10459 48195
rect 10517 48161 10551 48195
rect 10650 48161 10684 48195
rect 15945 48161 15979 48195
rect 8125 48093 8159 48127
rect 13001 48093 13035 48127
rect 13277 48093 13311 48127
rect 7481 48025 7515 48059
rect 1593 47957 1627 47991
rect 4905 47957 4939 47991
rect 7205 47957 7239 47991
rect 8677 47957 8711 47991
rect 9413 47957 9447 47991
rect 10149 47957 10183 47991
rect 10793 47957 10827 47991
rect 14381 47957 14415 47991
rect 15669 47957 15703 47991
rect 2881 47753 2915 47787
rect 4353 47753 4387 47787
rect 6745 47753 6779 47787
rect 8493 47753 8527 47787
rect 9137 47753 9171 47787
rect 9413 47753 9447 47787
rect 11069 47753 11103 47787
rect 13185 47753 13219 47787
rect 16681 47753 16715 47787
rect 4721 47685 4755 47719
rect 1777 47617 1811 47651
rect 15117 47617 15151 47651
rect 1501 47549 1535 47583
rect 5733 47549 5767 47583
rect 5917 47549 5951 47583
rect 6285 47549 6319 47583
rect 6929 47549 6963 47583
rect 8309 47549 8343 47583
rect 9689 47549 9723 47583
rect 10241 47549 10275 47583
rect 11805 47549 11839 47583
rect 11989 47549 12023 47583
rect 12357 47549 12391 47583
rect 15669 47549 15703 47583
rect 15853 47549 15887 47583
rect 15945 47549 15979 47583
rect 11529 47481 11563 47515
rect 12725 47481 12759 47515
rect 16405 47481 16439 47515
rect 5089 47413 5123 47447
rect 5457 47413 5491 47447
rect 7297 47413 7331 47447
rect 7757 47413 7791 47447
rect 9781 47413 9815 47447
rect 10701 47413 10735 47447
rect 13461 47413 13495 47447
rect 13829 47413 13863 47447
rect 15485 47413 15519 47447
rect 6285 47209 6319 47243
rect 7389 47209 7423 47243
rect 12817 47209 12851 47243
rect 14381 47209 14415 47243
rect 16405 47209 16439 47243
rect 4721 47141 4755 47175
rect 10333 47141 10367 47175
rect 16037 47141 16071 47175
rect 3525 47073 3559 47107
rect 3709 47073 3743 47107
rect 5181 47073 5215 47107
rect 5641 47073 5675 47107
rect 8033 47073 8067 47107
rect 8585 47073 8619 47107
rect 8769 47073 8803 47107
rect 9321 47073 9355 47107
rect 10977 47073 11011 47107
rect 16957 47073 16991 47107
rect 1685 47005 1719 47039
rect 3985 47005 4019 47039
rect 4997 47005 5031 47039
rect 8309 47005 8343 47039
rect 9781 47005 9815 47039
rect 12173 47005 12207 47039
rect 13001 47005 13035 47039
rect 13277 47005 13311 47039
rect 2053 46937 2087 46971
rect 5641 46937 5675 46971
rect 10241 46937 10275 46971
rect 11621 46937 11655 46971
rect 15669 46937 15703 46971
rect 17141 46937 17175 46971
rect 3525 46665 3559 46699
rect 4261 46665 4295 46699
rect 5641 46665 5675 46699
rect 7757 46665 7791 46699
rect 8493 46665 8527 46699
rect 9873 46665 9907 46699
rect 10609 46665 10643 46699
rect 11621 46665 11655 46699
rect 12633 46665 12667 46699
rect 17233 46665 17267 46699
rect 4629 46597 4663 46631
rect 1501 46529 1535 46563
rect 3157 46529 3191 46563
rect 5089 46529 5123 46563
rect 12725 46529 12759 46563
rect 14105 46529 14139 46563
rect 1777 46461 1811 46495
rect 5641 46461 5675 46495
rect 5917 46461 5951 46495
rect 6285 46461 6319 46495
rect 6929 46461 6963 46495
rect 9689 46461 9723 46495
rect 10149 46461 10183 46495
rect 11437 46461 11471 46495
rect 11897 46461 11931 46495
rect 13001 46461 13035 46495
rect 16037 46461 16071 46495
rect 17049 46461 17083 46495
rect 17509 46461 17543 46495
rect 8125 46393 8159 46427
rect 16589 46393 16623 46427
rect 3893 46325 3927 46359
rect 5457 46325 5491 46359
rect 8861 46325 8895 46359
rect 16221 46325 16255 46359
rect 16957 46325 16991 46359
rect 2053 46121 2087 46155
rect 5181 46121 5215 46155
rect 6101 46121 6135 46155
rect 7021 46121 7055 46155
rect 10609 46121 10643 46155
rect 12265 46121 12299 46155
rect 12633 46121 12667 46155
rect 17417 46121 17451 46155
rect 10241 46053 10275 46087
rect 10701 46053 10735 46087
rect 11069 46053 11103 46087
rect 12817 46053 12851 46087
rect 15669 46053 15703 46087
rect 6837 45985 6871 46019
rect 8033 45985 8067 46019
rect 8677 45985 8711 46019
rect 10517 45985 10551 46019
rect 12725 45985 12759 46019
rect 14657 45985 14691 46019
rect 16681 45985 16715 46019
rect 16957 45985 16991 46019
rect 17141 45985 17175 46019
rect 3801 45917 3835 45951
rect 4077 45917 4111 45951
rect 8585 45917 8619 45951
rect 10333 45917 10367 45951
rect 12449 45917 12483 45951
rect 13185 45917 13219 45951
rect 15301 45917 15335 45951
rect 16129 45917 16163 45951
rect 11897 45849 11931 45883
rect 16037 45849 16071 45883
rect 1593 45781 1627 45815
rect 5825 45781 5859 45815
rect 7297 45781 7331 45815
rect 8953 45781 8987 45815
rect 9873 45781 9907 45815
rect 11437 45781 11471 45815
rect 13461 45781 13495 45815
rect 13829 45781 13863 45815
rect 6745 45577 6779 45611
rect 7389 45577 7423 45611
rect 12909 45577 12943 45611
rect 4261 45509 4295 45543
rect 5089 45509 5123 45543
rect 7757 45509 7791 45543
rect 10885 45509 10919 45543
rect 11253 45509 11287 45543
rect 13277 45509 13311 45543
rect 16313 45509 16347 45543
rect 1501 45441 1535 45475
rect 3157 45441 3191 45475
rect 9505 45441 9539 45475
rect 15117 45441 15151 45475
rect 17325 45441 17359 45475
rect 18061 45441 18095 45475
rect 1777 45373 1811 45407
rect 4721 45373 4755 45407
rect 5641 45373 5675 45407
rect 5917 45373 5951 45407
rect 6285 45373 6319 45407
rect 6929 45373 6963 45407
rect 8493 45373 8527 45407
rect 8861 45373 8895 45407
rect 10149 45373 10183 45407
rect 10333 45373 10367 45407
rect 10609 45373 10643 45407
rect 11437 45373 11471 45407
rect 11805 45373 11839 45407
rect 12173 45373 12207 45407
rect 14197 45373 14231 45407
rect 14657 45373 14691 45407
rect 15485 45373 15519 45407
rect 15945 45373 15979 45407
rect 17601 45373 17635 45407
rect 17785 45373 17819 45407
rect 12633 45305 12667 45339
rect 16773 45305 16807 45339
rect 3801 45237 3835 45271
rect 5457 45237 5491 45271
rect 8125 45237 8159 45271
rect 13645 45237 13679 45271
rect 14013 45237 14047 45271
rect 14381 45237 14415 45271
rect 15669 45237 15703 45271
rect 2053 45033 2087 45067
rect 4261 45033 4295 45067
rect 8125 45033 8159 45067
rect 9781 45033 9815 45067
rect 10149 45033 10183 45067
rect 12173 45033 12207 45067
rect 12725 45033 12759 45067
rect 13001 45033 13035 45067
rect 15577 45033 15611 45067
rect 17509 45033 17543 45067
rect 6837 44965 6871 44999
rect 11529 44965 11563 44999
rect 4169 44897 4203 44931
rect 4721 44897 4755 44931
rect 6561 44897 6595 44931
rect 7527 44897 7561 44931
rect 7665 44897 7699 44931
rect 9045 44897 9079 44931
rect 9229 44897 9263 44931
rect 10609 44897 10643 44931
rect 10885 44897 10919 44931
rect 11345 44897 11379 44931
rect 13461 44897 13495 44931
rect 15209 44897 15243 44931
rect 15761 44897 15795 44931
rect 16037 44897 16071 44931
rect 16681 44897 16715 44931
rect 16957 44897 16991 44931
rect 5181 44829 5215 44863
rect 7389 44829 7423 44863
rect 9505 44829 9539 44863
rect 13185 44829 13219 44863
rect 5641 44761 5675 44795
rect 1593 44693 1627 44727
rect 6009 44693 6043 44727
rect 11805 44693 11839 44727
rect 14565 44693 14599 44727
rect 15761 44693 15795 44727
rect 1685 44489 1719 44523
rect 3525 44489 3559 44523
rect 7205 44489 7239 44523
rect 9413 44489 9447 44523
rect 11069 44489 11103 44523
rect 13277 44489 13311 44523
rect 14749 44489 14783 44523
rect 3893 44421 3927 44455
rect 6193 44421 6227 44455
rect 7389 44421 7423 44455
rect 8861 44421 8895 44455
rect 11529 44421 11563 44455
rect 15669 44421 15703 44455
rect 4905 44353 4939 44387
rect 5549 44353 5583 44387
rect 12725 44353 12759 44387
rect 16589 44353 16623 44387
rect 4261 44285 4295 44319
rect 5733 44285 5767 44319
rect 6285 44285 6319 44319
rect 7481 44285 7515 44319
rect 7941 44285 7975 44319
rect 8125 44285 8159 44319
rect 10241 44285 10275 44319
rect 10517 44285 10551 44319
rect 10701 44285 10735 44319
rect 11621 44285 11655 44319
rect 12265 44285 12299 44319
rect 12633 44285 12667 44319
rect 13921 44285 13955 44319
rect 14013 44285 14047 44319
rect 14381 44285 14415 44319
rect 16129 44285 16163 44319
rect 16497 44285 16531 44319
rect 16865 44285 16899 44319
rect 17601 44285 17635 44319
rect 5181 44217 5215 44251
rect 6837 44217 6871 44251
rect 9689 44217 9723 44251
rect 15025 44217 15059 44251
rect 15945 44217 15979 44251
rect 17877 44217 17911 44251
rect 6285 43945 6319 43979
rect 8309 43945 8343 43979
rect 12081 43945 12115 43979
rect 13001 43945 13035 43979
rect 15577 43945 15611 43979
rect 3157 43877 3191 43911
rect 4169 43877 4203 43911
rect 9413 43877 9447 43911
rect 15209 43877 15243 43911
rect 4905 43809 4939 43843
rect 6929 43809 6963 43843
rect 7297 43809 7331 43843
rect 7757 43809 7791 43843
rect 9965 43809 9999 43843
rect 10333 43809 10367 43843
rect 10977 43809 11011 43843
rect 12725 43809 12759 43843
rect 13461 43809 13495 43843
rect 15761 43809 15795 43843
rect 16037 43809 16071 43843
rect 16405 43809 16439 43843
rect 16957 43809 16991 43843
rect 1501 43741 1535 43775
rect 1777 43741 1811 43775
rect 4077 43741 4111 43775
rect 4997 43741 5031 43775
rect 9781 43741 9815 43775
rect 10425 43741 10459 43775
rect 11713 43741 11747 43775
rect 13185 43741 13219 43775
rect 16129 43741 16163 43775
rect 3893 43673 3927 43707
rect 5733 43673 5767 43707
rect 7757 43673 7791 43707
rect 3525 43605 3559 43639
rect 6561 43605 6595 43639
rect 8769 43605 8803 43639
rect 14565 43605 14599 43639
rect 17417 43605 17451 43639
rect 3525 43401 3559 43435
rect 3893 43401 3927 43435
rect 4169 43401 4203 43435
rect 5089 43401 5123 43435
rect 7389 43401 7423 43435
rect 7757 43401 7791 43435
rect 8309 43401 8343 43435
rect 9045 43401 9079 43435
rect 9505 43401 9539 43435
rect 11529 43401 11563 43435
rect 12357 43401 12391 43435
rect 13553 43401 13587 43435
rect 14197 43401 14231 43435
rect 15117 43401 15151 43435
rect 13921 43333 13955 43367
rect 1501 43265 1535 43299
rect 3157 43265 3191 43299
rect 6285 43265 6319 43299
rect 9873 43265 9907 43299
rect 13185 43265 13219 43299
rect 17417 43265 17451 43299
rect 1777 43197 1811 43231
rect 4077 43197 4111 43231
rect 4813 43197 4847 43231
rect 5917 43197 5951 43231
rect 6009 43197 6043 43231
rect 6377 43197 6411 43231
rect 6929 43197 6963 43231
rect 8585 43197 8619 43231
rect 9781 43197 9815 43231
rect 10057 43197 10091 43231
rect 10425 43197 10459 43231
rect 11989 43197 12023 43231
rect 12541 43197 12575 43231
rect 12909 43197 12943 43231
rect 14013 43197 14047 43231
rect 14473 43197 14507 43231
rect 16037 43197 16071 43231
rect 16681 43197 16715 43231
rect 17049 43197 17083 43231
rect 17325 43197 17359 43231
rect 5549 43061 5583 43095
rect 11253 43061 11287 43095
rect 15669 43061 15703 43095
rect 17877 43061 17911 43095
rect 2329 42857 2363 42891
rect 4997 42857 5031 42891
rect 6101 42857 6135 42891
rect 10517 42857 10551 42891
rect 11897 42857 11931 42891
rect 14289 42857 14323 42891
rect 16681 42857 16715 42891
rect 6653 42789 6687 42823
rect 3709 42721 3743 42755
rect 8217 42721 8251 42755
rect 8401 42721 8435 42755
rect 8769 42721 8803 42755
rect 9137 42721 9171 42755
rect 9689 42721 9723 42755
rect 10241 42721 10275 42755
rect 1961 42653 1995 42687
rect 3433 42653 3467 42687
rect 11529 42789 11563 42823
rect 10977 42721 11011 42755
rect 11069 42721 11103 42755
rect 12265 42721 12299 42755
rect 12909 42721 12943 42755
rect 13553 42721 13587 42755
rect 13829 42721 13863 42755
rect 13185 42653 13219 42687
rect 5733 42585 5767 42619
rect 8217 42585 8251 42619
rect 10517 42585 10551 42619
rect 10793 42585 10827 42619
rect 13921 42585 13955 42619
rect 14841 42721 14875 42755
rect 15209 42721 15243 42755
rect 15393 42721 15427 42755
rect 15945 42721 15979 42755
rect 16221 42721 16255 42755
rect 1593 42517 1627 42551
rect 7021 42517 7055 42551
rect 7757 42517 7791 42551
rect 10701 42517 10735 42551
rect 14289 42517 14323 42551
rect 14473 42517 14507 42551
rect 16129 42517 16163 42551
rect 17049 42517 17083 42551
rect 17417 42517 17451 42551
rect 2881 42313 2915 42347
rect 3525 42313 3559 42347
rect 4353 42313 4387 42347
rect 4813 42313 4847 42347
rect 7205 42313 7239 42347
rect 9505 42313 9539 42347
rect 9873 42313 9907 42347
rect 10241 42313 10275 42347
rect 10793 42313 10827 42347
rect 12173 42313 12207 42347
rect 13093 42313 13127 42347
rect 15025 42313 15059 42347
rect 15577 42313 15611 42347
rect 4997 42245 5031 42279
rect 7573 42245 7607 42279
rect 17233 42245 17267 42279
rect 1501 42177 1535 42211
rect 7757 42177 7791 42211
rect 7849 42177 7883 42211
rect 10609 42177 10643 42211
rect 17601 42177 17635 42211
rect 1777 42109 1811 42143
rect 5181 42109 5215 42143
rect 5641 42109 5675 42143
rect 5733 42109 5767 42143
rect 6101 42109 6135 42143
rect 6745 42109 6779 42143
rect 8585 42109 8619 42143
rect 8677 42109 8711 42143
rect 9137 42109 9171 42143
rect 9689 42109 9723 42143
rect 10701 42109 10735 42143
rect 11345 42109 11379 42143
rect 11713 42109 11747 42143
rect 13461 42109 13495 42143
rect 13645 42109 13679 42143
rect 14105 42109 14139 42143
rect 15853 42109 15887 42143
rect 16497 42109 16531 42143
rect 16865 42109 16899 42143
rect 17141 42109 17175 42143
rect 3893 42041 3927 42075
rect 14381 42041 14415 42075
rect 17969 42041 18003 42075
rect 12541 41973 12575 42007
rect 1961 41769 1995 41803
rect 3433 41769 3467 41803
rect 4353 41769 4387 41803
rect 7573 41769 7607 41803
rect 8309 41769 8343 41803
rect 10333 41769 10367 41803
rect 10701 41769 10735 41803
rect 14289 41769 14323 41803
rect 15117 41769 15151 41803
rect 16957 41769 16991 41803
rect 5917 41701 5951 41735
rect 8033 41701 8067 41735
rect 17325 41701 17359 41735
rect 5181 41633 5215 41667
rect 5641 41633 5675 41667
rect 7297 41633 7331 41667
rect 8493 41633 8527 41667
rect 9137 41633 9171 41667
rect 9505 41633 9539 41667
rect 9781 41633 9815 41667
rect 11437 41633 11471 41667
rect 11529 41633 11563 41667
rect 12449 41633 12483 41667
rect 13001 41633 13035 41667
rect 13461 41633 13495 41667
rect 15301 41633 15335 41667
rect 15577 41633 15611 41667
rect 15945 41633 15979 41667
rect 16681 41633 16715 41667
rect 4721 41565 4755 41599
rect 4997 41565 5031 41599
rect 12541 41565 12575 41599
rect 14657 41565 14691 41599
rect 15761 41565 15795 41599
rect 1593 41429 1627 41463
rect 6653 41429 6687 41463
rect 8585 41429 8619 41463
rect 12081 41429 12115 41463
rect 14013 41429 14047 41463
rect 3065 41225 3099 41259
rect 4629 41225 4663 41259
rect 6193 41225 6227 41259
rect 8769 41225 8803 41259
rect 14749 41225 14783 41259
rect 17969 41225 18003 41259
rect 5549 41157 5583 41191
rect 7481 41157 7515 41191
rect 9045 41157 9079 41191
rect 9413 41157 9447 41191
rect 9781 41157 9815 41191
rect 1501 41089 1535 41123
rect 4905 41089 4939 41123
rect 12633 41089 12667 41123
rect 13829 41089 13863 41123
rect 16773 41089 16807 41123
rect 1777 41021 1811 41055
rect 3893 41021 3927 41055
rect 5089 41021 5123 41055
rect 5641 41021 5675 41055
rect 6653 41021 6687 41055
rect 7021 41021 7055 41055
rect 7481 41021 7515 41055
rect 8585 41021 8619 41055
rect 9689 41021 9723 41055
rect 10057 41021 10091 41055
rect 10425 41021 10459 41055
rect 10977 41021 11011 41055
rect 11805 41021 11839 41055
rect 12173 41021 12207 41055
rect 12357 41021 12391 41055
rect 13001 41021 13035 41055
rect 13277 41021 13311 41055
rect 14197 41021 14231 41055
rect 16129 41021 16163 41055
rect 16221 41021 16255 41055
rect 16589 41021 16623 41055
rect 17325 41021 17359 41055
rect 11529 40953 11563 40987
rect 6561 40885 6595 40919
rect 8125 40885 8159 40919
rect 8493 40885 8527 40919
rect 15025 40885 15059 40919
rect 15485 40885 15519 40919
rect 17601 40885 17635 40919
rect 5089 40681 5123 40715
rect 5917 40681 5951 40715
rect 7021 40681 7055 40715
rect 7573 40681 7607 40715
rect 16405 40681 16439 40715
rect 16773 40681 16807 40715
rect 4721 40613 4755 40647
rect 8309 40613 8343 40647
rect 11529 40613 11563 40647
rect 13553 40613 13587 40647
rect 4905 40545 4939 40579
rect 6653 40545 6687 40579
rect 7389 40545 7423 40579
rect 8677 40545 8711 40579
rect 9045 40545 9079 40579
rect 9229 40545 9263 40579
rect 9689 40545 9723 40579
rect 10517 40545 10551 40579
rect 10793 40545 10827 40579
rect 10885 40545 10919 40579
rect 11069 40545 11103 40579
rect 12817 40545 12851 40579
rect 13093 40545 13127 40579
rect 13921 40545 13955 40579
rect 14565 40545 14599 40579
rect 15025 40545 15059 40579
rect 15393 40545 15427 40579
rect 15853 40545 15887 40579
rect 16865 40545 16899 40579
rect 8861 40477 8895 40511
rect 13277 40477 13311 40511
rect 14105 40477 14139 40511
rect 4353 40409 4387 40443
rect 6285 40409 6319 40443
rect 14197 40409 14231 40443
rect 17049 40409 17083 40443
rect 1593 40341 1627 40375
rect 1961 40341 1995 40375
rect 7941 40341 7975 40375
rect 10149 40341 10183 40375
rect 12081 40341 12115 40375
rect 17325 40341 17359 40375
rect 3801 40137 3835 40171
rect 11989 40137 12023 40171
rect 13737 40137 13771 40171
rect 14841 40137 14875 40171
rect 15485 40137 15519 40171
rect 17233 40137 17267 40171
rect 9781 40069 9815 40103
rect 14105 40069 14139 40103
rect 17785 40069 17819 40103
rect 5089 40001 5123 40035
rect 6561 40001 6595 40035
rect 3525 39933 3559 39967
rect 4261 39933 4295 39967
rect 4813 39933 4847 39967
rect 6285 39933 6319 39967
rect 6653 39933 6687 39967
rect 7205 39933 7239 39967
rect 7481 39933 7515 39967
rect 7849 39933 7883 39967
rect 9965 39933 9999 39967
rect 10241 39933 10275 39967
rect 11713 39933 11747 39967
rect 11897 39933 11931 39967
rect 12541 39933 12575 39967
rect 12633 39933 12667 39967
rect 13921 39933 13955 39967
rect 14381 39933 14415 39967
rect 16313 39933 16347 39967
rect 16405 39933 16439 39967
rect 16773 39933 16807 39967
rect 17325 39933 17359 39967
rect 6101 39865 6135 39899
rect 9413 39865 9447 39899
rect 15853 39865 15887 39899
rect 4353 39797 4387 39831
rect 5733 39797 5767 39831
rect 8493 39797 8527 39831
rect 8861 39797 8895 39831
rect 10885 39797 10919 39831
rect 11253 39797 11287 39831
rect 13369 39797 13403 39831
rect 4353 39593 4387 39627
rect 4629 39593 4663 39627
rect 5549 39593 5583 39627
rect 6285 39593 6319 39627
rect 8309 39593 8343 39627
rect 10057 39593 10091 39627
rect 11897 39593 11931 39627
rect 14565 39593 14599 39627
rect 17325 39593 17359 39627
rect 7849 39525 7883 39559
rect 14197 39525 14231 39559
rect 3249 39457 3283 39491
rect 3709 39457 3743 39491
rect 4629 39457 4663 39491
rect 5089 39457 5123 39491
rect 7389 39457 7423 39491
rect 7665 39457 7699 39491
rect 8769 39457 8803 39491
rect 10885 39457 10919 39491
rect 11345 39457 11379 39491
rect 12817 39457 12851 39491
rect 15577 39457 15611 39491
rect 15945 39457 15979 39491
rect 16313 39457 16347 39491
rect 16865 39457 16899 39491
rect 3341 39389 3375 39423
rect 11161 39389 11195 39423
rect 12541 39389 12575 39423
rect 15485 39389 15519 39423
rect 6653 39253 6687 39287
rect 8677 39253 8711 39287
rect 14933 39253 14967 39287
rect 15669 39253 15703 39287
rect 2697 39049 2731 39083
rect 3065 39049 3099 39083
rect 3433 39049 3467 39083
rect 3801 39049 3835 39083
rect 5457 39049 5491 39083
rect 6929 39049 6963 39083
rect 8401 39049 8435 39083
rect 13645 39049 13679 39083
rect 14381 39049 14415 39083
rect 15945 39049 15979 39083
rect 18245 39049 18279 39083
rect 6285 38981 6319 39015
rect 16221 38981 16255 39015
rect 4169 38913 4203 38947
rect 4261 38913 4295 38947
rect 10609 38913 10643 38947
rect 13001 38913 13035 38947
rect 15669 38913 15703 38947
rect 4997 38845 5031 38879
rect 5089 38845 5123 38879
rect 6837 38845 6871 38879
rect 7481 38845 7515 38879
rect 7573 38845 7607 38879
rect 8493 38845 8527 38879
rect 8861 38845 8895 38879
rect 9321 38845 9355 38879
rect 10057 38845 10091 38879
rect 10425 38845 10459 38879
rect 10793 38845 10827 38879
rect 11069 38845 11103 38879
rect 11989 38845 12023 38879
rect 12173 38845 12207 38879
rect 12817 38845 12851 38879
rect 13185 38845 13219 38879
rect 14197 38845 14231 38879
rect 14657 38845 14691 38879
rect 15117 38845 15151 38879
rect 16313 38845 16347 38879
rect 16497 38845 16531 38879
rect 16865 38845 16899 38879
rect 17417 38845 17451 38879
rect 2329 38777 2363 38811
rect 6009 38777 6043 38811
rect 11713 38777 11747 38811
rect 14105 38777 14139 38811
rect 17877 38777 17911 38811
rect 6653 38709 6687 38743
rect 3893 38505 3927 38539
rect 5365 38505 5399 38539
rect 6561 38505 6595 38539
rect 7021 38505 7055 38539
rect 7941 38505 7975 38539
rect 11805 38505 11839 38539
rect 13461 38505 13495 38539
rect 14013 38505 14047 38539
rect 14473 38505 14507 38539
rect 16405 38505 16439 38539
rect 16773 38505 16807 38539
rect 17049 38505 17083 38539
rect 3157 38437 3191 38471
rect 7573 38437 7607 38471
rect 10057 38437 10091 38471
rect 10609 38437 10643 38471
rect 11529 38437 11563 38471
rect 12173 38437 12207 38471
rect 1777 38369 1811 38403
rect 4261 38369 4295 38403
rect 6837 38369 6871 38403
rect 8033 38369 8067 38403
rect 8677 38369 8711 38403
rect 8769 38369 8803 38403
rect 9321 38369 9355 38403
rect 1501 38301 1535 38335
rect 3985 38301 4019 38335
rect 10793 38369 10827 38403
rect 11253 38369 11287 38403
rect 13001 38369 13035 38403
rect 13277 38369 13311 38403
rect 14749 38369 14783 38403
rect 14933 38369 14967 38403
rect 15577 38369 15611 38403
rect 15853 38369 15887 38403
rect 16865 38369 16899 38403
rect 10241 38301 10275 38335
rect 17325 38301 17359 38335
rect 10057 38233 10091 38267
rect 12909 38233 12943 38267
rect 13093 38233 13127 38267
rect 3525 38165 3559 38199
rect 6193 38165 6227 38199
rect 9229 38165 9263 38199
rect 9873 38165 9907 38199
rect 14657 38165 14691 38199
rect 3065 37961 3099 37995
rect 3525 37961 3559 37995
rect 9137 37961 9171 37995
rect 13829 37961 13863 37995
rect 14381 37961 14415 37995
rect 15117 37961 15151 37995
rect 15945 37961 15979 37995
rect 17785 37961 17819 37995
rect 7389 37893 7423 37927
rect 9689 37825 9723 37859
rect 12633 37825 12667 37859
rect 16865 37825 16899 37859
rect 1501 37757 1535 37791
rect 1777 37757 1811 37791
rect 4077 37757 4111 37791
rect 4353 37757 4387 37791
rect 6745 37757 6779 37791
rect 6929 37757 6963 37791
rect 7481 37757 7515 37791
rect 8493 37757 8527 37791
rect 10425 37757 10459 37791
rect 11989 37757 12023 37791
rect 12357 37757 12391 37791
rect 12725 37757 12759 37791
rect 14197 37757 14231 37791
rect 16037 37757 16071 37791
rect 16405 37757 16439 37791
rect 16773 37757 16807 37791
rect 17325 37757 17359 37791
rect 5733 37689 5767 37723
rect 6101 37689 6135 37723
rect 9505 37689 9539 37723
rect 9873 37689 9907 37723
rect 10057 37689 10091 37723
rect 14657 37689 14691 37723
rect 15485 37689 15519 37723
rect 3801 37621 3835 37655
rect 6469 37621 6503 37655
rect 8125 37621 8159 37655
rect 8677 37621 8711 37655
rect 9965 37621 9999 37655
rect 10793 37621 10827 37655
rect 11161 37621 11195 37655
rect 11897 37621 11931 37655
rect 13553 37621 13587 37655
rect 4997 37417 5031 37451
rect 6653 37417 6687 37451
rect 7297 37417 7331 37451
rect 7757 37417 7791 37451
rect 11437 37417 11471 37451
rect 13737 37417 13771 37451
rect 17417 37417 17451 37451
rect 6285 37349 6319 37383
rect 8493 37349 8527 37383
rect 12541 37349 12575 37383
rect 1593 37281 1627 37315
rect 1961 37281 1995 37315
rect 6837 37281 6871 37315
rect 8125 37281 8159 37315
rect 8769 37281 8803 37315
rect 9137 37281 9171 37315
rect 9321 37281 9355 37315
rect 9689 37281 9723 37315
rect 10057 37281 10091 37315
rect 10793 37281 10827 37315
rect 11253 37281 11287 37315
rect 12081 37281 12115 37315
rect 12725 37281 12759 37315
rect 14473 37281 14507 37315
rect 15025 37281 15059 37315
rect 15577 37281 15611 37315
rect 15853 37281 15887 37315
rect 16405 37281 16439 37315
rect 16957 37281 16991 37315
rect 3617 37213 3651 37247
rect 3893 37213 3927 37247
rect 14289 37213 14323 37247
rect 15117 37213 15151 37247
rect 16129 37213 16163 37247
rect 17141 37213 17175 37247
rect 7021 37145 7055 37179
rect 2329 37077 2363 37111
rect 3157 37077 3191 37111
rect 3433 37077 3467 37111
rect 5641 37077 5675 37111
rect 11069 37077 11103 37111
rect 4445 36873 4479 36907
rect 8493 36873 8527 36907
rect 8953 36873 8987 36907
rect 10241 36873 10275 36907
rect 10885 36873 10919 36907
rect 12173 36873 12207 36907
rect 12817 36873 12851 36907
rect 13553 36873 13587 36907
rect 15025 36873 15059 36907
rect 15485 36873 15519 36907
rect 18061 36873 18095 36907
rect 3709 36805 3743 36839
rect 4997 36805 5031 36839
rect 9229 36805 9263 36839
rect 9965 36805 9999 36839
rect 12541 36805 12575 36839
rect 14473 36805 14507 36839
rect 14749 36805 14783 36839
rect 4813 36737 4847 36771
rect 7205 36737 7239 36771
rect 13645 36737 13679 36771
rect 14381 36737 14415 36771
rect 5181 36669 5215 36703
rect 5549 36669 5583 36703
rect 5733 36669 5767 36703
rect 6285 36669 6319 36703
rect 7665 36669 7699 36703
rect 7987 36669 8021 36703
rect 8125 36669 8159 36703
rect 10701 36669 10735 36703
rect 12633 36669 12667 36703
rect 13093 36669 13127 36703
rect 15301 36669 15335 36703
rect 15761 36669 15795 36703
rect 16865 36669 16899 36703
rect 17233 36669 17267 36703
rect 17509 36669 17543 36703
rect 13921 36601 13955 36635
rect 14013 36601 14047 36635
rect 14473 36601 14507 36635
rect 16589 36601 16623 36635
rect 17785 36601 17819 36635
rect 1685 36533 1719 36567
rect 3249 36533 3283 36567
rect 6653 36533 6687 36567
rect 7021 36533 7055 36567
rect 11621 36533 11655 36567
rect 13829 36533 13863 36567
rect 16129 36533 16163 36567
rect 4813 36329 4847 36363
rect 6653 36329 6687 36363
rect 8585 36329 8619 36363
rect 9321 36329 9355 36363
rect 10609 36329 10643 36363
rect 12173 36329 12207 36363
rect 12725 36329 12759 36363
rect 13461 36329 13495 36363
rect 14105 36329 14139 36363
rect 14473 36329 14507 36363
rect 16405 36329 16439 36363
rect 17049 36329 17083 36363
rect 17417 36329 17451 36363
rect 4905 36261 4939 36295
rect 6285 36261 6319 36295
rect 8033 36261 8067 36295
rect 11529 36261 11563 36295
rect 5365 36193 5399 36227
rect 7021 36193 7055 36227
rect 7205 36193 7239 36227
rect 7573 36193 7607 36227
rect 9229 36193 9263 36227
rect 11345 36193 11379 36227
rect 13093 36193 13127 36227
rect 14749 36193 14783 36227
rect 14933 36193 14967 36227
rect 15301 36193 15335 36227
rect 16037 36193 16071 36227
rect 16865 36193 16899 36227
rect 1685 35989 1719 36023
rect 15945 35989 15979 36023
rect 16681 35989 16715 36023
rect 3065 35785 3099 35819
rect 4997 35785 5031 35819
rect 6377 35785 6411 35819
rect 7481 35785 7515 35819
rect 7849 35785 7883 35819
rect 8953 35785 8987 35819
rect 9321 35785 9355 35819
rect 10517 35785 10551 35819
rect 11069 35785 11103 35819
rect 12541 35785 12575 35819
rect 13093 35785 13127 35819
rect 14105 35785 14139 35819
rect 14749 35785 14783 35819
rect 15577 35785 15611 35819
rect 15853 35785 15887 35819
rect 16589 35785 16623 35819
rect 18153 35785 18187 35819
rect 8585 35717 8619 35751
rect 10149 35717 10183 35751
rect 14381 35717 14415 35751
rect 17509 35717 17543 35751
rect 1501 35649 1535 35683
rect 1777 35581 1811 35615
rect 6009 35581 6043 35615
rect 6745 35581 6779 35615
rect 7665 35581 7699 35615
rect 8125 35581 8159 35615
rect 9965 35581 9999 35615
rect 10885 35581 10919 35615
rect 11253 35581 11287 35615
rect 11713 35581 11747 35615
rect 11989 35581 12023 35615
rect 13185 35581 13219 35615
rect 14197 35581 14231 35615
rect 15393 35581 15427 35615
rect 16681 35581 16715 35615
rect 17233 35581 17267 35615
rect 17601 35581 17635 35615
rect 18429 35581 18463 35615
rect 7205 35445 7239 35479
rect 13369 35445 13403 35479
rect 13737 35445 13771 35479
rect 15025 35445 15059 35479
rect 6009 35241 6043 35275
rect 14197 35241 14231 35275
rect 14657 35241 14691 35275
rect 17417 35241 17451 35275
rect 10609 35173 10643 35207
rect 2605 35105 2639 35139
rect 7389 35105 7423 35139
rect 7527 35105 7561 35139
rect 7665 35105 7699 35139
rect 10701 35105 10735 35139
rect 13737 35105 13771 35139
rect 14749 35105 14783 35139
rect 16221 35105 16255 35139
rect 16589 35105 16623 35139
rect 16865 35105 16899 35139
rect 2329 35037 2363 35071
rect 3985 35037 4019 35071
rect 6837 35037 6871 35071
rect 15945 35037 15979 35071
rect 17141 35037 17175 35071
rect 4445 34969 4479 35003
rect 13921 34969 13955 35003
rect 14933 34969 14967 35003
rect 1593 34901 1627 34935
rect 4813 34901 4847 34935
rect 6377 34901 6411 34935
rect 9965 34901 9999 34935
rect 5825 34697 5859 34731
rect 6193 34697 6227 34731
rect 14749 34697 14783 34731
rect 15577 34697 15611 34731
rect 16221 34697 16255 34731
rect 2329 34629 2363 34663
rect 15853 34629 15887 34663
rect 17509 34629 17543 34663
rect 4537 34561 4571 34595
rect 5457 34561 5491 34595
rect 16865 34561 16899 34595
rect 18061 34561 18095 34595
rect 2697 34493 2731 34527
rect 3893 34493 3927 34527
rect 4905 34493 4939 34527
rect 5181 34493 5215 34527
rect 6285 34493 6319 34527
rect 6745 34493 6779 34527
rect 7481 34493 7515 34527
rect 7941 34493 7975 34527
rect 8493 34493 8527 34527
rect 10609 34493 10643 34527
rect 13829 34493 13863 34527
rect 15393 34493 15427 34527
rect 17233 34493 17267 34527
rect 17509 34493 17543 34527
rect 7205 34357 7239 34391
rect 6009 34153 6043 34187
rect 14197 34153 14231 34187
rect 15577 34153 15611 34187
rect 17417 34153 17451 34187
rect 6377 34085 6411 34119
rect 3525 34017 3559 34051
rect 6837 34017 6871 34051
rect 7389 34017 7423 34051
rect 7665 34017 7699 34051
rect 9597 34017 9631 34051
rect 9689 34017 9723 34051
rect 10057 34017 10091 34051
rect 14197 34017 14231 34051
rect 14841 34017 14875 34051
rect 15945 34017 15979 34051
rect 16497 34017 16531 34051
rect 16865 34017 16899 34051
rect 3249 33949 3283 33983
rect 4905 33949 4939 33983
rect 9781 33949 9815 33983
rect 14933 33949 14967 33983
rect 16221 33949 16255 33983
rect 17141 33949 17175 33983
rect 6929 33881 6963 33915
rect 3341 33609 3375 33643
rect 6653 33609 6687 33643
rect 8309 33609 8343 33643
rect 9045 33609 9079 33643
rect 9413 33609 9447 33643
rect 10425 33609 10459 33643
rect 14841 33609 14875 33643
rect 15577 33609 15611 33643
rect 15853 33609 15887 33643
rect 17509 33541 17543 33575
rect 6101 33473 6135 33507
rect 18429 33473 18463 33507
rect 4077 33405 4111 33439
rect 4353 33405 4387 33439
rect 6561 33405 6595 33439
rect 6929 33405 6963 33439
rect 7297 33405 7331 33439
rect 7849 33405 7883 33439
rect 9873 33405 9907 33439
rect 15669 33405 15703 33439
rect 16681 33405 16715 33439
rect 17049 33405 17083 33439
rect 17601 33405 17635 33439
rect 2053 33337 2087 33371
rect 2881 33337 2915 33371
rect 5733 33337 5767 33371
rect 6469 33337 6503 33371
rect 10701 33337 10735 33371
rect 1685 33269 1719 33303
rect 3801 33269 3835 33303
rect 10057 33269 10091 33303
rect 14105 33269 14139 33303
rect 14473 33269 14507 33303
rect 16221 33269 16255 33303
rect 16589 33269 16623 33303
rect 18061 33269 18095 33303
rect 2973 33065 3007 33099
rect 6285 33065 6319 33099
rect 6653 33065 6687 33099
rect 7113 33065 7147 33099
rect 7481 33065 7515 33099
rect 15393 33065 15427 33099
rect 15853 33065 15887 33099
rect 17785 33065 17819 33099
rect 17141 32997 17175 33031
rect 17417 32997 17451 33031
rect 4353 32929 4387 32963
rect 4721 32929 4755 32963
rect 5089 32929 5123 32963
rect 5457 32929 5491 32963
rect 5917 32929 5951 32963
rect 9597 32929 9631 32963
rect 9965 32929 9999 32963
rect 10149 32929 10183 32963
rect 10609 32929 10643 32963
rect 14013 32929 14047 32963
rect 14657 32929 14691 32963
rect 14841 32929 14875 32963
rect 16037 32929 16071 32963
rect 16405 32929 16439 32963
rect 16865 32929 16899 32963
rect 1409 32861 1443 32895
rect 1685 32861 1719 32895
rect 4537 32861 4571 32895
rect 9873 32861 9907 32895
rect 14289 32793 14323 32827
rect 3893 32725 3927 32759
rect 9137 32725 9171 32759
rect 11069 32725 11103 32759
rect 11437 32725 11471 32759
rect 2881 32521 2915 32555
rect 3525 32521 3559 32555
rect 5089 32521 5123 32555
rect 8033 32521 8067 32555
rect 8401 32521 8435 32555
rect 9045 32521 9079 32555
rect 14473 32521 14507 32555
rect 16129 32521 16163 32555
rect 18429 32521 18463 32555
rect 9321 32453 9355 32487
rect 1777 32385 1811 32419
rect 4537 32385 4571 32419
rect 4905 32385 4939 32419
rect 10149 32385 10183 32419
rect 11069 32385 11103 32419
rect 1501 32317 1535 32351
rect 4997 32317 5031 32351
rect 5365 32317 5399 32351
rect 5825 32317 5859 32351
rect 6377 32317 6411 32351
rect 8217 32317 8251 32351
rect 10609 32317 10643 32351
rect 11161 32317 11195 32351
rect 11621 32317 11655 32351
rect 11805 32317 11839 32351
rect 15485 32317 15519 32351
rect 16681 32317 16715 32351
rect 17233 32317 17267 32351
rect 17509 32317 17543 32351
rect 18061 32317 18095 32351
rect 3893 32249 3927 32283
rect 10517 32249 10551 32283
rect 14013 32249 14047 32283
rect 15117 32249 15151 32283
rect 15301 32249 15335 32283
rect 17785 32249 17819 32283
rect 13645 32181 13679 32215
rect 15577 32181 15611 32215
rect 16589 32181 16623 32215
rect 5365 31977 5399 32011
rect 5917 31977 5951 32011
rect 7665 31977 7699 32011
rect 9413 31977 9447 32011
rect 9873 31977 9907 32011
rect 12633 31977 12667 32011
rect 15577 31977 15611 32011
rect 3157 31909 3191 31943
rect 4537 31909 4571 31943
rect 5089 31909 5123 31943
rect 16037 31909 16071 31943
rect 16405 31909 16439 31943
rect 16497 31909 16531 31943
rect 16865 31909 16899 31943
rect 17233 31909 17267 31943
rect 1777 31841 1811 31875
rect 5825 31841 5859 31875
rect 6101 31841 6135 31875
rect 7757 31841 7791 31875
rect 8217 31841 8251 31875
rect 10241 31841 10275 31875
rect 11069 31841 11103 31875
rect 11437 31841 11471 31875
rect 12449 31841 12483 31875
rect 14565 31841 14599 31875
rect 14657 31841 14691 31875
rect 14841 31841 14875 31875
rect 15301 31841 15335 31875
rect 16313 31841 16347 31875
rect 1501 31773 1535 31807
rect 8585 31773 8619 31807
rect 16129 31773 16163 31807
rect 17509 31773 17543 31807
rect 10517 31705 10551 31739
rect 1961 31433 1995 31467
rect 5825 31433 5859 31467
rect 6469 31433 6503 31467
rect 7481 31433 7515 31467
rect 8677 31433 8711 31467
rect 14933 31433 14967 31467
rect 16497 31433 16531 31467
rect 2329 31365 2363 31399
rect 14289 31365 14323 31399
rect 8125 31297 8159 31331
rect 9137 31297 9171 31331
rect 15853 31297 15887 31331
rect 6285 31229 6319 31263
rect 7113 31229 7147 31263
rect 7849 31229 7883 31263
rect 8033 31229 8067 31263
rect 9505 31229 9539 31263
rect 9873 31229 9907 31263
rect 10333 31229 10367 31263
rect 10701 31229 10735 31263
rect 11805 31229 11839 31263
rect 12265 31229 12299 31263
rect 15485 31229 15519 31263
rect 16681 31229 16715 31263
rect 17233 31229 17267 31263
rect 17509 31229 17543 31263
rect 1593 31161 1627 31195
rect 12817 31161 12851 31195
rect 15301 31161 15335 31195
rect 17785 31161 17819 31195
rect 6101 31093 6135 31127
rect 9965 31093 9999 31127
rect 11621 31093 11655 31127
rect 12081 31093 12115 31127
rect 14657 31093 14691 31127
rect 16129 31093 16163 31127
rect 4721 30889 4755 30923
rect 8033 30889 8067 30923
rect 9873 30889 9907 30923
rect 10609 30889 10643 30923
rect 16037 30889 16071 30923
rect 16313 30889 16347 30923
rect 17509 30889 17543 30923
rect 3341 30821 3375 30855
rect 5917 30821 5951 30855
rect 10333 30821 10367 30855
rect 11805 30821 11839 30855
rect 15853 30821 15887 30855
rect 16497 30821 16531 30855
rect 16865 30821 16899 30855
rect 1961 30753 1995 30787
rect 5365 30753 5399 30787
rect 5641 30753 5675 30787
rect 1685 30685 1719 30719
rect 4997 30685 5031 30719
rect 15393 30617 15427 30651
rect 16405 30753 16439 30787
rect 16129 30685 16163 30719
rect 7665 30549 7699 30583
rect 12725 30549 12759 30583
rect 15853 30549 15887 30583
rect 17141 30549 17175 30583
rect 4629 30345 4663 30379
rect 15577 30345 15611 30379
rect 7573 30277 7607 30311
rect 12909 30277 12943 30311
rect 14749 30277 14783 30311
rect 15117 30277 15151 30311
rect 15853 30277 15887 30311
rect 16497 30277 16531 30311
rect 5181 30209 5215 30243
rect 9689 30209 9723 30243
rect 17785 30209 17819 30243
rect 5089 30141 5123 30175
rect 5457 30141 5491 30175
rect 5825 30141 5859 30175
rect 6561 30141 6595 30175
rect 7389 30141 7423 30175
rect 7849 30141 7883 30175
rect 8401 30141 8435 30175
rect 8861 30141 8895 30175
rect 9505 30141 9539 30175
rect 10333 30141 10367 30175
rect 13093 30141 13127 30175
rect 13277 30141 13311 30175
rect 13461 30141 13495 30175
rect 15669 30141 15703 30175
rect 16129 30141 16163 30175
rect 16681 30141 16715 30175
rect 17049 30141 17083 30175
rect 17509 30141 17543 30175
rect 18061 30141 18095 30175
rect 4997 30073 5031 30107
rect 1685 30005 1719 30039
rect 2145 30005 2179 30039
rect 6837 30005 6871 30039
rect 8585 30005 8619 30039
rect 12081 30005 12115 30039
rect 12541 30005 12575 30039
rect 1685 29801 1719 29835
rect 4537 29801 4571 29835
rect 5181 29801 5215 29835
rect 5549 29801 5583 29835
rect 7021 29801 7055 29835
rect 13369 29801 13403 29835
rect 15301 29801 15335 29835
rect 17141 29801 17175 29835
rect 3709 29733 3743 29767
rect 4445 29733 4479 29767
rect 5917 29733 5951 29767
rect 8217 29733 8251 29767
rect 15945 29733 15979 29767
rect 2053 29665 2087 29699
rect 2329 29665 2363 29699
rect 4721 29665 4755 29699
rect 6837 29665 6871 29699
rect 8309 29665 8343 29699
rect 9137 29665 9171 29699
rect 9321 29665 9355 29699
rect 10885 29665 10919 29699
rect 12449 29665 12483 29699
rect 13277 29665 13311 29699
rect 14381 29665 14415 29699
rect 16037 29665 16071 29699
rect 7757 29597 7791 29631
rect 13185 29597 13219 29631
rect 15761 29597 15795 29631
rect 9413 29461 9447 29495
rect 10701 29461 10735 29495
rect 12265 29461 12299 29495
rect 14565 29461 14599 29495
rect 16221 29461 16255 29495
rect 16773 29461 16807 29495
rect 17509 29461 17543 29495
rect 7481 29257 7515 29291
rect 9505 29257 9539 29291
rect 10149 29257 10183 29291
rect 10701 29257 10735 29291
rect 14381 29257 14415 29291
rect 16129 29257 16163 29291
rect 1501 29121 1535 29155
rect 5457 29121 5491 29155
rect 6837 29121 6871 29155
rect 9045 29121 9079 29155
rect 13829 29121 13863 29155
rect 15117 29121 15151 29155
rect 15301 29121 15335 29155
rect 1777 29053 1811 29087
rect 5365 29053 5399 29087
rect 7665 29053 7699 29087
rect 8309 29053 8343 29087
rect 8493 29053 8527 29087
rect 10333 29053 10367 29087
rect 12633 29053 12667 29087
rect 13001 29053 13035 29087
rect 13645 29053 13679 29087
rect 15393 29053 15427 29087
rect 16681 29053 16715 29087
rect 17141 29053 17175 29087
rect 17509 29053 17543 29087
rect 17785 29053 17819 29087
rect 3157 28985 3191 29019
rect 4629 28985 4663 29019
rect 4997 28985 5031 29019
rect 5641 28985 5675 29019
rect 5733 28985 5767 29019
rect 5825 28985 5859 29019
rect 6193 28985 6227 29019
rect 11805 28985 11839 29019
rect 15853 28985 15887 29019
rect 3433 28917 3467 28951
rect 7941 28917 7975 28951
rect 11437 28917 11471 28951
rect 12173 28917 12207 28951
rect 12541 28917 12575 28951
rect 16589 28917 16623 28951
rect 2237 28713 2271 28747
rect 2605 28713 2639 28747
rect 3433 28713 3467 28747
rect 6285 28713 6319 28747
rect 7113 28713 7147 28747
rect 7757 28713 7791 28747
rect 10333 28713 10367 28747
rect 12265 28713 12299 28747
rect 12725 28713 12759 28747
rect 13921 28713 13955 28747
rect 15853 28713 15887 28747
rect 17785 28713 17819 28747
rect 1409 28645 1443 28679
rect 15117 28645 15151 28679
rect 15485 28645 15519 28679
rect 17141 28645 17175 28679
rect 1593 28577 1627 28611
rect 3617 28577 3651 28611
rect 5273 28577 5307 28611
rect 5917 28577 5951 28611
rect 6929 28577 6963 28611
rect 8033 28577 8067 28611
rect 8493 28577 8527 28611
rect 8861 28577 8895 28611
rect 10149 28577 10183 28611
rect 10609 28577 10643 28611
rect 11345 28577 11379 28611
rect 12449 28577 12483 28611
rect 12909 28577 12943 28611
rect 13277 28577 13311 28611
rect 14657 28577 14691 28611
rect 16497 28577 16531 28611
rect 16865 28577 16899 28611
rect 1961 28509 1995 28543
rect 16221 28509 16255 28543
rect 4629 28441 4663 28475
rect 8769 28441 8803 28475
rect 11529 28441 11563 28475
rect 11897 28373 11931 28407
rect 17417 28373 17451 28407
rect 1961 28169 1995 28203
rect 2421 28169 2455 28203
rect 3525 28169 3559 28203
rect 7665 28169 7699 28203
rect 9045 28169 9079 28203
rect 9413 28169 9447 28203
rect 16129 28169 16163 28203
rect 7297 28101 7331 28135
rect 1685 28033 1719 28067
rect 6653 28033 6687 28067
rect 8309 28033 8343 28067
rect 8769 28033 8803 28067
rect 12081 28033 12115 28067
rect 14657 28033 14691 28067
rect 15301 28033 15335 28067
rect 17785 28033 17819 28067
rect 3893 27965 3927 27999
rect 4721 27965 4755 27999
rect 5825 27965 5859 27999
rect 6193 27965 6227 27999
rect 8585 27965 8619 27999
rect 10885 27965 10919 27999
rect 11897 27965 11931 27999
rect 12909 27965 12943 27999
rect 13185 27965 13219 27999
rect 13461 27965 13495 27999
rect 13645 27965 13679 27999
rect 13921 27965 13955 27999
rect 14381 27965 14415 27999
rect 15393 27965 15427 27999
rect 16681 27965 16715 27999
rect 17233 27965 17267 27999
rect 17509 27965 17543 27999
rect 7757 27897 7791 27931
rect 15853 27897 15887 27931
rect 16497 27897 16531 27931
rect 18061 27897 18095 27931
rect 4353 27829 4387 27863
rect 5273 27829 5307 27863
rect 5733 27829 5767 27863
rect 10149 27829 10183 27863
rect 11253 27829 11287 27863
rect 12449 27829 12483 27863
rect 12817 27829 12851 27863
rect 15025 27829 15059 27863
rect 5733 27625 5767 27659
rect 7021 27625 7055 27659
rect 8401 27625 8435 27659
rect 8769 27625 8803 27659
rect 12173 27625 12207 27659
rect 15393 27625 15427 27659
rect 17417 27625 17451 27659
rect 3709 27557 3743 27591
rect 5273 27557 5307 27591
rect 6653 27557 6687 27591
rect 13277 27557 13311 27591
rect 16037 27557 16071 27591
rect 1961 27489 1995 27523
rect 4261 27489 4295 27523
rect 4721 27489 4755 27523
rect 4997 27489 5031 27523
rect 7297 27489 7331 27523
rect 8033 27489 8067 27523
rect 10333 27489 10367 27523
rect 11345 27489 11379 27523
rect 12725 27489 12759 27523
rect 14105 27489 14139 27523
rect 14565 27489 14599 27523
rect 16681 27489 16715 27523
rect 16957 27489 16991 27523
rect 1685 27421 1719 27455
rect 4077 27421 4111 27455
rect 14657 27421 14691 27455
rect 16129 27421 16163 27455
rect 17141 27421 17175 27455
rect 11529 27353 11563 27387
rect 17785 27353 17819 27387
rect 3249 27285 3283 27319
rect 6101 27285 6135 27319
rect 7389 27285 7423 27319
rect 10517 27285 10551 27319
rect 11897 27285 11931 27319
rect 13553 27285 13587 27319
rect 13921 27285 13955 27319
rect 1777 27081 1811 27115
rect 3525 27081 3559 27115
rect 3893 27081 3927 27115
rect 6469 27081 6503 27115
rect 10425 27081 10459 27115
rect 12173 27081 12207 27115
rect 12725 27081 12759 27115
rect 13553 27081 13587 27115
rect 15577 27081 15611 27115
rect 7849 27013 7883 27047
rect 8401 27013 8435 27047
rect 11713 27013 11747 27047
rect 15853 27013 15887 27047
rect 17509 27013 17543 27047
rect 2789 26945 2823 26979
rect 5457 26945 5491 26979
rect 7205 26945 7239 26979
rect 8769 26945 8803 26979
rect 11253 26945 11287 26979
rect 16865 26945 16899 26979
rect 18061 26945 18095 26979
rect 2329 26877 2363 26911
rect 2697 26877 2731 26911
rect 3157 26877 3191 26911
rect 4077 26877 4111 26911
rect 4353 26877 4387 26911
rect 6101 26877 6135 26911
rect 6745 26877 6779 26911
rect 7481 26877 7515 26911
rect 7849 26877 7883 26911
rect 10701 26877 10735 26911
rect 11989 26877 12023 26911
rect 13921 26877 13955 26911
rect 14197 26877 14231 26911
rect 15669 26877 15703 26911
rect 17049 26877 17083 26911
rect 17601 26877 17635 26911
rect 18429 26877 18463 26911
rect 11897 26809 11931 26843
rect 13185 26809 13219 26843
rect 14381 26809 14415 26843
rect 6561 26741 6595 26775
rect 10885 26741 10919 26775
rect 11621 26741 11655 26775
rect 14657 26741 14691 26775
rect 16129 26741 16163 26775
rect 16589 26741 16623 26775
rect 5733 26537 5767 26571
rect 6653 26537 6687 26571
rect 8493 26537 8527 26571
rect 8677 26537 8711 26571
rect 11529 26537 11563 26571
rect 16037 26537 16071 26571
rect 17417 26537 17451 26571
rect 3617 26469 3651 26503
rect 5181 26469 5215 26503
rect 7757 26469 7791 26503
rect 16129 26469 16163 26503
rect 1593 26401 1627 26435
rect 1869 26401 1903 26435
rect 4077 26401 4111 26435
rect 4445 26401 4479 26435
rect 4905 26401 4939 26435
rect 7573 26401 7607 26435
rect 8769 26401 8803 26435
rect 9321 26401 9355 26435
rect 11345 26401 11379 26435
rect 13369 26401 13403 26435
rect 13553 26401 13587 26435
rect 14105 26401 14139 26435
rect 16681 26401 16715 26435
rect 16957 26401 16991 26435
rect 3249 26333 3283 26367
rect 9413 26333 9447 26367
rect 12173 26333 12207 26367
rect 14381 26333 14415 26367
rect 17141 26333 17175 26367
rect 3985 26265 4019 26299
rect 8125 26265 8159 26299
rect 11161 26265 11195 26299
rect 11897 26265 11931 26299
rect 12817 26265 12851 26299
rect 10057 26197 10091 26231
rect 1685 25993 1719 26027
rect 2053 25993 2087 26027
rect 2513 25993 2547 26027
rect 3433 25993 3467 26027
rect 3801 25993 3835 26027
rect 4169 25993 4203 26027
rect 7113 25993 7147 26027
rect 7665 25993 7699 26027
rect 9137 25993 9171 26027
rect 12817 25993 12851 26027
rect 15577 25993 15611 26027
rect 15853 25993 15887 26027
rect 18061 25993 18095 26027
rect 5733 25925 5767 25959
rect 8033 25925 8067 25959
rect 17509 25925 17543 25959
rect 6469 25857 6503 25891
rect 9873 25857 9907 25891
rect 12449 25857 12483 25891
rect 16865 25857 16899 25891
rect 18429 25857 18463 25891
rect 4077 25789 4111 25823
rect 4629 25789 4663 25823
rect 5181 25789 5215 25823
rect 5825 25789 5859 25823
rect 6377 25789 6411 25823
rect 8217 25789 8251 25823
rect 8401 25789 8435 25823
rect 8585 25789 8619 25823
rect 9505 25789 9539 25823
rect 9781 25789 9815 25823
rect 10149 25789 10183 25823
rect 10517 25789 10551 25823
rect 5549 25721 5583 25755
rect 11897 25721 11931 25755
rect 13001 25789 13035 25823
rect 13369 25789 13403 25823
rect 13461 25789 13495 25823
rect 14013 25789 14047 25823
rect 15669 25789 15703 25823
rect 16129 25789 16163 25823
rect 17049 25789 17083 25823
rect 17509 25789 17543 25823
rect 14473 25721 14507 25755
rect 11437 25653 11471 25687
rect 12173 25653 12207 25687
rect 12449 25653 12483 25687
rect 12633 25653 12667 25687
rect 16589 25653 16623 25687
rect 5917 25449 5951 25483
rect 8677 25449 8711 25483
rect 8953 25449 8987 25483
rect 9505 25449 9539 25483
rect 9873 25449 9907 25483
rect 12173 25449 12207 25483
rect 13645 25449 13679 25483
rect 15393 25449 15427 25483
rect 6653 25381 6687 25415
rect 4077 25313 4111 25347
rect 4629 25313 4663 25347
rect 5733 25313 5767 25347
rect 7297 25313 7331 25347
rect 7481 25313 7515 25347
rect 7941 25313 7975 25347
rect 9321 25313 9355 25347
rect 10149 25313 10183 25347
rect 10333 25313 10367 25347
rect 10885 25313 10919 25347
rect 12725 25313 12759 25347
rect 12909 25313 12943 25347
rect 13277 25313 13311 25347
rect 6285 25245 6319 25279
rect 11161 25245 11195 25279
rect 3341 25177 3375 25211
rect 7941 25177 7975 25211
rect 10425 25177 10459 25211
rect 15209 25313 15243 25347
rect 15577 25313 15611 25347
rect 15945 25313 15979 25347
rect 13829 25245 13863 25279
rect 16773 25245 16807 25279
rect 1593 25109 1627 25143
rect 3709 25109 3743 25143
rect 4629 25109 4663 25143
rect 13553 25109 13587 25143
rect 13645 25109 13679 25143
rect 17049 25109 17083 25143
rect 17417 25109 17451 25143
rect 5457 24905 5491 24939
rect 9045 24905 9079 24939
rect 15117 24905 15151 24939
rect 3893 24837 3927 24871
rect 17509 24837 17543 24871
rect 1685 24769 1719 24803
rect 3525 24769 3559 24803
rect 6469 24769 6503 24803
rect 8033 24769 8067 24803
rect 9505 24769 9539 24803
rect 10149 24769 10183 24803
rect 14749 24769 14783 24803
rect 15577 24769 15611 24803
rect 16589 24769 16623 24803
rect 16773 24769 16807 24803
rect 1409 24701 1443 24735
rect 4077 24701 4111 24735
rect 4353 24701 4387 24735
rect 6745 24701 6779 24735
rect 7481 24701 7515 24735
rect 8125 24701 8159 24735
rect 8493 24701 8527 24735
rect 10241 24701 10275 24735
rect 10517 24701 10551 24735
rect 13829 24701 13863 24735
rect 14197 24701 14231 24735
rect 15669 24701 15703 24735
rect 16129 24701 16163 24735
rect 17049 24701 17083 24735
rect 17509 24701 17543 24735
rect 3065 24633 3099 24667
rect 7297 24633 7331 24667
rect 13185 24633 13219 24667
rect 6009 24565 6043 24599
rect 6561 24565 6595 24599
rect 11621 24565 11655 24599
rect 12541 24565 12575 24599
rect 12909 24565 12943 24599
rect 13921 24565 13955 24599
rect 15853 24565 15887 24599
rect 1685 24361 1719 24395
rect 4997 24361 5031 24395
rect 5917 24361 5951 24395
rect 7113 24361 7147 24395
rect 7849 24361 7883 24395
rect 8309 24361 8343 24395
rect 10333 24361 10367 24395
rect 13829 24361 13863 24395
rect 14197 24361 14231 24395
rect 16681 24361 16715 24395
rect 17417 24361 17451 24395
rect 4537 24293 4571 24327
rect 11529 24293 11563 24327
rect 13461 24293 13495 24327
rect 2789 24225 2823 24259
rect 5181 24225 5215 24259
rect 5733 24225 5767 24259
rect 7021 24225 7055 24259
rect 9137 24225 9171 24259
rect 9597 24225 9631 24259
rect 10057 24225 10091 24259
rect 10793 24225 10827 24259
rect 11253 24225 11287 24259
rect 12909 24225 12943 24259
rect 14381 24225 14415 24259
rect 17049 24225 17083 24259
rect 2513 24157 2547 24191
rect 8401 24157 8435 24191
rect 15025 24157 15059 24191
rect 4905 24089 4939 24123
rect 6285 24089 6319 24123
rect 8677 24089 8711 24123
rect 10609 24089 10643 24123
rect 4077 24021 4111 24055
rect 5457 24021 5491 24055
rect 6653 24021 6687 24055
rect 11345 23817 11379 23851
rect 11713 23817 11747 23851
rect 14657 23817 14691 23851
rect 10149 23749 10183 23783
rect 18061 23749 18095 23783
rect 1777 23681 1811 23715
rect 5641 23681 5675 23715
rect 6745 23681 6779 23715
rect 10701 23681 10735 23715
rect 16773 23681 16807 23715
rect 17325 23681 17359 23715
rect 17785 23681 17819 23715
rect 1501 23613 1535 23647
rect 4445 23613 4479 23647
rect 4905 23613 4939 23647
rect 6561 23613 6595 23647
rect 7113 23613 7147 23647
rect 7297 23613 7331 23647
rect 7665 23613 7699 23647
rect 8033 23613 8067 23647
rect 9689 23613 9723 23647
rect 10425 23613 10459 23647
rect 12081 23613 12115 23647
rect 12909 23613 12943 23647
rect 13645 23613 13679 23647
rect 14013 23613 14047 23647
rect 14381 23613 14415 23647
rect 15761 23613 15795 23647
rect 16221 23613 16255 23647
rect 17601 23613 17635 23647
rect 3157 23545 3191 23579
rect 4813 23545 4847 23579
rect 5181 23545 5215 23579
rect 5273 23545 5307 23579
rect 6009 23545 6043 23579
rect 6377 23545 6411 23579
rect 9505 23545 9539 23579
rect 12541 23545 12575 23579
rect 13553 23545 13587 23579
rect 5089 23477 5123 23511
rect 8769 23477 8803 23511
rect 9045 23477 9079 23511
rect 15945 23477 15979 23511
rect 16589 23477 16623 23511
rect 1685 23273 1719 23307
rect 2605 23273 2639 23307
rect 2973 23273 3007 23307
rect 3709 23273 3743 23307
rect 6561 23273 6595 23307
rect 8493 23273 8527 23307
rect 8861 23273 8895 23307
rect 11069 23273 11103 23307
rect 13645 23273 13679 23307
rect 7941 23205 7975 23239
rect 15853 23205 15887 23239
rect 3893 23137 3927 23171
rect 3985 23137 4019 23171
rect 6837 23137 6871 23171
rect 7481 23137 7515 23171
rect 7665 23137 7699 23171
rect 9873 23137 9907 23171
rect 10241 23137 10275 23171
rect 10609 23137 10643 23171
rect 12449 23137 12483 23171
rect 12909 23137 12943 23171
rect 14381 23137 14415 23171
rect 14565 23137 14599 23171
rect 14749 23137 14783 23171
rect 16589 23137 16623 23171
rect 16957 23137 16991 23171
rect 17049 23137 17083 23171
rect 4261 23069 4295 23103
rect 6009 23069 6043 23103
rect 10793 23069 10827 23103
rect 13277 23069 13311 23103
rect 16497 23069 16531 23103
rect 1961 23001 1995 23035
rect 14197 23001 14231 23035
rect 5365 22933 5399 22967
rect 9505 22933 9539 22967
rect 12633 22933 12667 22967
rect 16037 22933 16071 22967
rect 17417 22933 17451 22967
rect 4261 22729 4295 22763
rect 6561 22729 6595 22763
rect 7941 22729 7975 22763
rect 9137 22729 9171 22763
rect 11069 22729 11103 22763
rect 11437 22729 11471 22763
rect 12909 22729 12943 22763
rect 15577 22729 15611 22763
rect 16497 22729 16531 22763
rect 9413 22661 9447 22695
rect 12541 22661 12575 22695
rect 13185 22661 13219 22695
rect 13645 22661 13679 22695
rect 15025 22661 15059 22695
rect 17509 22661 17543 22695
rect 4721 22593 4755 22627
rect 5457 22593 5491 22627
rect 8401 22593 8435 22627
rect 14289 22593 14323 22627
rect 14657 22593 14691 22627
rect 15301 22593 15335 22627
rect 16129 22593 16163 22627
rect 18061 22593 18095 22627
rect 4997 22525 5031 22559
rect 5181 22525 5215 22559
rect 8125 22525 8159 22559
rect 8769 22525 8803 22559
rect 9689 22525 9723 22559
rect 10425 22525 10459 22559
rect 10517 22525 10551 22559
rect 12357 22525 12391 22559
rect 13829 22525 13863 22559
rect 14197 22525 14231 22559
rect 15393 22525 15427 22559
rect 16681 22525 16715 22559
rect 17049 22525 17083 22559
rect 17601 22525 17635 22559
rect 18429 22525 18463 22559
rect 3801 22389 3835 22423
rect 4813 22389 4847 22423
rect 7113 22389 7147 22423
rect 7481 22389 7515 22423
rect 9781 22389 9815 22423
rect 12173 22389 12207 22423
rect 4537 22185 4571 22219
rect 4905 22185 4939 22219
rect 5917 22185 5951 22219
rect 6469 22185 6503 22219
rect 8493 22185 8527 22219
rect 3985 22117 4019 22151
rect 7573 22117 7607 22151
rect 9689 22117 9723 22151
rect 1869 22049 1903 22083
rect 2145 22049 2179 22083
rect 5365 22049 5399 22083
rect 5733 22049 5767 22083
rect 7021 22049 7055 22083
rect 7665 22049 7699 22083
rect 9597 22049 9631 22083
rect 10517 22049 10551 22083
rect 12909 22049 12943 22083
rect 14657 22049 14691 22083
rect 15025 22049 15059 22083
rect 15117 22049 15151 22083
rect 15577 22049 15611 22083
rect 16589 22049 16623 22083
rect 16865 22049 16899 22083
rect 8125 21981 8159 22015
rect 10241 21981 10275 22015
rect 10701 21981 10735 22015
rect 16129 21981 16163 22015
rect 17417 21981 17451 22015
rect 5181 21913 5215 21947
rect 13093 21913 13127 21947
rect 14473 21913 14507 21947
rect 16865 21913 16899 21947
rect 3433 21845 3467 21879
rect 7389 21845 7423 21879
rect 13461 21845 13495 21879
rect 13921 21845 13955 21879
rect 15945 21845 15979 21879
rect 1961 21641 1995 21675
rect 8033 21641 8067 21675
rect 8401 21641 8435 21675
rect 9965 21641 9999 21675
rect 10241 21641 10275 21675
rect 12173 21641 12207 21675
rect 12541 21641 12575 21675
rect 15669 21641 15703 21675
rect 2237 21573 2271 21607
rect 9505 21573 9539 21607
rect 13737 21573 13771 21607
rect 15945 21573 15979 21607
rect 6653 21505 6687 21539
rect 14381 21505 14415 21539
rect 14657 21505 14691 21539
rect 18061 21505 18095 21539
rect 4905 21437 4939 21471
rect 5273 21437 5307 21471
rect 6561 21437 6595 21471
rect 7297 21437 7331 21471
rect 8217 21437 8251 21471
rect 8677 21437 8711 21471
rect 11621 21437 11655 21471
rect 12633 21437 12667 21471
rect 12909 21437 12943 21471
rect 13645 21437 13679 21471
rect 13921 21437 13955 21471
rect 15761 21437 15795 21471
rect 16221 21437 16255 21471
rect 17325 21437 17359 21471
rect 17601 21437 17635 21471
rect 17785 21437 17819 21471
rect 5825 21369 5859 21403
rect 13093 21369 13127 21403
rect 16773 21369 16807 21403
rect 6193 21301 6227 21335
rect 6377 21301 6411 21335
rect 7757 21301 7791 21335
rect 11805 21301 11839 21335
rect 12817 21301 12851 21335
rect 12909 21301 12943 21335
rect 13553 21301 13587 21335
rect 15025 21301 15059 21335
rect 16589 21301 16623 21335
rect 3893 21097 3927 21131
rect 6285 21097 6319 21131
rect 8217 21097 8251 21131
rect 13185 21097 13219 21131
rect 13829 21097 13863 21131
rect 14197 21097 14231 21131
rect 17785 21097 17819 21131
rect 5917 21029 5951 21063
rect 6653 21029 6687 21063
rect 8769 21029 8803 21063
rect 15209 21029 15243 21063
rect 15945 21029 15979 21063
rect 17141 21029 17175 21063
rect 1409 20961 1443 20995
rect 1685 20961 1719 20995
rect 3801 20961 3835 20995
rect 4077 20961 4111 20995
rect 5825 20961 5859 20995
rect 7113 20961 7147 20995
rect 7481 20961 7515 20995
rect 7665 20961 7699 20995
rect 7941 20961 7975 20995
rect 8861 20961 8895 20995
rect 13277 20961 13311 20995
rect 15117 20961 15151 20995
rect 16037 20961 16071 20995
rect 16405 20961 16439 20995
rect 16865 20961 16899 20995
rect 2973 20757 3007 20791
rect 4353 20757 4387 20791
rect 12633 20757 12667 20791
rect 13461 20757 13495 20791
rect 15577 20757 15611 20791
rect 17417 20757 17451 20791
rect 1685 20553 1719 20587
rect 3617 20553 3651 20587
rect 6101 20553 6135 20587
rect 8769 20553 8803 20587
rect 9045 20553 9079 20587
rect 13369 20553 13403 20587
rect 14749 20553 14783 20587
rect 15117 20553 15151 20587
rect 15577 20553 15611 20587
rect 16497 20553 16531 20587
rect 1961 20485 1995 20519
rect 6469 20485 6503 20519
rect 9413 20485 9447 20519
rect 17509 20485 17543 20519
rect 4353 20417 4387 20451
rect 7757 20417 7791 20451
rect 10149 20417 10183 20451
rect 12357 20417 12391 20451
rect 16773 20417 16807 20451
rect 3249 20349 3283 20383
rect 3893 20349 3927 20383
rect 4077 20349 4111 20383
rect 6837 20349 6871 20383
rect 7205 20349 7239 20383
rect 7573 20349 7607 20383
rect 8585 20349 8619 20383
rect 9873 20349 9907 20383
rect 12265 20349 12299 20383
rect 12541 20349 12575 20383
rect 12633 20349 12667 20383
rect 14197 20349 14231 20383
rect 15669 20349 15703 20383
rect 16129 20349 16163 20383
rect 17233 20349 17267 20383
rect 17509 20349 17543 20383
rect 11897 20281 11931 20315
rect 12725 20281 12759 20315
rect 13093 20281 13127 20315
rect 3709 20213 3743 20247
rect 5457 20213 5491 20247
rect 8033 20213 8067 20247
rect 8401 20213 8435 20247
rect 11437 20213 11471 20247
rect 13829 20213 13863 20247
rect 14381 20213 14415 20247
rect 15853 20213 15887 20247
rect 1593 20009 1627 20043
rect 5273 20009 5307 20043
rect 6377 20009 6411 20043
rect 7665 20009 7699 20043
rect 12173 20009 12207 20043
rect 16313 20009 16347 20043
rect 17509 20009 17543 20043
rect 3433 19873 3467 19907
rect 6653 19873 6687 19907
rect 6929 19873 6963 19907
rect 13377 19873 13411 19907
rect 15393 19873 15427 19907
rect 15761 19873 15795 19907
rect 15853 19873 15887 19907
rect 17233 19873 17267 19907
rect 3157 19805 3191 19839
rect 6837 19805 6871 19839
rect 12541 19805 12575 19839
rect 12633 19805 12667 19839
rect 13461 19805 13495 19839
rect 14749 19737 14783 19771
rect 15209 19737 15243 19771
rect 4721 19669 4755 19703
rect 6469 19669 6503 19703
rect 7113 19669 7147 19703
rect 9873 19669 9907 19703
rect 13829 19669 13863 19703
rect 14197 19669 14231 19703
rect 16865 19669 16899 19703
rect 3433 19465 3467 19499
rect 3709 19465 3743 19499
rect 6561 19465 6595 19499
rect 7113 19465 7147 19499
rect 13737 19465 13771 19499
rect 16589 19397 16623 19431
rect 1409 19329 1443 19363
rect 13001 19329 13035 19363
rect 17785 19329 17819 19363
rect 1685 19261 1719 19295
rect 4813 19261 4847 19295
rect 5089 19261 5123 19295
rect 5188 19261 5222 19295
rect 5457 19261 5491 19295
rect 7849 19261 7883 19295
rect 8125 19261 8159 19295
rect 10609 19261 10643 19295
rect 11345 19261 11379 19295
rect 12909 19261 12943 19295
rect 13277 19261 13311 19295
rect 13461 19261 13495 19295
rect 15025 19261 15059 19295
rect 15301 19261 15335 19295
rect 15853 19261 15887 19295
rect 16313 19261 16347 19295
rect 17325 19261 17359 19295
rect 17601 19261 17635 19295
rect 3065 19193 3099 19227
rect 7573 19193 7607 19227
rect 11437 19193 11471 19227
rect 12265 19193 12299 19227
rect 14197 19193 14231 19227
rect 16773 19193 16807 19227
rect 4905 19125 4939 19159
rect 7665 19125 7699 19159
rect 11805 19125 11839 19159
rect 12173 19125 12207 19159
rect 14657 19125 14691 19159
rect 15485 19125 15519 19159
rect 1593 18921 1627 18955
rect 4997 18921 5031 18955
rect 6469 18921 6503 18955
rect 12633 18921 12667 18955
rect 13001 18921 13035 18955
rect 10793 18785 10827 18819
rect 11345 18785 11379 18819
rect 12449 18785 12483 18819
rect 14197 18785 14231 18819
rect 14565 18785 14599 18819
rect 16037 18785 16071 18819
rect 16497 18785 16531 18819
rect 11529 18717 11563 18751
rect 11805 18717 11839 18751
rect 14657 18717 14691 18751
rect 15393 18717 15427 18751
rect 15853 18717 15887 18751
rect 14013 18649 14047 18683
rect 16589 18649 16623 18683
rect 5365 18581 5399 18615
rect 12265 18581 12299 18615
rect 13277 18581 13311 18615
rect 3801 18377 3835 18411
rect 8033 18377 8067 18411
rect 10885 18377 10919 18411
rect 14657 18377 14691 18411
rect 12173 18309 12207 18343
rect 12633 18309 12667 18343
rect 13645 18309 13679 18343
rect 4169 18241 4203 18275
rect 15945 18241 15979 18275
rect 4445 18173 4479 18207
rect 6377 18173 6411 18207
rect 6653 18173 6687 18207
rect 6929 18173 6963 18207
rect 10517 18173 10551 18207
rect 11437 18173 11471 18207
rect 11805 18173 11839 18207
rect 12081 18173 12115 18207
rect 13829 18173 13863 18207
rect 14197 18173 14231 18207
rect 14289 18173 14323 18207
rect 15669 18173 15703 18207
rect 16497 18173 16531 18207
rect 16865 18173 16899 18207
rect 5825 18105 5859 18139
rect 6469 18105 6503 18139
rect 13277 18105 13311 18139
rect 1685 18037 1719 18071
rect 6101 18037 6135 18071
rect 6377 18037 6411 18071
rect 15117 18037 15151 18071
rect 16221 18037 16255 18071
rect 4169 17833 4203 17867
rect 10793 17833 10827 17867
rect 11805 17833 11839 17867
rect 12265 17833 12299 17867
rect 16497 17833 16531 17867
rect 8953 17765 8987 17799
rect 15761 17765 15795 17799
rect 1501 17697 1535 17731
rect 1777 17697 1811 17731
rect 7297 17697 7331 17731
rect 11345 17697 11379 17731
rect 13645 17697 13679 17731
rect 14013 17697 14047 17731
rect 15117 17697 15151 17731
rect 3157 17629 3191 17663
rect 7573 17629 7607 17663
rect 13737 17629 13771 17663
rect 14105 17629 14139 17663
rect 12909 17561 12943 17595
rect 11529 17493 11563 17527
rect 13093 17493 13127 17527
rect 14473 17493 14507 17527
rect 14933 17493 14967 17527
rect 16129 17493 16163 17527
rect 16773 17493 16807 17527
rect 9413 17289 9447 17323
rect 11621 17289 11655 17323
rect 15025 17221 15059 17255
rect 15577 17221 15611 17255
rect 1501 17153 1535 17187
rect 1777 17153 1811 17187
rect 4721 17153 4755 17187
rect 6377 17153 6411 17187
rect 7297 17153 7331 17187
rect 9965 17153 9999 17187
rect 12817 17153 12851 17187
rect 14749 17153 14783 17187
rect 4997 17085 5031 17119
rect 9689 17085 9723 17119
rect 12449 17085 12483 17119
rect 12633 17085 12667 17119
rect 12909 17085 12943 17119
rect 13461 17085 13495 17119
rect 15761 17085 15795 17119
rect 16129 17085 16163 17119
rect 16221 17085 16255 17119
rect 3157 17017 3191 17051
rect 4537 17017 4571 17051
rect 14381 17017 14415 17051
rect 7757 16949 7791 16983
rect 11069 16949 11103 16983
rect 11989 16949 12023 16983
rect 13921 16949 13955 16983
rect 1685 16745 1719 16779
rect 1961 16745 1995 16779
rect 4721 16745 4755 16779
rect 12265 16745 12299 16779
rect 12633 16745 12667 16779
rect 13093 16745 13127 16779
rect 16129 16745 16163 16779
rect 2329 16677 2363 16711
rect 3065 16609 3099 16643
rect 4445 16609 4479 16643
rect 9689 16609 9723 16643
rect 14105 16609 14139 16643
rect 14289 16609 14323 16643
rect 14473 16609 14507 16643
rect 16129 16609 16163 16643
rect 2789 16541 2823 16575
rect 15669 16541 15703 16575
rect 13921 16473 13955 16507
rect 15301 16473 15335 16507
rect 11161 16405 11195 16439
rect 13461 16405 13495 16439
rect 3433 16201 3467 16235
rect 3893 16201 3927 16235
rect 10609 16201 10643 16235
rect 12817 16201 12851 16235
rect 14013 16201 14047 16235
rect 14381 16201 14415 16235
rect 15577 16133 15611 16167
rect 1777 16065 1811 16099
rect 4353 16065 4387 16099
rect 11253 16065 11287 16099
rect 12081 16065 12115 16099
rect 13737 16065 13771 16099
rect 1501 15997 1535 16031
rect 3157 15997 3191 16031
rect 4077 15997 4111 16031
rect 11161 15997 11195 16031
rect 11989 15997 12023 16031
rect 13093 15997 13127 16031
rect 15761 15997 15795 16031
rect 15945 15997 15979 16031
rect 16129 15997 16163 16031
rect 10977 15929 11011 15963
rect 5641 15861 5675 15895
rect 15025 15861 15059 15895
rect 16681 15861 16715 15895
rect 1593 15657 1627 15691
rect 2881 15657 2915 15691
rect 3433 15657 3467 15691
rect 8861 15657 8895 15691
rect 13461 15657 13495 15691
rect 13829 15657 13863 15691
rect 15393 15657 15427 15691
rect 11437 15589 11471 15623
rect 3525 15521 3559 15555
rect 3801 15521 3835 15555
rect 7297 15521 7331 15555
rect 10057 15521 10091 15555
rect 13001 15521 13035 15555
rect 14473 15521 14507 15555
rect 14841 15521 14875 15555
rect 16129 15521 16163 15555
rect 16497 15521 16531 15555
rect 7573 15453 7607 15487
rect 9781 15453 9815 15487
rect 14933 15453 14967 15487
rect 14289 15385 14323 15419
rect 15945 15385 15979 15419
rect 2053 15317 2087 15351
rect 5089 15317 5123 15351
rect 11805 15317 11839 15351
rect 13185 15317 13219 15351
rect 15669 15317 15703 15351
rect 16865 15317 16899 15351
rect 3617 15113 3651 15147
rect 4261 15113 4295 15147
rect 4721 15113 4755 15147
rect 6469 15113 6503 15147
rect 7389 15113 7423 15147
rect 7665 15113 7699 15147
rect 10885 15113 10919 15147
rect 13001 15113 13035 15147
rect 13737 15113 13771 15147
rect 15117 15113 15151 15147
rect 15945 15113 15979 15147
rect 11253 15045 11287 15079
rect 16405 15045 16439 15079
rect 5181 14977 5215 15011
rect 11529 14977 11563 15011
rect 12357 14977 12391 15011
rect 4905 14909 4939 14943
rect 11713 14909 11747 14943
rect 12173 14909 12207 14943
rect 14197 14909 14231 14943
rect 14473 14909 14507 14943
rect 15577 14909 15611 14943
rect 16589 14909 16623 14943
rect 16773 14909 16807 14943
rect 16957 14909 16991 14943
rect 17417 14909 17451 14943
rect 14105 14841 14139 14875
rect 9873 14773 9907 14807
rect 10241 14773 10275 14807
rect 14381 14773 14415 14807
rect 14473 14773 14507 14807
rect 14749 14773 14783 14807
rect 4905 14569 4939 14603
rect 12265 14569 12299 14603
rect 15393 14569 15427 14603
rect 11529 14501 11563 14535
rect 2329 14433 2363 14467
rect 2605 14433 2639 14467
rect 10885 14433 10919 14467
rect 3985 14365 4019 14399
rect 12725 14501 12759 14535
rect 14473 14433 14507 14467
rect 14657 14433 14691 14467
rect 14841 14433 14875 14467
rect 16405 14433 16439 14467
rect 16773 14433 16807 14467
rect 16865 14433 16899 14467
rect 15853 14365 15887 14399
rect 14289 14297 14323 14331
rect 16221 14297 16255 14331
rect 12081 14229 12115 14263
rect 12265 14229 12299 14263
rect 13001 14229 13035 14263
rect 13829 14229 13863 14263
rect 2421 14025 2455 14059
rect 5641 14025 5675 14059
rect 7297 14025 7331 14059
rect 11345 14025 11379 14059
rect 11621 14025 11655 14059
rect 14105 14025 14139 14059
rect 15485 14025 15519 14059
rect 16405 14025 16439 14059
rect 2697 13957 2731 13991
rect 6009 13889 6043 13923
rect 14473 13957 14507 13991
rect 16773 13957 16807 13991
rect 11897 13889 11931 13923
rect 5733 13821 5767 13855
rect 10793 13821 10827 13855
rect 11069 13821 11103 13855
rect 11345 13821 11379 13855
rect 12081 13821 12115 13855
rect 12541 13821 12575 13855
rect 12817 13821 12851 13855
rect 13277 13821 13311 13855
rect 13369 13821 13403 13855
rect 15025 13821 15059 13855
rect 15301 13821 15335 13855
rect 16037 13821 16071 13855
rect 16957 13821 16991 13855
rect 17141 13821 17175 13855
rect 17325 13821 17359 13855
rect 10333 13685 10367 13719
rect 11253 13685 11287 13719
rect 1685 13481 1719 13515
rect 4905 13481 4939 13515
rect 5733 13481 5767 13515
rect 12173 13481 12207 13515
rect 16497 13481 16531 13515
rect 16865 13481 16899 13515
rect 11529 13413 11563 13447
rect 2973 13345 3007 13379
rect 3249 13345 3283 13379
rect 7573 13345 7607 13379
rect 9229 13345 9263 13379
rect 10333 13345 10367 13379
rect 10885 13345 10919 13379
rect 11345 13345 11379 13379
rect 12541 13345 12575 13379
rect 12817 13345 12851 13379
rect 14473 13345 14507 13379
rect 15485 13345 15519 13379
rect 15669 13345 15703 13379
rect 4629 13277 4663 13311
rect 7849 13277 7883 13311
rect 10241 13277 10275 13311
rect 13277 13277 13311 13311
rect 13921 13277 13955 13311
rect 14749 13277 14783 13311
rect 12633 13209 12667 13243
rect 15025 13209 15059 13243
rect 9781 13141 9815 13175
rect 13645 13141 13679 13175
rect 1593 12937 1627 12971
rect 2053 12937 2087 12971
rect 3341 12937 3375 12971
rect 3801 12937 3835 12971
rect 5641 12937 5675 12971
rect 7665 12937 7699 12971
rect 14197 12937 14231 12971
rect 16589 12937 16623 12971
rect 3065 12869 3099 12903
rect 7941 12869 7975 12903
rect 10057 12869 10091 12903
rect 10425 12869 10459 12903
rect 15577 12869 15611 12903
rect 4353 12801 4387 12835
rect 9505 12801 9539 12835
rect 11805 12801 11839 12835
rect 12541 12801 12575 12835
rect 14565 12801 14599 12835
rect 16221 12801 16255 12835
rect 4077 12733 4111 12767
rect 10609 12733 10643 12767
rect 11253 12733 11287 12767
rect 11437 12733 11471 12767
rect 12909 12733 12943 12767
rect 13093 12733 13127 12767
rect 13461 12733 13495 12767
rect 15117 12733 15151 12767
rect 15761 12733 15795 12767
rect 16129 12733 16163 12767
rect 17325 12733 17359 12767
rect 13737 12665 13771 12699
rect 2329 12597 2363 12631
rect 12173 12597 12207 12631
rect 16957 12597 16991 12631
rect 13001 12393 13035 12427
rect 14933 12393 14967 12427
rect 3065 12325 3099 12359
rect 8493 12325 8527 12359
rect 10517 12325 10551 12359
rect 12265 12325 12299 12359
rect 1685 12257 1719 12291
rect 4537 12257 4571 12291
rect 7113 12257 7147 12291
rect 10425 12257 10459 12291
rect 11345 12257 11379 12291
rect 13277 12257 13311 12291
rect 13737 12257 13771 12291
rect 14197 12257 14231 12291
rect 14473 12257 14507 12291
rect 16589 12257 16623 12291
rect 16773 12257 16807 12291
rect 16957 12257 16991 12291
rect 1409 12189 1443 12223
rect 4261 12189 4295 12223
rect 6837 12189 6871 12223
rect 10057 12189 10091 12223
rect 11069 12189 11103 12223
rect 11529 12189 11563 12223
rect 13829 12189 13863 12223
rect 15669 12189 15703 12223
rect 16405 12121 16439 12155
rect 4077 12053 4111 12087
rect 5825 12053 5859 12087
rect 11805 12053 11839 12087
rect 12725 12053 12759 12087
rect 15945 12053 15979 12087
rect 2973 11849 3007 11883
rect 3801 11849 3835 11883
rect 5917 11849 5951 11883
rect 8493 11849 8527 11883
rect 10517 11849 10551 11883
rect 14657 11849 14691 11883
rect 16957 11849 16991 11883
rect 13645 11781 13679 11815
rect 16497 11781 16531 11815
rect 1685 11713 1719 11747
rect 11069 11713 11103 11747
rect 12909 11713 12943 11747
rect 1409 11645 1443 11679
rect 4353 11645 4387 11679
rect 4629 11645 4663 11679
rect 7113 11645 7147 11679
rect 7389 11645 7423 11679
rect 10149 11645 10183 11679
rect 11253 11645 11287 11679
rect 11345 11645 11379 11679
rect 11713 11645 11747 11679
rect 12265 11645 12299 11679
rect 13829 11645 13863 11679
rect 14197 11645 14231 11679
rect 14289 11645 14323 11679
rect 15761 11645 15795 11679
rect 15945 11645 15979 11679
rect 16405 11645 16439 11679
rect 3433 11509 3467 11543
rect 6561 11509 6595 11543
rect 6929 11509 6963 11543
rect 10885 11509 10919 11543
rect 13277 11509 13311 11543
rect 15117 11509 15151 11543
rect 17325 11509 17359 11543
rect 8125 11305 8159 11339
rect 12265 11305 12299 11339
rect 14565 11305 14599 11339
rect 16129 11305 16163 11339
rect 16589 11305 16623 11339
rect 5825 11237 5859 11271
rect 9965 11237 9999 11271
rect 11805 11237 11839 11271
rect 1777 11169 1811 11203
rect 4445 11169 4479 11203
rect 10057 11169 10091 11203
rect 10701 11169 10735 11203
rect 10793 11169 10827 11203
rect 11345 11169 11379 11203
rect 12449 11169 12483 11203
rect 12817 11169 12851 11203
rect 13185 11169 13219 11203
rect 13829 11169 13863 11203
rect 14933 11169 14967 11203
rect 15669 11169 15703 11203
rect 15761 11169 15795 11203
rect 1501 11101 1535 11135
rect 4169 11101 4203 11135
rect 14197 11101 14231 11135
rect 14841 11101 14875 11135
rect 7205 11033 7239 11067
rect 7573 11033 7607 11067
rect 9597 11033 9631 11067
rect 3065 10965 3099 10999
rect 4077 10965 4111 10999
rect 10149 10965 10183 10999
rect 13645 10965 13679 10999
rect 3341 10761 3375 10795
rect 3801 10761 3835 10795
rect 5917 10761 5951 10795
rect 9137 10761 9171 10795
rect 11621 10761 11655 10795
rect 12081 10761 12115 10795
rect 12541 10761 12575 10795
rect 14749 10761 14783 10795
rect 16589 10693 16623 10727
rect 1685 10625 1719 10659
rect 3065 10625 3099 10659
rect 4629 10625 4663 10659
rect 8769 10625 8803 10659
rect 13921 10625 13955 10659
rect 15577 10625 15611 10659
rect 15853 10625 15887 10659
rect 1409 10557 1443 10591
rect 4353 10557 4387 10591
rect 8033 10557 8067 10591
rect 8217 10557 8251 10591
rect 8350 10557 8384 10591
rect 9689 10557 9723 10591
rect 9965 10557 9999 10591
rect 11345 10557 11379 10591
rect 13185 10557 13219 10591
rect 13553 10557 13587 10591
rect 13829 10557 13863 10591
rect 14197 10557 14231 10591
rect 16037 10557 16071 10591
rect 16497 10557 16531 10591
rect 7573 10489 7607 10523
rect 9413 10489 9447 10523
rect 7941 10421 7975 10455
rect 15025 10421 15059 10455
rect 4353 10217 4387 10251
rect 11345 10217 11379 10251
rect 12265 10217 12299 10251
rect 12725 10217 12759 10251
rect 14841 10217 14875 10251
rect 16405 10217 16439 10251
rect 16773 10217 16807 10251
rect 3157 10149 3191 10183
rect 4077 10149 4111 10183
rect 4721 10149 4755 10183
rect 7941 10149 7975 10183
rect 8493 10149 8527 10183
rect 1777 10081 1811 10115
rect 8033 10081 8067 10115
rect 9597 10081 9631 10115
rect 12909 10081 12943 10115
rect 14013 10081 14047 10115
rect 14473 10081 14507 10115
rect 15301 10081 15335 10115
rect 15577 10081 15611 10115
rect 1501 10013 1535 10047
rect 9321 10013 9355 10047
rect 7757 9877 7791 9911
rect 10885 9877 10919 9911
rect 11897 9877 11931 9911
rect 13093 9877 13127 9911
rect 13369 9877 13403 9911
rect 13829 9877 13863 9911
rect 16037 9877 16071 9911
rect 2053 9673 2087 9707
rect 2329 9673 2363 9707
rect 8125 9673 8159 9707
rect 11253 9673 11287 9707
rect 12909 9673 12943 9707
rect 13277 9673 13311 9707
rect 13461 9673 13495 9707
rect 1685 9605 1719 9639
rect 9413 9605 9447 9639
rect 14565 9605 14599 9639
rect 16589 9605 16623 9639
rect 9045 9537 9079 9571
rect 10701 9537 10735 9571
rect 14197 9537 14231 9571
rect 17693 9537 17727 9571
rect 7849 9469 7883 9503
rect 11437 9469 11471 9503
rect 11529 9469 11563 9503
rect 12173 9469 12207 9503
rect 12449 9469 12483 9503
rect 13737 9469 13771 9503
rect 14841 9469 14875 9503
rect 15485 9469 15519 9503
rect 17233 9469 17267 9503
rect 17601 9469 17635 9503
rect 13645 9401 13679 9435
rect 15853 9401 15887 9435
rect 16773 9401 16807 9435
rect 8585 9333 8619 9367
rect 10057 9333 10091 9367
rect 11069 9333 11103 9367
rect 16313 9333 16347 9367
rect 1593 9129 1627 9163
rect 1961 9129 1995 9163
rect 11805 9129 11839 9163
rect 13829 9129 13863 9163
rect 14197 9129 14231 9163
rect 11161 9061 11195 9095
rect 11529 9061 11563 9095
rect 15669 9061 15703 9095
rect 16221 9061 16255 9095
rect 9505 8993 9539 9027
rect 9781 8993 9815 9027
rect 12633 8993 12667 9027
rect 13001 8993 13035 9027
rect 13277 8993 13311 9027
rect 14841 8993 14875 9027
rect 15209 8993 15243 9027
rect 16313 8993 16347 9027
rect 15301 8925 15335 8959
rect 13277 8857 13311 8891
rect 14657 8857 14691 8891
rect 16037 8789 16071 8823
rect 9505 8585 9539 8619
rect 11345 8585 11379 8619
rect 11529 8585 11563 8619
rect 13185 8585 13219 8619
rect 14473 8585 14507 8619
rect 15117 8585 15151 8619
rect 16589 8585 16623 8619
rect 13921 8517 13955 8551
rect 15577 8517 15611 8551
rect 8769 8449 8803 8483
rect 10609 8449 10643 8483
rect 10977 8449 11011 8483
rect 9137 8381 9171 8415
rect 10517 8381 10551 8415
rect 11529 8381 11563 8415
rect 12081 8381 12115 8415
rect 12357 8381 12391 8415
rect 12725 8381 12759 8415
rect 15761 8381 15795 8415
rect 15945 8381 15979 8415
rect 16129 8381 16163 8415
rect 13553 8313 13587 8347
rect 16957 8313 16991 8347
rect 11529 8041 11563 8075
rect 14197 8041 14231 8075
rect 11161 7973 11195 8007
rect 8769 7905 8803 7939
rect 9045 7905 9079 7939
rect 13277 7905 13311 7939
rect 13461 7905 13495 7939
rect 14289 7905 14323 7939
rect 14841 7905 14875 7939
rect 15485 7905 15519 7939
rect 15853 7905 15887 7939
rect 12449 7837 12483 7871
rect 13001 7837 13035 7871
rect 15025 7837 15059 7871
rect 16405 7837 16439 7871
rect 13737 7769 13771 7803
rect 10333 7701 10367 7735
rect 9137 7497 9171 7531
rect 10885 7497 10919 7531
rect 12541 7497 12575 7531
rect 12817 7497 12851 7531
rect 8769 7429 8803 7463
rect 10609 7361 10643 7395
rect 12081 7361 12115 7395
rect 13093 7361 13127 7395
rect 15025 7361 15059 7395
rect 16497 7361 16531 7395
rect 5641 7293 5675 7327
rect 5917 7293 5951 7327
rect 11161 7293 11195 7327
rect 11989 7293 12023 7327
rect 13369 7293 13403 7327
rect 13829 7293 13863 7327
rect 14105 7293 14139 7327
rect 15393 7293 15427 7327
rect 15761 7293 15795 7327
rect 16221 7293 16255 7327
rect 7297 7225 7331 7259
rect 11253 7225 11287 7259
rect 14473 7225 14507 7259
rect 5549 7157 5583 7191
rect 5733 6953 5767 6987
rect 12725 6953 12759 6987
rect 13093 6953 13127 6987
rect 10149 6817 10183 6851
rect 11529 6817 11563 6851
rect 13185 6817 13219 6851
rect 13737 6817 13771 6851
rect 14381 6817 14415 6851
rect 14841 6817 14875 6851
rect 16589 6817 16623 6851
rect 16957 6817 16991 6851
rect 9873 6749 9907 6783
rect 13921 6749 13955 6783
rect 17049 6749 17083 6783
rect 12173 6681 12207 6715
rect 15761 6681 15795 6715
rect 16405 6681 16439 6715
rect 17417 6681 17451 6715
rect 15393 6613 15427 6647
rect 9965 6409 9999 6443
rect 10241 6409 10275 6443
rect 10885 6409 10919 6443
rect 11345 6409 11379 6443
rect 13185 6409 13219 6443
rect 15025 6409 15059 6443
rect 15853 6409 15887 6443
rect 16221 6409 16255 6443
rect 16589 6409 16623 6443
rect 13645 6341 13679 6375
rect 14749 6341 14783 6375
rect 17049 6341 17083 6375
rect 11621 6273 11655 6307
rect 12449 6273 12483 6307
rect 11529 6205 11563 6239
rect 12357 6205 12391 6239
rect 13829 6205 13863 6239
rect 14013 6205 14047 6239
rect 14197 6205 14231 6239
rect 17233 6205 17267 6239
rect 17417 6205 17451 6239
rect 17601 6205 17635 6239
rect 12909 6069 12943 6103
rect 11713 5865 11747 5899
rect 12173 5865 12207 5899
rect 13829 5865 13863 5899
rect 14289 5865 14323 5899
rect 16037 5865 16071 5899
rect 17417 5865 17451 5899
rect 8953 5797 8987 5831
rect 13185 5797 13219 5831
rect 13553 5797 13587 5831
rect 15301 5797 15335 5831
rect 2145 5729 2179 5763
rect 2421 5729 2455 5763
rect 3801 5729 3835 5763
rect 7573 5729 7607 5763
rect 9781 5729 9815 5763
rect 10057 5729 10091 5763
rect 12541 5729 12575 5763
rect 14657 5729 14691 5763
rect 16589 5729 16623 5763
rect 16957 5729 16991 5763
rect 17049 5729 17083 5763
rect 7297 5661 7331 5695
rect 11437 5661 11471 5695
rect 16405 5593 16439 5627
rect 2513 5321 2547 5355
rect 7757 5321 7791 5355
rect 10241 5321 10275 5355
rect 12541 5321 12575 5355
rect 13185 5321 13219 5355
rect 16957 5321 16991 5355
rect 13461 5253 13495 5287
rect 15577 5253 15611 5287
rect 16681 5253 16715 5287
rect 14013 5185 14047 5219
rect 15117 5185 15151 5219
rect 16221 5185 16255 5219
rect 2145 5117 2179 5151
rect 13921 5117 13955 5151
rect 14197 5117 14231 5151
rect 15761 5117 15795 5151
rect 16129 5117 16163 5151
rect 7297 4981 7331 5015
rect 9873 4981 9907 5015
rect 14657 4981 14691 5015
rect 1685 4777 1719 4811
rect 13737 4777 13771 4811
rect 14105 4777 14139 4811
rect 16773 4777 16807 4811
rect 15393 4709 15427 4743
rect 15761 4709 15795 4743
rect 14473 4641 14507 4675
rect 14749 4641 14783 4675
rect 15945 4641 15979 4675
rect 14289 4505 14323 4539
rect 14197 4233 14231 4267
rect 14565 4233 14599 4267
rect 15853 4233 15887 4267
rect 1409 4097 1443 4131
rect 1685 4097 1719 4131
rect 3065 4097 3099 4131
rect 10241 4097 10275 4131
rect 11897 4097 11931 4131
rect 10517 4029 10551 4063
rect 10057 3893 10091 3927
rect 1685 3689 1719 3723
rect 10241 3689 10275 3723
rect 9229 2601 9263 2635
rect 10057 2465 10091 2499
rect 9781 2397 9815 2431
rect 9505 2261 9539 2295
rect 11345 2261 11379 2295
<< metal1 >>
rect 3786 78616 3792 78668
rect 3844 78656 3850 78668
rect 4798 78656 4804 78668
rect 3844 78628 4804 78656
rect 3844 78616 3850 78628
rect 4798 78616 4804 78628
rect 4856 78616 4862 78668
rect 1104 77818 18860 77840
rect 1104 77766 7648 77818
rect 7700 77766 7712 77818
rect 7764 77766 7776 77818
rect 7828 77766 7840 77818
rect 7892 77766 14315 77818
rect 14367 77766 14379 77818
rect 14431 77766 14443 77818
rect 14495 77766 14507 77818
rect 14559 77766 18860 77818
rect 1104 77744 18860 77766
rect 3234 77460 3240 77512
rect 3292 77500 3298 77512
rect 15930 77500 15936 77512
rect 3292 77472 15936 77500
rect 3292 77460 3298 77472
rect 15930 77460 15936 77472
rect 15988 77460 15994 77512
rect 3326 77392 3332 77444
rect 3384 77432 3390 77444
rect 16022 77432 16028 77444
rect 3384 77404 16028 77432
rect 3384 77392 3390 77404
rect 16022 77392 16028 77404
rect 16080 77392 16086 77444
rect 1104 77274 18860 77296
rect 1104 77222 4315 77274
rect 4367 77222 4379 77274
rect 4431 77222 4443 77274
rect 4495 77222 4507 77274
rect 4559 77222 10982 77274
rect 11034 77222 11046 77274
rect 11098 77222 11110 77274
rect 11162 77222 11174 77274
rect 11226 77222 17648 77274
rect 17700 77222 17712 77274
rect 17764 77222 17776 77274
rect 17828 77222 17840 77274
rect 17892 77222 18860 77274
rect 1104 77200 18860 77222
rect 1104 76730 18860 76752
rect 1104 76678 7648 76730
rect 7700 76678 7712 76730
rect 7764 76678 7776 76730
rect 7828 76678 7840 76730
rect 7892 76678 14315 76730
rect 14367 76678 14379 76730
rect 14431 76678 14443 76730
rect 14495 76678 14507 76730
rect 14559 76678 18860 76730
rect 1104 76656 18860 76678
rect 1104 76186 18860 76208
rect 1104 76134 4315 76186
rect 4367 76134 4379 76186
rect 4431 76134 4443 76186
rect 4495 76134 4507 76186
rect 4559 76134 10982 76186
rect 11034 76134 11046 76186
rect 11098 76134 11110 76186
rect 11162 76134 11174 76186
rect 11226 76134 17648 76186
rect 17700 76134 17712 76186
rect 17764 76134 17776 76186
rect 17828 76134 17840 76186
rect 17892 76134 18860 76186
rect 1104 76112 18860 76134
rect 1104 75642 18860 75664
rect 1104 75590 7648 75642
rect 7700 75590 7712 75642
rect 7764 75590 7776 75642
rect 7828 75590 7840 75642
rect 7892 75590 14315 75642
rect 14367 75590 14379 75642
rect 14431 75590 14443 75642
rect 14495 75590 14507 75642
rect 14559 75590 18860 75642
rect 1104 75568 18860 75590
rect 4154 75420 4160 75472
rect 4212 75460 4218 75472
rect 4341 75463 4399 75469
rect 4341 75460 4353 75463
rect 4212 75432 4353 75460
rect 4212 75420 4218 75432
rect 4341 75429 4353 75432
rect 4387 75429 4399 75463
rect 4341 75423 4399 75429
rect 5166 75392 5172 75404
rect 5127 75364 5172 75392
rect 5166 75352 5172 75364
rect 5224 75352 5230 75404
rect 7098 75392 7104 75404
rect 7059 75364 7104 75392
rect 7098 75352 7104 75364
rect 7156 75352 7162 75404
rect 4890 75324 4896 75336
rect 4851 75296 4896 75324
rect 4890 75284 4896 75296
rect 4948 75284 4954 75336
rect 5353 75327 5411 75333
rect 5353 75293 5365 75327
rect 5399 75293 5411 75327
rect 5353 75287 5411 75293
rect 3970 75216 3976 75268
rect 4028 75256 4034 75268
rect 5368 75256 5396 75287
rect 4028 75228 5396 75256
rect 4028 75216 4034 75228
rect 2225 75191 2283 75197
rect 2225 75157 2237 75191
rect 2271 75188 2283 75191
rect 2958 75188 2964 75200
rect 2271 75160 2964 75188
rect 2271 75157 2283 75160
rect 2225 75151 2283 75157
rect 2958 75148 2964 75160
rect 3016 75148 3022 75200
rect 4154 75188 4160 75200
rect 4115 75160 4160 75188
rect 4154 75148 4160 75160
rect 4212 75148 4218 75200
rect 7282 75188 7288 75200
rect 7243 75160 7288 75188
rect 7282 75148 7288 75160
rect 7340 75148 7346 75200
rect 1104 75098 18860 75120
rect 1104 75046 4315 75098
rect 4367 75046 4379 75098
rect 4431 75046 4443 75098
rect 4495 75046 4507 75098
rect 4559 75046 10982 75098
rect 11034 75046 11046 75098
rect 11098 75046 11110 75098
rect 11162 75046 11174 75098
rect 11226 75046 17648 75098
rect 17700 75046 17712 75098
rect 17764 75046 17776 75098
rect 17828 75046 17840 75098
rect 17892 75046 18860 75098
rect 1104 75024 18860 75046
rect 3513 74987 3571 74993
rect 3513 74953 3525 74987
rect 3559 74984 3571 74987
rect 5166 74984 5172 74996
rect 3559 74956 5172 74984
rect 3559 74953 3571 74956
rect 3513 74947 3571 74953
rect 5166 74944 5172 74956
rect 5224 74984 5230 74996
rect 5813 74987 5871 74993
rect 5813 74984 5825 74987
rect 5224 74956 5825 74984
rect 5224 74944 5230 74956
rect 5813 74953 5825 74956
rect 5859 74953 5871 74987
rect 7006 74984 7012 74996
rect 6967 74956 7012 74984
rect 5813 74947 5871 74953
rect 7006 74944 7012 74956
rect 7064 74944 7070 74996
rect 2041 74919 2099 74925
rect 2041 74885 2053 74919
rect 2087 74916 2099 74919
rect 2087 74888 3188 74916
rect 2087 74885 2099 74888
rect 2041 74879 2099 74885
rect 2130 74848 2136 74860
rect 2091 74820 2136 74848
rect 2130 74808 2136 74820
rect 2188 74808 2194 74860
rect 2222 74740 2228 74792
rect 2280 74780 2286 74792
rect 2685 74783 2743 74789
rect 2685 74780 2697 74783
rect 2280 74752 2697 74780
rect 2280 74740 2286 74752
rect 2685 74749 2697 74752
rect 2731 74749 2743 74783
rect 2958 74780 2964 74792
rect 2871 74752 2964 74780
rect 2685 74743 2743 74749
rect 2958 74740 2964 74752
rect 3016 74740 3022 74792
rect 3160 74789 3188 74888
rect 3881 74851 3939 74857
rect 3881 74817 3893 74851
rect 3927 74848 3939 74851
rect 4890 74848 4896 74860
rect 3927 74820 4896 74848
rect 3927 74817 3939 74820
rect 3881 74811 3939 74817
rect 4890 74808 4896 74820
rect 4948 74808 4954 74860
rect 3145 74783 3203 74789
rect 3145 74749 3157 74783
rect 3191 74780 3203 74783
rect 3970 74780 3976 74792
rect 3191 74752 3976 74780
rect 3191 74749 3203 74752
rect 3145 74743 3203 74749
rect 3970 74740 3976 74752
rect 4028 74740 4034 74792
rect 4154 74740 4160 74792
rect 4212 74780 4218 74792
rect 4433 74783 4491 74789
rect 4433 74780 4445 74783
rect 4212 74752 4445 74780
rect 4212 74740 4218 74752
rect 4433 74749 4445 74752
rect 4479 74749 4491 74783
rect 4433 74743 4491 74749
rect 4709 74783 4767 74789
rect 4709 74749 4721 74783
rect 4755 74780 4767 74783
rect 4982 74780 4988 74792
rect 4755 74752 4988 74780
rect 4755 74749 4767 74752
rect 4709 74743 4767 74749
rect 2976 74712 3004 74740
rect 4062 74712 4068 74724
rect 2976 74684 4068 74712
rect 4062 74672 4068 74684
rect 4120 74672 4126 74724
rect 3970 74604 3976 74656
rect 4028 74644 4034 74656
rect 4249 74647 4307 74653
rect 4249 74644 4261 74647
rect 4028 74616 4261 74644
rect 4028 74604 4034 74616
rect 4249 74613 4261 74616
rect 4295 74613 4307 74647
rect 4448 74644 4476 74743
rect 4982 74740 4988 74752
rect 5040 74740 5046 74792
rect 6457 74783 6515 74789
rect 6457 74749 6469 74783
rect 6503 74780 6515 74783
rect 6730 74780 6736 74792
rect 6503 74752 6736 74780
rect 6503 74749 6515 74752
rect 6457 74743 6515 74749
rect 6730 74740 6736 74752
rect 6788 74780 6794 74792
rect 6917 74783 6975 74789
rect 6917 74780 6929 74783
rect 6788 74752 6929 74780
rect 6788 74740 6794 74752
rect 6917 74749 6929 74752
rect 6963 74749 6975 74783
rect 6917 74743 6975 74749
rect 7469 74783 7527 74789
rect 7469 74749 7481 74783
rect 7515 74749 7527 74783
rect 7469 74743 7527 74749
rect 6825 74715 6883 74721
rect 6825 74681 6837 74715
rect 6871 74712 6883 74715
rect 7374 74712 7380 74724
rect 6871 74684 7380 74712
rect 6871 74681 6883 74684
rect 6825 74675 6883 74681
rect 7374 74672 7380 74684
rect 7432 74712 7438 74724
rect 7484 74712 7512 74743
rect 7432 74684 7512 74712
rect 7432 74672 7438 74684
rect 5442 74644 5448 74656
rect 4448 74616 5448 74644
rect 4249 74607 4307 74613
rect 5442 74604 5448 74616
rect 5500 74604 5506 74656
rect 1104 74554 18860 74576
rect 1104 74502 7648 74554
rect 7700 74502 7712 74554
rect 7764 74502 7776 74554
rect 7828 74502 7840 74554
rect 7892 74502 14315 74554
rect 14367 74502 14379 74554
rect 14431 74502 14443 74554
rect 14495 74502 14507 74554
rect 14559 74502 18860 74554
rect 1104 74480 18860 74502
rect 4154 74400 4160 74452
rect 4212 74440 4218 74452
rect 4249 74443 4307 74449
rect 4249 74440 4261 74443
rect 4212 74412 4261 74440
rect 4212 74400 4218 74412
rect 4249 74409 4261 74412
rect 4295 74409 4307 74443
rect 4249 74403 4307 74409
rect 5534 74400 5540 74452
rect 5592 74440 5598 74452
rect 6086 74440 6092 74452
rect 5592 74412 6092 74440
rect 5592 74400 5598 74412
rect 6086 74400 6092 74412
rect 6144 74440 6150 74452
rect 6457 74443 6515 74449
rect 6457 74440 6469 74443
rect 6144 74412 6469 74440
rect 6144 74400 6150 74412
rect 6457 74409 6469 74412
rect 6503 74409 6515 74443
rect 6457 74403 6515 74409
rect 5169 74375 5227 74381
rect 5169 74341 5181 74375
rect 5215 74372 5227 74375
rect 5902 74372 5908 74384
rect 5215 74344 5908 74372
rect 5215 74341 5227 74344
rect 5169 74335 5227 74341
rect 5902 74332 5908 74344
rect 5960 74332 5966 74384
rect 7374 74332 7380 74384
rect 7432 74372 7438 74384
rect 7653 74375 7711 74381
rect 7653 74372 7665 74375
rect 7432 74344 7665 74372
rect 7432 74332 7438 74344
rect 7653 74341 7665 74344
rect 7699 74372 7711 74375
rect 8294 74372 8300 74384
rect 7699 74344 8300 74372
rect 7699 74341 7711 74344
rect 7653 74335 7711 74341
rect 8294 74332 8300 74344
rect 8352 74332 8358 74384
rect 2774 74264 2780 74316
rect 2832 74304 2838 74316
rect 2961 74307 3019 74313
rect 2961 74304 2973 74307
rect 2832 74276 2973 74304
rect 2832 74264 2838 74276
rect 2961 74273 2973 74276
rect 3007 74273 3019 74307
rect 5350 74304 5356 74316
rect 5311 74276 5356 74304
rect 2961 74267 3019 74273
rect 5350 74264 5356 74276
rect 5408 74264 5414 74316
rect 7742 74304 7748 74316
rect 7703 74276 7748 74304
rect 7742 74264 7748 74276
rect 7800 74264 7806 74316
rect 2130 74196 2136 74248
rect 2188 74236 2194 74248
rect 2682 74236 2688 74248
rect 2188 74208 2688 74236
rect 2188 74196 2194 74208
rect 2682 74196 2688 74208
rect 2740 74196 2746 74248
rect 4982 74236 4988 74248
rect 4895 74208 4988 74236
rect 4982 74196 4988 74208
rect 5040 74236 5046 74248
rect 7760 74236 7788 74264
rect 5040 74208 7788 74236
rect 5040 74196 5046 74208
rect 4709 74171 4767 74177
rect 4709 74137 4721 74171
rect 4755 74168 4767 74171
rect 5074 74168 5080 74180
rect 4755 74140 5080 74168
rect 4755 74137 4767 74140
rect 4709 74131 4767 74137
rect 5074 74128 5080 74140
rect 5132 74128 5138 74180
rect 6454 74128 6460 74180
rect 6512 74168 6518 74180
rect 7009 74171 7067 74177
rect 7009 74168 7021 74171
rect 6512 74140 7021 74168
rect 6512 74128 6518 74140
rect 7009 74137 7021 74140
rect 7055 74168 7067 74171
rect 7098 74168 7104 74180
rect 7055 74140 7104 74168
rect 7055 74137 7067 74140
rect 7009 74131 7067 74137
rect 7098 74128 7104 74140
rect 7156 74128 7162 74180
rect 2222 74100 2228 74112
rect 2183 74072 2228 74100
rect 2222 74060 2228 74072
rect 2280 74060 2286 74112
rect 5442 74100 5448 74112
rect 5403 74072 5448 74100
rect 5442 74060 5448 74072
rect 5500 74060 5506 74112
rect 6181 74103 6239 74109
rect 6181 74069 6193 74103
rect 6227 74100 6239 74103
rect 6546 74100 6552 74112
rect 6227 74072 6552 74100
rect 6227 74069 6239 74072
rect 6181 74063 6239 74069
rect 6546 74060 6552 74072
rect 6604 74060 6610 74112
rect 10137 74103 10195 74109
rect 10137 74069 10149 74103
rect 10183 74100 10195 74103
rect 10594 74100 10600 74112
rect 10183 74072 10600 74100
rect 10183 74069 10195 74072
rect 10137 74063 10195 74069
rect 10594 74060 10600 74072
rect 10652 74060 10658 74112
rect 1104 74010 18860 74032
rect 1104 73958 4315 74010
rect 4367 73958 4379 74010
rect 4431 73958 4443 74010
rect 4495 73958 4507 74010
rect 4559 73958 10982 74010
rect 11034 73958 11046 74010
rect 11098 73958 11110 74010
rect 11162 73958 11174 74010
rect 11226 73958 17648 74010
rect 17700 73958 17712 74010
rect 17764 73958 17776 74010
rect 17828 73958 17840 74010
rect 17892 73958 18860 74010
rect 1104 73936 18860 73958
rect 2130 73896 2136 73908
rect 2091 73868 2136 73896
rect 2130 73856 2136 73868
rect 2188 73856 2194 73908
rect 2222 73856 2228 73908
rect 2280 73896 2286 73908
rect 2869 73899 2927 73905
rect 2869 73896 2881 73899
rect 2280 73868 2881 73896
rect 2280 73856 2286 73868
rect 2869 73865 2881 73868
rect 2915 73865 2927 73899
rect 2869 73859 2927 73865
rect 3513 73831 3571 73837
rect 3513 73797 3525 73831
rect 3559 73828 3571 73831
rect 5902 73828 5908 73840
rect 3559 73800 5908 73828
rect 3559 73797 3571 73800
rect 3513 73791 3571 73797
rect 2501 73695 2559 73701
rect 2501 73661 2513 73695
rect 2547 73692 2559 73695
rect 2774 73692 2780 73704
rect 2547 73664 2780 73692
rect 2547 73661 2559 73664
rect 2501 73655 2559 73661
rect 2774 73652 2780 73664
rect 2832 73652 2838 73704
rect 2593 73627 2651 73633
rect 2593 73593 2605 73627
rect 2639 73624 2651 73627
rect 3528 73624 3556 73791
rect 5902 73788 5908 73800
rect 5960 73788 5966 73840
rect 3881 73763 3939 73769
rect 3881 73729 3893 73763
rect 3927 73760 3939 73763
rect 6086 73760 6092 73772
rect 3927 73732 5304 73760
rect 6047 73732 6092 73760
rect 3927 73729 3939 73732
rect 3881 73723 3939 73729
rect 5276 73704 5304 73732
rect 6086 73720 6092 73732
rect 6144 73720 6150 73772
rect 6365 73763 6423 73769
rect 6365 73729 6377 73763
rect 6411 73760 6423 73763
rect 6546 73760 6552 73772
rect 6411 73732 6552 73760
rect 6411 73729 6423 73732
rect 6365 73723 6423 73729
rect 6546 73720 6552 73732
rect 6604 73720 6610 73772
rect 10686 73760 10692 73772
rect 10647 73732 10692 73760
rect 10686 73720 10692 73732
rect 10744 73720 10750 73772
rect 4338 73652 4344 73704
rect 4396 73692 4402 73704
rect 4801 73695 4859 73701
rect 4801 73692 4813 73695
rect 4396 73664 4813 73692
rect 4396 73652 4402 73664
rect 4801 73661 4813 73664
rect 4847 73661 4859 73695
rect 5074 73692 5080 73704
rect 5035 73664 5080 73692
rect 4801 73655 4859 73661
rect 5074 73652 5080 73664
rect 5132 73652 5138 73704
rect 5258 73692 5264 73704
rect 5219 73664 5264 73692
rect 5258 73652 5264 73664
rect 5316 73652 5322 73704
rect 5350 73652 5356 73704
rect 5408 73692 5414 73704
rect 5629 73695 5687 73701
rect 5629 73692 5641 73695
rect 5408 73664 5641 73692
rect 5408 73652 5414 73664
rect 5629 73661 5641 73664
rect 5675 73692 5687 73695
rect 7190 73692 7196 73704
rect 5675 73664 7196 73692
rect 5675 73661 5687 73664
rect 5629 73655 5687 73661
rect 7190 73652 7196 73664
rect 7248 73652 7254 73704
rect 9306 73652 9312 73704
rect 9364 73692 9370 73704
rect 9493 73695 9551 73701
rect 9493 73692 9505 73695
rect 9364 73664 9505 73692
rect 9364 73652 9370 73664
rect 9493 73661 9505 73664
rect 9539 73692 9551 73695
rect 10045 73695 10103 73701
rect 10045 73692 10057 73695
rect 9539 73664 10057 73692
rect 9539 73661 9551 73664
rect 9493 73655 9551 73661
rect 10045 73661 10057 73664
rect 10091 73661 10103 73695
rect 10594 73692 10600 73704
rect 10555 73664 10600 73692
rect 10045 73655 10103 73661
rect 10594 73652 10600 73664
rect 10652 73652 10658 73704
rect 10781 73695 10839 73701
rect 10781 73661 10793 73695
rect 10827 73692 10839 73695
rect 11330 73692 11336 73704
rect 10827 73664 11336 73692
rect 10827 73661 10839 73664
rect 10781 73655 10839 73661
rect 4246 73624 4252 73636
rect 2639 73596 3556 73624
rect 4207 73596 4252 73624
rect 2639 73593 2651 73596
rect 2593 73587 2651 73593
rect 4246 73584 4252 73596
rect 4304 73584 4310 73636
rect 7374 73584 7380 73636
rect 7432 73624 7438 73636
rect 7742 73624 7748 73636
rect 7432 73596 7748 73624
rect 7432 73584 7438 73596
rect 7742 73584 7748 73596
rect 7800 73624 7806 73636
rect 8021 73627 8079 73633
rect 8021 73624 8033 73627
rect 7800 73596 8033 73624
rect 7800 73584 7806 73596
rect 8021 73593 8033 73596
rect 8067 73593 8079 73627
rect 8021 73587 8079 73593
rect 9953 73627 10011 73633
rect 9953 73593 9965 73627
rect 9999 73624 10011 73627
rect 10796 73624 10824 73655
rect 11330 73652 11336 73664
rect 11388 73652 11394 73704
rect 9999 73596 10824 73624
rect 9999 73593 10011 73596
rect 9953 73587 10011 73593
rect 5902 73556 5908 73568
rect 5863 73528 5908 73556
rect 5902 73516 5908 73528
rect 5960 73516 5966 73568
rect 5994 73516 6000 73568
rect 6052 73556 6058 73568
rect 7469 73559 7527 73565
rect 7469 73556 7481 73559
rect 6052 73528 7481 73556
rect 6052 73516 6058 73528
rect 7469 73525 7481 73528
rect 7515 73525 7527 73559
rect 7469 73519 7527 73525
rect 1104 73466 18860 73488
rect 1104 73414 7648 73466
rect 7700 73414 7712 73466
rect 7764 73414 7776 73466
rect 7828 73414 7840 73466
rect 7892 73414 14315 73466
rect 14367 73414 14379 73466
rect 14431 73414 14443 73466
rect 14495 73414 14507 73466
rect 14559 73414 18860 73466
rect 1104 73392 18860 73414
rect 2685 73355 2743 73361
rect 2685 73321 2697 73355
rect 2731 73352 2743 73355
rect 2774 73352 2780 73364
rect 2731 73324 2780 73352
rect 2731 73321 2743 73324
rect 2685 73315 2743 73321
rect 2774 73312 2780 73324
rect 2832 73352 2838 73364
rect 9306 73352 9312 73364
rect 2832 73324 7604 73352
rect 9267 73324 9312 73352
rect 2832 73312 2838 73324
rect 2866 73244 2872 73296
rect 2924 73284 2930 73296
rect 2961 73287 3019 73293
rect 2961 73284 2973 73287
rect 2924 73256 2973 73284
rect 2924 73244 2930 73256
rect 2961 73253 2973 73256
rect 3007 73253 3019 73287
rect 4798 73284 4804 73296
rect 4759 73256 4804 73284
rect 2961 73247 3019 73253
rect 4798 73244 4804 73256
rect 4856 73244 4862 73296
rect 6178 73244 6184 73296
rect 6236 73284 6242 73296
rect 7282 73284 7288 73296
rect 6236 73256 7288 73284
rect 6236 73244 6242 73256
rect 7282 73244 7288 73256
rect 7340 73284 7346 73296
rect 7340 73256 7420 73284
rect 7340 73244 7346 73256
rect 3789 73219 3847 73225
rect 3789 73216 3801 73219
rect 2700 73188 3801 73216
rect 2700 73160 2728 73188
rect 3789 73185 3801 73188
rect 3835 73216 3847 73219
rect 4338 73216 4344 73228
rect 3835 73188 4108 73216
rect 4299 73188 4344 73216
rect 3835 73185 3847 73188
rect 3789 73179 3847 73185
rect 2682 73108 2688 73160
rect 2740 73108 2746 73160
rect 3510 73148 3516 73160
rect 3471 73120 3516 73148
rect 3510 73108 3516 73120
rect 3568 73108 3574 73160
rect 3970 73148 3976 73160
rect 3883 73120 3976 73148
rect 3970 73108 3976 73120
rect 4028 73108 4034 73160
rect 4080 73148 4108 73188
rect 4338 73176 4344 73188
rect 4396 73176 4402 73228
rect 5353 73219 5411 73225
rect 5353 73185 5365 73219
rect 5399 73216 5411 73219
rect 5442 73216 5448 73228
rect 5399 73188 5448 73216
rect 5399 73185 5411 73188
rect 5353 73179 5411 73185
rect 5442 73176 5448 73188
rect 5500 73176 5506 73228
rect 5629 73219 5687 73225
rect 5629 73185 5641 73219
rect 5675 73216 5687 73219
rect 5994 73216 6000 73228
rect 5675 73188 6000 73216
rect 5675 73185 5687 73188
rect 5629 73179 5687 73185
rect 5994 73176 6000 73188
rect 6052 73176 6058 73228
rect 7392 73225 7420 73256
rect 6917 73219 6975 73225
rect 6917 73185 6929 73219
rect 6963 73185 6975 73219
rect 6917 73179 6975 73185
rect 7377 73219 7435 73225
rect 7377 73185 7389 73219
rect 7423 73185 7435 73219
rect 7377 73179 7435 73185
rect 4982 73148 4988 73160
rect 4080 73120 4988 73148
rect 4982 73108 4988 73120
rect 5040 73108 5046 73160
rect 5258 73108 5264 73160
rect 5316 73148 5322 73160
rect 5810 73148 5816 73160
rect 5316 73120 5816 73148
rect 5316 73108 5322 73120
rect 5810 73108 5816 73120
rect 5868 73108 5874 73160
rect 6730 73108 6736 73160
rect 6788 73148 6794 73160
rect 6932 73148 6960 73179
rect 6788 73120 6960 73148
rect 7576 73148 7604 73324
rect 9306 73312 9312 73324
rect 9364 73312 9370 73364
rect 8941 73219 8999 73225
rect 8941 73185 8953 73219
rect 8987 73216 8999 73219
rect 9214 73216 9220 73228
rect 8987 73188 9220 73216
rect 8987 73185 8999 73188
rect 8941 73179 8999 73185
rect 9214 73176 9220 73188
rect 9272 73176 9278 73228
rect 9490 73216 9496 73228
rect 9324 73188 9496 73216
rect 9033 73151 9091 73157
rect 9033 73148 9045 73151
rect 7576 73120 9045 73148
rect 6788 73108 6794 73120
rect 9033 73117 9045 73120
rect 9079 73148 9091 73151
rect 9324 73148 9352 73188
rect 9490 73176 9496 73188
rect 9548 73176 9554 73228
rect 9677 73219 9735 73225
rect 9677 73216 9689 73219
rect 9600 73188 9689 73216
rect 9600 73148 9628 73188
rect 9677 73185 9689 73188
rect 9723 73185 9735 73219
rect 10042 73216 10048 73228
rect 10003 73188 10048 73216
rect 9677 73179 9735 73185
rect 10042 73176 10048 73188
rect 10100 73176 10106 73228
rect 9079 73120 9352 73148
rect 9508 73120 9628 73148
rect 10873 73151 10931 73157
rect 9079 73117 9091 73120
rect 9033 73111 9091 73117
rect 3050 73040 3056 73092
rect 3108 73080 3114 73092
rect 3988 73080 4016 73108
rect 5074 73080 5080 73092
rect 3108 73052 5080 73080
rect 3108 73040 3114 73052
rect 5074 73040 5080 73052
rect 5132 73040 5138 73092
rect 6914 73080 6920 73092
rect 6875 73052 6920 73080
rect 6914 73040 6920 73052
rect 6972 73040 6978 73092
rect 8294 73040 8300 73092
rect 8352 73080 8358 73092
rect 9306 73080 9312 73092
rect 8352 73052 9312 73080
rect 8352 73040 8358 73052
rect 9306 73040 9312 73052
rect 9364 73080 9370 73092
rect 9508 73080 9536 73120
rect 10873 73117 10885 73151
rect 10919 73148 10931 73151
rect 11606 73148 11612 73160
rect 10919 73120 11612 73148
rect 10919 73117 10931 73120
rect 10873 73111 10931 73117
rect 11606 73108 11612 73120
rect 11664 73108 11670 73160
rect 9364 73052 9536 73080
rect 9364 73040 9370 73052
rect 4706 73012 4712 73024
rect 4667 72984 4712 73012
rect 4706 72972 4712 72984
rect 4764 72972 4770 73024
rect 6454 73012 6460 73024
rect 6415 72984 6460 73012
rect 6454 72972 6460 72984
rect 6512 72972 6518 73024
rect 8205 73015 8263 73021
rect 8205 72981 8217 73015
rect 8251 73012 8263 73015
rect 8570 73012 8576 73024
rect 8251 72984 8576 73012
rect 8251 72981 8263 72984
rect 8205 72975 8263 72981
rect 8570 72972 8576 72984
rect 8628 72972 8634 73024
rect 10870 72972 10876 73024
rect 10928 73012 10934 73024
rect 11149 73015 11207 73021
rect 11149 73012 11161 73015
rect 10928 72984 11161 73012
rect 10928 72972 10934 72984
rect 11149 72981 11161 72984
rect 11195 72981 11207 73015
rect 11149 72975 11207 72981
rect 1104 72922 18860 72944
rect 1104 72870 4315 72922
rect 4367 72870 4379 72922
rect 4431 72870 4443 72922
rect 4495 72870 4507 72922
rect 4559 72870 10982 72922
rect 11034 72870 11046 72922
rect 11098 72870 11110 72922
rect 11162 72870 11174 72922
rect 11226 72870 17648 72922
rect 17700 72870 17712 72922
rect 17764 72870 17776 72922
rect 17828 72870 17840 72922
rect 17892 72870 18860 72922
rect 1104 72848 18860 72870
rect 2682 72808 2688 72820
rect 2643 72780 2688 72808
rect 2682 72768 2688 72780
rect 2740 72768 2746 72820
rect 3050 72808 3056 72820
rect 3011 72780 3056 72808
rect 3050 72768 3056 72780
rect 3108 72768 3114 72820
rect 3878 72808 3884 72820
rect 3839 72780 3884 72808
rect 3878 72768 3884 72780
rect 3936 72768 3942 72820
rect 7006 72768 7012 72820
rect 7064 72808 7070 72820
rect 7745 72811 7803 72817
rect 7745 72808 7757 72811
rect 7064 72780 7757 72808
rect 7064 72768 7070 72780
rect 7745 72777 7757 72780
rect 7791 72777 7803 72811
rect 7745 72771 7803 72777
rect 8294 72768 8300 72820
rect 8352 72808 8358 72820
rect 8389 72811 8447 72817
rect 8389 72808 8401 72811
rect 8352 72780 8401 72808
rect 8352 72768 8358 72780
rect 8389 72777 8401 72780
rect 8435 72777 8447 72811
rect 8389 72771 8447 72777
rect 8570 72700 8576 72752
rect 8628 72740 8634 72752
rect 10870 72740 10876 72752
rect 8628 72712 10876 72740
rect 8628 72700 8634 72712
rect 10870 72700 10876 72712
rect 10928 72700 10934 72752
rect 11149 72743 11207 72749
rect 11149 72709 11161 72743
rect 11195 72740 11207 72743
rect 11330 72740 11336 72752
rect 11195 72712 11336 72740
rect 11195 72709 11207 72712
rect 11149 72703 11207 72709
rect 11330 72700 11336 72712
rect 11388 72700 11394 72752
rect 4525 72675 4583 72681
rect 4525 72641 4537 72675
rect 4571 72672 4583 72675
rect 4614 72672 4620 72684
rect 4571 72644 4620 72672
rect 4571 72641 4583 72644
rect 4525 72635 4583 72641
rect 4614 72632 4620 72644
rect 4672 72632 4678 72684
rect 4706 72632 4712 72684
rect 4764 72672 4770 72684
rect 5077 72675 5135 72681
rect 5077 72672 5089 72675
rect 4764 72644 5089 72672
rect 4764 72632 4770 72644
rect 5077 72641 5089 72644
rect 5123 72672 5135 72675
rect 5442 72672 5448 72684
rect 5123 72644 5448 72672
rect 5123 72641 5135 72644
rect 5077 72635 5135 72641
rect 5442 72632 5448 72644
rect 5500 72632 5506 72684
rect 6086 72632 6092 72684
rect 6144 72672 6150 72684
rect 6365 72675 6423 72681
rect 6365 72672 6377 72675
rect 6144 72644 6377 72672
rect 6144 72632 6150 72644
rect 6365 72641 6377 72644
rect 6411 72641 6423 72675
rect 10318 72672 10324 72684
rect 10231 72644 10324 72672
rect 6365 72635 6423 72641
rect 10318 72632 10324 72644
rect 10376 72672 10382 72684
rect 10376 72644 11836 72672
rect 10376 72632 10382 72644
rect 11808 72616 11836 72644
rect 5258 72564 5264 72616
rect 5316 72604 5322 72616
rect 5353 72607 5411 72613
rect 5353 72604 5365 72607
rect 5316 72576 5365 72604
rect 5316 72564 5322 72576
rect 5353 72573 5365 72576
rect 5399 72573 5411 72607
rect 5353 72567 5411 72573
rect 5537 72607 5595 72613
rect 5537 72573 5549 72607
rect 5583 72604 5595 72607
rect 5583 72576 5856 72604
rect 5583 72573 5595 72576
rect 5537 72567 5595 72573
rect 4433 72539 4491 72545
rect 4433 72505 4445 72539
rect 4479 72536 4491 72539
rect 5552 72536 5580 72567
rect 4479 72508 5580 72536
rect 4479 72505 4491 72508
rect 4433 72499 4491 72505
rect 5828 72480 5856 72576
rect 6454 72564 6460 72616
rect 6512 72604 6518 72616
rect 6641 72607 6699 72613
rect 6641 72604 6653 72607
rect 6512 72576 6653 72604
rect 6512 72564 6518 72576
rect 6641 72573 6653 72576
rect 6687 72604 6699 72607
rect 8018 72604 8024 72616
rect 6687 72576 8024 72604
rect 6687 72573 6699 72576
rect 6641 72567 6699 72573
rect 8018 72564 8024 72576
rect 8076 72564 8082 72616
rect 10870 72604 10876 72616
rect 10831 72576 10876 72604
rect 10870 72564 10876 72576
rect 10928 72564 10934 72616
rect 11425 72607 11483 72613
rect 11425 72573 11437 72607
rect 11471 72604 11483 72607
rect 11606 72604 11612 72616
rect 11471 72576 11612 72604
rect 11471 72573 11483 72576
rect 11425 72567 11483 72573
rect 11606 72564 11612 72576
rect 11664 72564 11670 72616
rect 11790 72604 11796 72616
rect 11751 72576 11796 72604
rect 11790 72564 11796 72576
rect 11848 72564 11854 72616
rect 11974 72604 11980 72616
rect 11935 72576 11980 72604
rect 11974 72564 11980 72576
rect 12032 72604 12038 72616
rect 12342 72604 12348 72616
rect 12032 72576 12348 72604
rect 12032 72564 12038 72576
rect 12342 72564 12348 72576
rect 12400 72564 12406 72616
rect 8849 72539 8907 72545
rect 8849 72505 8861 72539
rect 8895 72536 8907 72539
rect 10042 72536 10048 72548
rect 8895 72508 10048 72536
rect 8895 72505 8907 72508
rect 8849 72499 8907 72505
rect 10042 72496 10048 72508
rect 10100 72496 10106 72548
rect 12713 72539 12771 72545
rect 12713 72536 12725 72539
rect 12544 72508 12725 72536
rect 12544 72480 12572 72508
rect 12713 72505 12725 72508
rect 12759 72505 12771 72539
rect 12713 72499 12771 72505
rect 3421 72471 3479 72477
rect 3421 72437 3433 72471
rect 3467 72468 3479 72471
rect 3510 72468 3516 72480
rect 3467 72440 3516 72468
rect 3467 72437 3479 72440
rect 3421 72431 3479 72437
rect 3510 72428 3516 72440
rect 3568 72468 3574 72480
rect 4062 72468 4068 72480
rect 3568 72440 4068 72468
rect 3568 72428 3574 72440
rect 4062 72428 4068 72440
rect 4120 72428 4126 72480
rect 5810 72468 5816 72480
rect 5771 72440 5816 72468
rect 5810 72428 5816 72440
rect 5868 72428 5874 72480
rect 6178 72468 6184 72480
rect 6139 72440 6184 72468
rect 6178 72428 6184 72440
rect 6236 72428 6242 72480
rect 9214 72468 9220 72480
rect 9175 72440 9220 72468
rect 9214 72428 9220 72440
rect 9272 72428 9278 72480
rect 9674 72428 9680 72480
rect 9732 72468 9738 72480
rect 9953 72471 10011 72477
rect 9953 72468 9965 72471
rect 9732 72440 9965 72468
rect 9732 72428 9738 72440
rect 9953 72437 9965 72440
rect 9999 72468 10011 72471
rect 10502 72468 10508 72480
rect 9999 72440 10508 72468
rect 9999 72437 10011 72440
rect 9953 72431 10011 72437
rect 10502 72428 10508 72440
rect 10560 72428 10566 72480
rect 10689 72471 10747 72477
rect 10689 72437 10701 72471
rect 10735 72468 10747 72471
rect 12526 72468 12532 72480
rect 10735 72440 12532 72468
rect 10735 72437 10747 72440
rect 10689 72431 10747 72437
rect 12526 72428 12532 72440
rect 12584 72428 12590 72480
rect 1104 72378 18860 72400
rect 1104 72326 7648 72378
rect 7700 72326 7712 72378
rect 7764 72326 7776 72378
rect 7828 72326 7840 72378
rect 7892 72326 14315 72378
rect 14367 72326 14379 72378
rect 14431 72326 14443 72378
rect 14495 72326 14507 72378
rect 14559 72326 18860 72378
rect 1104 72304 18860 72326
rect 4982 72264 4988 72276
rect 4943 72236 4988 72264
rect 4982 72224 4988 72236
rect 5040 72224 5046 72276
rect 5534 72264 5540 72276
rect 5495 72236 5540 72264
rect 5534 72224 5540 72236
rect 5592 72224 5598 72276
rect 6086 72224 6092 72276
rect 6144 72264 6150 72276
rect 6181 72267 6239 72273
rect 6181 72264 6193 72267
rect 6144 72236 6193 72264
rect 6144 72224 6150 72236
rect 6181 72233 6193 72236
rect 6227 72233 6239 72267
rect 6181 72227 6239 72233
rect 10873 72267 10931 72273
rect 10873 72233 10885 72267
rect 10919 72264 10931 72267
rect 11974 72264 11980 72276
rect 10919 72236 11980 72264
rect 10919 72233 10931 72236
rect 10873 72227 10931 72233
rect 11974 72224 11980 72236
rect 12032 72224 12038 72276
rect 2774 72088 2780 72140
rect 2832 72128 2838 72140
rect 3234 72128 3240 72140
rect 2832 72100 3240 72128
rect 2832 72088 2838 72100
rect 3234 72088 3240 72100
rect 3292 72128 3298 72140
rect 3605 72131 3663 72137
rect 3605 72128 3617 72131
rect 3292 72100 3617 72128
rect 3292 72088 3298 72100
rect 3605 72097 3617 72100
rect 3651 72097 3663 72131
rect 3605 72091 3663 72097
rect 3694 72088 3700 72140
rect 3752 72128 3758 72140
rect 3881 72131 3939 72137
rect 3881 72128 3893 72131
rect 3752 72100 3893 72128
rect 3752 72088 3758 72100
rect 3881 72097 3893 72100
rect 3927 72097 3939 72131
rect 3881 72091 3939 72097
rect 6546 72088 6552 72140
rect 6604 72128 6610 72140
rect 6822 72128 6828 72140
rect 6604 72100 6828 72128
rect 6604 72088 6610 72100
rect 6822 72088 6828 72100
rect 6880 72128 6886 72140
rect 7098 72128 7104 72140
rect 6880 72100 7104 72128
rect 6880 72088 6886 72100
rect 7098 72088 7104 72100
rect 7156 72088 7162 72140
rect 8665 72131 8723 72137
rect 8665 72097 8677 72131
rect 8711 72128 8723 72131
rect 9214 72128 9220 72140
rect 8711 72100 9220 72128
rect 8711 72097 8723 72100
rect 8665 72091 8723 72097
rect 9214 72088 9220 72100
rect 9272 72088 9278 72140
rect 9306 72088 9312 72140
rect 9364 72128 9370 72140
rect 9674 72128 9680 72140
rect 9364 72100 9409 72128
rect 9635 72100 9680 72128
rect 9364 72088 9370 72100
rect 9674 72088 9680 72100
rect 9732 72088 9738 72140
rect 8110 72020 8116 72072
rect 8168 72060 8174 72072
rect 8570 72060 8576 72072
rect 8168 72032 8576 72060
rect 8168 72020 8174 72032
rect 8570 72020 8576 72032
rect 8628 72020 8634 72072
rect 8846 72060 8852 72072
rect 8807 72032 8852 72060
rect 8846 72020 8852 72032
rect 8904 72020 8910 72072
rect 5902 71952 5908 72004
rect 5960 71992 5966 72004
rect 6549 71995 6607 72001
rect 6549 71992 6561 71995
rect 5960 71964 6561 71992
rect 5960 71952 5966 71964
rect 6549 71961 6561 71964
rect 6595 71992 6607 71995
rect 6730 71992 6736 72004
rect 6595 71964 6736 71992
rect 6595 71961 6607 71964
rect 6549 71955 6607 71961
rect 6730 71952 6736 71964
rect 6788 71952 6794 72004
rect 7190 71952 7196 72004
rect 7248 71992 7254 72004
rect 7285 71995 7343 72001
rect 7285 71992 7297 71995
rect 7248 71964 7297 71992
rect 7248 71952 7254 71964
rect 7285 71961 7297 71964
rect 7331 71992 7343 71995
rect 8938 71992 8944 72004
rect 7331 71964 8944 71992
rect 7331 71961 7343 71964
rect 7285 71955 7343 71961
rect 8938 71952 8944 71964
rect 8996 71952 9002 72004
rect 7745 71927 7803 71933
rect 7745 71893 7757 71927
rect 7791 71924 7803 71927
rect 8202 71924 8208 71936
rect 7791 71896 8208 71924
rect 7791 71893 7803 71896
rect 7745 71887 7803 71893
rect 8202 71884 8208 71896
rect 8260 71884 8266 71936
rect 11241 71927 11299 71933
rect 11241 71893 11253 71927
rect 11287 71924 11299 71927
rect 11330 71924 11336 71936
rect 11287 71896 11336 71924
rect 11287 71893 11299 71896
rect 11241 71887 11299 71893
rect 11330 71884 11336 71896
rect 11388 71884 11394 71936
rect 1104 71834 18860 71856
rect 1104 71782 4315 71834
rect 4367 71782 4379 71834
rect 4431 71782 4443 71834
rect 4495 71782 4507 71834
rect 4559 71782 10982 71834
rect 11034 71782 11046 71834
rect 11098 71782 11110 71834
rect 11162 71782 11174 71834
rect 11226 71782 17648 71834
rect 17700 71782 17712 71834
rect 17764 71782 17776 71834
rect 17828 71782 17840 71834
rect 17892 71782 18860 71834
rect 1104 71760 18860 71782
rect 3234 71720 3240 71732
rect 3195 71692 3240 71720
rect 3234 71680 3240 71692
rect 3292 71680 3298 71732
rect 4617 71723 4675 71729
rect 4617 71689 4629 71723
rect 4663 71720 4675 71723
rect 5258 71720 5264 71732
rect 4663 71692 5264 71720
rect 4663 71689 4675 71692
rect 4617 71683 4675 71689
rect 5258 71680 5264 71692
rect 5316 71720 5322 71732
rect 6181 71723 6239 71729
rect 6181 71720 6193 71723
rect 5316 71692 6193 71720
rect 5316 71680 5322 71692
rect 6181 71689 6193 71692
rect 6227 71689 6239 71723
rect 6822 71720 6828 71732
rect 6783 71692 6828 71720
rect 6181 71683 6239 71689
rect 6822 71680 6828 71692
rect 6880 71680 6886 71732
rect 8662 71680 8668 71732
rect 8720 71720 8726 71732
rect 9125 71723 9183 71729
rect 9125 71720 9137 71723
rect 8720 71692 9137 71720
rect 8720 71680 8726 71692
rect 9125 71689 9137 71692
rect 9171 71720 9183 71723
rect 9306 71720 9312 71732
rect 9171 71692 9312 71720
rect 9171 71689 9183 71692
rect 9125 71683 9183 71689
rect 9306 71680 9312 71692
rect 9364 71680 9370 71732
rect 17494 71720 17500 71732
rect 17455 71692 17500 71720
rect 17494 71680 17500 71692
rect 17552 71680 17558 71732
rect 4801 71587 4859 71593
rect 4801 71553 4813 71587
rect 4847 71584 4859 71587
rect 5442 71584 5448 71596
rect 4847 71556 5448 71584
rect 4847 71553 4859 71556
rect 4801 71547 4859 71553
rect 5442 71544 5448 71556
rect 5500 71584 5506 71596
rect 6086 71584 6092 71596
rect 5500 71556 6092 71584
rect 5500 71544 5506 71556
rect 6086 71544 6092 71556
rect 6144 71584 6150 71596
rect 6546 71584 6552 71596
rect 6144 71556 6552 71584
rect 6144 71544 6150 71556
rect 6546 71544 6552 71556
rect 6604 71544 6610 71596
rect 7193 71587 7251 71593
rect 7193 71553 7205 71587
rect 7239 71584 7251 71587
rect 10594 71584 10600 71596
rect 7239 71556 8616 71584
rect 10555 71556 10600 71584
rect 7239 71553 7251 71556
rect 7193 71547 7251 71553
rect 5074 71516 5080 71528
rect 5035 71488 5080 71516
rect 5074 71476 5080 71488
rect 5132 71476 5138 71528
rect 7653 71519 7711 71525
rect 7653 71485 7665 71519
rect 7699 71485 7711 71519
rect 8202 71516 8208 71528
rect 8115 71488 8208 71516
rect 7653 71479 7711 71485
rect 3694 71380 3700 71392
rect 3655 71352 3700 71380
rect 3694 71340 3700 71352
rect 3752 71340 3758 71392
rect 7466 71380 7472 71392
rect 7427 71352 7472 71380
rect 7466 71340 7472 71352
rect 7524 71380 7530 71392
rect 7668 71380 7696 71479
rect 8202 71476 8208 71488
rect 8260 71516 8266 71528
rect 8386 71516 8392 71528
rect 8260 71488 8392 71516
rect 8260 71476 8266 71488
rect 8386 71476 8392 71488
rect 8444 71476 8450 71528
rect 8588 71525 8616 71556
rect 10594 71544 10600 71556
rect 10652 71544 10658 71596
rect 11330 71584 11336 71596
rect 11164 71556 11336 71584
rect 8573 71519 8631 71525
rect 8573 71485 8585 71519
rect 8619 71516 8631 71519
rect 8846 71516 8852 71528
rect 8619 71488 8852 71516
rect 8619 71485 8631 71488
rect 8573 71479 8631 71485
rect 8846 71476 8852 71488
rect 8904 71476 8910 71528
rect 11164 71525 11192 71556
rect 11330 71544 11336 71556
rect 11388 71584 11394 71596
rect 12897 71587 12955 71593
rect 12897 71584 12909 71587
rect 11388 71556 12909 71584
rect 11388 71544 11394 71556
rect 12897 71553 12909 71556
rect 12943 71553 12955 71587
rect 12897 71547 12955 71553
rect 11149 71519 11207 71525
rect 11149 71485 11161 71519
rect 11195 71485 11207 71519
rect 11149 71479 11207 71485
rect 11241 71519 11299 71525
rect 11241 71485 11253 71519
rect 11287 71516 11299 71519
rect 11287 71488 11376 71516
rect 11287 71485 11299 71488
rect 11241 71479 11299 71485
rect 11348 71460 11376 71488
rect 11422 71476 11428 71528
rect 11480 71516 11486 71528
rect 11698 71516 11704 71528
rect 11480 71488 11525 71516
rect 11659 71488 11704 71516
rect 11480 71476 11486 71488
rect 11698 71476 11704 71488
rect 11756 71476 11762 71528
rect 11882 71516 11888 71528
rect 11843 71488 11888 71516
rect 11882 71476 11888 71488
rect 11940 71476 11946 71528
rect 12802 71516 12808 71528
rect 12715 71488 12808 71516
rect 12802 71476 12808 71488
rect 12860 71516 12866 71528
rect 12989 71519 13047 71525
rect 12989 71516 13001 71519
rect 12860 71488 13001 71516
rect 12860 71476 12866 71488
rect 12989 71485 13001 71488
rect 13035 71485 13047 71519
rect 16114 71516 16120 71528
rect 16075 71488 16120 71516
rect 12989 71479 13047 71485
rect 16114 71476 16120 71488
rect 16172 71476 16178 71528
rect 16393 71519 16451 71525
rect 16393 71516 16405 71519
rect 16224 71488 16405 71516
rect 8754 71448 8760 71460
rect 8715 71420 8760 71448
rect 8754 71408 8760 71420
rect 8812 71408 8818 71460
rect 10505 71451 10563 71457
rect 10505 71417 10517 71451
rect 10551 71448 10563 71451
rect 11330 71448 11336 71460
rect 10551 71420 11336 71448
rect 10551 71417 10563 71420
rect 10505 71411 10563 71417
rect 11330 71408 11336 71420
rect 11388 71408 11394 71460
rect 7524 71352 7696 71380
rect 7524 71340 7530 71352
rect 9214 71340 9220 71392
rect 9272 71380 9278 71392
rect 9401 71383 9459 71389
rect 9401 71380 9413 71383
rect 9272 71352 9413 71380
rect 9272 71340 9278 71352
rect 9401 71349 9413 71352
rect 9447 71349 9459 71383
rect 9401 71343 9459 71349
rect 10137 71383 10195 71389
rect 10137 71349 10149 71383
rect 10183 71380 10195 71383
rect 11698 71380 11704 71392
rect 10183 71352 11704 71380
rect 10183 71349 10195 71352
rect 10137 71343 10195 71349
rect 11698 71340 11704 71352
rect 11756 71340 11762 71392
rect 16022 71380 16028 71392
rect 15983 71352 16028 71380
rect 16022 71340 16028 71352
rect 16080 71380 16086 71392
rect 16224 71380 16252 71488
rect 16393 71485 16405 71488
rect 16439 71485 16451 71519
rect 16393 71479 16451 71485
rect 16080 71352 16252 71380
rect 16080 71340 16086 71352
rect 1104 71290 18860 71312
rect 1104 71238 7648 71290
rect 7700 71238 7712 71290
rect 7764 71238 7776 71290
rect 7828 71238 7840 71290
rect 7892 71238 14315 71290
rect 14367 71238 14379 71290
rect 14431 71238 14443 71290
rect 14495 71238 14507 71290
rect 14559 71238 18860 71290
rect 1104 71216 18860 71238
rect 5442 71176 5448 71188
rect 5403 71148 5448 71176
rect 5442 71136 5448 71148
rect 5500 71136 5506 71188
rect 8205 71179 8263 71185
rect 8205 71145 8217 71179
rect 8251 71176 8263 71179
rect 8570 71176 8576 71188
rect 8251 71148 8576 71176
rect 8251 71145 8263 71148
rect 8205 71139 8263 71145
rect 8570 71136 8576 71148
rect 8628 71176 8634 71188
rect 9582 71176 9588 71188
rect 8628 71148 9588 71176
rect 8628 71136 8634 71148
rect 9582 71136 9588 71148
rect 9640 71136 9646 71188
rect 11057 71179 11115 71185
rect 11057 71145 11069 71179
rect 11103 71176 11115 71179
rect 11882 71176 11888 71188
rect 11103 71148 11888 71176
rect 11103 71145 11115 71148
rect 11057 71139 11115 71145
rect 11882 71136 11888 71148
rect 11940 71136 11946 71188
rect 10689 71111 10747 71117
rect 10689 71077 10701 71111
rect 10735 71108 10747 71111
rect 10778 71108 10784 71120
rect 10735 71080 10784 71108
rect 10735 71077 10747 71080
rect 10689 71071 10747 71077
rect 10778 71068 10784 71080
rect 10836 71108 10842 71120
rect 11422 71108 11428 71120
rect 10836 71080 11428 71108
rect 10836 71068 10842 71080
rect 11422 71068 11428 71080
rect 11480 71068 11486 71120
rect 4341 71043 4399 71049
rect 4341 71009 4353 71043
rect 4387 71040 4399 71043
rect 4522 71040 4528 71052
rect 4387 71012 4528 71040
rect 4387 71009 4399 71012
rect 4341 71003 4399 71009
rect 4522 71000 4528 71012
rect 4580 71000 4586 71052
rect 4706 71040 4712 71052
rect 4667 71012 4712 71040
rect 4706 71000 4712 71012
rect 4764 71000 4770 71052
rect 5074 71000 5080 71052
rect 5132 71040 5138 71052
rect 5169 71043 5227 71049
rect 5169 71040 5181 71043
rect 5132 71012 5181 71040
rect 5132 71000 5138 71012
rect 5169 71009 5181 71012
rect 5215 71040 5227 71043
rect 6730 71040 6736 71052
rect 5215 71012 6736 71040
rect 5215 71009 5227 71012
rect 5169 71003 5227 71009
rect 6730 71000 6736 71012
rect 6788 71040 6794 71052
rect 7469 71043 7527 71049
rect 7469 71040 7481 71043
rect 6788 71012 7481 71040
rect 6788 71000 6794 71012
rect 7469 71009 7481 71012
rect 7515 71040 7527 71043
rect 8110 71040 8116 71052
rect 7515 71012 8116 71040
rect 7515 71009 7527 71012
rect 7469 71003 7527 71009
rect 8110 71000 8116 71012
rect 8168 71000 8174 71052
rect 8754 71000 8760 71052
rect 8812 71040 8818 71052
rect 8941 71043 8999 71049
rect 8941 71040 8953 71043
rect 8812 71012 8953 71040
rect 8812 71000 8818 71012
rect 8941 71009 8953 71012
rect 8987 71009 8999 71043
rect 8941 71003 8999 71009
rect 6822 70972 6828 70984
rect 6783 70944 6828 70972
rect 6822 70932 6828 70944
rect 6880 70932 6886 70984
rect 9582 70972 9588 70984
rect 9543 70944 9588 70972
rect 9582 70932 9588 70944
rect 9640 70932 9646 70984
rect 4154 70904 4160 70916
rect 4115 70876 4160 70904
rect 4154 70864 4160 70876
rect 4212 70864 4218 70916
rect 8386 70796 8392 70848
rect 8444 70836 8450 70848
rect 8481 70839 8539 70845
rect 8481 70836 8493 70839
rect 8444 70808 8493 70836
rect 8444 70796 8450 70808
rect 8481 70805 8493 70808
rect 8527 70805 8539 70839
rect 8481 70799 8539 70805
rect 9953 70839 10011 70845
rect 9953 70805 9965 70839
rect 9999 70836 10011 70839
rect 10134 70836 10140 70848
rect 9999 70808 10140 70836
rect 9999 70805 10011 70808
rect 9953 70799 10011 70805
rect 10134 70796 10140 70808
rect 10192 70796 10198 70848
rect 10226 70796 10232 70848
rect 10284 70836 10290 70848
rect 11885 70839 11943 70845
rect 10284 70808 10329 70836
rect 10284 70796 10290 70808
rect 11885 70805 11897 70839
rect 11931 70836 11943 70839
rect 11974 70836 11980 70848
rect 11931 70808 11980 70836
rect 11931 70805 11943 70808
rect 11885 70799 11943 70805
rect 11974 70796 11980 70808
rect 12032 70796 12038 70848
rect 16114 70836 16120 70848
rect 16075 70808 16120 70836
rect 16114 70796 16120 70808
rect 16172 70796 16178 70848
rect 1104 70746 18860 70768
rect 1104 70694 4315 70746
rect 4367 70694 4379 70746
rect 4431 70694 4443 70746
rect 4495 70694 4507 70746
rect 4559 70694 10982 70746
rect 11034 70694 11046 70746
rect 11098 70694 11110 70746
rect 11162 70694 11174 70746
rect 11226 70694 17648 70746
rect 17700 70694 17712 70746
rect 17764 70694 17776 70746
rect 17828 70694 17840 70746
rect 17892 70694 18860 70746
rect 1104 70672 18860 70694
rect 1486 70592 1492 70644
rect 1544 70632 1550 70644
rect 2041 70635 2099 70641
rect 2041 70632 2053 70635
rect 1544 70604 2053 70632
rect 1544 70592 1550 70604
rect 2041 70601 2053 70604
rect 2087 70632 2099 70635
rect 2774 70632 2780 70644
rect 2087 70604 2780 70632
rect 2087 70601 2099 70604
rect 2041 70595 2099 70601
rect 2774 70592 2780 70604
rect 2832 70592 2838 70644
rect 4341 70635 4399 70641
rect 4341 70601 4353 70635
rect 4387 70632 4399 70635
rect 4706 70632 4712 70644
rect 4387 70604 4712 70632
rect 4387 70601 4399 70604
rect 4341 70595 4399 70601
rect 4706 70592 4712 70604
rect 4764 70592 4770 70644
rect 5534 70592 5540 70644
rect 5592 70632 5598 70644
rect 5905 70635 5963 70641
rect 5905 70632 5917 70635
rect 5592 70604 5917 70632
rect 5592 70592 5598 70604
rect 5905 70601 5917 70604
rect 5951 70601 5963 70635
rect 5905 70595 5963 70601
rect 7101 70635 7159 70641
rect 7101 70601 7113 70635
rect 7147 70632 7159 70635
rect 8570 70632 8576 70644
rect 7147 70604 8576 70632
rect 7147 70601 7159 70604
rect 7101 70595 7159 70601
rect 8570 70592 8576 70604
rect 8628 70592 8634 70644
rect 10318 70592 10324 70644
rect 10376 70632 10382 70644
rect 10778 70632 10784 70644
rect 10376 70604 10784 70632
rect 10376 70592 10382 70604
rect 10778 70592 10784 70604
rect 10836 70592 10842 70644
rect 11698 70592 11704 70644
rect 11756 70632 11762 70644
rect 11885 70635 11943 70641
rect 11885 70632 11897 70635
rect 11756 70604 11897 70632
rect 11756 70592 11762 70604
rect 11885 70601 11897 70604
rect 11931 70601 11943 70635
rect 11885 70595 11943 70601
rect 9493 70567 9551 70573
rect 9493 70533 9505 70567
rect 9539 70564 9551 70567
rect 9677 70567 9735 70573
rect 9677 70564 9689 70567
rect 9539 70536 9689 70564
rect 9539 70533 9551 70536
rect 9493 70527 9551 70533
rect 9677 70533 9689 70536
rect 9723 70564 9735 70567
rect 9723 70536 10456 70564
rect 9723 70533 9735 70536
rect 9677 70527 9735 70533
rect 5718 70496 5724 70508
rect 5631 70468 5724 70496
rect 5718 70456 5724 70468
rect 5776 70496 5782 70508
rect 7834 70496 7840 70508
rect 5776 70468 6592 70496
rect 7795 70468 7840 70496
rect 5776 70456 5782 70468
rect 5902 70428 5908 70440
rect 5863 70400 5908 70428
rect 5902 70388 5908 70400
rect 5960 70388 5966 70440
rect 6564 70437 6592 70468
rect 7834 70456 7840 70468
rect 7892 70456 7898 70508
rect 8110 70456 8116 70508
rect 8168 70496 8174 70508
rect 8297 70499 8355 70505
rect 8297 70496 8309 70499
rect 8168 70468 8309 70496
rect 8168 70456 8174 70468
rect 8297 70465 8309 70468
rect 8343 70496 8355 70499
rect 9033 70499 9091 70505
rect 9033 70496 9045 70499
rect 8343 70468 9045 70496
rect 8343 70465 8355 70468
rect 8297 70459 8355 70465
rect 9033 70465 9045 70468
rect 9079 70465 9091 70499
rect 10226 70496 10232 70508
rect 9033 70459 9091 70465
rect 9968 70468 10232 70496
rect 6549 70431 6607 70437
rect 6549 70397 6561 70431
rect 6595 70428 6607 70431
rect 6822 70428 6828 70440
rect 6595 70400 6828 70428
rect 6595 70397 6607 70400
rect 6549 70391 6607 70397
rect 6822 70388 6828 70400
rect 6880 70388 6886 70440
rect 8205 70431 8263 70437
rect 8205 70397 8217 70431
rect 8251 70428 8263 70431
rect 8386 70428 8392 70440
rect 8251 70400 8392 70428
rect 8251 70397 8263 70400
rect 8205 70391 8263 70397
rect 8386 70388 8392 70400
rect 8444 70388 8450 70440
rect 8570 70428 8576 70440
rect 8531 70400 8576 70428
rect 8570 70388 8576 70400
rect 8628 70388 8634 70440
rect 8665 70431 8723 70437
rect 8665 70397 8677 70431
rect 8711 70397 8723 70431
rect 8665 70391 8723 70397
rect 8680 70360 8708 70391
rect 9766 70388 9772 70440
rect 9824 70428 9830 70440
rect 9968 70437 9996 70468
rect 10226 70456 10232 70468
rect 10284 70456 10290 70508
rect 10428 70496 10456 70536
rect 10778 70496 10784 70508
rect 10428 70468 10548 70496
rect 10739 70468 10784 70496
rect 9953 70431 10011 70437
rect 9953 70428 9965 70431
rect 9824 70400 9965 70428
rect 9824 70388 9830 70400
rect 9953 70397 9965 70400
rect 9999 70397 10011 70431
rect 10134 70428 10140 70440
rect 10095 70400 10140 70428
rect 9953 70391 10011 70397
rect 10134 70388 10140 70400
rect 10192 70428 10198 70440
rect 10410 70428 10416 70440
rect 10192 70400 10416 70428
rect 10192 70388 10198 70400
rect 10410 70388 10416 70400
rect 10468 70388 10474 70440
rect 10520 70437 10548 70468
rect 10778 70456 10784 70468
rect 10836 70456 10842 70508
rect 10505 70431 10563 70437
rect 10505 70397 10517 70431
rect 10551 70397 10563 70431
rect 10505 70391 10563 70397
rect 11698 70388 11704 70440
rect 11756 70428 11762 70440
rect 11974 70428 11980 70440
rect 11756 70400 11980 70428
rect 11756 70388 11762 70400
rect 11974 70388 11980 70400
rect 12032 70388 12038 70440
rect 12066 70388 12072 70440
rect 12124 70428 12130 70440
rect 12161 70431 12219 70437
rect 12161 70428 12173 70431
rect 12124 70400 12173 70428
rect 12124 70388 12130 70400
rect 12161 70397 12173 70400
rect 12207 70397 12219 70431
rect 12161 70391 12219 70397
rect 12529 70431 12587 70437
rect 12529 70397 12541 70431
rect 12575 70397 12587 70431
rect 12529 70391 12587 70397
rect 12544 70360 12572 70391
rect 7484 70332 8708 70360
rect 11808 70332 12572 70360
rect 7484 70304 7512 70332
rect 11808 70304 11836 70332
rect 1673 70295 1731 70301
rect 1673 70261 1685 70295
rect 1719 70292 1731 70295
rect 1762 70292 1768 70304
rect 1719 70264 1768 70292
rect 1719 70261 1731 70264
rect 1673 70255 1731 70261
rect 1762 70252 1768 70264
rect 1820 70252 1826 70304
rect 4062 70252 4068 70304
rect 4120 70292 4126 70304
rect 4614 70292 4620 70304
rect 4120 70264 4620 70292
rect 4120 70252 4126 70264
rect 4614 70252 4620 70264
rect 4672 70252 4678 70304
rect 7466 70292 7472 70304
rect 7427 70264 7472 70292
rect 7466 70252 7472 70264
rect 7524 70252 7530 70304
rect 8018 70252 8024 70304
rect 8076 70292 8082 70304
rect 9582 70292 9588 70304
rect 8076 70264 9588 70292
rect 8076 70252 8082 70264
rect 9582 70252 9588 70264
rect 9640 70252 9646 70304
rect 9677 70295 9735 70301
rect 9677 70261 9689 70295
rect 9723 70292 9735 70295
rect 10134 70292 10140 70304
rect 9723 70264 10140 70292
rect 9723 70261 9735 70264
rect 9677 70255 9735 70261
rect 10134 70252 10140 70264
rect 10192 70252 10198 70304
rect 11701 70295 11759 70301
rect 11701 70261 11713 70295
rect 11747 70292 11759 70295
rect 11790 70292 11796 70304
rect 11747 70264 11796 70292
rect 11747 70261 11759 70264
rect 11701 70255 11759 70261
rect 11790 70252 11796 70264
rect 11848 70252 11854 70304
rect 1104 70202 18860 70224
rect 1104 70150 7648 70202
rect 7700 70150 7712 70202
rect 7764 70150 7776 70202
rect 7828 70150 7840 70202
rect 7892 70150 14315 70202
rect 14367 70150 14379 70202
rect 14431 70150 14443 70202
rect 14495 70150 14507 70202
rect 14559 70150 18860 70202
rect 1104 70128 18860 70150
rect 6641 70091 6699 70097
rect 6641 70057 6653 70091
rect 6687 70088 6699 70091
rect 6730 70088 6736 70100
rect 6687 70060 6736 70088
rect 6687 70057 6699 70060
rect 6641 70051 6699 70057
rect 6730 70048 6736 70060
rect 6788 70048 6794 70100
rect 8754 70088 8760 70100
rect 8715 70060 8760 70088
rect 8754 70048 8760 70060
rect 8812 70048 8818 70100
rect 9950 70020 9956 70032
rect 9508 69992 9956 70020
rect 1486 69952 1492 69964
rect 1447 69924 1492 69952
rect 1486 69912 1492 69924
rect 1544 69912 1550 69964
rect 4798 69912 4804 69964
rect 4856 69952 4862 69964
rect 5077 69955 5135 69961
rect 5077 69952 5089 69955
rect 4856 69924 5089 69952
rect 4856 69912 4862 69924
rect 5077 69921 5089 69924
rect 5123 69921 5135 69955
rect 5077 69915 5135 69921
rect 7101 69955 7159 69961
rect 7101 69921 7113 69955
rect 7147 69952 7159 69955
rect 7374 69952 7380 69964
rect 7147 69924 7380 69952
rect 7147 69921 7159 69924
rect 7101 69915 7159 69921
rect 7374 69912 7380 69924
rect 7432 69952 7438 69964
rect 8202 69952 8208 69964
rect 7432 69924 8208 69952
rect 7432 69912 7438 69924
rect 8202 69912 8208 69924
rect 8260 69912 8266 69964
rect 9508 69961 9536 69992
rect 9950 69980 9956 69992
rect 10008 70020 10014 70032
rect 11057 70023 11115 70029
rect 11057 70020 11069 70023
rect 10008 69992 11069 70020
rect 10008 69980 10014 69992
rect 11057 69989 11069 69992
rect 11103 69989 11115 70023
rect 11057 69983 11115 69989
rect 9493 69955 9551 69961
rect 9493 69921 9505 69955
rect 9539 69921 9551 69955
rect 9674 69952 9680 69964
rect 9635 69924 9680 69952
rect 9493 69915 9551 69921
rect 9674 69912 9680 69924
rect 9732 69912 9738 69964
rect 10045 69955 10103 69961
rect 10045 69952 10057 69955
rect 9876 69924 10057 69952
rect 1762 69884 1768 69896
rect 1723 69856 1768 69884
rect 1762 69844 1768 69856
rect 1820 69844 1826 69896
rect 6546 69844 6552 69896
rect 6604 69884 6610 69896
rect 6825 69887 6883 69893
rect 6825 69884 6837 69887
rect 6604 69856 6837 69884
rect 6604 69844 6610 69856
rect 6825 69853 6837 69856
rect 6871 69853 6883 69887
rect 9766 69884 9772 69896
rect 9727 69856 9772 69884
rect 6825 69847 6883 69853
rect 9766 69844 9772 69856
rect 9824 69844 9830 69896
rect 9876 69828 9904 69924
rect 10045 69921 10057 69924
rect 10091 69952 10103 69955
rect 10134 69952 10140 69964
rect 10091 69924 10140 69952
rect 10091 69921 10103 69924
rect 10045 69915 10103 69921
rect 10134 69912 10140 69924
rect 10192 69912 10198 69964
rect 10410 69912 10416 69964
rect 10468 69952 10474 69964
rect 10597 69955 10655 69961
rect 10597 69952 10609 69955
rect 10468 69924 10609 69952
rect 10468 69912 10474 69924
rect 10597 69921 10609 69924
rect 10643 69921 10655 69955
rect 10597 69915 10655 69921
rect 9858 69776 9864 69828
rect 9916 69776 9922 69828
rect 11974 69776 11980 69828
rect 12032 69816 12038 69828
rect 12161 69819 12219 69825
rect 12161 69816 12173 69819
rect 12032 69788 12173 69816
rect 12032 69776 12038 69788
rect 12161 69785 12173 69788
rect 12207 69785 12219 69819
rect 12161 69779 12219 69785
rect 2498 69708 2504 69760
rect 2556 69748 2562 69760
rect 2869 69751 2927 69757
rect 2869 69748 2881 69751
rect 2556 69720 2881 69748
rect 2556 69708 2562 69720
rect 2869 69717 2881 69720
rect 2915 69717 2927 69751
rect 2869 69711 2927 69717
rect 4157 69751 4215 69757
rect 4157 69717 4169 69751
rect 4203 69748 4215 69751
rect 4614 69748 4620 69760
rect 4203 69720 4620 69748
rect 4203 69717 4215 69720
rect 4157 69711 4215 69717
rect 4614 69708 4620 69720
rect 4672 69708 4678 69760
rect 5258 69748 5264 69760
rect 5219 69720 5264 69748
rect 5258 69708 5264 69720
rect 5316 69748 5322 69760
rect 5813 69751 5871 69757
rect 5813 69748 5825 69751
rect 5316 69720 5825 69748
rect 5316 69708 5322 69720
rect 5813 69717 5825 69720
rect 5859 69748 5871 69751
rect 5902 69748 5908 69760
rect 5859 69720 5908 69748
rect 5859 69717 5871 69720
rect 5813 69711 5871 69717
rect 5902 69708 5908 69720
rect 5960 69708 5966 69760
rect 8386 69748 8392 69760
rect 8347 69720 8392 69748
rect 8386 69708 8392 69720
rect 8444 69708 8450 69760
rect 9217 69751 9275 69757
rect 9217 69717 9229 69751
rect 9263 69748 9275 69751
rect 10410 69748 10416 69760
rect 9263 69720 10416 69748
rect 9263 69717 9275 69720
rect 9217 69711 9275 69717
rect 10410 69708 10416 69720
rect 10468 69708 10474 69760
rect 11885 69751 11943 69757
rect 11885 69717 11897 69751
rect 11931 69748 11943 69751
rect 12066 69748 12072 69760
rect 11931 69720 12072 69748
rect 11931 69717 11943 69720
rect 11885 69711 11943 69717
rect 12066 69708 12072 69720
rect 12124 69708 12130 69760
rect 1104 69658 18860 69680
rect 1104 69606 4315 69658
rect 4367 69606 4379 69658
rect 4431 69606 4443 69658
rect 4495 69606 4507 69658
rect 4559 69606 10982 69658
rect 11034 69606 11046 69658
rect 11098 69606 11110 69658
rect 11162 69606 11174 69658
rect 11226 69606 17648 69658
rect 17700 69606 17712 69658
rect 17764 69606 17776 69658
rect 17828 69606 17840 69658
rect 17892 69606 18860 69658
rect 1104 69584 18860 69606
rect 5721 69547 5779 69553
rect 5721 69513 5733 69547
rect 5767 69544 5779 69547
rect 5810 69544 5816 69556
rect 5767 69516 5816 69544
rect 5767 69513 5779 69516
rect 5721 69507 5779 69513
rect 5810 69504 5816 69516
rect 5868 69504 5874 69556
rect 9490 69504 9496 69556
rect 9548 69544 9554 69556
rect 9861 69547 9919 69553
rect 9861 69544 9873 69547
rect 9548 69516 9873 69544
rect 9548 69504 9554 69516
rect 9861 69513 9873 69516
rect 9907 69513 9919 69547
rect 9861 69507 9919 69513
rect 4154 69476 4160 69488
rect 4115 69448 4160 69476
rect 4154 69436 4160 69448
rect 4212 69436 4218 69488
rect 5828 69476 5856 69504
rect 6730 69476 6736 69488
rect 5828 69448 6736 69476
rect 6730 69436 6736 69448
rect 6788 69476 6794 69488
rect 6788 69448 6868 69476
rect 6788 69436 6794 69448
rect 1765 69411 1823 69417
rect 1765 69377 1777 69411
rect 1811 69408 1823 69411
rect 2498 69408 2504 69420
rect 1811 69380 2504 69408
rect 1811 69377 1823 69380
rect 1765 69371 1823 69377
rect 2498 69368 2504 69380
rect 2556 69368 2562 69420
rect 5810 69408 5816 69420
rect 5771 69380 5816 69408
rect 5810 69368 5816 69380
rect 5868 69368 5874 69420
rect 6840 69417 6868 69448
rect 12066 69436 12072 69488
rect 12124 69476 12130 69488
rect 12124 69448 12296 69476
rect 12124 69436 12130 69448
rect 6825 69411 6883 69417
rect 6825 69377 6837 69411
rect 6871 69377 6883 69411
rect 6825 69371 6883 69377
rect 7466 69368 7472 69420
rect 7524 69408 7530 69420
rect 7653 69411 7711 69417
rect 7653 69408 7665 69411
rect 7524 69380 7665 69408
rect 7524 69368 7530 69380
rect 7653 69377 7665 69380
rect 7699 69377 7711 69411
rect 7653 69371 7711 69377
rect 9125 69411 9183 69417
rect 9125 69377 9137 69411
rect 9171 69408 9183 69411
rect 9171 69380 10180 69408
rect 9171 69377 9183 69380
rect 9125 69371 9183 69377
rect 10152 69352 10180 69380
rect 11882 69368 11888 69420
rect 11940 69408 11946 69420
rect 12161 69411 12219 69417
rect 12161 69408 12173 69411
rect 11940 69380 12173 69408
rect 11940 69368 11946 69380
rect 12161 69377 12173 69380
rect 12207 69377 12219 69411
rect 12161 69371 12219 69377
rect 2317 69343 2375 69349
rect 2317 69309 2329 69343
rect 2363 69340 2375 69343
rect 2590 69340 2596 69352
rect 2363 69312 2596 69340
rect 2363 69309 2375 69312
rect 2317 69303 2375 69309
rect 2590 69300 2596 69312
rect 2648 69300 2654 69352
rect 4062 69340 4068 69352
rect 3804 69312 4068 69340
rect 1762 69232 1768 69284
rect 1820 69272 1826 69284
rect 2133 69275 2191 69281
rect 2133 69272 2145 69275
rect 1820 69244 2145 69272
rect 1820 69232 1826 69244
rect 2133 69241 2145 69244
rect 2179 69272 2191 69275
rect 2179 69244 3464 69272
rect 2179 69241 2191 69244
rect 2133 69235 2191 69241
rect 2222 69164 2228 69216
rect 2280 69204 2286 69216
rect 2409 69207 2467 69213
rect 2409 69204 2421 69207
rect 2280 69176 2421 69204
rect 2280 69164 2286 69176
rect 2409 69173 2421 69176
rect 2455 69173 2467 69207
rect 2409 69167 2467 69173
rect 2590 69164 2596 69216
rect 2648 69204 2654 69216
rect 3050 69204 3056 69216
rect 2648 69176 3056 69204
rect 2648 69164 2654 69176
rect 3050 69164 3056 69176
rect 3108 69164 3114 69216
rect 3436 69213 3464 69244
rect 3421 69207 3479 69213
rect 3421 69173 3433 69207
rect 3467 69204 3479 69207
rect 3602 69204 3608 69216
rect 3467 69176 3608 69204
rect 3467 69173 3479 69176
rect 3421 69167 3479 69173
rect 3602 69164 3608 69176
rect 3660 69164 3666 69216
rect 3694 69164 3700 69216
rect 3752 69204 3758 69216
rect 3804 69213 3832 69312
rect 4062 69300 4068 69312
rect 4120 69300 4126 69352
rect 4614 69340 4620 69352
rect 4575 69312 4620 69340
rect 4614 69300 4620 69312
rect 4672 69300 4678 69352
rect 6362 69340 6368 69352
rect 6323 69312 6368 69340
rect 6362 69300 6368 69312
rect 6420 69300 6426 69352
rect 6638 69340 6644 69352
rect 6599 69312 6644 69340
rect 6638 69300 6644 69312
rect 6696 69300 6702 69352
rect 7190 69300 7196 69352
rect 7248 69340 7254 69352
rect 7561 69343 7619 69349
rect 7561 69340 7573 69343
rect 7248 69312 7573 69340
rect 7248 69300 7254 69312
rect 7561 69309 7573 69312
rect 7607 69340 7619 69343
rect 8202 69340 8208 69352
rect 7607 69312 8208 69340
rect 7607 69309 7619 69312
rect 7561 69303 7619 69309
rect 8202 69300 8208 69312
rect 8260 69300 8266 69352
rect 9950 69340 9956 69352
rect 9911 69312 9956 69340
rect 9950 69300 9956 69312
rect 10008 69300 10014 69352
rect 10134 69340 10140 69352
rect 10095 69312 10140 69340
rect 10134 69300 10140 69312
rect 10192 69300 10198 69352
rect 10505 69343 10563 69349
rect 10505 69340 10517 69343
rect 10244 69312 10517 69340
rect 8757 69275 8815 69281
rect 8757 69241 8769 69275
rect 8803 69272 8815 69275
rect 9674 69272 9680 69284
rect 8803 69244 9680 69272
rect 8803 69241 8815 69244
rect 8757 69235 8815 69241
rect 9674 69232 9680 69244
rect 9732 69232 9738 69284
rect 3789 69207 3847 69213
rect 3789 69204 3801 69207
rect 3752 69176 3801 69204
rect 3752 69164 3758 69176
rect 3789 69173 3801 69176
rect 3835 69173 3847 69207
rect 3789 69167 3847 69173
rect 4798 69164 4804 69216
rect 4856 69204 4862 69216
rect 5077 69207 5135 69213
rect 5077 69204 5089 69207
rect 4856 69176 5089 69204
rect 4856 69164 4862 69176
rect 5077 69173 5089 69176
rect 5123 69173 5135 69207
rect 5077 69167 5135 69173
rect 7193 69207 7251 69213
rect 7193 69173 7205 69207
rect 7239 69204 7251 69207
rect 7374 69204 7380 69216
rect 7239 69176 7380 69204
rect 7239 69173 7251 69176
rect 7193 69167 7251 69173
rect 7374 69164 7380 69176
rect 7432 69164 7438 69216
rect 9490 69204 9496 69216
rect 9451 69176 9496 69204
rect 9490 69164 9496 69176
rect 9548 69204 9554 69216
rect 10244 69204 10272 69312
rect 10505 69309 10517 69312
rect 10551 69309 10563 69343
rect 10505 69303 10563 69309
rect 11241 69343 11299 69349
rect 11241 69309 11253 69343
rect 11287 69309 11299 69343
rect 11241 69303 11299 69309
rect 11256 69272 11284 69303
rect 11974 69300 11980 69352
rect 12032 69340 12038 69352
rect 12069 69343 12127 69349
rect 12069 69340 12081 69343
rect 12032 69312 12081 69340
rect 12032 69300 12038 69312
rect 12069 69309 12081 69312
rect 12115 69309 12127 69343
rect 12268 69340 12296 69448
rect 12437 69343 12495 69349
rect 12437 69340 12449 69343
rect 12268 69312 12449 69340
rect 12069 69303 12127 69309
rect 12437 69309 12449 69312
rect 12483 69309 12495 69343
rect 12437 69303 12495 69309
rect 12805 69343 12863 69349
rect 12805 69309 12817 69343
rect 12851 69309 12863 69343
rect 12805 69303 12863 69309
rect 11609 69275 11667 69281
rect 11609 69272 11621 69275
rect 11256 69244 11621 69272
rect 11609 69241 11621 69244
rect 11655 69272 11667 69275
rect 11790 69272 11796 69284
rect 11655 69244 11796 69272
rect 11655 69241 11667 69244
rect 11609 69235 11667 69241
rect 11790 69232 11796 69244
rect 11848 69272 11854 69284
rect 12342 69272 12348 69284
rect 11848 69244 12348 69272
rect 11848 69232 11854 69244
rect 12342 69232 12348 69244
rect 12400 69232 12406 69284
rect 9548 69176 10272 69204
rect 9548 69164 9554 69176
rect 11054 69164 11060 69216
rect 11112 69204 11118 69216
rect 11885 69207 11943 69213
rect 11885 69204 11897 69207
rect 11112 69176 11897 69204
rect 11112 69164 11118 69176
rect 11885 69173 11897 69176
rect 11931 69204 11943 69207
rect 12820 69204 12848 69303
rect 11931 69176 12848 69204
rect 11931 69173 11943 69176
rect 11885 69167 11943 69173
rect 1104 69114 18860 69136
rect 1104 69062 7648 69114
rect 7700 69062 7712 69114
rect 7764 69062 7776 69114
rect 7828 69062 7840 69114
rect 7892 69062 14315 69114
rect 14367 69062 14379 69114
rect 14431 69062 14443 69114
rect 14495 69062 14507 69114
rect 14559 69062 18860 69114
rect 1104 69040 18860 69062
rect 5534 69000 5540 69012
rect 5447 68972 5540 69000
rect 5534 68960 5540 68972
rect 5592 69000 5598 69012
rect 5994 69000 6000 69012
rect 5592 68972 6000 69000
rect 5592 68960 5598 68972
rect 5994 68960 6000 68972
rect 6052 68960 6058 69012
rect 6273 69003 6331 69009
rect 6273 68969 6285 69003
rect 6319 69000 6331 69003
rect 6638 69000 6644 69012
rect 6319 68972 6644 69000
rect 6319 68969 6331 68972
rect 6273 68963 6331 68969
rect 6638 68960 6644 68972
rect 6696 68960 6702 69012
rect 3510 68932 3516 68944
rect 3471 68904 3516 68932
rect 3510 68892 3516 68904
rect 3568 68892 3574 68944
rect 9490 68892 9496 68944
rect 9548 68932 9554 68944
rect 13817 68935 13875 68941
rect 9548 68904 9812 68932
rect 9548 68892 9554 68904
rect 2222 68864 2228 68876
rect 2183 68836 2228 68864
rect 2222 68824 2228 68836
rect 2280 68824 2286 68876
rect 2498 68864 2504 68876
rect 2459 68836 2504 68864
rect 2498 68824 2504 68836
rect 2556 68824 2562 68876
rect 3878 68824 3884 68876
rect 3936 68864 3942 68876
rect 4341 68867 4399 68873
rect 4341 68864 4353 68867
rect 3936 68836 4353 68864
rect 3936 68824 3942 68836
rect 4341 68833 4353 68836
rect 4387 68833 4399 68867
rect 5350 68864 5356 68876
rect 5311 68836 5356 68864
rect 4341 68827 4399 68833
rect 5350 68824 5356 68836
rect 5408 68824 5414 68876
rect 8018 68864 8024 68876
rect 7979 68836 8024 68864
rect 8018 68824 8024 68836
rect 8076 68824 8082 68876
rect 8389 68867 8447 68873
rect 8389 68833 8401 68867
rect 8435 68864 8447 68867
rect 8570 68864 8576 68876
rect 8435 68836 8576 68864
rect 8435 68833 8447 68836
rect 8389 68827 8447 68833
rect 8570 68824 8576 68836
rect 8628 68824 8634 68876
rect 9784 68873 9812 68904
rect 13817 68901 13829 68935
rect 13863 68932 13875 68935
rect 14090 68932 14096 68944
rect 13863 68904 14096 68932
rect 13863 68901 13875 68904
rect 13817 68895 13875 68901
rect 14090 68892 14096 68904
rect 14148 68892 14154 68944
rect 9677 68867 9735 68873
rect 9677 68833 9689 68867
rect 9723 68833 9735 68867
rect 9677 68827 9735 68833
rect 9769 68867 9827 68873
rect 9769 68833 9781 68867
rect 9815 68833 9827 68867
rect 9769 68827 9827 68833
rect 10413 68867 10471 68873
rect 10413 68833 10425 68867
rect 10459 68833 10471 68867
rect 10413 68827 10471 68833
rect 1670 68796 1676 68808
rect 1631 68768 1676 68796
rect 1670 68756 1676 68768
rect 1728 68756 1734 68808
rect 2685 68799 2743 68805
rect 2685 68765 2697 68799
rect 2731 68796 2743 68799
rect 2774 68796 2780 68808
rect 2731 68768 2780 68796
rect 2731 68765 2743 68768
rect 2685 68759 2743 68765
rect 2774 68756 2780 68768
rect 2832 68756 2838 68808
rect 4062 68756 4068 68808
rect 4120 68796 4126 68808
rect 4525 68799 4583 68805
rect 4120 68768 4165 68796
rect 4120 68756 4126 68768
rect 4525 68765 4537 68799
rect 4571 68796 4583 68799
rect 4982 68796 4988 68808
rect 4571 68768 4988 68796
rect 4571 68765 4583 68768
rect 4525 68759 4583 68765
rect 4982 68756 4988 68768
rect 5040 68756 5046 68808
rect 7006 68756 7012 68808
rect 7064 68796 7070 68808
rect 7377 68799 7435 68805
rect 7377 68796 7389 68799
rect 7064 68768 7389 68796
rect 7064 68756 7070 68768
rect 7377 68765 7389 68768
rect 7423 68765 7435 68799
rect 7377 68759 7435 68765
rect 7929 68799 7987 68805
rect 7929 68765 7941 68799
rect 7975 68765 7987 68799
rect 8294 68796 8300 68808
rect 8255 68768 8300 68796
rect 7929 68759 7987 68765
rect 4893 68731 4951 68737
rect 4893 68697 4905 68731
rect 4939 68728 4951 68731
rect 5074 68728 5080 68740
rect 4939 68700 5080 68728
rect 4939 68697 4951 68700
rect 4893 68691 4951 68697
rect 5074 68688 5080 68700
rect 5132 68688 5138 68740
rect 5905 68731 5963 68737
rect 5905 68697 5917 68731
rect 5951 68728 5963 68731
rect 6362 68728 6368 68740
rect 5951 68700 6368 68728
rect 5951 68697 5963 68700
rect 5905 68691 5963 68697
rect 6362 68688 6368 68700
rect 6420 68728 6426 68740
rect 6914 68728 6920 68740
rect 6420 68700 6920 68728
rect 6420 68688 6426 68700
rect 6914 68688 6920 68700
rect 6972 68688 6978 68740
rect 7944 68728 7972 68759
rect 8294 68756 8300 68768
rect 8352 68756 8358 68808
rect 8018 68728 8024 68740
rect 7944 68700 8024 68728
rect 8018 68688 8024 68700
rect 8076 68688 8082 68740
rect 8941 68731 8999 68737
rect 8941 68697 8953 68731
rect 8987 68728 8999 68731
rect 9692 68728 9720 68827
rect 10042 68796 10048 68808
rect 10003 68768 10048 68796
rect 10042 68756 10048 68768
rect 10100 68756 10106 68808
rect 10428 68796 10456 68827
rect 10502 68824 10508 68876
rect 10560 68864 10566 68876
rect 10689 68867 10747 68873
rect 10689 68864 10701 68867
rect 10560 68836 10701 68864
rect 10560 68824 10566 68836
rect 10689 68833 10701 68836
rect 10735 68833 10747 68867
rect 12434 68864 12440 68876
rect 12395 68836 12440 68864
rect 10689 68827 10747 68833
rect 12434 68824 12440 68836
rect 12492 68824 12498 68876
rect 13906 68824 13912 68876
rect 13964 68864 13970 68876
rect 14001 68867 14059 68873
rect 14001 68864 14013 68867
rect 13964 68836 14013 68864
rect 13964 68824 13970 68836
rect 14001 68833 14013 68836
rect 14047 68833 14059 68867
rect 14001 68827 14059 68833
rect 14369 68799 14427 68805
rect 10428 68768 10732 68796
rect 10704 68740 10732 68768
rect 14369 68765 14381 68799
rect 14415 68796 14427 68799
rect 15010 68796 15016 68808
rect 14415 68768 15016 68796
rect 14415 68765 14427 68768
rect 14369 68759 14427 68765
rect 15010 68756 15016 68768
rect 15068 68756 15074 68808
rect 15930 68756 15936 68808
rect 15988 68796 15994 68808
rect 16114 68796 16120 68808
rect 15988 68768 16120 68796
rect 15988 68756 15994 68768
rect 16114 68756 16120 68768
rect 16172 68756 16178 68808
rect 9950 68728 9956 68740
rect 8987 68700 9956 68728
rect 8987 68697 8999 68700
rect 8941 68691 8999 68697
rect 9950 68688 9956 68700
rect 10008 68688 10014 68740
rect 10686 68688 10692 68740
rect 10744 68688 10750 68740
rect 1762 68620 1768 68672
rect 1820 68660 1826 68672
rect 2130 68660 2136 68672
rect 1820 68632 2136 68660
rect 1820 68620 1826 68632
rect 2130 68620 2136 68632
rect 2188 68660 2194 68672
rect 2961 68663 3019 68669
rect 2961 68660 2973 68663
rect 2188 68632 2973 68660
rect 2188 68620 2194 68632
rect 2961 68629 2973 68632
rect 3007 68629 3019 68663
rect 2961 68623 3019 68629
rect 3421 68663 3479 68669
rect 3421 68629 3433 68663
rect 3467 68660 3479 68663
rect 3602 68660 3608 68672
rect 3467 68632 3608 68660
rect 3467 68629 3479 68632
rect 3421 68623 3479 68629
rect 3602 68620 3608 68632
rect 3660 68620 3666 68672
rect 6086 68620 6092 68672
rect 6144 68660 6150 68672
rect 6546 68660 6552 68672
rect 6144 68632 6552 68660
rect 6144 68620 6150 68632
rect 6546 68620 6552 68632
rect 6604 68620 6610 68672
rect 7285 68663 7343 68669
rect 7285 68629 7297 68663
rect 7331 68660 7343 68663
rect 7374 68660 7380 68672
rect 7331 68632 7380 68660
rect 7331 68629 7343 68632
rect 7285 68623 7343 68629
rect 7374 68620 7380 68632
rect 7432 68620 7438 68672
rect 9214 68660 9220 68672
rect 9175 68632 9220 68660
rect 9214 68620 9220 68632
rect 9272 68660 9278 68672
rect 9858 68660 9864 68672
rect 9272 68632 9864 68660
rect 9272 68620 9278 68632
rect 9858 68620 9864 68632
rect 9916 68620 9922 68672
rect 11241 68663 11299 68669
rect 11241 68629 11253 68663
rect 11287 68660 11299 68663
rect 11422 68660 11428 68672
rect 11287 68632 11428 68660
rect 11287 68629 11299 68632
rect 11241 68623 11299 68629
rect 11422 68620 11428 68632
rect 11480 68620 11486 68672
rect 11606 68660 11612 68672
rect 11567 68632 11612 68660
rect 11606 68620 11612 68632
rect 11664 68620 11670 68672
rect 12066 68660 12072 68672
rect 12027 68632 12072 68660
rect 12066 68620 12072 68632
rect 12124 68620 12130 68672
rect 12618 68660 12624 68672
rect 12579 68632 12624 68660
rect 12618 68620 12624 68632
rect 12676 68620 12682 68672
rect 12802 68620 12808 68672
rect 12860 68660 12866 68672
rect 12897 68663 12955 68669
rect 12897 68660 12909 68663
rect 12860 68632 12909 68660
rect 12860 68620 12866 68632
rect 12897 68629 12909 68632
rect 12943 68629 12955 68663
rect 13354 68660 13360 68672
rect 13315 68632 13360 68660
rect 12897 68623 12955 68629
rect 13354 68620 13360 68632
rect 13412 68620 13418 68672
rect 16114 68660 16120 68672
rect 16075 68632 16120 68660
rect 16114 68620 16120 68632
rect 16172 68620 16178 68672
rect 1104 68570 18860 68592
rect 1104 68518 4315 68570
rect 4367 68518 4379 68570
rect 4431 68518 4443 68570
rect 4495 68518 4507 68570
rect 4559 68518 10982 68570
rect 11034 68518 11046 68570
rect 11098 68518 11110 68570
rect 11162 68518 11174 68570
rect 11226 68518 17648 68570
rect 17700 68518 17712 68570
rect 17764 68518 17776 68570
rect 17828 68518 17840 68570
rect 17892 68518 18860 68570
rect 1104 68496 18860 68518
rect 6730 68456 6736 68468
rect 6691 68428 6736 68456
rect 6730 68416 6736 68428
rect 6788 68416 6794 68468
rect 7469 68459 7527 68465
rect 7469 68425 7481 68459
rect 7515 68456 7527 68459
rect 8570 68456 8576 68468
rect 7515 68428 8576 68456
rect 7515 68425 7527 68428
rect 7469 68419 7527 68425
rect 8570 68416 8576 68428
rect 8628 68416 8634 68468
rect 17494 68456 17500 68468
rect 17455 68428 17500 68456
rect 17494 68416 17500 68428
rect 17552 68416 17558 68468
rect 7101 68391 7159 68397
rect 7101 68357 7113 68391
rect 7147 68388 7159 68391
rect 7926 68388 7932 68400
rect 7147 68360 7932 68388
rect 7147 68357 7159 68360
rect 7101 68351 7159 68357
rect 7926 68348 7932 68360
rect 7984 68348 7990 68400
rect 9950 68348 9956 68400
rect 10008 68388 10014 68400
rect 10318 68388 10324 68400
rect 10008 68360 10324 68388
rect 10008 68348 10014 68360
rect 10318 68348 10324 68360
rect 10376 68348 10382 68400
rect 10778 68348 10784 68400
rect 10836 68388 10842 68400
rect 11238 68388 11244 68400
rect 10836 68360 11244 68388
rect 10836 68348 10842 68360
rect 11238 68348 11244 68360
rect 11296 68348 11302 68400
rect 11330 68348 11336 68400
rect 11388 68388 11394 68400
rect 11388 68360 11744 68388
rect 11388 68348 11394 68360
rect 1486 68320 1492 68332
rect 1447 68292 1492 68320
rect 1486 68280 1492 68292
rect 1544 68280 1550 68332
rect 1762 68320 1768 68332
rect 1723 68292 1768 68320
rect 1762 68280 1768 68292
rect 1820 68280 1826 68332
rect 3881 68323 3939 68329
rect 3881 68289 3893 68323
rect 3927 68320 3939 68323
rect 4982 68320 4988 68332
rect 3927 68292 4988 68320
rect 3927 68289 3939 68292
rect 3881 68283 3939 68289
rect 4982 68280 4988 68292
rect 5040 68280 5046 68332
rect 9125 68323 9183 68329
rect 9125 68289 9137 68323
rect 9171 68320 9183 68323
rect 10686 68320 10692 68332
rect 9171 68292 10692 68320
rect 9171 68289 9183 68292
rect 9125 68283 9183 68289
rect 10686 68280 10692 68292
rect 10744 68280 10750 68332
rect 11606 68320 11612 68332
rect 11072 68292 11612 68320
rect 4065 68255 4123 68261
rect 4065 68252 4077 68255
rect 3712 68224 4077 68252
rect 2774 68144 2780 68196
rect 2832 68184 2838 68196
rect 3421 68187 3479 68193
rect 3421 68184 3433 68187
rect 2832 68156 3433 68184
rect 2832 68144 2838 68156
rect 3421 68153 3433 68156
rect 3467 68153 3479 68187
rect 3421 68147 3479 68153
rect 3712 68128 3740 68224
rect 4065 68221 4077 68224
rect 4111 68221 4123 68255
rect 4065 68215 4123 68221
rect 4341 68255 4399 68261
rect 4341 68221 4353 68255
rect 4387 68252 4399 68255
rect 5074 68252 5080 68264
rect 4387 68224 5080 68252
rect 4387 68221 4399 68224
rect 4341 68215 4399 68221
rect 5074 68212 5080 68224
rect 5132 68212 5138 68264
rect 5626 68212 5632 68264
rect 5684 68252 5690 68264
rect 6457 68255 6515 68261
rect 6457 68252 6469 68255
rect 5684 68224 6469 68252
rect 5684 68212 5690 68224
rect 6457 68221 6469 68224
rect 6503 68252 6515 68255
rect 6549 68255 6607 68261
rect 6549 68252 6561 68255
rect 6503 68224 6561 68252
rect 6503 68221 6515 68224
rect 6457 68215 6515 68221
rect 6549 68221 6561 68224
rect 6595 68221 6607 68255
rect 6549 68215 6607 68221
rect 7374 68212 7380 68264
rect 7432 68252 7438 68264
rect 11072 68261 11100 68292
rect 11606 68280 11612 68292
rect 11664 68280 11670 68332
rect 11716 68329 11744 68360
rect 11701 68323 11759 68329
rect 11701 68289 11713 68323
rect 11747 68289 11759 68323
rect 11701 68283 11759 68289
rect 16025 68323 16083 68329
rect 16025 68289 16037 68323
rect 16071 68320 16083 68323
rect 16071 68292 16436 68320
rect 16071 68289 16083 68292
rect 16025 68283 16083 68289
rect 16408 68264 16436 68292
rect 7653 68255 7711 68261
rect 7653 68252 7665 68255
rect 7432 68224 7665 68252
rect 7432 68212 7438 68224
rect 7653 68221 7665 68224
rect 7699 68221 7711 68255
rect 7653 68215 7711 68221
rect 9769 68255 9827 68261
rect 9769 68221 9781 68255
rect 9815 68221 9827 68255
rect 9769 68215 9827 68221
rect 11057 68255 11115 68261
rect 11057 68221 11069 68255
rect 11103 68221 11115 68255
rect 11057 68215 11115 68221
rect 5350 68144 5356 68196
rect 5408 68184 5414 68196
rect 5997 68187 6055 68193
rect 5997 68184 6009 68187
rect 5408 68156 6009 68184
rect 5408 68144 5414 68156
rect 5997 68153 6009 68156
rect 6043 68153 6055 68187
rect 5997 68147 6055 68153
rect 8478 68144 8484 68196
rect 8536 68184 8542 68196
rect 8846 68184 8852 68196
rect 8536 68156 8852 68184
rect 8536 68144 8542 68156
rect 8846 68144 8852 68156
rect 8904 68144 8910 68196
rect 9784 68184 9812 68215
rect 11146 68212 11152 68264
rect 11204 68252 11210 68264
rect 11422 68252 11428 68264
rect 11204 68224 11428 68252
rect 11204 68212 11210 68224
rect 11422 68212 11428 68224
rect 11480 68212 11486 68264
rect 11517 68255 11575 68261
rect 11517 68221 11529 68255
rect 11563 68252 11575 68255
rect 12618 68252 12624 68264
rect 11563 68224 12624 68252
rect 11563 68221 11575 68224
rect 11517 68215 11575 68221
rect 10134 68184 10140 68196
rect 9784 68156 10140 68184
rect 10134 68144 10140 68156
rect 10192 68184 10198 68196
rect 10321 68187 10379 68193
rect 10321 68184 10333 68187
rect 10192 68156 10333 68184
rect 10192 68144 10198 68156
rect 10321 68153 10333 68156
rect 10367 68184 10379 68187
rect 10778 68184 10784 68196
rect 10367 68156 10784 68184
rect 10367 68153 10379 68156
rect 10321 68147 10379 68153
rect 10778 68144 10784 68156
rect 10836 68144 10842 68196
rect 2866 68116 2872 68128
rect 2827 68088 2872 68116
rect 2866 68076 2872 68088
rect 2924 68076 2930 68128
rect 3694 68076 3700 68128
rect 3752 68076 3758 68128
rect 3878 68076 3884 68128
rect 3936 68116 3942 68128
rect 5445 68119 5503 68125
rect 5445 68116 5457 68119
rect 3936 68088 5457 68116
rect 3936 68076 3942 68088
rect 5445 68085 5457 68088
rect 5491 68085 5503 68119
rect 8018 68116 8024 68128
rect 7979 68088 8024 68116
rect 5445 68079 5503 68085
rect 8018 68076 8024 68088
rect 8076 68076 8082 68128
rect 8386 68076 8392 68128
rect 8444 68116 8450 68128
rect 8665 68119 8723 68125
rect 8665 68116 8677 68119
rect 8444 68088 8677 68116
rect 8444 68076 8450 68088
rect 8665 68085 8677 68088
rect 8711 68085 8723 68119
rect 9490 68116 9496 68128
rect 9451 68088 9496 68116
rect 8665 68079 8723 68085
rect 9490 68076 9496 68088
rect 9548 68076 9554 68128
rect 9766 68076 9772 68128
rect 9824 68116 9830 68128
rect 9953 68119 10011 68125
rect 9953 68116 9965 68119
rect 9824 68088 9965 68116
rect 9824 68076 9830 68088
rect 9953 68085 9965 68088
rect 9999 68085 10011 68119
rect 9953 68079 10011 68085
rect 10689 68119 10747 68125
rect 10689 68085 10701 68119
rect 10735 68116 10747 68119
rect 11330 68116 11336 68128
rect 10735 68088 11336 68116
rect 10735 68085 10747 68088
rect 10689 68079 10747 68085
rect 11330 68076 11336 68088
rect 11388 68116 11394 68128
rect 11532 68116 11560 68215
rect 12618 68212 12624 68224
rect 12676 68212 12682 68264
rect 12802 68252 12808 68264
rect 12763 68224 12808 68252
rect 12802 68212 12808 68224
rect 12860 68212 12866 68264
rect 13170 68252 13176 68264
rect 13131 68224 13176 68252
rect 13170 68212 13176 68224
rect 13228 68212 13234 68264
rect 13354 68252 13360 68264
rect 13315 68224 13360 68252
rect 13354 68212 13360 68224
rect 13412 68212 13418 68264
rect 16114 68252 16120 68264
rect 16075 68224 16120 68252
rect 16114 68212 16120 68224
rect 16172 68212 16178 68264
rect 16390 68252 16396 68264
rect 16351 68224 16396 68252
rect 16390 68212 16396 68224
rect 16448 68212 16454 68264
rect 12434 68116 12440 68128
rect 11388 68088 11560 68116
rect 12395 68088 12440 68116
rect 11388 68076 11394 68088
rect 12434 68076 12440 68088
rect 12492 68076 12498 68128
rect 13906 68116 13912 68128
rect 13867 68088 13912 68116
rect 13906 68076 13912 68088
rect 13964 68076 13970 68128
rect 14090 68076 14096 68128
rect 14148 68116 14154 68128
rect 14277 68119 14335 68125
rect 14277 68116 14289 68119
rect 14148 68088 14289 68116
rect 14148 68076 14154 68088
rect 14277 68085 14289 68088
rect 14323 68116 14335 68119
rect 15102 68116 15108 68128
rect 14323 68088 15108 68116
rect 14323 68085 14335 68088
rect 14277 68079 14335 68085
rect 15102 68076 15108 68088
rect 15160 68076 15166 68128
rect 1104 68026 18860 68048
rect 1104 67974 7648 68026
rect 7700 67974 7712 68026
rect 7764 67974 7776 68026
rect 7828 67974 7840 68026
rect 7892 67974 14315 68026
rect 14367 67974 14379 68026
rect 14431 67974 14443 68026
rect 14495 67974 14507 68026
rect 14559 67974 18860 68026
rect 1104 67952 18860 67974
rect 1673 67915 1731 67921
rect 1673 67881 1685 67915
rect 1719 67912 1731 67915
rect 2222 67912 2228 67924
rect 1719 67884 2228 67912
rect 1719 67881 1731 67884
rect 1673 67875 1731 67881
rect 2222 67872 2228 67884
rect 2280 67872 2286 67924
rect 3513 67915 3571 67921
rect 3513 67881 3525 67915
rect 3559 67912 3571 67915
rect 3878 67912 3884 67924
rect 3559 67884 3884 67912
rect 3559 67881 3571 67884
rect 3513 67875 3571 67881
rect 3878 67872 3884 67884
rect 3936 67872 3942 67924
rect 4062 67912 4068 67924
rect 4023 67884 4068 67912
rect 4062 67872 4068 67884
rect 4120 67872 4126 67924
rect 4890 67912 4896 67924
rect 4851 67884 4896 67912
rect 4890 67872 4896 67884
rect 4948 67872 4954 67924
rect 7929 67915 7987 67921
rect 7929 67881 7941 67915
rect 7975 67912 7987 67915
rect 8294 67912 8300 67924
rect 7975 67884 8300 67912
rect 7975 67881 7987 67884
rect 7929 67875 7987 67881
rect 8294 67872 8300 67884
rect 8352 67872 8358 67924
rect 8386 67872 8392 67924
rect 8444 67912 8450 67924
rect 9769 67915 9827 67921
rect 9769 67912 9781 67915
rect 8444 67884 9781 67912
rect 8444 67872 8450 67884
rect 9769 67881 9781 67884
rect 9815 67912 9827 67915
rect 10410 67912 10416 67924
rect 9815 67884 10416 67912
rect 9815 67881 9827 67884
rect 9769 67875 9827 67881
rect 10410 67872 10416 67884
rect 10468 67872 10474 67924
rect 1486 67804 1492 67856
rect 1544 67844 1550 67856
rect 2498 67844 2504 67856
rect 1544 67816 2504 67844
rect 1544 67804 1550 67816
rect 2498 67804 2504 67816
rect 2556 67844 2562 67856
rect 3053 67847 3111 67853
rect 3053 67844 3065 67847
rect 2556 67816 3065 67844
rect 2556 67804 2562 67816
rect 3053 67813 3065 67816
rect 3099 67813 3111 67847
rect 7561 67847 7619 67853
rect 7561 67844 7573 67847
rect 3053 67807 3111 67813
rect 5460 67816 7573 67844
rect 2593 67779 2651 67785
rect 2593 67745 2605 67779
rect 2639 67776 2651 67779
rect 2866 67776 2872 67788
rect 2639 67748 2872 67776
rect 2639 67745 2651 67748
rect 2593 67739 2651 67745
rect 2866 67736 2872 67748
rect 2924 67736 2930 67788
rect 3326 67736 3332 67788
rect 3384 67776 3390 67788
rect 3605 67779 3663 67785
rect 3605 67776 3617 67779
rect 3384 67748 3617 67776
rect 3384 67736 3390 67748
rect 3605 67745 3617 67748
rect 3651 67745 3663 67779
rect 3605 67739 3663 67745
rect 3694 67736 3700 67788
rect 3752 67776 3758 67788
rect 4062 67776 4068 67788
rect 3752 67748 4068 67776
rect 3752 67736 3758 67748
rect 4062 67736 4068 67748
rect 4120 67736 4126 67788
rect 4801 67779 4859 67785
rect 4801 67776 4813 67779
rect 4724 67748 4813 67776
rect 1762 67708 1768 67720
rect 1723 67680 1768 67708
rect 1762 67668 1768 67680
rect 1820 67668 1826 67720
rect 2314 67708 2320 67720
rect 2275 67680 2320 67708
rect 2314 67668 2320 67680
rect 2372 67668 2378 67720
rect 2774 67668 2780 67720
rect 2832 67708 2838 67720
rect 2832 67680 2877 67708
rect 2832 67668 2838 67680
rect 4724 67652 4752 67748
rect 4801 67745 4813 67748
rect 4847 67745 4859 67779
rect 4801 67739 4859 67745
rect 4890 67736 4896 67788
rect 4948 67776 4954 67788
rect 5460 67785 5488 67816
rect 7561 67813 7573 67816
rect 7607 67844 7619 67847
rect 8110 67844 8116 67856
rect 7607 67816 8116 67844
rect 7607 67813 7619 67816
rect 7561 67807 7619 67813
rect 8110 67804 8116 67816
rect 8168 67804 8174 67856
rect 10134 67804 10140 67856
rect 10192 67844 10198 67856
rect 10229 67847 10287 67853
rect 10229 67844 10241 67847
rect 10192 67816 10241 67844
rect 10192 67804 10198 67816
rect 10229 67813 10241 67816
rect 10275 67844 10287 67847
rect 10318 67844 10324 67856
rect 10275 67816 10324 67844
rect 10275 67813 10287 67816
rect 10229 67807 10287 67813
rect 10318 67804 10324 67816
rect 10376 67804 10382 67856
rect 11146 67844 11152 67856
rect 10980 67816 11152 67844
rect 5445 67779 5503 67785
rect 5445 67776 5457 67779
rect 4948 67748 5457 67776
rect 4948 67736 4954 67748
rect 5445 67745 5457 67748
rect 5491 67745 5503 67779
rect 7466 67776 7472 67788
rect 7427 67748 7472 67776
rect 5445 67739 5503 67745
rect 7466 67736 7472 67748
rect 7524 67736 7530 67788
rect 8938 67736 8944 67788
rect 8996 67776 9002 67788
rect 9309 67779 9367 67785
rect 9309 67776 9321 67779
rect 8996 67748 9321 67776
rect 8996 67736 9002 67748
rect 9309 67745 9321 67748
rect 9355 67745 9367 67779
rect 9309 67739 9367 67745
rect 10597 67779 10655 67785
rect 10597 67745 10609 67779
rect 10643 67776 10655 67779
rect 10686 67776 10692 67788
rect 10643 67748 10692 67776
rect 10643 67745 10655 67748
rect 10597 67739 10655 67745
rect 10686 67736 10692 67748
rect 10744 67736 10750 67788
rect 10980 67785 11008 67816
rect 11146 67804 11152 67816
rect 11204 67844 11210 67856
rect 11606 67844 11612 67856
rect 11204 67816 11612 67844
rect 11204 67804 11210 67816
rect 11606 67804 11612 67816
rect 11664 67804 11670 67856
rect 10965 67779 11023 67785
rect 10965 67745 10977 67779
rect 11011 67745 11023 67779
rect 11330 67776 11336 67788
rect 11243 67748 11336 67776
rect 10965 67739 11023 67745
rect 11330 67736 11336 67748
rect 11388 67736 11394 67788
rect 12437 67779 12495 67785
rect 12437 67745 12449 67779
rect 12483 67745 12495 67779
rect 12437 67739 12495 67745
rect 12989 67779 13047 67785
rect 12989 67745 13001 67779
rect 13035 67745 13047 67779
rect 13170 67776 13176 67788
rect 13131 67748 13176 67776
rect 12989 67739 13047 67745
rect 5629 67711 5687 67717
rect 5629 67677 5641 67711
rect 5675 67677 5687 67711
rect 5629 67671 5687 67677
rect 3786 67640 3792 67652
rect 3747 67612 3792 67640
rect 3786 67600 3792 67612
rect 3844 67600 3850 67652
rect 4706 67640 4712 67652
rect 4667 67612 4712 67640
rect 4706 67600 4712 67612
rect 4764 67600 4770 67652
rect 5644 67640 5672 67671
rect 5460 67612 5672 67640
rect 9493 67643 9551 67649
rect 5166 67532 5172 67584
rect 5224 67572 5230 67584
rect 5460 67572 5488 67612
rect 9493 67609 9505 67643
rect 9539 67640 9551 67643
rect 9539 67612 9628 67640
rect 9539 67609 9551 67612
rect 9493 67603 9551 67609
rect 6178 67572 6184 67584
rect 5224 67544 5488 67572
rect 6139 67544 6184 67572
rect 5224 67532 5230 67544
rect 6178 67532 6184 67544
rect 6236 67532 6242 67584
rect 8018 67532 8024 67584
rect 8076 67572 8082 67584
rect 8205 67575 8263 67581
rect 8205 67572 8217 67575
rect 8076 67544 8217 67572
rect 8076 67532 8082 67544
rect 8205 67541 8217 67544
rect 8251 67541 8263 67575
rect 9600 67572 9628 67612
rect 11348 67584 11376 67736
rect 11517 67711 11575 67717
rect 11517 67677 11529 67711
rect 11563 67708 11575 67711
rect 12161 67711 12219 67717
rect 12161 67708 12173 67711
rect 11563 67680 12173 67708
rect 11563 67677 11575 67680
rect 11517 67671 11575 67677
rect 12161 67677 12173 67680
rect 12207 67708 12219 67711
rect 12452 67708 12480 67739
rect 12207 67680 12480 67708
rect 13004 67708 13032 67739
rect 13170 67736 13176 67748
rect 13228 67736 13234 67788
rect 15286 67736 15292 67788
rect 15344 67776 15350 67788
rect 15749 67779 15807 67785
rect 15749 67776 15761 67779
rect 15344 67748 15761 67776
rect 15344 67736 15350 67748
rect 15749 67745 15761 67748
rect 15795 67745 15807 67779
rect 15749 67739 15807 67745
rect 13722 67708 13728 67720
rect 13004 67680 13728 67708
rect 12207 67677 12219 67680
rect 12161 67671 12219 67677
rect 13722 67668 13728 67680
rect 13780 67668 13786 67720
rect 15473 67711 15531 67717
rect 15473 67677 15485 67711
rect 15519 67708 15531 67711
rect 15930 67708 15936 67720
rect 15519 67680 15936 67708
rect 15519 67677 15531 67680
rect 15473 67671 15531 67677
rect 15930 67668 15936 67680
rect 15988 67668 15994 67720
rect 17126 67708 17132 67720
rect 17087 67680 17132 67708
rect 17126 67668 17132 67680
rect 17184 67668 17190 67720
rect 9858 67572 9864 67584
rect 9600 67544 9864 67572
rect 8205 67535 8263 67541
rect 9858 67532 9864 67544
rect 9916 67572 9922 67584
rect 10870 67572 10876 67584
rect 9916 67544 10876 67572
rect 9916 67532 9922 67544
rect 10870 67532 10876 67544
rect 10928 67532 10934 67584
rect 11330 67532 11336 67584
rect 11388 67532 11394 67584
rect 12529 67575 12587 67581
rect 12529 67541 12541 67575
rect 12575 67572 12587 67575
rect 13078 67572 13084 67584
rect 12575 67544 13084 67572
rect 12575 67541 12587 67544
rect 12529 67535 12587 67541
rect 13078 67532 13084 67544
rect 13136 67532 13142 67584
rect 1104 67482 18860 67504
rect 1104 67430 4315 67482
rect 4367 67430 4379 67482
rect 4431 67430 4443 67482
rect 4495 67430 4507 67482
rect 4559 67430 10982 67482
rect 11034 67430 11046 67482
rect 11098 67430 11110 67482
rect 11162 67430 11174 67482
rect 11226 67430 17648 67482
rect 17700 67430 17712 67482
rect 17764 67430 17776 67482
rect 17828 67430 17840 67482
rect 17892 67430 18860 67482
rect 1104 67408 18860 67430
rect 2866 67368 2872 67380
rect 2827 67340 2872 67368
rect 2866 67328 2872 67340
rect 2924 67328 2930 67380
rect 4890 67368 4896 67380
rect 4851 67340 4896 67368
rect 4890 67328 4896 67340
rect 4948 67328 4954 67380
rect 6730 67368 6736 67380
rect 6691 67340 6736 67368
rect 6730 67328 6736 67340
rect 6788 67328 6794 67380
rect 6914 67328 6920 67380
rect 6972 67368 6978 67380
rect 7285 67371 7343 67377
rect 7285 67368 7297 67371
rect 6972 67340 7297 67368
rect 6972 67328 6978 67340
rect 7285 67337 7297 67340
rect 7331 67337 7343 67371
rect 7285 67331 7343 67337
rect 13170 67328 13176 67380
rect 13228 67368 13234 67380
rect 13633 67371 13691 67377
rect 13633 67368 13645 67371
rect 13228 67340 13645 67368
rect 13228 67328 13234 67340
rect 13633 67337 13645 67340
rect 13679 67337 13691 67371
rect 13633 67331 13691 67337
rect 3970 67192 3976 67244
rect 4028 67232 4034 67244
rect 5353 67235 5411 67241
rect 5353 67232 5365 67235
rect 4028 67204 5365 67232
rect 4028 67192 4034 67204
rect 5353 67201 5365 67204
rect 5399 67201 5411 67235
rect 5353 67195 5411 67201
rect 6365 67235 6423 67241
rect 6365 67201 6377 67235
rect 6411 67232 6423 67235
rect 6748 67232 6776 67328
rect 14366 67300 14372 67312
rect 14327 67272 14372 67300
rect 14366 67260 14372 67272
rect 14424 67260 14430 67312
rect 8205 67235 8263 67241
rect 8205 67232 8217 67235
rect 6411 67204 6776 67232
rect 7208 67204 8217 67232
rect 6411 67201 6423 67204
rect 6365 67195 6423 67201
rect 7208 67176 7236 67204
rect 8205 67201 8217 67204
rect 8251 67201 8263 67235
rect 10502 67232 10508 67244
rect 10463 67204 10508 67232
rect 8205 67195 8263 67201
rect 10502 67192 10508 67204
rect 10560 67192 10566 67244
rect 11974 67192 11980 67244
rect 12032 67232 12038 67244
rect 16025 67235 16083 67241
rect 12032 67204 12572 67232
rect 12032 67192 12038 67204
rect 1854 67164 1860 67176
rect 1815 67136 1860 67164
rect 1854 67124 1860 67136
rect 1912 67124 1918 67176
rect 4246 67164 4252 67176
rect 4159 67136 4252 67164
rect 4246 67124 4252 67136
rect 4304 67164 4310 67176
rect 5626 67164 5632 67176
rect 4304 67136 5632 67164
rect 4304 67124 4310 67136
rect 5626 67124 5632 67136
rect 5684 67124 5690 67176
rect 5902 67164 5908 67176
rect 5863 67136 5908 67164
rect 5902 67124 5908 67136
rect 5960 67124 5966 67176
rect 6178 67164 6184 67176
rect 6091 67136 6184 67164
rect 6178 67124 6184 67136
rect 6236 67124 6242 67176
rect 7190 67164 7196 67176
rect 7151 67136 7196 67164
rect 7190 67124 7196 67136
rect 7248 67124 7254 67176
rect 7929 67167 7987 67173
rect 7929 67133 7941 67167
rect 7975 67164 7987 67167
rect 8018 67164 8024 67176
rect 7975 67136 8024 67164
rect 7975 67133 7987 67136
rect 7929 67127 7987 67133
rect 2225 67099 2283 67105
rect 2225 67065 2237 67099
rect 2271 67096 2283 67099
rect 6196 67096 6224 67124
rect 6822 67096 6828 67108
rect 2271 67068 3372 67096
rect 2271 67065 2283 67068
rect 2225 67059 2283 67065
rect 3344 67040 3372 67068
rect 4448 67068 5212 67096
rect 6196 67068 6828 67096
rect 2593 67031 2651 67037
rect 2593 66997 2605 67031
rect 2639 67028 2651 67031
rect 2774 67028 2780 67040
rect 2639 67000 2780 67028
rect 2639 66997 2651 67000
rect 2593 66991 2651 66997
rect 2774 66988 2780 67000
rect 2832 66988 2838 67040
rect 3326 66988 3332 67040
rect 3384 67028 3390 67040
rect 4448 67037 4476 67068
rect 5184 67040 5212 67068
rect 6822 67056 6828 67068
rect 6880 67056 6886 67108
rect 7101 67099 7159 67105
rect 7101 67065 7113 67099
rect 7147 67096 7159 67099
rect 7944 67096 7972 67127
rect 8018 67124 8024 67136
rect 8076 67124 8082 67176
rect 9674 67164 9680 67176
rect 9635 67136 9680 67164
rect 9674 67124 9680 67136
rect 9732 67124 9738 67176
rect 10045 67167 10103 67173
rect 10045 67133 10057 67167
rect 10091 67133 10103 67167
rect 10410 67164 10416 67176
rect 10371 67136 10416 67164
rect 10045 67127 10103 67133
rect 7147 67068 7972 67096
rect 7147 67065 7159 67068
rect 7101 67059 7159 67065
rect 3605 67031 3663 67037
rect 3605 67028 3617 67031
rect 3384 67000 3617 67028
rect 3384 66988 3390 67000
rect 3605 66997 3617 67000
rect 3651 66997 3663 67031
rect 3605 66991 3663 66997
rect 4433 67031 4491 67037
rect 4433 66997 4445 67031
rect 4479 66997 4491 67031
rect 5166 67028 5172 67040
rect 5127 67000 5172 67028
rect 4433 66991 4491 66997
rect 5166 66988 5172 67000
rect 5224 66988 5230 67040
rect 7466 66988 7472 67040
rect 7524 67028 7530 67040
rect 8570 67028 8576 67040
rect 7524 67000 8576 67028
rect 7524 66988 7530 67000
rect 8570 66988 8576 67000
rect 8628 66988 8634 67040
rect 8938 66988 8944 67040
rect 8996 67028 9002 67040
rect 9033 67031 9091 67037
rect 9033 67028 9045 67031
rect 8996 67000 9045 67028
rect 8996 66988 9002 67000
rect 9033 66997 9045 67000
rect 9079 66997 9091 67031
rect 9490 67028 9496 67040
rect 9451 67000 9496 67028
rect 9033 66991 9091 66997
rect 9490 66988 9496 67000
rect 9548 67028 9554 67040
rect 10060 67028 10088 67127
rect 10410 67124 10416 67136
rect 10468 67124 10474 67176
rect 12158 67164 12164 67176
rect 12119 67136 12164 67164
rect 12158 67124 12164 67136
rect 12216 67124 12222 67176
rect 12544 67173 12572 67204
rect 16025 67201 16037 67235
rect 16071 67232 16083 67235
rect 16071 67204 16436 67232
rect 16071 67201 16083 67204
rect 16025 67195 16083 67201
rect 12529 67167 12587 67173
rect 12529 67133 12541 67167
rect 12575 67133 12587 67167
rect 12529 67127 12587 67133
rect 12897 67167 12955 67173
rect 12897 67133 12909 67167
rect 12943 67133 12955 67167
rect 12897 67127 12955 67133
rect 12250 67056 12256 67108
rect 12308 67096 12314 67108
rect 12434 67096 12440 67108
rect 12308 67068 12440 67096
rect 12308 67056 12314 67068
rect 12434 67056 12440 67068
rect 12492 67096 12498 67108
rect 12912 67096 12940 67127
rect 12986 67124 12992 67176
rect 13044 67164 13050 67176
rect 14185 67167 14243 67173
rect 14185 67164 14197 67167
rect 13044 67136 14197 67164
rect 13044 67124 13050 67136
rect 14185 67133 14197 67136
rect 14231 67164 14243 67167
rect 14645 67167 14703 67173
rect 14645 67164 14657 67167
rect 14231 67136 14657 67164
rect 14231 67133 14243 67136
rect 14185 67127 14243 67133
rect 14645 67133 14657 67136
rect 14691 67133 14703 67167
rect 14645 67127 14703 67133
rect 15105 67167 15163 67173
rect 15105 67133 15117 67167
rect 15151 67164 15163 67167
rect 15378 67164 15384 67176
rect 15151 67136 15384 67164
rect 15151 67133 15163 67136
rect 15105 67127 15163 67133
rect 15378 67124 15384 67136
rect 15436 67164 15442 67176
rect 15930 67164 15936 67176
rect 15436 67136 15936 67164
rect 15436 67124 15442 67136
rect 15930 67124 15936 67136
rect 15988 67164 15994 67176
rect 16408 67173 16436 67204
rect 16117 67167 16175 67173
rect 16117 67164 16129 67167
rect 15988 67136 16129 67164
rect 15988 67124 15994 67136
rect 16117 67133 16129 67136
rect 16163 67133 16175 67167
rect 16117 67127 16175 67133
rect 16393 67167 16451 67173
rect 16393 67133 16405 67167
rect 16439 67164 16451 67167
rect 16482 67164 16488 67176
rect 16439 67136 16488 67164
rect 16439 67133 16451 67136
rect 16393 67127 16451 67133
rect 16482 67124 16488 67136
rect 16540 67124 16546 67176
rect 13262 67096 13268 67108
rect 12492 67068 12940 67096
rect 13223 67068 13268 67096
rect 12492 67056 12498 67068
rect 13262 67056 13268 67068
rect 13320 67056 13326 67108
rect 9548 67000 10088 67028
rect 11241 67031 11299 67037
rect 9548 66988 9554 67000
rect 11241 66997 11253 67031
rect 11287 67028 11299 67031
rect 11330 67028 11336 67040
rect 11287 67000 11336 67028
rect 11287 66997 11299 67000
rect 11241 66991 11299 66997
rect 11330 66988 11336 67000
rect 11388 66988 11394 67040
rect 11606 67028 11612 67040
rect 11567 67000 11612 67028
rect 11606 66988 11612 67000
rect 11664 66988 11670 67040
rect 11974 67028 11980 67040
rect 11935 67000 11980 67028
rect 11974 66988 11980 67000
rect 12032 66988 12038 67040
rect 13814 66988 13820 67040
rect 13872 67028 13878 67040
rect 14001 67031 14059 67037
rect 14001 67028 14013 67031
rect 13872 67000 14013 67028
rect 13872 66988 13878 67000
rect 14001 66997 14013 67000
rect 14047 66997 14059 67031
rect 14001 66991 14059 66997
rect 15286 66988 15292 67040
rect 15344 67028 15350 67040
rect 15473 67031 15531 67037
rect 15473 67028 15485 67031
rect 15344 67000 15485 67028
rect 15344 66988 15350 67000
rect 15473 66997 15485 67000
rect 15519 66997 15531 67031
rect 17494 67028 17500 67040
rect 17455 67000 17500 67028
rect 15473 66991 15531 66997
rect 17494 66988 17500 67000
rect 17552 66988 17558 67040
rect 1104 66938 18860 66960
rect 1104 66886 7648 66938
rect 7700 66886 7712 66938
rect 7764 66886 7776 66938
rect 7828 66886 7840 66938
rect 7892 66886 14315 66938
rect 14367 66886 14379 66938
rect 14431 66886 14443 66938
rect 14495 66886 14507 66938
rect 14559 66886 18860 66938
rect 1104 66864 18860 66886
rect 2041 66827 2099 66833
rect 2041 66793 2053 66827
rect 2087 66824 2099 66827
rect 2314 66824 2320 66836
rect 2087 66796 2320 66824
rect 2087 66793 2099 66796
rect 2041 66787 2099 66793
rect 2314 66784 2320 66796
rect 2372 66824 2378 66836
rect 2501 66827 2559 66833
rect 2501 66824 2513 66827
rect 2372 66796 2513 66824
rect 2372 66784 2378 66796
rect 2501 66793 2513 66796
rect 2547 66793 2559 66827
rect 2501 66787 2559 66793
rect 2866 66784 2872 66836
rect 2924 66824 2930 66836
rect 3789 66827 3847 66833
rect 3789 66824 3801 66827
rect 2924 66796 3801 66824
rect 2924 66784 2930 66796
rect 3789 66793 3801 66796
rect 3835 66824 3847 66827
rect 4246 66824 4252 66836
rect 3835 66796 4252 66824
rect 3835 66793 3847 66796
rect 3789 66787 3847 66793
rect 4246 66784 4252 66796
rect 4304 66784 4310 66836
rect 8570 66784 8576 66836
rect 8628 66824 8634 66836
rect 9309 66827 9367 66833
rect 9309 66824 9321 66827
rect 8628 66796 9321 66824
rect 8628 66784 8634 66796
rect 9309 66793 9321 66796
rect 9355 66824 9367 66827
rect 9674 66824 9680 66836
rect 9355 66796 9680 66824
rect 9355 66793 9367 66796
rect 9309 66787 9367 66793
rect 9674 66784 9680 66796
rect 9732 66784 9738 66836
rect 15930 66784 15936 66836
rect 15988 66824 15994 66836
rect 16945 66827 17003 66833
rect 16945 66824 16957 66827
rect 15988 66796 16957 66824
rect 15988 66784 15994 66796
rect 16945 66793 16957 66796
rect 16991 66793 17003 66827
rect 16945 66787 17003 66793
rect 2130 66716 2136 66768
rect 2188 66756 2194 66768
rect 2225 66759 2283 66765
rect 2225 66756 2237 66759
rect 2188 66728 2237 66756
rect 2188 66716 2194 66728
rect 2225 66725 2237 66728
rect 2271 66725 2283 66759
rect 2225 66719 2283 66725
rect 11974 66716 11980 66768
rect 12032 66756 12038 66768
rect 12032 66728 13216 66756
rect 12032 66716 12038 66728
rect 2409 66691 2467 66697
rect 2409 66657 2421 66691
rect 2455 66688 2467 66691
rect 2590 66688 2596 66700
rect 2455 66660 2596 66688
rect 2455 66657 2467 66660
rect 2409 66651 2467 66657
rect 2590 66648 2596 66660
rect 2648 66648 2654 66700
rect 3326 66648 3332 66700
rect 3384 66688 3390 66700
rect 3605 66691 3663 66697
rect 3605 66688 3617 66691
rect 3384 66660 3617 66688
rect 3384 66648 3390 66660
rect 3605 66657 3617 66660
rect 3651 66657 3663 66691
rect 5258 66688 5264 66700
rect 5219 66660 5264 66688
rect 3605 66651 3663 66657
rect 5258 66648 5264 66660
rect 5316 66648 5322 66700
rect 5626 66648 5632 66700
rect 5684 66688 5690 66700
rect 5813 66691 5871 66697
rect 5813 66688 5825 66691
rect 5684 66660 5825 66688
rect 5684 66648 5690 66660
rect 5813 66657 5825 66660
rect 5859 66688 5871 66691
rect 6546 66688 6552 66700
rect 5859 66660 6552 66688
rect 5859 66657 5871 66660
rect 5813 66651 5871 66657
rect 6546 66648 6552 66660
rect 6604 66648 6610 66700
rect 6730 66648 6736 66700
rect 6788 66688 6794 66700
rect 7098 66688 7104 66700
rect 6788 66660 7104 66688
rect 6788 66648 6794 66660
rect 7098 66648 7104 66660
rect 7156 66648 7162 66700
rect 7466 66688 7472 66700
rect 7427 66660 7472 66688
rect 7466 66648 7472 66660
rect 7524 66688 7530 66700
rect 8202 66688 8208 66700
rect 7524 66660 8208 66688
rect 7524 66648 7530 66660
rect 8202 66648 8208 66660
rect 8260 66648 8266 66700
rect 8481 66691 8539 66697
rect 8481 66657 8493 66691
rect 8527 66688 8539 66691
rect 9122 66688 9128 66700
rect 8527 66660 9128 66688
rect 8527 66657 8539 66660
rect 8481 66651 8539 66657
rect 9122 66648 9128 66660
rect 9180 66648 9186 66700
rect 9582 66688 9588 66700
rect 9543 66660 9588 66688
rect 9582 66648 9588 66660
rect 9640 66648 9646 66700
rect 9858 66688 9864 66700
rect 9819 66660 9864 66688
rect 9858 66648 9864 66660
rect 9916 66648 9922 66700
rect 10229 66691 10287 66697
rect 10229 66657 10241 66691
rect 10275 66657 10287 66691
rect 10229 66651 10287 66657
rect 5537 66623 5595 66629
rect 5537 66589 5549 66623
rect 5583 66620 5595 66623
rect 5902 66620 5908 66632
rect 5583 66592 5908 66620
rect 5583 66589 5595 66592
rect 5537 66583 5595 66589
rect 5902 66580 5908 66592
rect 5960 66620 5966 66632
rect 6181 66623 6239 66629
rect 6181 66620 6193 66623
rect 5960 66592 6193 66620
rect 5960 66580 5966 66592
rect 6181 66589 6193 66592
rect 6227 66589 6239 66623
rect 9674 66620 9680 66632
rect 9635 66592 9680 66620
rect 6181 66583 6239 66589
rect 9674 66580 9680 66592
rect 9732 66580 9738 66632
rect 5074 66512 5080 66564
rect 5132 66552 5138 66564
rect 5994 66552 6000 66564
rect 5132 66524 6000 66552
rect 5132 66512 5138 66524
rect 5994 66512 6000 66524
rect 6052 66512 6058 66564
rect 8665 66555 8723 66561
rect 8665 66521 8677 66555
rect 8711 66552 8723 66555
rect 9214 66552 9220 66564
rect 8711 66524 9220 66552
rect 8711 66521 8723 66524
rect 8665 66515 8723 66521
rect 9214 66512 9220 66524
rect 9272 66552 9278 66564
rect 10244 66552 10272 66651
rect 12434 66648 12440 66700
rect 12492 66688 12498 66700
rect 12894 66688 12900 66700
rect 12492 66660 12537 66688
rect 12855 66660 12900 66688
rect 12492 66648 12498 66660
rect 12894 66648 12900 66660
rect 12952 66648 12958 66700
rect 13188 66697 13216 66728
rect 13173 66691 13231 66697
rect 13173 66657 13185 66691
rect 13219 66657 13231 66691
rect 13173 66651 13231 66657
rect 14366 66648 14372 66700
rect 14424 66688 14430 66700
rect 15013 66691 15071 66697
rect 15013 66688 15025 66691
rect 14424 66660 15025 66688
rect 14424 66648 14430 66660
rect 15013 66657 15025 66660
rect 15059 66688 15071 66691
rect 16114 66688 16120 66700
rect 15059 66660 16120 66688
rect 15059 66657 15071 66660
rect 15013 66651 15071 66657
rect 16114 66648 16120 66660
rect 16172 66648 16178 66700
rect 11885 66623 11943 66629
rect 11885 66589 11897 66623
rect 11931 66620 11943 66623
rect 12158 66620 12164 66632
rect 11931 66592 12164 66620
rect 11931 66589 11943 66592
rect 11885 66583 11943 66589
rect 12158 66580 12164 66592
rect 12216 66580 12222 66632
rect 12526 66580 12532 66632
rect 12584 66620 12590 66632
rect 12986 66620 12992 66632
rect 12584 66592 12992 66620
rect 12584 66580 12590 66592
rect 12986 66580 12992 66592
rect 13044 66580 13050 66632
rect 15194 66580 15200 66632
rect 15252 66620 15258 66632
rect 15289 66623 15347 66629
rect 15289 66620 15301 66623
rect 15252 66592 15301 66620
rect 15252 66580 15258 66592
rect 15289 66589 15301 66592
rect 15335 66589 15347 66623
rect 16666 66620 16672 66632
rect 16627 66592 16672 66620
rect 15289 66583 15347 66589
rect 16666 66580 16672 66592
rect 16724 66580 16730 66632
rect 10410 66552 10416 66564
rect 9272 66524 10416 66552
rect 9272 66512 9278 66524
rect 10410 66512 10416 66524
rect 10468 66512 10474 66564
rect 1673 66487 1731 66493
rect 1673 66453 1685 66487
rect 1719 66484 1731 66487
rect 1854 66484 1860 66496
rect 1719 66456 1860 66484
rect 1719 66453 1731 66456
rect 1673 66447 1731 66453
rect 1854 66444 1860 66456
rect 1912 66444 1918 66496
rect 4985 66487 5043 66493
rect 4985 66453 4997 66487
rect 5031 66484 5043 66487
rect 5166 66484 5172 66496
rect 5031 66456 5172 66484
rect 5031 66453 5043 66456
rect 4985 66447 5043 66453
rect 5166 66444 5172 66456
rect 5224 66444 5230 66496
rect 6641 66487 6699 66493
rect 6641 66453 6653 66487
rect 6687 66484 6699 66487
rect 6822 66484 6828 66496
rect 6687 66456 6828 66484
rect 6687 66453 6699 66456
rect 6641 66447 6699 66453
rect 6822 66444 6828 66456
rect 6880 66444 6886 66496
rect 7101 66487 7159 66493
rect 7101 66453 7113 66487
rect 7147 66484 7159 66487
rect 7282 66484 7288 66496
rect 7147 66456 7288 66484
rect 7147 66453 7159 66456
rect 7101 66447 7159 66453
rect 7282 66444 7288 66456
rect 7340 66444 7346 66496
rect 7653 66487 7711 66493
rect 7653 66453 7665 66487
rect 7699 66484 7711 66487
rect 8202 66484 8208 66496
rect 7699 66456 8208 66484
rect 7699 66453 7711 66456
rect 7653 66447 7711 66453
rect 8202 66444 8208 66456
rect 8260 66444 8266 66496
rect 10686 66444 10692 66496
rect 10744 66484 10750 66496
rect 11057 66487 11115 66493
rect 11057 66484 11069 66487
rect 10744 66456 11069 66484
rect 10744 66444 10750 66456
rect 11057 66453 11069 66456
rect 11103 66453 11115 66487
rect 12250 66484 12256 66496
rect 12211 66456 12256 66484
rect 11057 66447 11115 66453
rect 12250 66444 12256 66456
rect 12308 66444 12314 66496
rect 12526 66484 12532 66496
rect 12487 66456 12532 66484
rect 12526 66444 12532 66456
rect 12584 66444 12590 66496
rect 1104 66394 18860 66416
rect 1104 66342 4315 66394
rect 4367 66342 4379 66394
rect 4431 66342 4443 66394
rect 4495 66342 4507 66394
rect 4559 66342 10982 66394
rect 11034 66342 11046 66394
rect 11098 66342 11110 66394
rect 11162 66342 11174 66394
rect 11226 66342 17648 66394
rect 17700 66342 17712 66394
rect 17764 66342 17776 66394
rect 17828 66342 17840 66394
rect 17892 66342 18860 66394
rect 1104 66320 18860 66342
rect 1765 66283 1823 66289
rect 1765 66249 1777 66283
rect 1811 66280 1823 66283
rect 2501 66283 2559 66289
rect 2501 66280 2513 66283
rect 1811 66252 2513 66280
rect 1811 66249 1823 66252
rect 1765 66243 1823 66249
rect 2501 66249 2513 66252
rect 2547 66280 2559 66283
rect 2590 66280 2596 66292
rect 2547 66252 2596 66280
rect 2547 66249 2559 66252
rect 2501 66243 2559 66249
rect 2590 66240 2596 66252
rect 2648 66240 2654 66292
rect 2866 66280 2872 66292
rect 2827 66252 2872 66280
rect 2866 66240 2872 66252
rect 2924 66240 2930 66292
rect 5166 66240 5172 66292
rect 5224 66280 5230 66292
rect 6825 66283 6883 66289
rect 5224 66252 5488 66280
rect 5224 66240 5230 66252
rect 3418 66172 3424 66224
rect 3476 66212 3482 66224
rect 4985 66215 5043 66221
rect 4985 66212 4997 66215
rect 3476 66184 4997 66212
rect 3476 66172 3482 66184
rect 4985 66181 4997 66184
rect 5031 66181 5043 66215
rect 5460 66212 5488 66252
rect 6825 66249 6837 66283
rect 6871 66280 6883 66283
rect 7466 66280 7472 66292
rect 6871 66252 7472 66280
rect 6871 66249 6883 66252
rect 6825 66243 6883 66249
rect 7466 66240 7472 66252
rect 7524 66240 7530 66292
rect 9490 66240 9496 66292
rect 9548 66280 9554 66292
rect 10042 66280 10048 66292
rect 9548 66252 10048 66280
rect 9548 66240 9554 66252
rect 10042 66240 10048 66252
rect 10100 66240 10106 66292
rect 13998 66240 14004 66292
rect 14056 66280 14062 66292
rect 14366 66280 14372 66292
rect 14056 66252 14372 66280
rect 14056 66240 14062 66252
rect 14366 66240 14372 66252
rect 14424 66240 14430 66292
rect 5460 66184 5764 66212
rect 4985 66175 5043 66181
rect 4433 66147 4491 66153
rect 4433 66113 4445 66147
rect 4479 66144 4491 66147
rect 5626 66144 5632 66156
rect 4479 66116 5632 66144
rect 4479 66113 4491 66116
rect 4433 66107 4491 66113
rect 5626 66104 5632 66116
rect 5684 66104 5690 66156
rect 5736 66153 5764 66184
rect 9214 66172 9220 66224
rect 9272 66212 9278 66224
rect 9858 66212 9864 66224
rect 9272 66184 9864 66212
rect 9272 66172 9278 66184
rect 9858 66172 9864 66184
rect 9916 66172 9922 66224
rect 10134 66212 10140 66224
rect 10060 66184 10140 66212
rect 5721 66147 5779 66153
rect 5721 66113 5733 66147
rect 5767 66113 5779 66147
rect 5721 66107 5779 66113
rect 6457 66147 6515 66153
rect 6457 66113 6469 66147
rect 6503 66144 6515 66147
rect 6503 66116 8156 66144
rect 6503 66113 6515 66116
rect 6457 66107 6515 66113
rect 1581 66079 1639 66085
rect 1581 66045 1593 66079
rect 1627 66076 1639 66079
rect 1627 66048 1900 66076
rect 1627 66045 1639 66048
rect 1581 66039 1639 66045
rect 1872 65952 1900 66048
rect 2866 66036 2872 66088
rect 2924 66076 2930 66088
rect 2961 66079 3019 66085
rect 2961 66076 2973 66079
rect 2924 66048 2973 66076
rect 2924 66036 2930 66048
rect 2961 66045 2973 66048
rect 3007 66076 3019 66079
rect 3602 66076 3608 66088
rect 3007 66048 3608 66076
rect 3007 66045 3019 66048
rect 2961 66039 3019 66045
rect 3602 66036 3608 66048
rect 3660 66036 3666 66088
rect 5074 66076 5080 66088
rect 5035 66048 5080 66076
rect 5074 66036 5080 66048
rect 5132 66036 5138 66088
rect 5537 66079 5595 66085
rect 5537 66045 5549 66079
rect 5583 66076 5595 66079
rect 6472 66076 6500 66107
rect 8128 66088 8156 66116
rect 7282 66076 7288 66088
rect 5583 66048 6500 66076
rect 7243 66048 7288 66076
rect 5583 66045 5595 66048
rect 5537 66039 5595 66045
rect 4801 66011 4859 66017
rect 4801 65977 4813 66011
rect 4847 66008 4859 66011
rect 5552 66008 5580 66039
rect 7282 66036 7288 66048
rect 7340 66036 7346 66088
rect 7561 66079 7619 66085
rect 7561 66045 7573 66079
rect 7607 66045 7619 66079
rect 8110 66076 8116 66088
rect 8071 66048 8116 66076
rect 7561 66039 7619 66045
rect 4847 65980 5580 66008
rect 4847 65977 4859 65980
rect 4801 65971 4859 65977
rect 6822 65968 6828 66020
rect 6880 66008 6886 66020
rect 7576 66008 7604 66039
rect 8110 66036 8116 66048
rect 8168 66036 8174 66088
rect 8570 66076 8576 66088
rect 8483 66048 8576 66076
rect 8570 66036 8576 66048
rect 8628 66076 8634 66088
rect 9582 66076 9588 66088
rect 8628 66048 9588 66076
rect 8628 66036 8634 66048
rect 9582 66036 9588 66048
rect 9640 66036 9646 66088
rect 10060 66076 10088 66184
rect 10134 66172 10140 66184
rect 10192 66172 10198 66224
rect 11054 66172 11060 66224
rect 11112 66212 11118 66224
rect 11517 66215 11575 66221
rect 11517 66212 11529 66215
rect 11112 66184 11529 66212
rect 11112 66172 11118 66184
rect 11517 66181 11529 66184
rect 11563 66212 11575 66215
rect 11606 66212 11612 66224
rect 11563 66184 11612 66212
rect 11563 66181 11575 66184
rect 11517 66175 11575 66181
rect 11606 66172 11612 66184
rect 11664 66172 11670 66224
rect 12434 66172 12440 66224
rect 12492 66212 12498 66224
rect 13633 66215 13691 66221
rect 13633 66212 13645 66215
rect 12492 66184 13645 66212
rect 12492 66172 12498 66184
rect 13633 66181 13645 66184
rect 13679 66181 13691 66215
rect 13633 66175 13691 66181
rect 12989 66147 13047 66153
rect 12989 66113 13001 66147
rect 13035 66144 13047 66147
rect 13354 66144 13360 66156
rect 13035 66116 13360 66144
rect 13035 66113 13047 66116
rect 12989 66107 13047 66113
rect 13354 66104 13360 66116
rect 13412 66104 13418 66156
rect 15105 66147 15163 66153
rect 15105 66113 15117 66147
rect 15151 66144 15163 66147
rect 15470 66144 15476 66156
rect 15151 66116 15476 66144
rect 15151 66113 15163 66116
rect 15105 66107 15163 66113
rect 15470 66104 15476 66116
rect 15528 66144 15534 66156
rect 15565 66147 15623 66153
rect 15565 66144 15577 66147
rect 15528 66116 15577 66144
rect 15528 66104 15534 66116
rect 15565 66113 15577 66116
rect 15611 66113 15623 66147
rect 15565 66107 15623 66113
rect 10129 66079 10187 66085
rect 10129 66076 10141 66079
rect 9692 66048 10141 66076
rect 8202 66008 8208 66020
rect 6880 65980 8208 66008
rect 6880 65968 6886 65980
rect 8202 65968 8208 65980
rect 8260 65968 8266 66020
rect 9692 65952 9720 66048
rect 10129 66045 10141 66048
rect 10175 66076 10187 66079
rect 10597 66079 10655 66085
rect 10597 66076 10609 66079
rect 10175 66048 10609 66076
rect 10175 66045 10187 66048
rect 10129 66039 10187 66045
rect 10597 66045 10609 66048
rect 10643 66045 10655 66079
rect 11333 66079 11391 66085
rect 11333 66076 11345 66079
rect 10597 66039 10655 66045
rect 11256 66048 11345 66076
rect 11256 65952 11284 66048
rect 11333 66045 11345 66048
rect 11379 66076 11391 66079
rect 11974 66076 11980 66088
rect 11379 66048 11980 66076
rect 11379 66045 11391 66048
rect 11333 66039 11391 66045
rect 11974 66036 11980 66048
rect 12032 66076 12038 66088
rect 12069 66079 12127 66085
rect 12069 66076 12081 66079
rect 12032 66048 12081 66076
rect 12032 66036 12038 66048
rect 12069 66045 12081 66048
rect 12115 66045 12127 66079
rect 12069 66039 12127 66045
rect 12526 66036 12532 66088
rect 12584 66076 12590 66088
rect 12621 66079 12679 66085
rect 12621 66076 12633 66079
rect 12584 66048 12633 66076
rect 12584 66036 12590 66048
rect 12621 66045 12633 66048
rect 12667 66045 12679 66079
rect 13262 66076 13268 66088
rect 13223 66048 13268 66076
rect 12621 66039 12679 66045
rect 13262 66036 13268 66048
rect 13320 66036 13326 66088
rect 15289 66079 15347 66085
rect 15289 66045 15301 66079
rect 15335 66076 15347 66079
rect 15378 66076 15384 66088
rect 15335 66048 15384 66076
rect 15335 66045 15347 66048
rect 15289 66039 15347 66045
rect 15378 66036 15384 66048
rect 15436 66036 15442 66088
rect 11790 65968 11796 66020
rect 11848 66008 11854 66020
rect 12802 66008 12808 66020
rect 11848 65980 12808 66008
rect 11848 65968 11854 65980
rect 12802 65968 12808 65980
rect 12860 65968 12866 66020
rect 1854 65900 1860 65952
rect 1912 65940 1918 65952
rect 2041 65943 2099 65949
rect 2041 65940 2053 65943
rect 1912 65912 2053 65940
rect 1912 65900 1918 65912
rect 2041 65909 2053 65912
rect 2087 65909 2099 65943
rect 2041 65903 2099 65909
rect 2774 65900 2780 65952
rect 2832 65940 2838 65952
rect 3145 65943 3203 65949
rect 3145 65940 3157 65943
rect 2832 65912 3157 65940
rect 2832 65900 2838 65912
rect 3145 65909 3157 65912
rect 3191 65909 3203 65943
rect 3145 65903 3203 65909
rect 3326 65900 3332 65952
rect 3384 65940 3390 65952
rect 3605 65943 3663 65949
rect 3605 65940 3617 65943
rect 3384 65912 3617 65940
rect 3384 65900 3390 65912
rect 3605 65909 3617 65912
rect 3651 65909 3663 65943
rect 3605 65903 3663 65909
rect 4614 65900 4620 65952
rect 4672 65940 4678 65952
rect 4890 65940 4896 65952
rect 4672 65912 4896 65940
rect 4672 65900 4678 65912
rect 4890 65900 4896 65912
rect 4948 65900 4954 65952
rect 7466 65900 7472 65952
rect 7524 65940 7530 65952
rect 7837 65943 7895 65949
rect 7837 65940 7849 65943
rect 7524 65912 7849 65940
rect 7524 65900 7530 65912
rect 7837 65909 7849 65912
rect 7883 65909 7895 65943
rect 9122 65940 9128 65952
rect 9083 65912 9128 65940
rect 7837 65903 7895 65909
rect 9122 65900 9128 65912
rect 9180 65900 9186 65952
rect 9214 65900 9220 65952
rect 9272 65940 9278 65952
rect 9401 65943 9459 65949
rect 9401 65940 9413 65943
rect 9272 65912 9413 65940
rect 9272 65900 9278 65912
rect 9401 65909 9413 65912
rect 9447 65909 9459 65943
rect 9401 65903 9459 65909
rect 9674 65900 9680 65952
rect 9732 65900 9738 65952
rect 9766 65900 9772 65952
rect 9824 65940 9830 65952
rect 9953 65943 10011 65949
rect 9953 65940 9965 65943
rect 9824 65912 9965 65940
rect 9824 65900 9830 65912
rect 9953 65909 9965 65912
rect 9999 65940 10011 65943
rect 10042 65940 10048 65952
rect 9999 65912 10048 65940
rect 9999 65909 10011 65912
rect 9953 65903 10011 65909
rect 10042 65900 10048 65912
rect 10100 65900 10106 65952
rect 10318 65940 10324 65952
rect 10279 65912 10324 65940
rect 10318 65900 10324 65912
rect 10376 65900 10382 65952
rect 11238 65940 11244 65952
rect 11199 65912 11244 65940
rect 11238 65900 11244 65912
rect 11296 65900 11302 65952
rect 11330 65900 11336 65952
rect 11388 65940 11394 65952
rect 11606 65940 11612 65952
rect 11388 65912 11612 65940
rect 11388 65900 11394 65912
rect 11606 65900 11612 65912
rect 11664 65900 11670 65952
rect 12529 65943 12587 65949
rect 12529 65909 12541 65943
rect 12575 65940 12587 65943
rect 12894 65940 12900 65952
rect 12575 65912 12900 65940
rect 12575 65909 12587 65912
rect 12529 65903 12587 65909
rect 12894 65900 12900 65912
rect 12952 65900 12958 65952
rect 14734 65940 14740 65952
rect 14695 65912 14740 65940
rect 14734 65900 14740 65912
rect 14792 65940 14798 65952
rect 15102 65940 15108 65952
rect 14792 65912 15108 65940
rect 14792 65900 14798 65912
rect 15102 65900 15108 65912
rect 15160 65900 15166 65952
rect 16574 65900 16580 65952
rect 16632 65940 16638 65952
rect 16669 65943 16727 65949
rect 16669 65940 16681 65943
rect 16632 65912 16681 65940
rect 16632 65900 16638 65912
rect 16669 65909 16681 65912
rect 16715 65909 16727 65943
rect 16669 65903 16727 65909
rect 1104 65850 18860 65872
rect 1104 65798 7648 65850
rect 7700 65798 7712 65850
rect 7764 65798 7776 65850
rect 7828 65798 7840 65850
rect 7892 65798 14315 65850
rect 14367 65798 14379 65850
rect 14431 65798 14443 65850
rect 14495 65798 14507 65850
rect 14559 65798 18860 65850
rect 1104 65776 18860 65798
rect 2130 65696 2136 65748
rect 2188 65736 2194 65748
rect 2314 65736 2320 65748
rect 2188 65708 2320 65736
rect 2188 65696 2194 65708
rect 2314 65696 2320 65708
rect 2372 65736 2378 65748
rect 2593 65739 2651 65745
rect 2593 65736 2605 65739
rect 2372 65708 2605 65736
rect 2372 65696 2378 65708
rect 2593 65705 2605 65708
rect 2639 65705 2651 65739
rect 2593 65699 2651 65705
rect 7101 65739 7159 65745
rect 7101 65705 7113 65739
rect 7147 65736 7159 65739
rect 8570 65736 8576 65748
rect 7147 65708 8576 65736
rect 7147 65705 7159 65708
rect 7101 65699 7159 65705
rect 8570 65696 8576 65708
rect 8628 65696 8634 65748
rect 8754 65696 8760 65748
rect 8812 65736 8818 65748
rect 8812 65708 9168 65736
rect 8812 65696 8818 65708
rect 9140 65680 9168 65708
rect 10134 65696 10140 65748
rect 10192 65736 10198 65748
rect 11057 65739 11115 65745
rect 11057 65736 11069 65739
rect 10192 65708 11069 65736
rect 10192 65696 10198 65708
rect 11057 65705 11069 65708
rect 11103 65705 11115 65739
rect 11057 65699 11115 65705
rect 12526 65696 12532 65748
rect 12584 65736 12590 65748
rect 12989 65739 13047 65745
rect 12989 65736 13001 65739
rect 12584 65708 13001 65736
rect 12584 65696 12590 65708
rect 12989 65705 13001 65708
rect 13035 65705 13047 65739
rect 12989 65699 13047 65705
rect 13906 65696 13912 65748
rect 13964 65736 13970 65748
rect 14737 65739 14795 65745
rect 14737 65736 14749 65739
rect 13964 65708 14749 65736
rect 13964 65696 13970 65708
rect 14737 65705 14749 65708
rect 14783 65705 14795 65739
rect 15378 65736 15384 65748
rect 15339 65708 15384 65736
rect 14737 65699 14795 65705
rect 15378 65696 15384 65708
rect 15436 65696 15442 65748
rect 16114 65736 16120 65748
rect 16075 65708 16120 65736
rect 16114 65696 16120 65708
rect 16172 65696 16178 65748
rect 2498 65628 2504 65680
rect 2556 65668 2562 65680
rect 2866 65668 2872 65680
rect 2556 65640 2872 65668
rect 2556 65628 2562 65640
rect 2866 65628 2872 65640
rect 2924 65668 2930 65680
rect 2961 65671 3019 65677
rect 2961 65668 2973 65671
rect 2924 65640 2973 65668
rect 2924 65628 2930 65640
rect 2961 65637 2973 65640
rect 3007 65668 3019 65671
rect 3007 65640 4200 65668
rect 3007 65637 3019 65640
rect 2961 65631 3019 65637
rect 3145 65603 3203 65609
rect 3145 65569 3157 65603
rect 3191 65600 3203 65603
rect 3326 65600 3332 65612
rect 3191 65572 3332 65600
rect 3191 65569 3203 65572
rect 3145 65563 3203 65569
rect 3326 65560 3332 65572
rect 3384 65560 3390 65612
rect 4172 65609 4200 65640
rect 9122 65628 9128 65680
rect 9180 65628 9186 65680
rect 10965 65671 11023 65677
rect 10965 65668 10977 65671
rect 10888 65640 10977 65668
rect 4157 65603 4215 65609
rect 4157 65569 4169 65603
rect 4203 65569 4215 65603
rect 4798 65600 4804 65612
rect 4157 65563 4215 65569
rect 4356 65572 4804 65600
rect 4356 65532 4384 65572
rect 4798 65560 4804 65572
rect 4856 65560 4862 65612
rect 6641 65603 6699 65609
rect 6641 65569 6653 65603
rect 6687 65600 6699 65603
rect 7466 65600 7472 65612
rect 6687 65572 7472 65600
rect 6687 65569 6699 65572
rect 6641 65563 6699 65569
rect 7466 65560 7472 65572
rect 7524 65560 7530 65612
rect 7926 65600 7932 65612
rect 7887 65572 7932 65600
rect 7926 65560 7932 65572
rect 7984 65560 7990 65612
rect 8205 65603 8263 65609
rect 8205 65569 8217 65603
rect 8251 65569 8263 65603
rect 8205 65563 8263 65569
rect 3988 65504 4384 65532
rect 4433 65535 4491 65541
rect 3988 65476 4016 65504
rect 4433 65501 4445 65535
rect 4479 65532 4491 65535
rect 5442 65532 5448 65544
rect 4479 65504 5448 65532
rect 4479 65501 4491 65504
rect 4433 65495 4491 65501
rect 5442 65492 5448 65504
rect 5500 65492 5506 65544
rect 8021 65535 8079 65541
rect 8021 65501 8033 65535
rect 8067 65532 8079 65535
rect 8110 65532 8116 65544
rect 8067 65504 8116 65532
rect 8067 65501 8079 65504
rect 8021 65495 8079 65501
rect 8110 65492 8116 65504
rect 8168 65492 8174 65544
rect 3329 65467 3387 65473
rect 3329 65433 3341 65467
rect 3375 65464 3387 65467
rect 3970 65464 3976 65476
rect 3375 65436 3976 65464
rect 3375 65433 3387 65436
rect 3329 65427 3387 65433
rect 3970 65424 3976 65436
rect 4028 65424 4034 65476
rect 7466 65424 7472 65476
rect 7524 65464 7530 65476
rect 8220 65464 8248 65563
rect 8386 65560 8392 65612
rect 8444 65600 8450 65612
rect 8665 65603 8723 65609
rect 8665 65600 8677 65603
rect 8444 65572 8677 65600
rect 8444 65560 8450 65572
rect 8665 65569 8677 65572
rect 8711 65569 8723 65603
rect 8665 65563 8723 65569
rect 8754 65560 8760 65612
rect 8812 65600 8818 65612
rect 9033 65603 9091 65609
rect 9033 65600 9045 65603
rect 8812 65572 9045 65600
rect 8812 65560 8818 65572
rect 9033 65569 9045 65572
rect 9079 65569 9091 65603
rect 9033 65563 9091 65569
rect 10686 65560 10692 65612
rect 10744 65600 10750 65612
rect 10888 65600 10916 65640
rect 10965 65637 10977 65640
rect 11011 65637 11023 65671
rect 10965 65631 11023 65637
rect 11149 65671 11207 65677
rect 11149 65637 11161 65671
rect 11195 65668 11207 65671
rect 11330 65668 11336 65680
rect 11195 65640 11336 65668
rect 11195 65637 11207 65640
rect 11149 65631 11207 65637
rect 11330 65628 11336 65640
rect 11388 65628 11394 65680
rect 12713 65671 12771 65677
rect 12713 65637 12725 65671
rect 12759 65668 12771 65671
rect 13262 65668 13268 65680
rect 12759 65640 13268 65668
rect 12759 65637 12771 65640
rect 12713 65631 12771 65637
rect 13262 65628 13268 65640
rect 13320 65628 13326 65680
rect 12250 65600 12256 65612
rect 10744 65572 10916 65600
rect 11348 65572 12256 65600
rect 10744 65560 10750 65572
rect 10594 65492 10600 65544
rect 10652 65532 10658 65544
rect 10781 65535 10839 65541
rect 10781 65532 10793 65535
rect 10652 65504 10793 65532
rect 10652 65492 10658 65504
rect 10781 65501 10793 65504
rect 10827 65532 10839 65535
rect 11348 65532 11376 65572
rect 12250 65560 12256 65572
rect 12308 65560 12314 65612
rect 13170 65560 13176 65612
rect 13228 65600 13234 65612
rect 13357 65603 13415 65609
rect 13357 65600 13369 65603
rect 13228 65572 13369 65600
rect 13228 65560 13234 65572
rect 13357 65569 13369 65572
rect 13403 65600 13415 65603
rect 13998 65600 14004 65612
rect 13403 65572 14004 65600
rect 13403 65569 13415 65572
rect 13357 65563 13415 65569
rect 13998 65560 14004 65572
rect 14056 65560 14062 65612
rect 11514 65532 11520 65544
rect 10827 65504 11376 65532
rect 11427 65504 11520 65532
rect 10827 65501 10839 65504
rect 10781 65495 10839 65501
rect 11514 65492 11520 65504
rect 11572 65532 11578 65544
rect 11974 65532 11980 65544
rect 11572 65504 11980 65532
rect 11572 65492 11578 65504
rect 11974 65492 11980 65504
rect 12032 65492 12038 65544
rect 13630 65532 13636 65544
rect 13591 65504 13636 65532
rect 13630 65492 13636 65504
rect 13688 65492 13694 65544
rect 7524 65436 8248 65464
rect 9677 65467 9735 65473
rect 7524 65424 7530 65436
rect 9677 65433 9689 65467
rect 9723 65464 9735 65467
rect 10410 65464 10416 65476
rect 9723 65436 10416 65464
rect 9723 65433 9735 65436
rect 9677 65427 9735 65433
rect 10410 65424 10416 65436
rect 10468 65424 10474 65476
rect 2222 65396 2228 65408
rect 2183 65368 2228 65396
rect 2222 65356 2228 65368
rect 2280 65356 2286 65408
rect 3694 65396 3700 65408
rect 3655 65368 3700 65396
rect 3694 65356 3700 65368
rect 3752 65356 3758 65408
rect 4065 65399 4123 65405
rect 4065 65365 4077 65399
rect 4111 65396 4123 65399
rect 5074 65396 5080 65408
rect 4111 65368 5080 65396
rect 4111 65365 4123 65368
rect 4065 65359 4123 65365
rect 5074 65356 5080 65368
rect 5132 65356 5138 65408
rect 5534 65396 5540 65408
rect 5495 65368 5540 65396
rect 5534 65356 5540 65368
rect 5592 65356 5598 65408
rect 6086 65396 6092 65408
rect 6047 65368 6092 65396
rect 6086 65356 6092 65368
rect 6144 65356 6150 65408
rect 9950 65356 9956 65408
rect 10008 65396 10014 65408
rect 10137 65399 10195 65405
rect 10137 65396 10149 65399
rect 10008 65368 10149 65396
rect 10008 65356 10014 65368
rect 10137 65365 10149 65368
rect 10183 65365 10195 65399
rect 10137 65359 10195 65365
rect 11885 65399 11943 65405
rect 11885 65365 11897 65399
rect 11931 65396 11943 65399
rect 12250 65396 12256 65408
rect 11931 65368 12256 65396
rect 11931 65365 11943 65368
rect 11885 65359 11943 65365
rect 12250 65356 12256 65368
rect 12308 65356 12314 65408
rect 1104 65306 18860 65328
rect 1104 65254 4315 65306
rect 4367 65254 4379 65306
rect 4431 65254 4443 65306
rect 4495 65254 4507 65306
rect 4559 65254 10982 65306
rect 11034 65254 11046 65306
rect 11098 65254 11110 65306
rect 11162 65254 11174 65306
rect 11226 65254 17648 65306
rect 17700 65254 17712 65306
rect 17764 65254 17776 65306
rect 17828 65254 17840 65306
rect 17892 65254 18860 65306
rect 1104 65232 18860 65254
rect 3237 65195 3295 65201
rect 3237 65161 3249 65195
rect 3283 65192 3295 65195
rect 3326 65192 3332 65204
rect 3283 65164 3332 65192
rect 3283 65161 3295 65164
rect 3237 65155 3295 65161
rect 3326 65152 3332 65164
rect 3384 65152 3390 65204
rect 5258 65192 5264 65204
rect 5219 65164 5264 65192
rect 5258 65152 5264 65164
rect 5316 65152 5322 65204
rect 6086 65192 6092 65204
rect 5644 65164 6092 65192
rect 4062 65084 4068 65136
rect 4120 65124 4126 65136
rect 5644 65124 5672 65164
rect 6086 65152 6092 65164
rect 6144 65152 6150 65204
rect 6914 65152 6920 65204
rect 6972 65192 6978 65204
rect 7009 65195 7067 65201
rect 7009 65192 7021 65195
rect 6972 65164 7021 65192
rect 6972 65152 6978 65164
rect 7009 65161 7021 65164
rect 7055 65161 7067 65195
rect 7926 65192 7932 65204
rect 7887 65164 7932 65192
rect 7009 65155 7067 65161
rect 7926 65152 7932 65164
rect 7984 65152 7990 65204
rect 9493 65195 9551 65201
rect 9493 65161 9505 65195
rect 9539 65192 9551 65195
rect 9582 65192 9588 65204
rect 9539 65164 9588 65192
rect 9539 65161 9551 65164
rect 9493 65155 9551 65161
rect 9582 65152 9588 65164
rect 9640 65152 9646 65204
rect 10594 65152 10600 65204
rect 10652 65192 10658 65204
rect 11333 65195 11391 65201
rect 11333 65192 11345 65195
rect 10652 65164 11345 65192
rect 10652 65152 10658 65164
rect 11333 65161 11345 65164
rect 11379 65161 11391 65195
rect 13170 65192 13176 65204
rect 13131 65164 13176 65192
rect 11333 65155 11391 65161
rect 13170 65152 13176 65164
rect 13228 65152 13234 65204
rect 17494 65192 17500 65204
rect 17455 65164 17500 65192
rect 17494 65152 17500 65164
rect 17552 65152 17558 65204
rect 4120 65096 5672 65124
rect 4120 65084 4126 65096
rect 2590 65016 2596 65068
rect 2648 65056 2654 65068
rect 2685 65059 2743 65065
rect 2685 65056 2697 65059
rect 2648 65028 2697 65056
rect 2648 65016 2654 65028
rect 2685 65025 2697 65028
rect 2731 65025 2743 65059
rect 2685 65019 2743 65025
rect 3694 65016 3700 65068
rect 3752 65056 3758 65068
rect 5534 65056 5540 65068
rect 3752 65028 5540 65056
rect 3752 65016 3758 65028
rect 1762 64948 1768 65000
rect 1820 64988 1826 65000
rect 2222 64988 2228 65000
rect 1820 64960 2228 64988
rect 1820 64948 1826 64960
rect 2222 64948 2228 64960
rect 2280 64948 2286 65000
rect 4356 64997 4384 65028
rect 5534 65016 5540 65028
rect 5592 65016 5598 65068
rect 5644 65065 5672 65096
rect 10152 65096 10824 65124
rect 5629 65059 5687 65065
rect 5629 65025 5641 65059
rect 5675 65025 5687 65059
rect 5629 65019 5687 65025
rect 5810 65016 5816 65068
rect 5868 65056 5874 65068
rect 5905 65059 5963 65065
rect 5905 65056 5917 65059
rect 5868 65028 5917 65056
rect 5868 65016 5874 65028
rect 5905 65025 5917 65028
rect 5951 65025 5963 65059
rect 5905 65019 5963 65025
rect 2409 64991 2467 64997
rect 2409 64957 2421 64991
rect 2455 64957 2467 64991
rect 2409 64951 2467 64957
rect 4341 64991 4399 64997
rect 4341 64957 4353 64991
rect 4387 64957 4399 64991
rect 4341 64951 4399 64957
rect 4617 64991 4675 64997
rect 4617 64957 4629 64991
rect 4663 64957 4675 64991
rect 4617 64951 4675 64957
rect 2133 64923 2191 64929
rect 2133 64889 2145 64923
rect 2179 64920 2191 64923
rect 2424 64920 2452 64951
rect 2498 64920 2504 64932
rect 2179 64892 2504 64920
rect 2179 64889 2191 64892
rect 2133 64883 2191 64889
rect 2498 64880 2504 64892
rect 2556 64880 2562 64932
rect 3881 64923 3939 64929
rect 3881 64889 3893 64923
rect 3927 64920 3939 64923
rect 4632 64920 4660 64951
rect 4706 64948 4712 65000
rect 4764 64988 4770 65000
rect 4801 64991 4859 64997
rect 4801 64988 4813 64991
rect 4764 64960 4813 64988
rect 4764 64948 4770 64960
rect 4801 64957 4813 64960
rect 4847 64957 4859 64991
rect 4801 64951 4859 64957
rect 8294 64948 8300 65000
rect 8352 64988 8358 65000
rect 8573 64991 8631 64997
rect 8573 64988 8585 64991
rect 8352 64960 8585 64988
rect 8352 64948 8358 64960
rect 8573 64957 8585 64960
rect 8619 64957 8631 64991
rect 8573 64951 8631 64957
rect 4890 64920 4896 64932
rect 3927 64892 4896 64920
rect 3927 64889 3939 64892
rect 3881 64883 3939 64889
rect 4890 64880 4896 64892
rect 4948 64880 4954 64932
rect 8588 64920 8616 64951
rect 8938 64948 8944 65000
rect 8996 64988 9002 65000
rect 9950 64988 9956 65000
rect 8996 64960 9956 64988
rect 8996 64948 9002 64960
rect 9950 64948 9956 64960
rect 10008 64988 10014 65000
rect 10152 64997 10180 65096
rect 10594 65056 10600 65068
rect 10555 65028 10600 65056
rect 10594 65016 10600 65028
rect 10652 65016 10658 65068
rect 10137 64991 10195 64997
rect 10137 64988 10149 64991
rect 10008 64960 10149 64988
rect 10008 64948 10014 64960
rect 10137 64957 10149 64960
rect 10183 64957 10195 64991
rect 10686 64988 10692 65000
rect 10647 64960 10692 64988
rect 10137 64951 10195 64957
rect 10686 64948 10692 64960
rect 10744 64948 10750 65000
rect 8846 64920 8852 64932
rect 8588 64892 8852 64920
rect 8846 64880 8852 64892
rect 8904 64920 8910 64932
rect 9033 64923 9091 64929
rect 9033 64920 9045 64923
rect 8904 64892 9045 64920
rect 8904 64880 8910 64892
rect 9033 64889 9045 64892
rect 9079 64889 9091 64923
rect 9033 64883 9091 64889
rect 10045 64923 10103 64929
rect 10045 64889 10057 64923
rect 10091 64920 10103 64923
rect 10704 64920 10732 64948
rect 10091 64892 10732 64920
rect 10796 64920 10824 65096
rect 16025 65059 16083 65065
rect 16025 65025 16037 65059
rect 16071 65056 16083 65059
rect 16071 65028 16436 65056
rect 16071 65025 16083 65028
rect 16025 65019 16083 65025
rect 16408 65000 16436 65028
rect 12342 64988 12348 65000
rect 12303 64960 12348 64988
rect 12342 64948 12348 64960
rect 12400 64948 12406 65000
rect 12437 64991 12495 64997
rect 12437 64957 12449 64991
rect 12483 64988 12495 64991
rect 13265 64991 13323 64997
rect 13265 64988 13277 64991
rect 12483 64960 13277 64988
rect 12483 64957 12495 64960
rect 12437 64951 12495 64957
rect 13265 64957 13277 64960
rect 13311 64988 13323 64991
rect 13998 64988 14004 65000
rect 13311 64960 14004 64988
rect 13311 64957 13323 64960
rect 13265 64951 13323 64957
rect 13998 64948 14004 64960
rect 14056 64988 14062 65000
rect 14093 64991 14151 64997
rect 14093 64988 14105 64991
rect 14056 64960 14105 64988
rect 14056 64948 14062 64960
rect 14093 64957 14105 64960
rect 14139 64957 14151 64991
rect 16114 64988 16120 65000
rect 16075 64960 16120 64988
rect 14093 64951 14151 64957
rect 16114 64948 16120 64960
rect 16172 64948 16178 65000
rect 16390 64988 16396 65000
rect 16351 64960 16396 64988
rect 16390 64948 16396 64960
rect 16448 64948 16454 65000
rect 12710 64920 12716 64932
rect 10796 64892 12716 64920
rect 10091 64889 10103 64892
rect 10045 64883 10103 64889
rect 12710 64880 12716 64892
rect 12768 64920 12774 64932
rect 12894 64920 12900 64932
rect 12768 64892 12900 64920
rect 12768 64880 12774 64892
rect 12894 64880 12900 64892
rect 12952 64880 12958 64932
rect 13630 64880 13636 64932
rect 13688 64920 13694 64932
rect 13817 64923 13875 64929
rect 13817 64920 13829 64923
rect 13688 64892 13829 64920
rect 13688 64880 13694 64892
rect 13817 64889 13829 64892
rect 13863 64920 13875 64923
rect 15102 64920 15108 64932
rect 13863 64892 15108 64920
rect 13863 64889 13875 64892
rect 13817 64883 13875 64889
rect 15102 64880 15108 64892
rect 15160 64880 15166 64932
rect 1765 64855 1823 64861
rect 1765 64821 1777 64855
rect 1811 64852 1823 64855
rect 2866 64852 2872 64864
rect 1811 64824 2872 64852
rect 1811 64821 1823 64824
rect 1765 64815 1823 64821
rect 2866 64812 2872 64824
rect 2924 64812 2930 64864
rect 7466 64812 7472 64864
rect 7524 64852 7530 64864
rect 7561 64855 7619 64861
rect 7561 64852 7573 64855
rect 7524 64824 7573 64852
rect 7524 64812 7530 64824
rect 7561 64821 7573 64824
rect 7607 64821 7619 64855
rect 7561 64815 7619 64821
rect 8389 64855 8447 64861
rect 8389 64821 8401 64855
rect 8435 64852 8447 64855
rect 8478 64852 8484 64864
rect 8435 64824 8484 64852
rect 8435 64821 8447 64824
rect 8389 64815 8447 64821
rect 8478 64812 8484 64824
rect 8536 64852 8542 64864
rect 8754 64852 8760 64864
rect 8536 64824 8760 64852
rect 8536 64812 8542 64824
rect 8754 64812 8760 64824
rect 8812 64812 8818 64864
rect 10134 64812 10140 64864
rect 10192 64852 10198 64864
rect 11149 64855 11207 64861
rect 11149 64852 11161 64855
rect 10192 64824 11161 64852
rect 10192 64812 10198 64824
rect 11149 64821 11161 64824
rect 11195 64821 11207 64855
rect 11149 64815 11207 64821
rect 11333 64855 11391 64861
rect 11333 64821 11345 64855
rect 11379 64852 11391 64855
rect 11609 64855 11667 64861
rect 11609 64852 11621 64855
rect 11379 64824 11621 64852
rect 11379 64821 11391 64824
rect 11333 64815 11391 64821
rect 11609 64821 11621 64824
rect 11655 64852 11667 64855
rect 13449 64855 13507 64861
rect 13449 64852 13461 64855
rect 11655 64824 13461 64852
rect 11655 64821 11667 64824
rect 11609 64815 11667 64821
rect 13449 64821 13461 64824
rect 13495 64821 13507 64855
rect 13449 64815 13507 64821
rect 1104 64762 18860 64784
rect 1104 64710 7648 64762
rect 7700 64710 7712 64762
rect 7764 64710 7776 64762
rect 7828 64710 7840 64762
rect 7892 64710 14315 64762
rect 14367 64710 14379 64762
rect 14431 64710 14443 64762
rect 14495 64710 14507 64762
rect 14559 64710 18860 64762
rect 1104 64688 18860 64710
rect 3418 64608 3424 64660
rect 3476 64648 3482 64660
rect 4062 64648 4068 64660
rect 3476 64620 4068 64648
rect 3476 64608 3482 64620
rect 4062 64608 4068 64620
rect 4120 64608 4126 64660
rect 6638 64648 6644 64660
rect 6551 64620 6644 64648
rect 6638 64608 6644 64620
rect 6696 64648 6702 64660
rect 8386 64648 8392 64660
rect 6696 64620 8392 64648
rect 6696 64608 6702 64620
rect 8386 64608 8392 64620
rect 8444 64608 8450 64660
rect 9858 64608 9864 64660
rect 9916 64648 9922 64660
rect 9953 64651 10011 64657
rect 9953 64648 9965 64651
rect 9916 64620 9965 64648
rect 9916 64608 9922 64620
rect 9953 64617 9965 64620
rect 9999 64617 10011 64651
rect 9953 64611 10011 64617
rect 7101 64583 7159 64589
rect 7101 64549 7113 64583
rect 7147 64580 7159 64583
rect 8478 64580 8484 64592
rect 7147 64552 8484 64580
rect 7147 64549 7159 64552
rect 7101 64543 7159 64549
rect 8478 64540 8484 64552
rect 8536 64540 8542 64592
rect 9600 64552 10732 64580
rect 9600 64524 9628 64552
rect 2777 64515 2835 64521
rect 2777 64481 2789 64515
rect 2823 64512 2835 64515
rect 2866 64512 2872 64524
rect 2823 64484 2872 64512
rect 2823 64481 2835 64484
rect 2777 64475 2835 64481
rect 2866 64472 2872 64484
rect 2924 64512 2930 64524
rect 3878 64512 3884 64524
rect 2924 64484 3884 64512
rect 2924 64472 2930 64484
rect 3878 64472 3884 64484
rect 3936 64472 3942 64524
rect 3970 64472 3976 64524
rect 4028 64512 4034 64524
rect 4614 64512 4620 64524
rect 4028 64484 4620 64512
rect 4028 64472 4034 64484
rect 4614 64472 4620 64484
rect 4672 64512 4678 64524
rect 5261 64515 5319 64521
rect 5261 64512 5273 64515
rect 4672 64484 5273 64512
rect 4672 64472 4678 64484
rect 5261 64481 5273 64484
rect 5307 64481 5319 64515
rect 5261 64475 5319 64481
rect 7282 64472 7288 64524
rect 7340 64512 7346 64524
rect 7561 64515 7619 64521
rect 7561 64512 7573 64515
rect 7340 64484 7573 64512
rect 7340 64472 7346 64484
rect 7561 64481 7573 64484
rect 7607 64481 7619 64515
rect 8294 64512 8300 64524
rect 7561 64475 7619 64481
rect 7668 64484 8300 64512
rect 3050 64444 3056 64456
rect 3011 64416 3056 64444
rect 3050 64404 3056 64416
rect 3108 64404 3114 64456
rect 6362 64404 6368 64456
rect 6420 64444 6426 64456
rect 7668 64444 7696 64484
rect 8294 64472 8300 64484
rect 8352 64512 8358 64524
rect 8389 64515 8447 64521
rect 8389 64512 8401 64515
rect 8352 64484 8401 64512
rect 8352 64472 8358 64484
rect 8389 64481 8401 64484
rect 8435 64481 8447 64515
rect 8389 64475 8447 64481
rect 6420 64416 7696 64444
rect 7837 64447 7895 64453
rect 6420 64404 6426 64416
rect 7837 64413 7849 64447
rect 7883 64444 7895 64447
rect 8202 64444 8208 64456
rect 7883 64416 8208 64444
rect 7883 64413 7895 64416
rect 7837 64407 7895 64413
rect 8202 64404 8208 64416
rect 8260 64404 8266 64456
rect 8404 64444 8432 64475
rect 8570 64472 8576 64524
rect 8628 64512 8634 64524
rect 8849 64515 8907 64521
rect 8849 64512 8861 64515
rect 8628 64484 8861 64512
rect 8628 64472 8634 64484
rect 8849 64481 8861 64484
rect 8895 64512 8907 64515
rect 9582 64512 9588 64524
rect 8895 64484 9588 64512
rect 8895 64481 8907 64484
rect 8849 64475 8907 64481
rect 9582 64472 9588 64484
rect 9640 64472 9646 64524
rect 10134 64512 10140 64524
rect 10095 64484 10140 64512
rect 10134 64472 10140 64484
rect 10192 64472 10198 64524
rect 10318 64512 10324 64524
rect 10279 64484 10324 64512
rect 10318 64472 10324 64484
rect 10376 64472 10382 64524
rect 10704 64521 10732 64552
rect 10689 64515 10747 64521
rect 10689 64481 10701 64515
rect 10735 64481 10747 64515
rect 10689 64475 10747 64481
rect 10778 64472 10784 64524
rect 10836 64512 10842 64524
rect 11241 64515 11299 64521
rect 11241 64512 11253 64515
rect 10836 64484 11253 64512
rect 10836 64472 10842 64484
rect 11241 64481 11253 64484
rect 11287 64481 11299 64515
rect 11241 64475 11299 64481
rect 13078 64472 13084 64524
rect 13136 64512 13142 64524
rect 13265 64515 13323 64521
rect 13265 64512 13277 64515
rect 13136 64484 13277 64512
rect 13136 64472 13142 64484
rect 13265 64481 13277 64484
rect 13311 64481 13323 64515
rect 13265 64475 13323 64481
rect 15102 64472 15108 64524
rect 15160 64512 15166 64524
rect 15473 64515 15531 64521
rect 15473 64512 15485 64515
rect 15160 64484 15485 64512
rect 15160 64472 15166 64484
rect 15473 64481 15485 64484
rect 15519 64512 15531 64515
rect 16114 64512 16120 64524
rect 15519 64484 16120 64512
rect 15519 64481 15531 64484
rect 15473 64475 15531 64481
rect 16114 64472 16120 64484
rect 16172 64472 16178 64524
rect 8662 64444 8668 64456
rect 8404 64416 8668 64444
rect 8662 64404 8668 64416
rect 8720 64404 8726 64456
rect 10336 64444 10364 64472
rect 11330 64444 11336 64456
rect 10336 64416 11336 64444
rect 11330 64404 11336 64416
rect 11388 64444 11394 64456
rect 11609 64447 11667 64453
rect 11609 64444 11621 64447
rect 11388 64416 11621 64444
rect 11388 64404 11394 64416
rect 11609 64413 11621 64416
rect 11655 64413 11667 64447
rect 12986 64444 12992 64456
rect 12947 64416 12992 64444
rect 11609 64407 11667 64413
rect 12986 64404 12992 64416
rect 13044 64404 13050 64456
rect 14366 64444 14372 64456
rect 14327 64416 14372 64444
rect 14366 64404 14372 64416
rect 14424 64404 14430 64456
rect 15654 64404 15660 64456
rect 15712 64444 15718 64456
rect 15749 64447 15807 64453
rect 15749 64444 15761 64447
rect 15712 64416 15761 64444
rect 15712 64404 15718 64416
rect 15749 64413 15761 64416
rect 15795 64413 15807 64447
rect 16850 64444 16856 64456
rect 16811 64416 16856 64444
rect 15749 64407 15807 64413
rect 16850 64404 16856 64416
rect 16908 64404 16914 64456
rect 2225 64379 2283 64385
rect 2225 64345 2237 64379
rect 2271 64376 2283 64379
rect 2682 64376 2688 64388
rect 2271 64348 2688 64376
rect 2271 64345 2283 64348
rect 2225 64339 2283 64345
rect 2682 64336 2688 64348
rect 2740 64336 2746 64388
rect 6273 64379 6331 64385
rect 6273 64345 6285 64379
rect 6319 64376 6331 64379
rect 7098 64376 7104 64388
rect 6319 64348 7104 64376
rect 6319 64345 6331 64348
rect 6273 64339 6331 64345
rect 7098 64336 7104 64348
rect 7156 64376 7162 64388
rect 8113 64379 8171 64385
rect 8113 64376 8125 64379
rect 7156 64348 8125 64376
rect 7156 64336 7162 64348
rect 8113 64345 8125 64348
rect 8159 64345 8171 64379
rect 8113 64339 8171 64345
rect 1673 64311 1731 64317
rect 1673 64277 1685 64311
rect 1719 64308 1731 64311
rect 1762 64308 1768 64320
rect 1719 64280 1768 64308
rect 1719 64277 1731 64280
rect 1673 64271 1731 64277
rect 1762 64268 1768 64280
rect 1820 64268 1826 64320
rect 2406 64268 2412 64320
rect 2464 64308 2470 64320
rect 2593 64311 2651 64317
rect 2593 64308 2605 64311
rect 2464 64280 2605 64308
rect 2464 64268 2470 64280
rect 2593 64277 2605 64280
rect 2639 64308 2651 64311
rect 4157 64311 4215 64317
rect 4157 64308 4169 64311
rect 2639 64280 4169 64308
rect 2639 64277 2651 64280
rect 2593 64271 2651 64277
rect 4157 64277 4169 64280
rect 4203 64277 4215 64311
rect 4157 64271 4215 64277
rect 4890 64268 4896 64320
rect 4948 64308 4954 64320
rect 4985 64311 5043 64317
rect 4985 64308 4997 64311
rect 4948 64280 4997 64308
rect 4948 64268 4954 64280
rect 4985 64277 4997 64280
rect 5031 64308 5043 64311
rect 5445 64311 5503 64317
rect 5445 64308 5457 64311
rect 5031 64280 5457 64308
rect 5031 64277 5043 64280
rect 4985 64271 5043 64277
rect 5445 64277 5457 64280
rect 5491 64277 5503 64311
rect 5810 64308 5816 64320
rect 5771 64280 5816 64308
rect 5445 64271 5503 64277
rect 5810 64268 5816 64280
rect 5868 64268 5874 64320
rect 9306 64308 9312 64320
rect 9267 64280 9312 64308
rect 9306 64268 9312 64280
rect 9364 64268 9370 64320
rect 9766 64308 9772 64320
rect 9727 64280 9772 64308
rect 9766 64268 9772 64280
rect 9824 64268 9830 64320
rect 1104 64218 18860 64240
rect 1104 64166 4315 64218
rect 4367 64166 4379 64218
rect 4431 64166 4443 64218
rect 4495 64166 4507 64218
rect 4559 64166 10982 64218
rect 11034 64166 11046 64218
rect 11098 64166 11110 64218
rect 11162 64166 11174 64218
rect 11226 64166 17648 64218
rect 17700 64166 17712 64218
rect 17764 64166 17776 64218
rect 17828 64166 17840 64218
rect 17892 64166 18860 64218
rect 1104 64144 18860 64166
rect 6362 64104 6368 64116
rect 6323 64076 6368 64104
rect 6362 64064 6368 64076
rect 6420 64064 6426 64116
rect 9493 64107 9551 64113
rect 9493 64073 9505 64107
rect 9539 64104 9551 64107
rect 10318 64104 10324 64116
rect 9539 64076 10324 64104
rect 9539 64073 9551 64076
rect 9493 64067 9551 64073
rect 10318 64064 10324 64076
rect 10376 64064 10382 64116
rect 15102 64104 15108 64116
rect 15063 64076 15108 64104
rect 15102 64064 15108 64076
rect 15160 64064 15166 64116
rect 2041 64039 2099 64045
rect 2041 64005 2053 64039
rect 2087 64036 2099 64039
rect 2774 64036 2780 64048
rect 2087 64008 2780 64036
rect 2087 64005 2099 64008
rect 2041 63999 2099 64005
rect 2774 63996 2780 64008
rect 2832 64036 2838 64048
rect 3881 64039 3939 64045
rect 2832 64008 3188 64036
rect 2832 63996 2838 64008
rect 2682 63900 2688 63912
rect 2643 63872 2688 63900
rect 2682 63860 2688 63872
rect 2740 63860 2746 63912
rect 3160 63909 3188 64008
rect 3881 64005 3893 64039
rect 3927 64036 3939 64039
rect 4062 64036 4068 64048
rect 3927 64008 4068 64036
rect 3927 64005 3939 64008
rect 3881 63999 3939 64005
rect 4062 63996 4068 64008
rect 4120 63996 4126 64048
rect 9306 63996 9312 64048
rect 9364 64036 9370 64048
rect 10502 64036 10508 64048
rect 9364 64008 10508 64036
rect 9364 63996 9370 64008
rect 10502 63996 10508 64008
rect 10560 63996 10566 64048
rect 11330 63996 11336 64048
rect 11388 63996 11394 64048
rect 4154 63928 4160 63980
rect 4212 63968 4218 63980
rect 4706 63968 4712 63980
rect 4212 63940 4712 63968
rect 4212 63928 4218 63940
rect 4706 63928 4712 63940
rect 4764 63928 4770 63980
rect 6086 63928 6092 63980
rect 6144 63968 6150 63980
rect 8386 63968 8392 63980
rect 6144 63940 7328 63968
rect 6144 63928 6150 63940
rect 2961 63903 3019 63909
rect 2961 63869 2973 63903
rect 3007 63869 3019 63903
rect 2961 63863 3019 63869
rect 3145 63903 3203 63909
rect 3145 63869 3157 63903
rect 3191 63900 3203 63903
rect 3602 63900 3608 63912
rect 3191 63872 3608 63900
rect 3191 63869 3203 63872
rect 3145 63863 3203 63869
rect 2130 63832 2136 63844
rect 2091 63804 2136 63832
rect 2130 63792 2136 63804
rect 2188 63792 2194 63844
rect 2406 63792 2412 63844
rect 2464 63832 2470 63844
rect 2976 63832 3004 63863
rect 3602 63860 3608 63872
rect 3660 63860 3666 63912
rect 4525 63903 4583 63909
rect 4525 63869 4537 63903
rect 4571 63900 4583 63903
rect 5258 63900 5264 63912
rect 4571 63872 5264 63900
rect 4571 63869 4583 63872
rect 4525 63863 4583 63869
rect 5258 63860 5264 63872
rect 5316 63860 5322 63912
rect 5445 63903 5503 63909
rect 5445 63869 5457 63903
rect 5491 63869 5503 63903
rect 7098 63900 7104 63912
rect 7059 63872 7104 63900
rect 5445 63863 5503 63869
rect 2464 63804 3004 63832
rect 2464 63792 2470 63804
rect 3050 63792 3056 63844
rect 3108 63832 3114 63844
rect 3513 63835 3571 63841
rect 3513 63832 3525 63835
rect 3108 63804 3525 63832
rect 3108 63792 3114 63804
rect 3513 63801 3525 63804
rect 3559 63832 3571 63835
rect 4062 63832 4068 63844
rect 3559 63804 4068 63832
rect 3559 63801 3571 63804
rect 3513 63795 3571 63801
rect 4062 63792 4068 63804
rect 4120 63792 4126 63844
rect 4890 63792 4896 63844
rect 4948 63832 4954 63844
rect 5460 63832 5488 63863
rect 7098 63860 7104 63872
rect 7156 63860 7162 63912
rect 7300 63909 7328 63940
rect 8128 63940 8392 63968
rect 7285 63903 7343 63909
rect 7285 63869 7297 63903
rect 7331 63869 7343 63903
rect 7926 63900 7932 63912
rect 7887 63872 7932 63900
rect 7285 63863 7343 63869
rect 7926 63860 7932 63872
rect 7984 63860 7990 63912
rect 8128 63909 8156 63940
rect 8386 63928 8392 63940
rect 8444 63928 8450 63980
rect 11057 63971 11115 63977
rect 11057 63968 11069 63971
rect 9784 63940 11069 63968
rect 9784 63912 9812 63940
rect 11057 63937 11069 63940
rect 11103 63968 11115 63971
rect 11348 63968 11376 63996
rect 11103 63940 12480 63968
rect 11103 63937 11115 63940
rect 11057 63931 11115 63937
rect 8113 63903 8171 63909
rect 8113 63869 8125 63903
rect 8159 63869 8171 63903
rect 8113 63863 8171 63869
rect 8202 63860 8208 63912
rect 8260 63900 8266 63912
rect 8478 63900 8484 63912
rect 8260 63872 8484 63900
rect 8260 63860 8266 63872
rect 8478 63860 8484 63872
rect 8536 63860 8542 63912
rect 9766 63900 9772 63912
rect 9727 63872 9772 63900
rect 9766 63860 9772 63872
rect 9824 63860 9830 63912
rect 10321 63903 10379 63909
rect 10321 63869 10333 63903
rect 10367 63869 10379 63903
rect 10502 63900 10508 63912
rect 10463 63872 10508 63900
rect 10321 63863 10379 63869
rect 7190 63832 7196 63844
rect 4948 63804 5488 63832
rect 7151 63804 7196 63832
rect 4948 63792 4954 63804
rect 7190 63792 7196 63804
rect 7248 63792 7254 63844
rect 1670 63764 1676 63776
rect 1631 63736 1676 63764
rect 1670 63724 1676 63736
rect 1728 63724 1734 63776
rect 4614 63724 4620 63776
rect 4672 63764 4678 63776
rect 4801 63767 4859 63773
rect 4801 63764 4813 63767
rect 4672 63736 4813 63764
rect 4672 63724 4678 63736
rect 4801 63733 4813 63736
rect 4847 63733 4859 63767
rect 5074 63764 5080 63776
rect 5035 63736 5080 63764
rect 4801 63727 4859 63733
rect 5074 63724 5080 63736
rect 5132 63724 5138 63776
rect 6733 63767 6791 63773
rect 6733 63733 6745 63767
rect 6779 63764 6791 63767
rect 7466 63764 7472 63776
rect 6779 63736 7472 63764
rect 6779 63733 6791 63736
rect 6733 63727 6791 63733
rect 7466 63724 7472 63736
rect 7524 63764 7530 63776
rect 7944 63764 7972 63860
rect 9125 63835 9183 63841
rect 9125 63801 9137 63835
rect 9171 63832 9183 63835
rect 9950 63832 9956 63844
rect 9171 63804 9956 63832
rect 9171 63801 9183 63804
rect 9125 63795 9183 63801
rect 9950 63792 9956 63804
rect 10008 63832 10014 63844
rect 10336 63832 10364 63863
rect 10502 63860 10508 63872
rect 10560 63860 10566 63912
rect 11333 63903 11391 63909
rect 11333 63869 11345 63903
rect 11379 63900 11391 63903
rect 11609 63903 11667 63909
rect 11609 63900 11621 63903
rect 11379 63872 11621 63900
rect 11379 63869 11391 63872
rect 11333 63863 11391 63869
rect 11609 63869 11621 63872
rect 11655 63869 11667 63903
rect 12066 63900 12072 63912
rect 12027 63872 12072 63900
rect 11609 63863 11667 63869
rect 12066 63860 12072 63872
rect 12124 63860 12130 63912
rect 12452 63909 12480 63940
rect 15378 63928 15384 63980
rect 15436 63928 15442 63980
rect 16025 63971 16083 63977
rect 16025 63937 16037 63971
rect 16071 63968 16083 63971
rect 16071 63940 16436 63968
rect 16071 63937 16083 63940
rect 16025 63931 16083 63937
rect 12437 63903 12495 63909
rect 12437 63869 12449 63903
rect 12483 63869 12495 63903
rect 13078 63900 13084 63912
rect 13039 63872 13084 63900
rect 12437 63863 12495 63869
rect 13078 63860 13084 63872
rect 13136 63860 13142 63912
rect 13541 63903 13599 63909
rect 13541 63869 13553 63903
rect 13587 63869 13599 63903
rect 13998 63900 14004 63912
rect 13959 63872 14004 63900
rect 13541 63863 13599 63869
rect 10008 63804 10364 63832
rect 10008 63792 10014 63804
rect 11054 63792 11060 63844
rect 11112 63832 11118 63844
rect 11112 63804 11744 63832
rect 11112 63792 11118 63804
rect 7524 63736 7972 63764
rect 7524 63724 7530 63736
rect 8478 63724 8484 63776
rect 8536 63764 8542 63776
rect 9398 63764 9404 63776
rect 8536 63736 9404 63764
rect 8536 63724 8542 63736
rect 9398 63724 9404 63736
rect 9456 63724 9462 63776
rect 9674 63724 9680 63776
rect 9732 63764 9738 63776
rect 9769 63767 9827 63773
rect 9769 63764 9781 63767
rect 9732 63736 9781 63764
rect 9732 63724 9738 63736
rect 9769 63733 9781 63736
rect 9815 63733 9827 63767
rect 9769 63727 9827 63733
rect 11146 63724 11152 63776
rect 11204 63764 11210 63776
rect 11716 63773 11744 63804
rect 12526 63792 12532 63844
rect 12584 63832 12590 63844
rect 13357 63835 13415 63841
rect 13357 63832 13369 63835
rect 12584 63804 13369 63832
rect 12584 63792 12590 63804
rect 13357 63801 13369 63804
rect 13403 63832 13415 63835
rect 13556 63832 13584 63863
rect 13998 63860 14004 63872
rect 14056 63900 14062 63912
rect 14553 63903 14611 63909
rect 14553 63900 14565 63903
rect 14056 63872 14565 63900
rect 14056 63860 14062 63872
rect 14553 63869 14565 63872
rect 14599 63869 14611 63903
rect 15396 63900 15424 63928
rect 15562 63900 15568 63912
rect 15396 63872 15568 63900
rect 14553 63863 14611 63869
rect 15562 63860 15568 63872
rect 15620 63900 15626 63912
rect 16408 63909 16436 63940
rect 16117 63903 16175 63909
rect 16117 63900 16129 63903
rect 15620 63872 16129 63900
rect 15620 63860 15626 63872
rect 16117 63869 16129 63872
rect 16163 63869 16175 63903
rect 16117 63863 16175 63869
rect 16393 63903 16451 63909
rect 16393 63869 16405 63903
rect 16439 63900 16451 63903
rect 16482 63900 16488 63912
rect 16439 63872 16488 63900
rect 16439 63869 16451 63872
rect 16393 63863 16451 63869
rect 16482 63860 16488 63872
rect 16540 63860 16546 63912
rect 13403 63804 13584 63832
rect 13403 63801 13415 63804
rect 13357 63795 13415 63801
rect 11333 63767 11391 63773
rect 11333 63764 11345 63767
rect 11204 63736 11345 63764
rect 11204 63724 11210 63736
rect 11333 63733 11345 63736
rect 11379 63764 11391 63767
rect 11425 63767 11483 63773
rect 11425 63764 11437 63767
rect 11379 63736 11437 63764
rect 11379 63733 11391 63736
rect 11333 63727 11391 63733
rect 11425 63733 11437 63736
rect 11471 63733 11483 63767
rect 11425 63727 11483 63733
rect 11701 63767 11759 63773
rect 11701 63733 11713 63767
rect 11747 63733 11759 63767
rect 11701 63727 11759 63733
rect 13262 63724 13268 63776
rect 13320 63764 13326 63776
rect 13633 63767 13691 63773
rect 13633 63764 13645 63767
rect 13320 63736 13645 63764
rect 13320 63724 13326 63736
rect 13633 63733 13645 63736
rect 13679 63733 13691 63767
rect 13633 63727 13691 63733
rect 15565 63767 15623 63773
rect 15565 63733 15577 63767
rect 15611 63764 15623 63767
rect 15654 63764 15660 63776
rect 15611 63736 15660 63764
rect 15611 63733 15623 63736
rect 15565 63727 15623 63733
rect 15654 63724 15660 63736
rect 15712 63724 15718 63776
rect 17494 63764 17500 63776
rect 17455 63736 17500 63764
rect 17494 63724 17500 63736
rect 17552 63724 17558 63776
rect 1104 63674 18860 63696
rect 1104 63622 7648 63674
rect 7700 63622 7712 63674
rect 7764 63622 7776 63674
rect 7828 63622 7840 63674
rect 7892 63622 14315 63674
rect 14367 63622 14379 63674
rect 14431 63622 14443 63674
rect 14495 63622 14507 63674
rect 14559 63622 18860 63674
rect 1104 63600 18860 63622
rect 5258 63520 5264 63572
rect 5316 63560 5322 63572
rect 5629 63563 5687 63569
rect 5629 63560 5641 63563
rect 5316 63532 5641 63560
rect 5316 63520 5322 63532
rect 5629 63529 5641 63532
rect 5675 63529 5687 63563
rect 5629 63523 5687 63529
rect 6086 63520 6092 63572
rect 6144 63560 6150 63572
rect 6181 63563 6239 63569
rect 6181 63560 6193 63563
rect 6144 63532 6193 63560
rect 6144 63520 6150 63532
rect 6181 63529 6193 63532
rect 6227 63560 6239 63563
rect 6362 63560 6368 63572
rect 6227 63532 6368 63560
rect 6227 63529 6239 63532
rect 6181 63523 6239 63529
rect 6362 63520 6368 63532
rect 6420 63520 6426 63572
rect 6638 63560 6644 63572
rect 6599 63532 6644 63560
rect 6638 63520 6644 63532
rect 6696 63520 6702 63572
rect 8570 63560 8576 63572
rect 8312 63532 8576 63560
rect 7929 63495 7987 63501
rect 7929 63461 7941 63495
rect 7975 63492 7987 63495
rect 8312 63492 8340 63532
rect 8570 63520 8576 63532
rect 8628 63520 8634 63572
rect 10134 63520 10140 63572
rect 10192 63560 10198 63572
rect 10502 63560 10508 63572
rect 10192 63532 10508 63560
rect 10192 63520 10198 63532
rect 10502 63520 10508 63532
rect 10560 63560 10566 63572
rect 10560 63532 11008 63560
rect 10560 63520 10566 63532
rect 9858 63492 9864 63504
rect 7975 63464 8340 63492
rect 9232 63464 9864 63492
rect 7975 63461 7987 63464
rect 7929 63455 7987 63461
rect 1489 63427 1547 63433
rect 1489 63393 1501 63427
rect 1535 63424 1547 63427
rect 1535 63396 2728 63424
rect 1535 63393 1547 63396
rect 1489 63387 1547 63393
rect 1762 63356 1768 63368
rect 1675 63328 1768 63356
rect 1762 63316 1768 63328
rect 1820 63356 1826 63368
rect 2130 63356 2136 63368
rect 1820 63328 2136 63356
rect 1820 63316 1826 63328
rect 2130 63316 2136 63328
rect 2188 63316 2194 63368
rect 2700 63300 2728 63396
rect 3878 63384 3884 63436
rect 3936 63424 3942 63436
rect 4249 63427 4307 63433
rect 4249 63424 4261 63427
rect 3936 63396 4261 63424
rect 3936 63384 3942 63396
rect 4249 63393 4261 63396
rect 4295 63393 4307 63427
rect 4249 63387 4307 63393
rect 7469 63427 7527 63433
rect 7469 63393 7481 63427
rect 7515 63393 7527 63427
rect 7469 63387 7527 63393
rect 7561 63427 7619 63433
rect 7561 63393 7573 63427
rect 7607 63424 7619 63427
rect 8018 63424 8024 63436
rect 7607 63396 8024 63424
rect 7607 63393 7619 63396
rect 7561 63387 7619 63393
rect 3970 63316 3976 63368
rect 4028 63356 4034 63368
rect 4522 63356 4528 63368
rect 4028 63328 4528 63356
rect 4028 63316 4034 63328
rect 4522 63316 4528 63328
rect 4580 63316 4586 63368
rect 7484 63356 7512 63387
rect 8018 63384 8024 63396
rect 8076 63384 8082 63436
rect 9232 63433 9260 63464
rect 9858 63452 9864 63464
rect 9916 63452 9922 63504
rect 10980 63492 11008 63532
rect 11606 63520 11612 63572
rect 11664 63560 11670 63572
rect 11701 63563 11759 63569
rect 11701 63560 11713 63563
rect 11664 63532 11713 63560
rect 11664 63520 11670 63532
rect 11701 63529 11713 63532
rect 11747 63560 11759 63563
rect 12066 63560 12072 63572
rect 11747 63532 12072 63560
rect 11747 63529 11759 63532
rect 11701 63523 11759 63529
rect 12066 63520 12072 63532
rect 12124 63520 12130 63572
rect 15562 63560 15568 63572
rect 15523 63532 15568 63560
rect 15562 63520 15568 63532
rect 15620 63560 15626 63572
rect 15746 63560 15752 63572
rect 15620 63532 15752 63560
rect 15620 63520 15626 63532
rect 15746 63520 15752 63532
rect 15804 63560 15810 63572
rect 16485 63563 16543 63569
rect 16485 63560 16497 63563
rect 15804 63532 16497 63560
rect 15804 63520 15810 63532
rect 16485 63529 16497 63532
rect 16531 63529 16543 63563
rect 16485 63523 16543 63529
rect 11149 63495 11207 63501
rect 11149 63492 11161 63495
rect 10980 63464 11161 63492
rect 11149 63461 11161 63464
rect 11195 63461 11207 63495
rect 11149 63455 11207 63461
rect 9217 63427 9275 63433
rect 9217 63393 9229 63427
rect 9263 63393 9275 63427
rect 9398 63424 9404 63436
rect 9359 63396 9404 63424
rect 9217 63387 9275 63393
rect 9398 63384 9404 63396
rect 9456 63424 9462 63436
rect 9582 63424 9588 63436
rect 9456 63396 9588 63424
rect 9456 63384 9462 63396
rect 9582 63384 9588 63396
rect 9640 63384 9646 63436
rect 9766 63424 9772 63436
rect 9727 63396 9772 63424
rect 9766 63384 9772 63396
rect 9824 63384 9830 63436
rect 10137 63427 10195 63433
rect 10137 63393 10149 63427
rect 10183 63393 10195 63427
rect 10686 63424 10692 63436
rect 10647 63396 10692 63424
rect 10137 63387 10195 63393
rect 7742 63356 7748 63368
rect 7484 63328 7748 63356
rect 7742 63316 7748 63328
rect 7800 63316 7806 63368
rect 9030 63316 9036 63368
rect 9088 63356 9094 63368
rect 10152 63356 10180 63387
rect 10686 63384 10692 63396
rect 10744 63384 10750 63436
rect 12437 63427 12495 63433
rect 12437 63393 12449 63427
rect 12483 63424 12495 63427
rect 12526 63424 12532 63436
rect 12483 63396 12532 63424
rect 12483 63393 12495 63396
rect 12437 63387 12495 63393
rect 12526 63384 12532 63396
rect 12584 63384 12590 63436
rect 13541 63427 13599 63433
rect 13541 63393 13553 63427
rect 13587 63424 13599 63427
rect 14734 63424 14740 63436
rect 13587 63396 14740 63424
rect 13587 63393 13599 63396
rect 13541 63387 13599 63393
rect 14734 63384 14740 63396
rect 14792 63424 14798 63436
rect 15102 63424 15108 63436
rect 14792 63396 15108 63424
rect 14792 63384 14798 63396
rect 15102 63384 15108 63396
rect 15160 63384 15166 63436
rect 15562 63384 15568 63436
rect 15620 63424 15626 63436
rect 16025 63427 16083 63433
rect 16025 63424 16037 63427
rect 15620 63396 16037 63424
rect 15620 63384 15626 63396
rect 16025 63393 16037 63396
rect 16071 63393 16083 63427
rect 16025 63387 16083 63393
rect 10962 63356 10968 63368
rect 9088 63328 10968 63356
rect 9088 63316 9094 63328
rect 10962 63316 10968 63328
rect 11020 63316 11026 63368
rect 11422 63316 11428 63368
rect 11480 63356 11486 63368
rect 11480 63328 13492 63356
rect 11480 63316 11486 63328
rect 2682 63248 2688 63300
rect 2740 63288 2746 63300
rect 3418 63288 3424 63300
rect 2740 63260 3424 63288
rect 2740 63248 2746 63260
rect 3418 63248 3424 63260
rect 3476 63248 3482 63300
rect 9214 63288 9220 63300
rect 9175 63260 9220 63288
rect 9214 63248 9220 63260
rect 9272 63248 9278 63300
rect 9674 63248 9680 63300
rect 9732 63288 9738 63300
rect 10226 63288 10232 63300
rect 9732 63260 10232 63288
rect 9732 63248 9738 63260
rect 10226 63248 10232 63260
rect 10284 63248 10290 63300
rect 1670 63180 1676 63232
rect 1728 63220 1734 63232
rect 2222 63220 2228 63232
rect 1728 63192 2228 63220
rect 1728 63180 1734 63192
rect 2222 63180 2228 63192
rect 2280 63220 2286 63232
rect 2869 63223 2927 63229
rect 2869 63220 2881 63223
rect 2280 63192 2881 63220
rect 2280 63180 2286 63192
rect 2869 63189 2881 63192
rect 2915 63189 2927 63223
rect 4062 63220 4068 63232
rect 4023 63192 4068 63220
rect 2869 63183 2927 63189
rect 4062 63180 4068 63192
rect 4120 63180 4126 63232
rect 8294 63220 8300 63232
rect 8207 63192 8300 63220
rect 8294 63180 8300 63192
rect 8352 63220 8358 63232
rect 9582 63220 9588 63232
rect 8352 63192 9588 63220
rect 8352 63180 8358 63192
rect 9582 63180 9588 63192
rect 9640 63180 9646 63232
rect 10042 63180 10048 63232
rect 10100 63220 10106 63232
rect 12621 63223 12679 63229
rect 12621 63220 12633 63223
rect 10100 63192 12633 63220
rect 10100 63180 10106 63192
rect 12621 63189 12633 63192
rect 12667 63189 12679 63223
rect 12986 63220 12992 63232
rect 12899 63192 12992 63220
rect 12621 63183 12679 63189
rect 12986 63180 12992 63192
rect 13044 63220 13050 63232
rect 13354 63220 13360 63232
rect 13044 63192 13360 63220
rect 13044 63180 13050 63192
rect 13354 63180 13360 63192
rect 13412 63180 13418 63232
rect 13464 63220 13492 63328
rect 13722 63316 13728 63368
rect 13780 63356 13786 63368
rect 13817 63359 13875 63365
rect 13817 63356 13829 63359
rect 13780 63328 13829 63356
rect 13780 63316 13786 63328
rect 13817 63325 13829 63328
rect 13863 63325 13875 63359
rect 13817 63319 13875 63325
rect 14826 63220 14832 63232
rect 13464 63192 14832 63220
rect 14826 63180 14832 63192
rect 14884 63220 14890 63232
rect 14921 63223 14979 63229
rect 14921 63220 14933 63223
rect 14884 63192 14933 63220
rect 14884 63180 14890 63192
rect 14921 63189 14933 63192
rect 14967 63189 14979 63223
rect 16206 63220 16212 63232
rect 16167 63192 16212 63220
rect 14921 63183 14979 63189
rect 16206 63180 16212 63192
rect 16264 63180 16270 63232
rect 1104 63130 18860 63152
rect 1104 63078 4315 63130
rect 4367 63078 4379 63130
rect 4431 63078 4443 63130
rect 4495 63078 4507 63130
rect 4559 63078 10982 63130
rect 11034 63078 11046 63130
rect 11098 63078 11110 63130
rect 11162 63078 11174 63130
rect 11226 63078 17648 63130
rect 17700 63078 17712 63130
rect 17764 63078 17776 63130
rect 17828 63078 17840 63130
rect 17892 63078 18860 63130
rect 1104 63056 18860 63078
rect 2590 62976 2596 63028
rect 2648 63016 2654 63028
rect 3145 63019 3203 63025
rect 3145 63016 3157 63019
rect 2648 62988 3157 63016
rect 2648 62976 2654 62988
rect 3145 62985 3157 62988
rect 3191 62985 3203 63019
rect 3145 62979 3203 62985
rect 3881 63019 3939 63025
rect 3881 62985 3893 63019
rect 3927 63016 3939 63019
rect 3970 63016 3976 63028
rect 3927 62988 3976 63016
rect 3927 62985 3939 62988
rect 3881 62979 3939 62985
rect 3970 62976 3976 62988
rect 4028 62976 4034 63028
rect 4154 62976 4160 63028
rect 4212 63016 4218 63028
rect 4341 63019 4399 63025
rect 4341 63016 4353 63019
rect 4212 62988 4353 63016
rect 4212 62976 4218 62988
rect 4341 62985 4353 62988
rect 4387 62985 4399 63019
rect 4341 62979 4399 62985
rect 4985 63019 5043 63025
rect 4985 62985 4997 63019
rect 5031 63016 5043 63019
rect 5442 63016 5448 63028
rect 5031 62988 5448 63016
rect 5031 62985 5043 62988
rect 4985 62979 5043 62985
rect 2041 62883 2099 62889
rect 2041 62849 2053 62883
rect 2087 62880 2099 62883
rect 2608 62880 2636 62976
rect 5000 62880 5028 62979
rect 5442 62976 5448 62988
rect 5500 62976 5506 63028
rect 8113 63019 8171 63025
rect 8113 62985 8125 63019
rect 8159 63016 8171 63019
rect 9398 63016 9404 63028
rect 8159 62988 9404 63016
rect 8159 62985 8171 62988
rect 8113 62979 8171 62985
rect 9398 62976 9404 62988
rect 9456 62976 9462 63028
rect 9950 63016 9956 63028
rect 9911 62988 9956 63016
rect 9950 62976 9956 62988
rect 10008 62976 10014 63028
rect 11425 63019 11483 63025
rect 11425 62985 11437 63019
rect 11471 63016 11483 63019
rect 12618 63016 12624 63028
rect 11471 62988 12624 63016
rect 11471 62985 11483 62988
rect 11425 62979 11483 62985
rect 8481 62951 8539 62957
rect 8481 62917 8493 62951
rect 8527 62948 8539 62951
rect 9030 62948 9036 62960
rect 8527 62920 9036 62948
rect 8527 62917 8539 62920
rect 8481 62911 8539 62917
rect 9030 62908 9036 62920
rect 9088 62908 9094 62960
rect 10686 62948 10692 62960
rect 9876 62920 10692 62948
rect 2087 62852 2636 62880
rect 4264 62852 5028 62880
rect 9125 62883 9183 62889
rect 2087 62849 2099 62852
rect 2041 62843 2099 62849
rect 2222 62772 2228 62824
rect 2280 62812 2286 62824
rect 2317 62815 2375 62821
rect 2317 62812 2329 62815
rect 2280 62784 2329 62812
rect 2280 62772 2286 62784
rect 2317 62781 2329 62784
rect 2363 62781 2375 62815
rect 2498 62812 2504 62824
rect 2459 62784 2504 62812
rect 2317 62775 2375 62781
rect 2498 62772 2504 62784
rect 2556 62812 2562 62824
rect 4264 62821 4292 62852
rect 9125 62849 9137 62883
rect 9171 62880 9183 62883
rect 9398 62880 9404 62892
rect 9171 62852 9404 62880
rect 9171 62849 9183 62852
rect 9125 62843 9183 62849
rect 2777 62815 2835 62821
rect 2777 62812 2789 62815
rect 2556 62784 2789 62812
rect 2556 62772 2562 62784
rect 2777 62781 2789 62784
rect 2823 62781 2835 62815
rect 2777 62775 2835 62781
rect 4249 62815 4307 62821
rect 4249 62781 4261 62815
rect 4295 62781 4307 62815
rect 4249 62775 4307 62781
rect 4798 62772 4804 62824
rect 4856 62812 4862 62824
rect 5626 62812 5632 62824
rect 4856 62784 5632 62812
rect 4856 62772 4862 62784
rect 5626 62772 5632 62784
rect 5684 62772 5690 62824
rect 5810 62772 5816 62824
rect 5868 62812 5874 62824
rect 6181 62815 6239 62821
rect 6181 62812 6193 62815
rect 5868 62784 6193 62812
rect 5868 62772 5874 62784
rect 6181 62781 6193 62784
rect 6227 62812 6239 62815
rect 6638 62812 6644 62824
rect 6227 62784 6644 62812
rect 6227 62781 6239 62784
rect 6181 62775 6239 62781
rect 6638 62772 6644 62784
rect 6696 62772 6702 62824
rect 6822 62772 6828 62824
rect 6880 62812 6886 62824
rect 7466 62812 7472 62824
rect 6880 62784 7472 62812
rect 6880 62772 6886 62784
rect 7466 62772 7472 62784
rect 7524 62772 7530 62824
rect 8573 62815 8631 62821
rect 8573 62781 8585 62815
rect 8619 62812 8631 62815
rect 9140 62812 9168 62843
rect 9398 62840 9404 62852
rect 9456 62840 9462 62892
rect 8619 62784 9168 62812
rect 8619 62781 8631 62784
rect 8573 62775 8631 62781
rect 1486 62744 1492 62756
rect 1447 62716 1492 62744
rect 1486 62704 1492 62716
rect 1544 62704 1550 62756
rect 4062 62744 4068 62756
rect 3975 62716 4068 62744
rect 4062 62704 4068 62716
rect 4120 62744 4126 62756
rect 4982 62744 4988 62756
rect 4120 62716 4988 62744
rect 4120 62704 4126 62716
rect 4982 62704 4988 62716
rect 5040 62704 5046 62756
rect 7742 62744 7748 62756
rect 7703 62716 7748 62744
rect 7742 62704 7748 62716
rect 7800 62704 7806 62756
rect 8386 62704 8392 62756
rect 8444 62744 8450 62756
rect 9401 62747 9459 62753
rect 9401 62744 9413 62747
rect 8444 62716 9413 62744
rect 8444 62704 8450 62716
rect 9401 62713 9413 62716
rect 9447 62744 9459 62747
rect 9876 62744 9904 62920
rect 10686 62908 10692 62920
rect 10744 62908 10750 62960
rect 11440 62880 11468 62979
rect 12618 62976 12624 62988
rect 12676 62976 12682 63028
rect 14734 63016 14740 63028
rect 14695 62988 14740 63016
rect 14734 62976 14740 62988
rect 14792 62976 14798 63028
rect 15010 63016 15016 63028
rect 14971 62988 15016 63016
rect 15010 62976 15016 62988
rect 15068 62976 15074 63028
rect 16942 63016 16948 63028
rect 16903 62988 16948 63016
rect 16942 62976 16948 62988
rect 17000 62976 17006 63028
rect 10060 62852 11468 62880
rect 12621 62883 12679 62889
rect 10060 62824 10088 62852
rect 12621 62849 12633 62883
rect 12667 62880 12679 62883
rect 15028 62880 15056 62976
rect 15657 62883 15715 62889
rect 15657 62880 15669 62883
rect 12667 62852 13032 62880
rect 15028 62852 15669 62880
rect 12667 62849 12679 62852
rect 12621 62843 12679 62849
rect 10042 62812 10048 62824
rect 9955 62784 10048 62812
rect 10042 62772 10048 62784
rect 10100 62772 10106 62824
rect 10226 62812 10232 62824
rect 10187 62784 10232 62812
rect 10226 62772 10232 62784
rect 10284 62772 10290 62824
rect 10686 62812 10692 62824
rect 10647 62784 10692 62812
rect 10686 62772 10692 62784
rect 10744 62812 10750 62824
rect 10962 62812 10968 62824
rect 10744 62784 10968 62812
rect 10744 62772 10750 62784
rect 10962 62772 10968 62784
rect 11020 62772 11026 62824
rect 13004 62821 13032 62852
rect 15657 62849 15669 62852
rect 15703 62849 15715 62883
rect 15657 62843 15715 62849
rect 12713 62815 12771 62821
rect 12713 62781 12725 62815
rect 12759 62781 12771 62815
rect 12713 62775 12771 62781
rect 12989 62815 13047 62821
rect 12989 62781 13001 62815
rect 13035 62812 13047 62815
rect 13078 62812 13084 62824
rect 13035 62784 13084 62812
rect 13035 62781 13047 62784
rect 12989 62775 13047 62781
rect 9447 62716 9904 62744
rect 9447 62713 9459 62716
rect 9401 62707 9459 62713
rect 4154 62636 4160 62688
rect 4212 62676 4218 62688
rect 4706 62676 4712 62688
rect 4212 62648 4712 62676
rect 4212 62636 4218 62648
rect 4706 62636 4712 62648
rect 4764 62636 4770 62688
rect 4798 62636 4804 62688
rect 4856 62676 4862 62688
rect 5261 62679 5319 62685
rect 5261 62676 5273 62679
rect 4856 62648 5273 62676
rect 4856 62636 4862 62648
rect 5261 62645 5273 62648
rect 5307 62645 5319 62679
rect 6546 62676 6552 62688
rect 6507 62648 6552 62676
rect 5261 62639 5319 62645
rect 6546 62636 6552 62648
rect 6604 62636 6610 62688
rect 7282 62676 7288 62688
rect 7243 62648 7288 62676
rect 7282 62636 7288 62648
rect 7340 62636 7346 62688
rect 8754 62676 8760 62688
rect 8715 62648 8760 62676
rect 8754 62636 8760 62648
rect 8812 62636 8818 62688
rect 12158 62636 12164 62688
rect 12216 62676 12222 62688
rect 12253 62679 12311 62685
rect 12253 62676 12265 62679
rect 12216 62648 12265 62676
rect 12216 62636 12222 62648
rect 12253 62645 12265 62648
rect 12299 62676 12311 62679
rect 12526 62676 12532 62688
rect 12299 62648 12532 62676
rect 12299 62645 12311 62648
rect 12253 62639 12311 62645
rect 12526 62636 12532 62648
rect 12584 62636 12590 62688
rect 12728 62676 12756 62775
rect 13078 62772 13084 62784
rect 13136 62772 13142 62824
rect 15010 62772 15016 62824
rect 15068 62812 15074 62824
rect 15381 62815 15439 62821
rect 15381 62812 15393 62815
rect 15068 62784 15393 62812
rect 15068 62772 15074 62784
rect 15381 62781 15393 62784
rect 15427 62812 15439 62815
rect 15746 62812 15752 62824
rect 15427 62784 15752 62812
rect 15427 62781 15439 62784
rect 15381 62775 15439 62781
rect 15746 62772 15752 62784
rect 15804 62772 15810 62824
rect 13354 62676 13360 62688
rect 12728 62648 13360 62676
rect 13354 62636 13360 62648
rect 13412 62636 13418 62688
rect 13814 62636 13820 62688
rect 13872 62676 13878 62688
rect 14093 62679 14151 62685
rect 14093 62676 14105 62679
rect 13872 62648 14105 62676
rect 13872 62636 13878 62648
rect 14093 62645 14105 62648
rect 14139 62645 14151 62679
rect 14093 62639 14151 62645
rect 1104 62586 18860 62608
rect 1104 62534 7648 62586
rect 7700 62534 7712 62586
rect 7764 62534 7776 62586
rect 7828 62534 7840 62586
rect 7892 62534 14315 62586
rect 14367 62534 14379 62586
rect 14431 62534 14443 62586
rect 14495 62534 14507 62586
rect 14559 62534 18860 62586
rect 1104 62512 18860 62534
rect 2406 62472 2412 62484
rect 2367 62444 2412 62472
rect 2406 62432 2412 62444
rect 2464 62432 2470 62484
rect 3878 62432 3884 62484
rect 3936 62472 3942 62484
rect 4617 62475 4675 62481
rect 4617 62472 4629 62475
rect 3936 62444 4629 62472
rect 3936 62432 3942 62444
rect 4617 62441 4629 62444
rect 4663 62472 4675 62475
rect 4798 62472 4804 62484
rect 4663 62444 4804 62472
rect 4663 62441 4675 62444
rect 4617 62435 4675 62441
rect 4798 62432 4804 62444
rect 4856 62432 4862 62484
rect 8941 62475 8999 62481
rect 8941 62441 8953 62475
rect 8987 62441 8999 62475
rect 8941 62435 8999 62441
rect 9677 62475 9735 62481
rect 9677 62441 9689 62475
rect 9723 62472 9735 62475
rect 9858 62472 9864 62484
rect 9723 62444 9864 62472
rect 9723 62441 9735 62444
rect 9677 62435 9735 62441
rect 1581 62339 1639 62345
rect 1581 62305 1593 62339
rect 1627 62336 1639 62339
rect 1670 62336 1676 62348
rect 1627 62308 1676 62336
rect 1627 62305 1639 62308
rect 1581 62299 1639 62305
rect 1670 62296 1676 62308
rect 1728 62296 1734 62348
rect 1765 62339 1823 62345
rect 1765 62305 1777 62339
rect 1811 62336 1823 62339
rect 2424 62336 2452 62432
rect 2866 62364 2872 62416
rect 2924 62404 2930 62416
rect 2961 62407 3019 62413
rect 2961 62404 2973 62407
rect 2924 62376 2973 62404
rect 2924 62364 2930 62376
rect 2961 62373 2973 62376
rect 3007 62373 3019 62407
rect 8956 62404 8984 62435
rect 9858 62432 9864 62444
rect 9916 62432 9922 62484
rect 10226 62472 10232 62484
rect 10187 62444 10232 62472
rect 10226 62432 10232 62444
rect 10284 62432 10290 62484
rect 12621 62475 12679 62481
rect 12621 62441 12633 62475
rect 12667 62472 12679 62475
rect 12710 62472 12716 62484
rect 12667 62444 12716 62472
rect 12667 62441 12679 62444
rect 12621 62435 12679 62441
rect 12710 62432 12716 62444
rect 12768 62432 12774 62484
rect 10244 62404 10272 62432
rect 8956 62376 10272 62404
rect 2961 62367 3019 62373
rect 1811 62308 2452 62336
rect 3789 62339 3847 62345
rect 1811 62305 1823 62308
rect 1765 62299 1823 62305
rect 3789 62305 3801 62339
rect 3835 62336 3847 62339
rect 8757 62339 8815 62345
rect 3835 62308 4384 62336
rect 3835 62305 3847 62308
rect 3789 62299 3847 62305
rect 2130 62268 2136 62280
rect 2043 62240 2136 62268
rect 2130 62228 2136 62240
rect 2188 62268 2194 62280
rect 2777 62271 2835 62277
rect 2777 62268 2789 62271
rect 2188 62240 2789 62268
rect 2188 62228 2194 62240
rect 2777 62237 2789 62240
rect 2823 62237 2835 62271
rect 2777 62231 2835 62237
rect 3418 62228 3424 62280
rect 3476 62268 3482 62280
rect 3513 62271 3571 62277
rect 3513 62268 3525 62271
rect 3476 62240 3525 62268
rect 3476 62228 3482 62240
rect 3513 62237 3525 62240
rect 3559 62237 3571 62271
rect 3970 62268 3976 62280
rect 3931 62240 3976 62268
rect 3513 62231 3571 62237
rect 3970 62228 3976 62240
rect 4028 62228 4034 62280
rect 2958 62160 2964 62212
rect 3016 62200 3022 62212
rect 4062 62200 4068 62212
rect 3016 62172 4068 62200
rect 3016 62160 3022 62172
rect 4062 62160 4068 62172
rect 4120 62160 4126 62212
rect 4356 62209 4384 62308
rect 8757 62305 8769 62339
rect 8803 62336 8815 62339
rect 8938 62336 8944 62348
rect 8803 62308 8944 62336
rect 8803 62305 8815 62308
rect 8757 62299 8815 62305
rect 8938 62296 8944 62308
rect 8996 62296 9002 62348
rect 9769 62339 9827 62345
rect 9769 62305 9781 62339
rect 9815 62336 9827 62339
rect 9858 62336 9864 62348
rect 9815 62308 9864 62336
rect 9815 62305 9827 62308
rect 9769 62299 9827 62305
rect 9858 62296 9864 62308
rect 9916 62296 9922 62348
rect 11330 62336 11336 62348
rect 11291 62308 11336 62336
rect 11330 62296 11336 62308
rect 11388 62296 11394 62348
rect 12434 62296 12440 62348
rect 12492 62336 12498 62348
rect 12897 62339 12955 62345
rect 12897 62336 12909 62339
rect 12492 62308 12909 62336
rect 12492 62296 12498 62308
rect 12897 62305 12909 62308
rect 12943 62305 12955 62339
rect 12897 62299 12955 62305
rect 13354 62296 13360 62348
rect 13412 62336 13418 62348
rect 13725 62339 13783 62345
rect 13725 62336 13737 62339
rect 13412 62308 13737 62336
rect 13412 62296 13418 62308
rect 13725 62305 13737 62308
rect 13771 62336 13783 62339
rect 14274 62336 14280 62348
rect 13771 62308 14280 62336
rect 13771 62305 13783 62308
rect 13725 62299 13783 62305
rect 14274 62296 14280 62308
rect 14332 62296 14338 62348
rect 11514 62268 11520 62280
rect 11475 62240 11520 62268
rect 11514 62228 11520 62240
rect 11572 62228 11578 62280
rect 13998 62268 14004 62280
rect 13959 62240 14004 62268
rect 13998 62228 14004 62240
rect 14056 62228 14062 62280
rect 15194 62268 15200 62280
rect 15155 62240 15200 62268
rect 15194 62228 15200 62240
rect 15252 62228 15258 62280
rect 15562 62228 15568 62280
rect 15620 62268 15626 62280
rect 16025 62271 16083 62277
rect 16025 62268 16037 62271
rect 15620 62240 16037 62268
rect 15620 62228 15626 62240
rect 16025 62237 16037 62240
rect 16071 62237 16083 62271
rect 16025 62231 16083 62237
rect 4341 62203 4399 62209
rect 4341 62169 4353 62203
rect 4387 62200 4399 62203
rect 4706 62200 4712 62212
rect 4387 62172 4712 62200
rect 4387 62169 4399 62172
rect 4341 62163 4399 62169
rect 4706 62160 4712 62172
rect 4764 62160 4770 62212
rect 9309 62203 9367 62209
rect 9309 62169 9321 62203
rect 9355 62200 9367 62203
rect 9766 62200 9772 62212
rect 9355 62172 9772 62200
rect 9355 62169 9367 62172
rect 9309 62163 9367 62169
rect 9766 62160 9772 62172
rect 9824 62200 9830 62212
rect 10134 62200 10140 62212
rect 9824 62172 10140 62200
rect 9824 62160 9830 62172
rect 10134 62160 10140 62172
rect 10192 62160 10198 62212
rect 9490 62092 9496 62144
rect 9548 62132 9554 62144
rect 9953 62135 10011 62141
rect 9953 62132 9965 62135
rect 9548 62104 9965 62132
rect 9548 62092 9554 62104
rect 9953 62101 9965 62104
rect 9999 62101 10011 62135
rect 10686 62132 10692 62144
rect 10647 62104 10692 62132
rect 9953 62095 10011 62101
rect 10686 62092 10692 62104
rect 10744 62092 10750 62144
rect 13633 62135 13691 62141
rect 13633 62101 13645 62135
rect 13679 62132 13691 62135
rect 13722 62132 13728 62144
rect 13679 62104 13728 62132
rect 13679 62101 13691 62104
rect 13633 62095 13691 62101
rect 13722 62092 13728 62104
rect 13780 62132 13786 62144
rect 15378 62132 15384 62144
rect 13780 62104 15384 62132
rect 13780 62092 13786 62104
rect 15378 62092 15384 62104
rect 15436 62092 15442 62144
rect 1104 62042 18860 62064
rect 1104 61990 4315 62042
rect 4367 61990 4379 62042
rect 4431 61990 4443 62042
rect 4495 61990 4507 62042
rect 4559 61990 10982 62042
rect 11034 61990 11046 62042
rect 11098 61990 11110 62042
rect 11162 61990 11174 62042
rect 11226 61990 17648 62042
rect 17700 61990 17712 62042
rect 17764 61990 17776 62042
rect 17828 61990 17840 62042
rect 17892 61990 18860 62042
rect 1104 61968 18860 61990
rect 3053 61931 3111 61937
rect 3053 61897 3065 61931
rect 3099 61928 3111 61931
rect 3145 61931 3203 61937
rect 3145 61928 3157 61931
rect 3099 61900 3157 61928
rect 3099 61897 3111 61900
rect 3053 61891 3111 61897
rect 3145 61897 3157 61900
rect 3191 61928 3203 61931
rect 3970 61928 3976 61940
rect 3191 61900 3976 61928
rect 3191 61897 3203 61900
rect 3145 61891 3203 61897
rect 3970 61888 3976 61900
rect 4028 61888 4034 61940
rect 6914 61888 6920 61940
rect 6972 61928 6978 61940
rect 7098 61928 7104 61940
rect 6972 61900 7104 61928
rect 6972 61888 6978 61900
rect 7098 61888 7104 61900
rect 7156 61888 7162 61940
rect 8754 61888 8760 61940
rect 8812 61928 8818 61940
rect 9401 61931 9459 61937
rect 9401 61928 9413 61931
rect 8812 61900 9413 61928
rect 8812 61888 8818 61900
rect 9401 61897 9413 61900
rect 9447 61897 9459 61931
rect 9401 61891 9459 61897
rect 11149 61931 11207 61937
rect 11149 61897 11161 61931
rect 11195 61928 11207 61931
rect 11330 61928 11336 61940
rect 11195 61900 11336 61928
rect 11195 61897 11207 61900
rect 11149 61891 11207 61897
rect 8849 61863 8907 61869
rect 8849 61829 8861 61863
rect 8895 61860 8907 61863
rect 8938 61860 8944 61872
rect 8895 61832 8944 61860
rect 8895 61829 8907 61832
rect 8849 61823 8907 61829
rect 8938 61820 8944 61832
rect 8996 61820 9002 61872
rect 2041 61795 2099 61801
rect 2041 61761 2053 61795
rect 2087 61792 2099 61795
rect 2130 61792 2136 61804
rect 2087 61764 2136 61792
rect 2087 61761 2099 61764
rect 2041 61755 2099 61761
rect 2130 61752 2136 61764
rect 2188 61752 2194 61804
rect 2498 61792 2504 61804
rect 2240 61764 2504 61792
rect 1670 61684 1676 61736
rect 1728 61724 1734 61736
rect 2240 61724 2268 61764
rect 2498 61752 2504 61764
rect 2556 61752 2562 61804
rect 2682 61752 2688 61804
rect 2740 61792 2746 61804
rect 3878 61792 3884 61804
rect 2740 61764 3884 61792
rect 2740 61752 2746 61764
rect 3878 61752 3884 61764
rect 3936 61792 3942 61804
rect 4065 61795 4123 61801
rect 4065 61792 4077 61795
rect 3936 61764 4077 61792
rect 3936 61752 3942 61764
rect 4065 61761 4077 61764
rect 4111 61761 4123 61795
rect 4065 61755 4123 61761
rect 8478 61752 8484 61804
rect 8536 61792 8542 61804
rect 9122 61792 9128 61804
rect 8536 61764 9128 61792
rect 8536 61752 8542 61764
rect 9122 61752 9128 61764
rect 9180 61752 9186 61804
rect 9416 61792 9444 61891
rect 11330 61888 11336 61900
rect 11388 61888 11394 61940
rect 11514 61888 11520 61940
rect 11572 61928 11578 61940
rect 11793 61931 11851 61937
rect 11793 61928 11805 61931
rect 11572 61900 11805 61928
rect 11572 61888 11578 61900
rect 11793 61897 11805 61900
rect 11839 61897 11851 61931
rect 14734 61928 14740 61940
rect 14695 61900 14740 61928
rect 11793 61891 11851 61897
rect 11808 61792 11836 61891
rect 14734 61888 14740 61900
rect 14792 61888 14798 61940
rect 12253 61863 12311 61869
rect 12253 61829 12265 61863
rect 12299 61860 12311 61863
rect 13262 61860 13268 61872
rect 12299 61832 13268 61860
rect 12299 61829 12311 61832
rect 12253 61823 12311 61829
rect 13262 61820 13268 61832
rect 13320 61820 13326 61872
rect 14274 61860 14280 61872
rect 14187 61832 14280 61860
rect 14274 61820 14280 61832
rect 14332 61860 14338 61872
rect 14642 61860 14648 61872
rect 14332 61832 14648 61860
rect 14332 61820 14338 61832
rect 14642 61820 14648 61832
rect 14700 61860 14706 61872
rect 15010 61860 15016 61872
rect 14700 61832 15016 61860
rect 14700 61820 14706 61832
rect 15010 61820 15016 61832
rect 15068 61820 15074 61872
rect 13541 61795 13599 61801
rect 9416 61764 10180 61792
rect 11808 61764 12756 61792
rect 1728 61696 2268 61724
rect 2317 61727 2375 61733
rect 1728 61684 1734 61696
rect 2317 61693 2329 61727
rect 2363 61693 2375 61727
rect 2317 61687 2375 61693
rect 4341 61727 4399 61733
rect 4341 61693 4353 61727
rect 4387 61724 4399 61727
rect 4706 61724 4712 61736
rect 4387 61696 4712 61724
rect 4387 61693 4399 61696
rect 4341 61687 4399 61693
rect 1486 61656 1492 61668
rect 1447 61628 1492 61656
rect 1486 61616 1492 61628
rect 1544 61616 1550 61668
rect 2332 61656 2360 61687
rect 4706 61684 4712 61696
rect 4764 61684 4770 61736
rect 10152 61733 10180 61764
rect 12728 61736 12756 61764
rect 13541 61761 13553 61795
rect 13587 61792 13599 61795
rect 13630 61792 13636 61804
rect 13587 61764 13636 61792
rect 13587 61761 13599 61764
rect 13541 61755 13599 61761
rect 13630 61752 13636 61764
rect 13688 61752 13694 61804
rect 15105 61795 15163 61801
rect 15105 61761 15117 61795
rect 15151 61792 15163 61795
rect 15151 61764 15608 61792
rect 15151 61761 15163 61764
rect 15105 61755 15163 61761
rect 15580 61736 15608 61764
rect 9953 61727 10011 61733
rect 9953 61693 9965 61727
rect 9999 61693 10011 61727
rect 9953 61687 10011 61693
rect 10137 61727 10195 61733
rect 10137 61693 10149 61727
rect 10183 61693 10195 61727
rect 10137 61687 10195 61693
rect 3050 61656 3056 61668
rect 2332 61628 3056 61656
rect 3050 61616 3056 61628
rect 3108 61656 3114 61668
rect 3697 61659 3755 61665
rect 3697 61656 3709 61659
rect 3108 61628 3709 61656
rect 3108 61616 3114 61628
rect 3697 61625 3709 61628
rect 3743 61625 3755 61659
rect 9968 61656 9996 61687
rect 10318 61684 10324 61736
rect 10376 61724 10382 61736
rect 10505 61727 10563 61733
rect 10505 61724 10517 61727
rect 10376 61696 10517 61724
rect 10376 61684 10382 61696
rect 10505 61693 10517 61696
rect 10551 61693 10563 61727
rect 10505 61687 10563 61693
rect 11517 61727 11575 61733
rect 11517 61693 11529 61727
rect 11563 61724 11575 61727
rect 12529 61727 12587 61733
rect 12529 61724 12541 61727
rect 11563 61696 12541 61724
rect 11563 61693 11575 61696
rect 11517 61687 11575 61693
rect 12529 61693 12541 61696
rect 12575 61693 12587 61727
rect 12710 61724 12716 61736
rect 12623 61696 12716 61724
rect 12529 61687 12587 61693
rect 10226 61656 10232 61668
rect 9968 61628 10232 61656
rect 3697 61619 3755 61625
rect 10226 61616 10232 61628
rect 10284 61616 10290 61668
rect 12544 61656 12572 61687
rect 12710 61684 12716 61696
rect 12768 61684 12774 61736
rect 13262 61724 13268 61736
rect 13223 61696 13268 61724
rect 13262 61684 13268 61696
rect 13320 61684 13326 61736
rect 14734 61684 14740 61736
rect 14792 61724 14798 61736
rect 15289 61727 15347 61733
rect 15289 61724 15301 61727
rect 14792 61696 15301 61724
rect 14792 61684 14798 61696
rect 15289 61693 15301 61696
rect 15335 61693 15347 61727
rect 15562 61724 15568 61736
rect 15523 61696 15568 61724
rect 15289 61687 15347 61693
rect 12618 61656 12624 61668
rect 12531 61628 12624 61656
rect 12618 61616 12624 61628
rect 12676 61656 12682 61668
rect 13722 61656 13728 61668
rect 12676 61628 13728 61656
rect 12676 61616 12682 61628
rect 13722 61616 13728 61628
rect 13780 61616 13786 61668
rect 3142 61588 3148 61600
rect 3103 61560 3148 61588
rect 3142 61548 3148 61560
rect 3200 61548 3206 61600
rect 3418 61588 3424 61600
rect 3379 61560 3424 61588
rect 3418 61548 3424 61560
rect 3476 61548 3482 61600
rect 5442 61588 5448 61600
rect 5403 61560 5448 61588
rect 5442 61548 5448 61560
rect 5500 61548 5506 61600
rect 8478 61588 8484 61600
rect 8439 61560 8484 61588
rect 8478 61548 8484 61560
rect 8536 61548 8542 61600
rect 9953 61591 10011 61597
rect 9953 61557 9965 61591
rect 9999 61588 10011 61591
rect 10134 61588 10140 61600
rect 9999 61560 10140 61588
rect 9999 61557 10011 61560
rect 9953 61551 10011 61557
rect 10134 61548 10140 61560
rect 10192 61548 10198 61600
rect 11514 61548 11520 61600
rect 11572 61588 11578 61600
rect 11698 61588 11704 61600
rect 11572 61560 11704 61588
rect 11572 61548 11578 61560
rect 11698 61548 11704 61560
rect 11756 61548 11762 61600
rect 13909 61591 13967 61597
rect 13909 61557 13921 61591
rect 13955 61588 13967 61591
rect 13998 61588 14004 61600
rect 13955 61560 14004 61588
rect 13955 61557 13967 61560
rect 13909 61551 13967 61557
rect 13998 61548 14004 61560
rect 14056 61588 14062 61600
rect 14918 61588 14924 61600
rect 14056 61560 14924 61588
rect 14056 61548 14062 61560
rect 14918 61548 14924 61560
rect 14976 61548 14982 61600
rect 15304 61588 15332 61687
rect 15562 61684 15568 61696
rect 15620 61684 15626 61736
rect 15930 61588 15936 61600
rect 15304 61560 15936 61588
rect 15930 61548 15936 61560
rect 15988 61548 15994 61600
rect 16666 61588 16672 61600
rect 16627 61560 16672 61588
rect 16666 61548 16672 61560
rect 16724 61548 16730 61600
rect 1104 61498 18860 61520
rect 1104 61446 7648 61498
rect 7700 61446 7712 61498
rect 7764 61446 7776 61498
rect 7828 61446 7840 61498
rect 7892 61446 14315 61498
rect 14367 61446 14379 61498
rect 14431 61446 14443 61498
rect 14495 61446 14507 61498
rect 14559 61446 18860 61498
rect 1104 61424 18860 61446
rect 3050 61384 3056 61396
rect 3011 61356 3056 61384
rect 3050 61344 3056 61356
rect 3108 61344 3114 61396
rect 3418 61344 3424 61396
rect 3476 61384 3482 61396
rect 4249 61387 4307 61393
rect 4249 61384 4261 61387
rect 3476 61356 4261 61384
rect 3476 61344 3482 61356
rect 4249 61353 4261 61356
rect 4295 61353 4307 61387
rect 4798 61384 4804 61396
rect 4759 61356 4804 61384
rect 4249 61347 4307 61353
rect 4798 61344 4804 61356
rect 4856 61344 4862 61396
rect 9766 61384 9772 61396
rect 9679 61356 9772 61384
rect 9766 61344 9772 61356
rect 9824 61384 9830 61396
rect 10226 61384 10232 61396
rect 9824 61356 10232 61384
rect 9824 61344 9830 61356
rect 10226 61344 10232 61356
rect 10284 61344 10290 61396
rect 3513 61319 3571 61325
rect 3513 61285 3525 61319
rect 3559 61316 3571 61319
rect 4706 61316 4712 61328
rect 3559 61288 4712 61316
rect 3559 61285 3571 61288
rect 3513 61279 3571 61285
rect 4706 61276 4712 61288
rect 4764 61276 4770 61328
rect 7374 61276 7380 61328
rect 7432 61316 7438 61328
rect 7558 61316 7564 61328
rect 7432 61288 7564 61316
rect 7432 61276 7438 61288
rect 7558 61276 7564 61288
rect 7616 61276 7622 61328
rect 8018 61276 8024 61328
rect 8076 61316 8082 61328
rect 13446 61316 13452 61328
rect 8076 61288 8984 61316
rect 8076 61276 8082 61288
rect 1210 61208 1216 61260
rect 1268 61248 1274 61260
rect 1489 61251 1547 61257
rect 1489 61248 1501 61251
rect 1268 61220 1501 61248
rect 1268 61208 1274 61220
rect 1489 61217 1501 61220
rect 1535 61248 1547 61251
rect 2682 61248 2688 61260
rect 1535 61220 2688 61248
rect 1535 61217 1547 61220
rect 1489 61211 1547 61217
rect 2682 61208 2688 61220
rect 2740 61208 2746 61260
rect 3694 61208 3700 61260
rect 3752 61248 3758 61260
rect 3973 61251 4031 61257
rect 3973 61248 3985 61251
rect 3752 61220 3985 61248
rect 3752 61208 3758 61220
rect 3973 61217 3985 61220
rect 4019 61217 4031 61251
rect 3973 61211 4031 61217
rect 4157 61251 4215 61257
rect 4157 61217 4169 61251
rect 4203 61248 4215 61251
rect 5442 61248 5448 61260
rect 4203 61220 5448 61248
rect 4203 61217 4215 61220
rect 4157 61211 4215 61217
rect 1762 61180 1768 61192
rect 1723 61152 1768 61180
rect 1762 61140 1768 61152
rect 1820 61180 1826 61192
rect 3789 61183 3847 61189
rect 3789 61180 3801 61183
rect 1820 61152 3801 61180
rect 1820 61140 1826 61152
rect 3789 61149 3801 61152
rect 3835 61149 3847 61183
rect 3789 61143 3847 61149
rect 3418 61072 3424 61124
rect 3476 61112 3482 61124
rect 4172 61112 4200 61211
rect 5442 61208 5448 61220
rect 5500 61208 5506 61260
rect 8294 61248 8300 61260
rect 8255 61220 8300 61248
rect 8294 61208 8300 61220
rect 8352 61208 8358 61260
rect 8754 61248 8760 61260
rect 8715 61220 8760 61248
rect 8754 61208 8760 61220
rect 8812 61208 8818 61260
rect 8956 61257 8984 61288
rect 13004 61288 13452 61316
rect 8941 61251 8999 61257
rect 8941 61217 8953 61251
rect 8987 61248 8999 61251
rect 9766 61248 9772 61260
rect 8987 61220 9772 61248
rect 8987 61217 8999 61220
rect 8941 61211 8999 61217
rect 9766 61208 9772 61220
rect 9824 61208 9830 61260
rect 9858 61208 9864 61260
rect 9916 61248 9922 61260
rect 10505 61251 10563 61257
rect 10505 61248 10517 61251
rect 9916 61220 10517 61248
rect 9916 61208 9922 61220
rect 10505 61217 10517 61220
rect 10551 61217 10563 61251
rect 11054 61248 11060 61260
rect 11015 61220 11060 61248
rect 10505 61211 10563 61217
rect 11054 61208 11060 61220
rect 11112 61248 11118 61260
rect 11422 61248 11428 61260
rect 11112 61220 11428 61248
rect 11112 61208 11118 61220
rect 11422 61208 11428 61220
rect 11480 61208 11486 61260
rect 13004 61257 13032 61288
rect 13446 61276 13452 61288
rect 13504 61276 13510 61328
rect 12989 61251 13047 61257
rect 12989 61217 13001 61251
rect 13035 61217 13047 61251
rect 13170 61248 13176 61260
rect 13131 61220 13176 61248
rect 12989 61211 13047 61217
rect 13170 61208 13176 61220
rect 13228 61208 13234 61260
rect 13814 61208 13820 61260
rect 13872 61248 13878 61260
rect 14642 61248 14648 61260
rect 13872 61220 14648 61248
rect 13872 61208 13878 61220
rect 14642 61208 14648 61220
rect 14700 61248 14706 61260
rect 14737 61251 14795 61257
rect 14737 61248 14749 61251
rect 14700 61220 14749 61248
rect 14700 61208 14706 61220
rect 14737 61217 14749 61220
rect 14783 61217 14795 61251
rect 14737 61211 14795 61217
rect 7190 61140 7196 61192
rect 7248 61180 7254 61192
rect 7374 61180 7380 61192
rect 7248 61152 7380 61180
rect 7248 61140 7254 61152
rect 7374 61140 7380 61152
rect 7432 61140 7438 61192
rect 3476 61084 4200 61112
rect 8312 61112 8340 61208
rect 8772 61180 8800 61208
rect 9030 61180 9036 61192
rect 8772 61152 9036 61180
rect 9030 61140 9036 61152
rect 9088 61140 9094 61192
rect 9490 61140 9496 61192
rect 9548 61180 9554 61192
rect 10042 61180 10048 61192
rect 9548 61152 10048 61180
rect 9548 61140 9554 61152
rect 10042 61140 10048 61152
rect 10100 61140 10106 61192
rect 10873 61183 10931 61189
rect 10873 61149 10885 61183
rect 10919 61180 10931 61183
rect 11330 61180 11336 61192
rect 10919 61152 11336 61180
rect 10919 61149 10931 61152
rect 10873 61143 10931 61149
rect 11330 61140 11336 61152
rect 11388 61140 11394 61192
rect 13449 61183 13507 61189
rect 13449 61149 13461 61183
rect 13495 61180 13507 61183
rect 13630 61180 13636 61192
rect 13495 61152 13636 61180
rect 13495 61149 13507 61152
rect 13449 61143 13507 61149
rect 13630 61140 13636 61152
rect 13688 61140 13694 61192
rect 15010 61180 15016 61192
rect 14971 61152 15016 61180
rect 15010 61140 15016 61152
rect 15068 61140 15074 61192
rect 8312 61084 8708 61112
rect 3476 61072 3482 61084
rect 8680 61056 8708 61084
rect 4062 61004 4068 61056
rect 4120 61044 4126 61056
rect 4614 61044 4620 61056
rect 4120 61016 4620 61044
rect 4120 61004 4126 61016
rect 4614 61004 4620 61016
rect 4672 61004 4678 61056
rect 8294 61044 8300 61056
rect 8255 61016 8300 61044
rect 8294 61004 8300 61016
rect 8352 61004 8358 61056
rect 8662 61004 8668 61056
rect 8720 61004 8726 61056
rect 10137 61047 10195 61053
rect 10137 61013 10149 61047
rect 10183 61044 10195 61047
rect 10226 61044 10232 61056
rect 10183 61016 10232 61044
rect 10183 61013 10195 61016
rect 10137 61007 10195 61013
rect 10226 61004 10232 61016
rect 10284 61004 10290 61056
rect 11977 61047 12035 61053
rect 11977 61013 11989 61047
rect 12023 61044 12035 61047
rect 12342 61044 12348 61056
rect 12023 61016 12348 61044
rect 12023 61013 12035 61016
rect 11977 61007 12035 61013
rect 12342 61004 12348 61016
rect 12400 61004 12406 61056
rect 16114 61044 16120 61056
rect 16075 61016 16120 61044
rect 16114 61004 16120 61016
rect 16172 61004 16178 61056
rect 1104 60954 18860 60976
rect 1104 60902 4315 60954
rect 4367 60902 4379 60954
rect 4431 60902 4443 60954
rect 4495 60902 4507 60954
rect 4559 60902 10982 60954
rect 11034 60902 11046 60954
rect 11098 60902 11110 60954
rect 11162 60902 11174 60954
rect 11226 60902 17648 60954
rect 17700 60902 17712 60954
rect 17764 60902 17776 60954
rect 17828 60902 17840 60954
rect 17892 60902 18860 60954
rect 1104 60880 18860 60902
rect 3418 60840 3424 60852
rect 3379 60812 3424 60840
rect 3418 60800 3424 60812
rect 3476 60800 3482 60852
rect 3694 60800 3700 60852
rect 3752 60840 3758 60852
rect 3789 60843 3847 60849
rect 3789 60840 3801 60843
rect 3752 60812 3801 60840
rect 3752 60800 3758 60812
rect 3789 60809 3801 60812
rect 3835 60840 3847 60843
rect 3835 60812 4016 60840
rect 3835 60809 3847 60812
rect 3789 60803 3847 60809
rect 1946 60664 1952 60716
rect 2004 60704 2010 60716
rect 2133 60707 2191 60713
rect 2133 60704 2145 60707
rect 2004 60676 2145 60704
rect 2004 60664 2010 60676
rect 2133 60673 2145 60676
rect 2179 60673 2191 60707
rect 3988 60704 4016 60812
rect 5258 60800 5264 60852
rect 5316 60840 5322 60852
rect 5534 60840 5540 60852
rect 5316 60812 5540 60840
rect 5316 60800 5322 60812
rect 5534 60800 5540 60812
rect 5592 60800 5598 60852
rect 8478 60800 8484 60852
rect 8536 60840 8542 60852
rect 9401 60843 9459 60849
rect 9401 60840 9413 60843
rect 8536 60812 9413 60840
rect 8536 60800 8542 60812
rect 9401 60809 9413 60812
rect 9447 60840 9459 60843
rect 9858 60840 9864 60852
rect 9447 60812 9864 60840
rect 9447 60809 9459 60812
rect 9401 60803 9459 60809
rect 9858 60800 9864 60812
rect 9916 60800 9922 60852
rect 10042 60800 10048 60852
rect 10100 60840 10106 60852
rect 10137 60843 10195 60849
rect 10137 60840 10149 60843
rect 10100 60812 10149 60840
rect 10100 60800 10106 60812
rect 10137 60809 10149 60812
rect 10183 60840 10195 60843
rect 11422 60840 11428 60852
rect 10183 60812 10732 60840
rect 11383 60812 11428 60840
rect 10183 60809 10195 60812
rect 10137 60803 10195 60809
rect 10413 60775 10471 60781
rect 10413 60741 10425 60775
rect 10459 60741 10471 60775
rect 10413 60735 10471 60741
rect 3988 60676 4108 60704
rect 2133 60667 2191 60673
rect 2682 60636 2688 60648
rect 2643 60608 2688 60636
rect 2682 60596 2688 60608
rect 2740 60596 2746 60648
rect 2866 60596 2872 60648
rect 2924 60636 2930 60648
rect 2961 60639 3019 60645
rect 2961 60636 2973 60639
rect 2924 60608 2973 60636
rect 2924 60596 2930 60608
rect 2961 60605 2973 60608
rect 3007 60605 3019 60639
rect 2961 60599 3019 60605
rect 3050 60596 3056 60648
rect 3108 60636 3114 60648
rect 3145 60639 3203 60645
rect 3145 60636 3157 60639
rect 3108 60608 3157 60636
rect 3108 60596 3114 60608
rect 3145 60605 3157 60608
rect 3191 60605 3203 60639
rect 3145 60599 3203 60605
rect 2041 60571 2099 60577
rect 2041 60537 2053 60571
rect 2087 60568 2099 60571
rect 3068 60568 3096 60596
rect 4080 60577 4108 60676
rect 8938 60664 8944 60716
rect 8996 60704 9002 60716
rect 9122 60704 9128 60716
rect 8996 60676 9128 60704
rect 8996 60664 9002 60676
rect 9122 60664 9128 60676
rect 9180 60664 9186 60716
rect 10428 60648 10456 60735
rect 4249 60639 4307 60645
rect 4249 60605 4261 60639
rect 4295 60636 4307 60639
rect 4614 60636 4620 60648
rect 4295 60608 4620 60636
rect 4295 60605 4307 60608
rect 4249 60599 4307 60605
rect 4614 60596 4620 60608
rect 4672 60636 4678 60648
rect 5261 60639 5319 60645
rect 5261 60636 5273 60639
rect 4672 60608 5273 60636
rect 4672 60596 4678 60608
rect 5261 60605 5273 60608
rect 5307 60605 5319 60639
rect 8294 60636 8300 60648
rect 8255 60608 8300 60636
rect 5261 60599 5319 60605
rect 8294 60596 8300 60608
rect 8352 60596 8358 60648
rect 10410 60596 10416 60648
rect 10468 60596 10474 60648
rect 10594 60636 10600 60648
rect 10555 60608 10600 60636
rect 10594 60596 10600 60608
rect 10652 60596 10658 60648
rect 10704 60636 10732 60812
rect 11422 60800 11428 60812
rect 11480 60800 11486 60852
rect 13170 60800 13176 60852
rect 13228 60840 13234 60852
rect 13725 60843 13783 60849
rect 13725 60840 13737 60843
rect 13228 60812 13737 60840
rect 13228 60800 13234 60812
rect 13725 60809 13737 60812
rect 13771 60809 13783 60843
rect 13725 60803 13783 60809
rect 11790 60772 11796 60784
rect 11440 60744 11796 60772
rect 11440 60716 11468 60744
rect 11790 60732 11796 60744
rect 11848 60732 11854 60784
rect 14642 60732 14648 60784
rect 14700 60772 14706 60784
rect 14700 60744 15148 60772
rect 14700 60732 14706 60744
rect 11422 60664 11428 60716
rect 11480 60664 11486 60716
rect 11974 60704 11980 60716
rect 11808 60676 11980 60704
rect 11808 60648 11836 60676
rect 11974 60664 11980 60676
rect 12032 60664 12038 60716
rect 12526 60704 12532 60716
rect 12487 60676 12532 60704
rect 12526 60664 12532 60676
rect 12584 60664 12590 60716
rect 15120 60704 15148 60744
rect 15473 60707 15531 60713
rect 15473 60704 15485 60707
rect 15120 60676 15485 60704
rect 15473 60673 15485 60676
rect 15519 60673 15531 60707
rect 15473 60667 15531 60673
rect 16025 60707 16083 60713
rect 16025 60673 16037 60707
rect 16071 60704 16083 60707
rect 16071 60676 16436 60704
rect 16071 60673 16083 60676
rect 16025 60667 16083 60673
rect 10873 60639 10931 60645
rect 10873 60636 10885 60639
rect 10704 60608 10885 60636
rect 10873 60605 10885 60608
rect 10919 60605 10931 60639
rect 10873 60599 10931 60605
rect 11790 60596 11796 60648
rect 11848 60596 11854 60648
rect 11885 60639 11943 60645
rect 11885 60605 11897 60639
rect 11931 60605 11943 60639
rect 11885 60599 11943 60605
rect 2087 60540 3096 60568
rect 4065 60571 4123 60577
rect 2087 60537 2099 60540
rect 2041 60531 2099 60537
rect 4065 60537 4077 60571
rect 4111 60568 4123 60571
rect 4893 60571 4951 60577
rect 4893 60568 4905 60571
rect 4111 60540 4905 60568
rect 4111 60537 4123 60540
rect 4065 60531 4123 60537
rect 4893 60537 4905 60540
rect 4939 60537 4951 60571
rect 4893 60531 4951 60537
rect 1670 60500 1676 60512
rect 1631 60472 1676 60500
rect 1670 60460 1676 60472
rect 1728 60460 1734 60512
rect 4338 60500 4344 60512
rect 4299 60472 4344 60500
rect 4338 60460 4344 60472
rect 4396 60460 4402 60512
rect 7837 60503 7895 60509
rect 7837 60469 7849 60503
rect 7883 60500 7895 60503
rect 8018 60500 8024 60512
rect 7883 60472 8024 60500
rect 7883 60469 7895 60472
rect 7837 60463 7895 60469
rect 8018 60460 8024 60472
rect 8076 60460 8082 60512
rect 8386 60500 8392 60512
rect 8347 60472 8392 60500
rect 8386 60460 8392 60472
rect 8444 60460 8450 60512
rect 9033 60503 9091 60509
rect 9033 60469 9045 60503
rect 9079 60500 9091 60503
rect 9122 60500 9128 60512
rect 9079 60472 9128 60500
rect 9079 60469 9091 60472
rect 9033 60463 9091 60469
rect 9122 60460 9128 60472
rect 9180 60460 9186 60512
rect 11793 60503 11851 60509
rect 11793 60469 11805 60503
rect 11839 60500 11851 60503
rect 11900 60500 11928 60599
rect 12434 60596 12440 60648
rect 12492 60636 12498 60648
rect 12710 60636 12716 60648
rect 12492 60608 12537 60636
rect 12671 60608 12716 60636
rect 12492 60596 12498 60608
rect 12710 60596 12716 60608
rect 12768 60596 12774 60648
rect 15488 60636 15516 60667
rect 16114 60636 16120 60648
rect 15488 60608 16120 60636
rect 16114 60596 16120 60608
rect 16172 60596 16178 60648
rect 16408 60645 16436 60676
rect 16393 60639 16451 60645
rect 16393 60605 16405 60639
rect 16439 60636 16451 60639
rect 16482 60636 16488 60648
rect 16439 60608 16488 60636
rect 16439 60605 16451 60608
rect 16393 60599 16451 60605
rect 16482 60596 16488 60608
rect 16540 60596 16546 60648
rect 11974 60500 11980 60512
rect 11839 60472 11980 60500
rect 11839 60469 11851 60472
rect 11793 60463 11851 60469
rect 11974 60460 11980 60472
rect 12032 60460 12038 60512
rect 13446 60500 13452 60512
rect 13407 60472 13452 60500
rect 13446 60460 13452 60472
rect 13504 60460 13510 60512
rect 14829 60503 14887 60509
rect 14829 60469 14841 60503
rect 14875 60500 14887 60503
rect 15010 60500 15016 60512
rect 14875 60472 15016 60500
rect 14875 60469 14887 60472
rect 14829 60463 14887 60469
rect 15010 60460 15016 60472
rect 15068 60460 15074 60512
rect 17494 60500 17500 60512
rect 17455 60472 17500 60500
rect 17494 60460 17500 60472
rect 17552 60460 17558 60512
rect 1104 60410 18860 60432
rect 1104 60358 7648 60410
rect 7700 60358 7712 60410
rect 7764 60358 7776 60410
rect 7828 60358 7840 60410
rect 7892 60358 14315 60410
rect 14367 60358 14379 60410
rect 14431 60358 14443 60410
rect 14495 60358 14507 60410
rect 14559 60358 18860 60410
rect 1104 60336 18860 60358
rect 2225 60299 2283 60305
rect 2225 60265 2237 60299
rect 2271 60296 2283 60299
rect 2682 60296 2688 60308
rect 2271 60268 2688 60296
rect 2271 60265 2283 60268
rect 2225 60259 2283 60265
rect 2682 60256 2688 60268
rect 2740 60256 2746 60308
rect 4614 60296 4620 60308
rect 4575 60268 4620 60296
rect 4614 60256 4620 60268
rect 4672 60256 4678 60308
rect 7101 60299 7159 60305
rect 7101 60265 7113 60299
rect 7147 60296 7159 60299
rect 7374 60296 7380 60308
rect 7147 60268 7380 60296
rect 7147 60265 7159 60268
rect 7101 60259 7159 60265
rect 7374 60256 7380 60268
rect 7432 60256 7438 60308
rect 8021 60299 8079 60305
rect 8021 60265 8033 60299
rect 8067 60296 8079 60299
rect 8294 60296 8300 60308
rect 8067 60268 8300 60296
rect 8067 60265 8079 60268
rect 8021 60259 8079 60265
rect 8294 60256 8300 60268
rect 8352 60256 8358 60308
rect 9766 60256 9772 60308
rect 9824 60296 9830 60308
rect 10137 60299 10195 60305
rect 10137 60296 10149 60299
rect 9824 60268 10149 60296
rect 9824 60256 9830 60268
rect 10137 60265 10149 60268
rect 10183 60265 10195 60299
rect 10137 60259 10195 60265
rect 10410 60256 10416 60308
rect 10468 60256 10474 60308
rect 11977 60299 12035 60305
rect 11977 60265 11989 60299
rect 12023 60296 12035 60299
rect 12710 60296 12716 60308
rect 12023 60268 12716 60296
rect 12023 60265 12035 60268
rect 11977 60259 12035 60265
rect 12710 60256 12716 60268
rect 12768 60256 12774 60308
rect 14001 60299 14059 60305
rect 14001 60265 14013 60299
rect 14047 60296 14059 60299
rect 14734 60296 14740 60308
rect 14047 60268 14740 60296
rect 14047 60265 14059 60268
rect 14001 60259 14059 60265
rect 2774 60120 2780 60172
rect 2832 60160 2838 60172
rect 3237 60163 3295 60169
rect 3237 60160 3249 60163
rect 2832 60132 3249 60160
rect 2832 60120 2838 60132
rect 3237 60129 3249 60132
rect 3283 60160 3295 60163
rect 6089 60163 6147 60169
rect 3283 60132 3740 60160
rect 3283 60129 3295 60132
rect 3237 60123 3295 60129
rect 3712 60104 3740 60132
rect 6089 60129 6101 60163
rect 6135 60160 6147 60163
rect 6365 60163 6423 60169
rect 6365 60160 6377 60163
rect 6135 60132 6377 60160
rect 6135 60129 6147 60132
rect 6089 60123 6147 60129
rect 6365 60129 6377 60132
rect 6411 60160 6423 60163
rect 6454 60160 6460 60172
rect 6411 60132 6460 60160
rect 6411 60129 6423 60132
rect 6365 60123 6423 60129
rect 6454 60120 6460 60132
rect 6512 60120 6518 60172
rect 8662 60120 8668 60172
rect 8720 60160 8726 60172
rect 8757 60163 8815 60169
rect 8757 60160 8769 60163
rect 8720 60132 8769 60160
rect 8720 60120 8726 60132
rect 8757 60129 8769 60132
rect 8803 60129 8815 60163
rect 10428 60160 10456 60256
rect 14016 60228 14044 60259
rect 14734 60256 14740 60268
rect 14792 60256 14798 60308
rect 16114 60296 16120 60308
rect 16075 60268 16120 60296
rect 16114 60256 16120 60268
rect 16172 60256 16178 60308
rect 12728 60200 14044 60228
rect 10870 60160 10876 60172
rect 10428 60132 10876 60160
rect 8757 60123 8815 60129
rect 10870 60120 10876 60132
rect 10928 60120 10934 60172
rect 12434 60120 12440 60172
rect 12492 60160 12498 60172
rect 12728 60169 12756 60200
rect 12713 60163 12771 60169
rect 12713 60160 12725 60163
rect 12492 60132 12725 60160
rect 12492 60120 12498 60132
rect 12713 60129 12725 60132
rect 12759 60129 12771 60163
rect 12713 60123 12771 60129
rect 12805 60163 12863 60169
rect 12805 60129 12817 60163
rect 12851 60129 12863 60163
rect 12805 60123 12863 60129
rect 2866 60052 2872 60104
rect 2924 60092 2930 60104
rect 2961 60095 3019 60101
rect 2961 60092 2973 60095
rect 2924 60064 2973 60092
rect 2924 60052 2930 60064
rect 2961 60061 2973 60064
rect 3007 60092 3019 60095
rect 3418 60092 3424 60104
rect 3007 60064 3424 60092
rect 3007 60061 3019 60064
rect 2961 60055 3019 60061
rect 3418 60052 3424 60064
rect 3476 60092 3482 60104
rect 3513 60095 3571 60101
rect 3513 60092 3525 60095
rect 3476 60064 3525 60092
rect 3476 60052 3482 60064
rect 3513 60061 3525 60064
rect 3559 60061 3571 60095
rect 3513 60055 3571 60061
rect 3694 60052 3700 60104
rect 3752 60052 3758 60104
rect 9398 60092 9404 60104
rect 9359 60064 9404 60092
rect 9398 60052 9404 60064
rect 9456 60052 9462 60104
rect 11517 60095 11575 60101
rect 11517 60061 11529 60095
rect 11563 60092 11575 60095
rect 11698 60092 11704 60104
rect 11563 60064 11704 60092
rect 11563 60061 11575 60064
rect 11517 60055 11575 60061
rect 11698 60052 11704 60064
rect 11756 60052 11762 60104
rect 6178 60024 6184 60036
rect 6139 59996 6184 60024
rect 6178 59984 6184 59996
rect 6236 59984 6242 60036
rect 12710 59984 12716 60036
rect 12768 60024 12774 60036
rect 12820 60024 12848 60123
rect 13170 60120 13176 60172
rect 13228 60160 13234 60172
rect 13228 60132 13273 60160
rect 13228 60120 13234 60132
rect 12986 60092 12992 60104
rect 12947 60064 12992 60092
rect 12986 60052 12992 60064
rect 13044 60052 13050 60104
rect 13998 60024 14004 60036
rect 12768 59996 14004 60024
rect 12768 59984 12774 59996
rect 13998 59984 14004 59996
rect 14056 59984 14062 60036
rect 1673 59959 1731 59965
rect 1673 59925 1685 59959
rect 1719 59956 1731 59959
rect 1762 59956 1768 59968
rect 1719 59928 1768 59956
rect 1719 59925 1731 59928
rect 1673 59919 1731 59925
rect 1762 59916 1768 59928
rect 1820 59956 1826 59968
rect 1946 59956 1952 59968
rect 1820 59928 1952 59956
rect 1820 59916 1826 59928
rect 1946 59916 1952 59928
rect 2004 59916 2010 59968
rect 2593 59959 2651 59965
rect 2593 59925 2605 59959
rect 2639 59956 2651 59959
rect 2682 59956 2688 59968
rect 2639 59928 2688 59956
rect 2639 59925 2651 59928
rect 2593 59919 2651 59925
rect 2682 59916 2688 59928
rect 2740 59916 2746 59968
rect 8294 59956 8300 59968
rect 8255 59928 8300 59956
rect 8294 59916 8300 59928
rect 8352 59956 8358 59968
rect 8570 59956 8576 59968
rect 8352 59928 8576 59956
rect 8352 59916 8358 59928
rect 8570 59916 8576 59928
rect 8628 59916 8634 59968
rect 10594 59956 10600 59968
rect 10555 59928 10600 59956
rect 10594 59916 10600 59928
rect 10652 59916 10658 59968
rect 11514 59916 11520 59968
rect 11572 59956 11578 59968
rect 14826 59956 14832 59968
rect 11572 59928 14832 59956
rect 11572 59916 11578 59928
rect 14826 59916 14832 59928
rect 14884 59916 14890 59968
rect 1104 59866 18860 59888
rect 1104 59814 4315 59866
rect 4367 59814 4379 59866
rect 4431 59814 4443 59866
rect 4495 59814 4507 59866
rect 4559 59814 10982 59866
rect 11034 59814 11046 59866
rect 11098 59814 11110 59866
rect 11162 59814 11174 59866
rect 11226 59814 17648 59866
rect 17700 59814 17712 59866
rect 17764 59814 17776 59866
rect 17828 59814 17840 59866
rect 17892 59814 18860 59866
rect 1104 59792 18860 59814
rect 3694 59752 3700 59764
rect 3655 59724 3700 59752
rect 3694 59712 3700 59724
rect 3752 59712 3758 59764
rect 4798 59712 4804 59764
rect 4856 59752 4862 59764
rect 4893 59755 4951 59761
rect 4893 59752 4905 59755
rect 4856 59724 4905 59752
rect 4856 59712 4862 59724
rect 4893 59721 4905 59724
rect 4939 59721 4951 59755
rect 5626 59752 5632 59764
rect 5587 59724 5632 59752
rect 4893 59715 4951 59721
rect 5626 59712 5632 59724
rect 5684 59712 5690 59764
rect 6270 59752 6276 59764
rect 6231 59724 6276 59752
rect 6270 59712 6276 59724
rect 6328 59712 6334 59764
rect 6730 59712 6736 59764
rect 6788 59752 6794 59764
rect 6825 59755 6883 59761
rect 6825 59752 6837 59755
rect 6788 59724 6837 59752
rect 6788 59712 6794 59724
rect 6825 59721 6837 59724
rect 6871 59721 6883 59755
rect 6825 59715 6883 59721
rect 1486 59644 1492 59696
rect 1544 59684 1550 59696
rect 1673 59687 1731 59693
rect 1673 59684 1685 59687
rect 1544 59656 1685 59684
rect 1544 59644 1550 59656
rect 1673 59653 1685 59656
rect 1719 59684 1731 59687
rect 2317 59687 2375 59693
rect 2317 59684 2329 59687
rect 1719 59656 2329 59684
rect 1719 59653 1731 59656
rect 1673 59647 1731 59653
rect 2317 59653 2329 59656
rect 2363 59653 2375 59687
rect 5644 59684 5672 59712
rect 6178 59684 6184 59696
rect 5644 59656 6184 59684
rect 2317 59647 2375 59653
rect 6178 59644 6184 59656
rect 6236 59644 6242 59696
rect 6840 59684 6868 59715
rect 9030 59712 9036 59764
rect 9088 59752 9094 59764
rect 9401 59755 9459 59761
rect 9401 59752 9413 59755
rect 9088 59724 9413 59752
rect 9088 59712 9094 59724
rect 9401 59721 9413 59724
rect 9447 59721 9459 59755
rect 9401 59715 9459 59721
rect 6840 59656 7512 59684
rect 6454 59616 6460 59628
rect 5092 59588 6460 59616
rect 2501 59551 2559 59557
rect 2501 59517 2513 59551
rect 2547 59548 2559 59551
rect 2682 59548 2688 59560
rect 2547 59520 2688 59548
rect 2547 59517 2559 59520
rect 2501 59511 2559 59517
rect 2682 59508 2688 59520
rect 2740 59508 2746 59560
rect 5092 59557 5120 59588
rect 6454 59576 6460 59588
rect 6512 59576 6518 59628
rect 6914 59576 6920 59628
rect 6972 59616 6978 59628
rect 7101 59619 7159 59625
rect 7101 59616 7113 59619
rect 6972 59588 7113 59616
rect 6972 59576 6978 59588
rect 7101 59585 7113 59588
rect 7147 59585 7159 59619
rect 7101 59579 7159 59585
rect 2869 59551 2927 59557
rect 2869 59517 2881 59551
rect 2915 59517 2927 59551
rect 2869 59511 2927 59517
rect 4433 59551 4491 59557
rect 4433 59517 4445 59551
rect 4479 59548 4491 59551
rect 5077 59551 5135 59557
rect 5077 59548 5089 59551
rect 4479 59520 5089 59548
rect 4479 59517 4491 59520
rect 4433 59511 4491 59517
rect 5077 59517 5089 59520
rect 5123 59517 5135 59551
rect 5077 59511 5135 59517
rect 5261 59551 5319 59557
rect 5261 59517 5273 59551
rect 5307 59548 5319 59551
rect 5810 59548 5816 59560
rect 5307 59520 5816 59548
rect 5307 59517 5319 59520
rect 5261 59511 5319 59517
rect 2884 59424 2912 59511
rect 2133 59415 2191 59421
rect 2133 59381 2145 59415
rect 2179 59412 2191 59415
rect 2866 59412 2872 59424
rect 2179 59384 2872 59412
rect 2179 59381 2191 59384
rect 2133 59375 2191 59381
rect 2866 59372 2872 59384
rect 2924 59372 2930 59424
rect 3329 59415 3387 59421
rect 3329 59381 3341 59415
rect 3375 59412 3387 59415
rect 3418 59412 3424 59424
rect 3375 59384 3424 59412
rect 3375 59381 3387 59384
rect 3329 59375 3387 59381
rect 3418 59372 3424 59384
rect 3476 59372 3482 59424
rect 4801 59415 4859 59421
rect 4801 59381 4813 59415
rect 4847 59412 4859 59415
rect 5276 59412 5304 59511
rect 5810 59508 5816 59520
rect 5868 59548 5874 59560
rect 5994 59548 6000 59560
rect 5868 59520 6000 59548
rect 5868 59508 5874 59520
rect 5994 59508 6000 59520
rect 6052 59508 6058 59560
rect 7282 59548 7288 59560
rect 7243 59520 7288 59548
rect 7282 59508 7288 59520
rect 7340 59508 7346 59560
rect 7377 59551 7435 59557
rect 7377 59517 7389 59551
rect 7423 59517 7435 59551
rect 7484 59548 7512 59656
rect 7745 59551 7803 59557
rect 7745 59548 7757 59551
rect 7484 59520 7757 59548
rect 7377 59511 7435 59517
rect 7745 59517 7757 59520
rect 7791 59517 7803 59551
rect 9416 59548 9444 59715
rect 10594 59712 10600 59764
rect 10652 59752 10658 59764
rect 12161 59755 12219 59761
rect 10652 59724 11008 59752
rect 10652 59712 10658 59724
rect 10045 59619 10103 59625
rect 10045 59585 10057 59619
rect 10091 59616 10103 59619
rect 10778 59616 10784 59628
rect 10091 59588 10640 59616
rect 10739 59588 10784 59616
rect 10091 59585 10103 59588
rect 10045 59579 10103 59585
rect 10137 59551 10195 59557
rect 10137 59548 10149 59551
rect 9416 59520 10149 59548
rect 7745 59511 7803 59517
rect 10137 59517 10149 59520
rect 10183 59548 10195 59551
rect 10410 59548 10416 59560
rect 10183 59520 10416 59548
rect 10183 59517 10195 59520
rect 10137 59511 10195 59517
rect 7190 59440 7196 59492
rect 7248 59480 7254 59492
rect 7392 59480 7420 59511
rect 10410 59508 10416 59520
rect 10468 59508 10474 59560
rect 10612 59548 10640 59588
rect 10778 59576 10784 59588
rect 10836 59576 10842 59628
rect 10686 59548 10692 59560
rect 10612 59520 10692 59548
rect 10686 59508 10692 59520
rect 10744 59508 10750 59560
rect 10873 59551 10931 59557
rect 10873 59517 10885 59551
rect 10919 59517 10931 59551
rect 10873 59511 10931 59517
rect 7248 59452 7420 59480
rect 7248 59440 7254 59452
rect 8478 59440 8484 59492
rect 8536 59480 8542 59492
rect 8938 59480 8944 59492
rect 8536 59452 8944 59480
rect 8536 59440 8542 59452
rect 8938 59440 8944 59452
rect 8996 59480 9002 59492
rect 9033 59483 9091 59489
rect 9033 59480 9045 59483
rect 8996 59452 9045 59480
rect 8996 59440 9002 59452
rect 9033 59449 9045 59452
rect 9079 59449 9091 59483
rect 9033 59443 9091 59449
rect 9766 59440 9772 59492
rect 9824 59480 9830 59492
rect 10888 59480 10916 59511
rect 9824 59452 10916 59480
rect 9824 59440 9830 59452
rect 8662 59412 8668 59424
rect 4847 59384 5304 59412
rect 8623 59384 8668 59412
rect 4847 59381 4859 59384
rect 4801 59375 4859 59381
rect 8662 59372 8668 59384
rect 8720 59372 8726 59424
rect 10686 59372 10692 59424
rect 10744 59412 10750 59424
rect 10980 59412 11008 59724
rect 12161 59721 12173 59755
rect 12207 59752 12219 59755
rect 13170 59752 13176 59764
rect 12207 59724 13176 59752
rect 12207 59721 12219 59724
rect 12161 59715 12219 59721
rect 13170 59712 13176 59724
rect 13228 59712 13234 59764
rect 13446 59752 13452 59764
rect 13407 59724 13452 59752
rect 13446 59712 13452 59724
rect 13504 59712 13510 59764
rect 13998 59752 14004 59764
rect 13959 59724 14004 59752
rect 13998 59712 14004 59724
rect 14056 59712 14062 59764
rect 14090 59712 14096 59764
rect 14148 59752 14154 59764
rect 17497 59755 17555 59761
rect 17497 59752 17509 59755
rect 14148 59724 17509 59752
rect 14148 59712 14154 59724
rect 17497 59721 17509 59724
rect 17543 59721 17555 59755
rect 17497 59715 17555 59721
rect 11793 59687 11851 59693
rect 11793 59653 11805 59687
rect 11839 59684 11851 59687
rect 13538 59684 13544 59696
rect 11839 59656 13544 59684
rect 11839 59653 11851 59656
rect 11793 59647 11851 59653
rect 13538 59644 13544 59656
rect 13596 59644 13602 59696
rect 14369 59619 14427 59625
rect 14369 59616 14381 59619
rect 12544 59588 14381 59616
rect 12544 59560 12572 59588
rect 14369 59585 14381 59588
rect 14415 59585 14427 59619
rect 14369 59579 14427 59585
rect 16025 59619 16083 59625
rect 16025 59585 16037 59619
rect 16071 59616 16083 59619
rect 16071 59588 16436 59616
rect 16071 59585 16083 59588
rect 16025 59579 16083 59585
rect 16408 59560 16436 59588
rect 12526 59548 12532 59560
rect 12487 59520 12532 59548
rect 12526 59508 12532 59520
rect 12584 59508 12590 59560
rect 12710 59548 12716 59560
rect 12671 59520 12716 59548
rect 12710 59508 12716 59520
rect 12768 59508 12774 59560
rect 12986 59548 12992 59560
rect 12947 59520 12992 59548
rect 12986 59508 12992 59520
rect 13044 59508 13050 59560
rect 13538 59548 13544 59560
rect 13499 59520 13544 59548
rect 13538 59508 13544 59520
rect 13596 59508 13602 59560
rect 15930 59508 15936 59560
rect 15988 59548 15994 59560
rect 16117 59551 16175 59557
rect 16117 59548 16129 59551
rect 15988 59520 16129 59548
rect 15988 59508 15994 59520
rect 16117 59517 16129 59520
rect 16163 59517 16175 59551
rect 16390 59548 16396 59560
rect 16351 59520 16396 59548
rect 16117 59511 16175 59517
rect 16390 59508 16396 59520
rect 16448 59508 16454 59560
rect 12342 59440 12348 59492
rect 12400 59480 12406 59492
rect 13004 59480 13032 59508
rect 12400 59452 13032 59480
rect 12400 59440 12406 59452
rect 10744 59384 11008 59412
rect 10744 59372 10750 59384
rect 13262 59372 13268 59424
rect 13320 59412 13326 59424
rect 13446 59412 13452 59424
rect 13320 59384 13452 59412
rect 13320 59372 13326 59384
rect 13446 59372 13452 59384
rect 13504 59372 13510 59424
rect 1104 59322 18860 59344
rect 1104 59270 7648 59322
rect 7700 59270 7712 59322
rect 7764 59270 7776 59322
rect 7828 59270 7840 59322
rect 7892 59270 14315 59322
rect 14367 59270 14379 59322
rect 14431 59270 14443 59322
rect 14495 59270 14507 59322
rect 14559 59270 18860 59322
rect 1104 59248 18860 59270
rect 2332 59180 2820 59208
rect 1578 59140 1584 59152
rect 1539 59112 1584 59140
rect 1578 59100 1584 59112
rect 1636 59100 1642 59152
rect 1762 59100 1768 59152
rect 1820 59140 1826 59152
rect 2332 59140 2360 59180
rect 1820 59112 2360 59140
rect 1820 59100 1826 59112
rect 1486 59072 1492 59084
rect 1447 59044 1492 59072
rect 1486 59032 1492 59044
rect 1544 59032 1550 59084
rect 2332 59081 2360 59112
rect 2317 59075 2375 59081
rect 2317 59041 2329 59075
rect 2363 59041 2375 59075
rect 2792 59072 2820 59180
rect 2866 59168 2872 59220
rect 2924 59208 2930 59220
rect 3513 59211 3571 59217
rect 3513 59208 3525 59211
rect 2924 59180 3525 59208
rect 2924 59168 2930 59180
rect 3513 59177 3525 59180
rect 3559 59177 3571 59211
rect 3513 59171 3571 59177
rect 3881 59211 3939 59217
rect 3881 59177 3893 59211
rect 3927 59208 3939 59211
rect 4798 59208 4804 59220
rect 3927 59180 4804 59208
rect 3927 59177 3939 59180
rect 3881 59171 3939 59177
rect 4798 59168 4804 59180
rect 4856 59168 4862 59220
rect 10321 59211 10379 59217
rect 10321 59177 10333 59211
rect 10367 59208 10379 59211
rect 10594 59208 10600 59220
rect 10367 59180 10600 59208
rect 10367 59177 10379 59180
rect 10321 59171 10379 59177
rect 10594 59168 10600 59180
rect 10652 59168 10658 59220
rect 10870 59208 10876 59220
rect 10831 59180 10876 59208
rect 10870 59168 10876 59180
rect 10928 59168 10934 59220
rect 11425 59211 11483 59217
rect 11425 59177 11437 59211
rect 11471 59208 11483 59211
rect 11606 59208 11612 59220
rect 11471 59180 11612 59208
rect 11471 59177 11483 59180
rect 11425 59171 11483 59177
rect 11606 59168 11612 59180
rect 11664 59168 11670 59220
rect 12253 59211 12311 59217
rect 12253 59177 12265 59211
rect 12299 59208 12311 59211
rect 12342 59208 12348 59220
rect 12299 59180 12348 59208
rect 12299 59177 12311 59180
rect 12253 59171 12311 59177
rect 12342 59168 12348 59180
rect 12400 59168 12406 59220
rect 13173 59211 13231 59217
rect 13173 59177 13185 59211
rect 13219 59208 13231 59211
rect 13814 59208 13820 59220
rect 13219 59180 13820 59208
rect 13219 59177 13231 59180
rect 13173 59171 13231 59177
rect 5442 59100 5448 59152
rect 5500 59140 5506 59152
rect 8386 59140 8392 59152
rect 5500 59112 5856 59140
rect 5500 59100 5506 59112
rect 3329 59075 3387 59081
rect 2792 59044 2912 59072
rect 2317 59035 2375 59041
rect 1670 58964 1676 59016
rect 1728 59004 1734 59016
rect 2222 59004 2228 59016
rect 1728 58976 2228 59004
rect 1728 58964 1734 58976
rect 2222 58964 2228 58976
rect 2280 59004 2286 59016
rect 2409 59007 2467 59013
rect 2409 59004 2421 59007
rect 2280 58976 2421 59004
rect 2280 58964 2286 58976
rect 2409 58973 2421 58976
rect 2455 58973 2467 59007
rect 2409 58967 2467 58973
rect 2884 58945 2912 59044
rect 3329 59041 3341 59075
rect 3375 59072 3387 59075
rect 4614 59072 4620 59084
rect 3375 59044 4620 59072
rect 3375 59041 3387 59044
rect 3329 59035 3387 59041
rect 4614 59032 4620 59044
rect 4672 59032 4678 59084
rect 4982 59032 4988 59084
rect 5040 59072 5046 59084
rect 5353 59075 5411 59081
rect 5353 59072 5365 59075
rect 5040 59044 5365 59072
rect 5040 59032 5046 59044
rect 5353 59041 5365 59044
rect 5399 59041 5411 59075
rect 5718 59072 5724 59084
rect 5679 59044 5724 59072
rect 5353 59035 5411 59041
rect 5718 59032 5724 59044
rect 5776 59032 5782 59084
rect 5828 59081 5856 59112
rect 7944 59112 8392 59140
rect 5813 59075 5871 59081
rect 5813 59041 5825 59075
rect 5859 59072 5871 59075
rect 6822 59072 6828 59084
rect 5859 59044 6828 59072
rect 5859 59041 5871 59044
rect 5813 59035 5871 59041
rect 6822 59032 6828 59044
rect 6880 59032 6886 59084
rect 7374 59032 7380 59084
rect 7432 59072 7438 59084
rect 7944 59081 7972 59112
rect 8386 59100 8392 59112
rect 8444 59100 8450 59152
rect 11885 59143 11943 59149
rect 11885 59109 11897 59143
rect 11931 59140 11943 59143
rect 12710 59140 12716 59152
rect 11931 59112 12716 59140
rect 11931 59109 11943 59112
rect 11885 59103 11943 59109
rect 12710 59100 12716 59112
rect 12768 59140 12774 59152
rect 13262 59140 13268 59152
rect 12768 59112 13268 59140
rect 12768 59100 12774 59112
rect 13262 59100 13268 59112
rect 13320 59100 13326 59152
rect 7469 59075 7527 59081
rect 7469 59072 7481 59075
rect 7432 59044 7481 59072
rect 7432 59032 7438 59044
rect 7469 59041 7481 59044
rect 7515 59072 7527 59075
rect 7929 59075 7987 59081
rect 7929 59072 7941 59075
rect 7515 59044 7941 59072
rect 7515 59041 7527 59044
rect 7469 59035 7527 59041
rect 7929 59041 7941 59044
rect 7975 59041 7987 59075
rect 8478 59072 8484 59084
rect 8439 59044 8484 59072
rect 7929 59035 7987 59041
rect 8478 59032 8484 59044
rect 8536 59032 8542 59084
rect 9033 59075 9091 59081
rect 9033 59041 9045 59075
rect 9079 59041 9091 59075
rect 9033 59035 9091 59041
rect 4801 59007 4859 59013
rect 4801 58973 4813 59007
rect 4847 59004 4859 59007
rect 5736 59004 5764 59032
rect 8662 59004 8668 59016
rect 4847 58976 5764 59004
rect 8623 58976 8668 59004
rect 4847 58973 4859 58976
rect 4801 58967 4859 58973
rect 8662 58964 8668 58976
rect 8720 58964 8726 59016
rect 9048 59004 9076 59035
rect 9122 59032 9128 59084
rect 9180 59072 9186 59084
rect 9217 59075 9275 59081
rect 9217 59072 9229 59075
rect 9180 59044 9229 59072
rect 9180 59032 9186 59044
rect 9217 59041 9229 59044
rect 9263 59041 9275 59075
rect 9766 59072 9772 59084
rect 9727 59044 9772 59072
rect 9217 59035 9275 59041
rect 9766 59032 9772 59044
rect 9824 59032 9830 59084
rect 11241 59075 11299 59081
rect 11241 59041 11253 59075
rect 11287 59072 11299 59075
rect 11606 59072 11612 59084
rect 11287 59044 11612 59072
rect 11287 59041 11299 59044
rect 11241 59035 11299 59041
rect 11606 59032 11612 59044
rect 11664 59072 11670 59084
rect 12158 59072 12164 59084
rect 11664 59044 12164 59072
rect 11664 59032 11670 59044
rect 12158 59032 12164 59044
rect 12216 59032 12222 59084
rect 13357 59075 13415 59081
rect 13357 59041 13369 59075
rect 13403 59041 13415 59075
rect 13357 59035 13415 59041
rect 9490 59004 9496 59016
rect 9048 58976 9496 59004
rect 9490 58964 9496 58976
rect 9548 58964 9554 59016
rect 2869 58939 2927 58945
rect 2869 58905 2881 58939
rect 2915 58936 2927 58939
rect 3237 58939 3295 58945
rect 3237 58936 3249 58939
rect 2915 58908 3249 58936
rect 2915 58905 2927 58908
rect 2869 58899 2927 58905
rect 3237 58905 3249 58908
rect 3283 58936 3295 58939
rect 4062 58936 4068 58948
rect 3283 58908 4068 58936
rect 3283 58905 3295 58908
rect 3237 58899 3295 58905
rect 4062 58896 4068 58908
rect 4120 58896 4126 58948
rect 5169 58939 5227 58945
rect 5169 58905 5181 58939
rect 5215 58936 5227 58939
rect 5994 58936 6000 58948
rect 5215 58908 6000 58936
rect 5215 58905 5227 58908
rect 5169 58899 5227 58905
rect 5994 58896 6000 58908
rect 6052 58936 6058 58948
rect 6181 58939 6239 58945
rect 6181 58936 6193 58939
rect 6052 58908 6193 58936
rect 6052 58896 6058 58908
rect 6181 58905 6193 58908
rect 6227 58905 6239 58939
rect 6181 58899 6239 58905
rect 12434 58896 12440 58948
rect 12492 58936 12498 58948
rect 13372 58936 13400 59035
rect 13464 59013 13492 59180
rect 13814 59168 13820 59180
rect 13872 59168 13878 59220
rect 13449 59007 13507 59013
rect 13449 58973 13461 59007
rect 13495 58973 13507 59007
rect 13449 58967 13507 58973
rect 13725 59007 13783 59013
rect 13725 58973 13737 59007
rect 13771 59004 13783 59007
rect 13906 59004 13912 59016
rect 13771 58976 13912 59004
rect 13771 58973 13783 58976
rect 13725 58967 13783 58973
rect 13906 58964 13912 58976
rect 13964 58964 13970 59016
rect 14826 59004 14832 59016
rect 14787 58976 14832 59004
rect 14826 58964 14832 58976
rect 14884 58964 14890 59016
rect 12492 58908 13400 58936
rect 12492 58896 12498 58908
rect 6638 58868 6644 58880
rect 6599 58840 6644 58868
rect 6638 58828 6644 58840
rect 6696 58828 6702 58880
rect 7101 58871 7159 58877
rect 7101 58837 7113 58871
rect 7147 58868 7159 58871
rect 7190 58868 7196 58880
rect 7147 58840 7196 58868
rect 7147 58837 7159 58840
rect 7101 58831 7159 58837
rect 7190 58828 7196 58840
rect 7248 58868 7254 58880
rect 7653 58871 7711 58877
rect 7653 58868 7665 58871
rect 7248 58840 7665 58868
rect 7248 58828 7254 58840
rect 7653 58837 7665 58840
rect 7699 58837 7711 58871
rect 8294 58868 8300 58880
rect 8255 58840 8300 58868
rect 7653 58831 7711 58837
rect 8294 58828 8300 58840
rect 8352 58828 8358 58880
rect 12802 58868 12808 58880
rect 12763 58840 12808 58868
rect 12802 58828 12808 58840
rect 12860 58828 12866 58880
rect 13372 58868 13400 58908
rect 14642 58868 14648 58880
rect 13372 58840 14648 58868
rect 14642 58828 14648 58840
rect 14700 58828 14706 58880
rect 15930 58828 15936 58880
rect 15988 58868 15994 58880
rect 16117 58871 16175 58877
rect 16117 58868 16129 58871
rect 15988 58840 16129 58868
rect 15988 58828 15994 58840
rect 16117 58837 16129 58840
rect 16163 58837 16175 58871
rect 16117 58831 16175 58837
rect 1104 58778 18860 58800
rect 1104 58726 4315 58778
rect 4367 58726 4379 58778
rect 4431 58726 4443 58778
rect 4495 58726 4507 58778
rect 4559 58726 10982 58778
rect 11034 58726 11046 58778
rect 11098 58726 11110 58778
rect 11162 58726 11174 58778
rect 11226 58726 17648 58778
rect 17700 58726 17712 58778
rect 17764 58726 17776 58778
rect 17828 58726 17840 58778
rect 17892 58726 18860 58778
rect 1104 58704 18860 58726
rect 2774 58624 2780 58676
rect 2832 58664 2838 58676
rect 2869 58667 2927 58673
rect 2869 58664 2881 58667
rect 2832 58636 2881 58664
rect 2832 58624 2838 58636
rect 2869 58633 2881 58636
rect 2915 58633 2927 58667
rect 4614 58664 4620 58676
rect 4575 58636 4620 58664
rect 2869 58627 2927 58633
rect 4614 58624 4620 58636
rect 4672 58624 4678 58676
rect 4982 58664 4988 58676
rect 4943 58636 4988 58664
rect 4982 58624 4988 58636
rect 5040 58624 5046 58676
rect 7653 58667 7711 58673
rect 7653 58633 7665 58667
rect 7699 58664 7711 58667
rect 8018 58664 8024 58676
rect 7699 58636 8024 58664
rect 7699 58633 7711 58636
rect 7653 58627 7711 58633
rect 8018 58624 8024 58636
rect 8076 58624 8082 58676
rect 14642 58664 14648 58676
rect 14603 58636 14648 58664
rect 14642 58624 14648 58636
rect 14700 58624 14706 58676
rect 4062 58556 4068 58608
rect 4120 58596 4126 58608
rect 5537 58599 5595 58605
rect 5537 58596 5549 58599
rect 4120 58568 5549 58596
rect 4120 58556 4126 58568
rect 5537 58565 5549 58568
rect 5583 58565 5595 58599
rect 5537 58559 5595 58565
rect 7285 58599 7343 58605
rect 7285 58565 7297 58599
rect 7331 58596 7343 58599
rect 9674 58596 9680 58608
rect 7331 58568 9680 58596
rect 7331 58565 7343 58568
rect 7285 58559 7343 58565
rect 1210 58488 1216 58540
rect 1268 58528 1274 58540
rect 1489 58531 1547 58537
rect 1489 58528 1501 58531
rect 1268 58500 1501 58528
rect 1268 58488 1274 58500
rect 1489 58497 1501 58500
rect 1535 58497 1547 58531
rect 1762 58528 1768 58540
rect 1723 58500 1768 58528
rect 1489 58491 1547 58497
rect 1504 58324 1532 58491
rect 1762 58488 1768 58500
rect 1820 58488 1826 58540
rect 6822 58528 6828 58540
rect 5736 58500 6828 58528
rect 3513 58463 3571 58469
rect 3513 58429 3525 58463
rect 3559 58460 3571 58463
rect 4065 58463 4123 58469
rect 4065 58460 4077 58463
rect 3559 58432 4077 58460
rect 3559 58429 3571 58432
rect 3513 58423 3571 58429
rect 4065 58429 4077 58432
rect 4111 58460 4123 58463
rect 4614 58460 4620 58472
rect 4111 58432 4620 58460
rect 4111 58429 4123 58432
rect 4065 58423 4123 58429
rect 4614 58420 4620 58432
rect 4672 58420 4678 58472
rect 5736 58469 5764 58500
rect 6822 58488 6828 58500
rect 6880 58488 6886 58540
rect 8680 58537 8708 58568
rect 9674 58556 9680 58568
rect 9732 58556 9738 58608
rect 10410 58596 10416 58608
rect 10371 58568 10416 58596
rect 10410 58556 10416 58568
rect 10468 58556 10474 58608
rect 11238 58556 11244 58608
rect 11296 58596 11302 58608
rect 11422 58596 11428 58608
rect 11296 58568 11428 58596
rect 11296 58556 11302 58568
rect 11422 58556 11428 58568
rect 11480 58556 11486 58608
rect 8665 58531 8723 58537
rect 8665 58497 8677 58531
rect 8711 58497 8723 58531
rect 8665 58491 8723 58497
rect 11793 58531 11851 58537
rect 11793 58497 11805 58531
rect 11839 58528 11851 58531
rect 12158 58528 12164 58540
rect 11839 58500 12164 58528
rect 11839 58497 11851 58500
rect 11793 58491 11851 58497
rect 12158 58488 12164 58500
rect 12216 58528 12222 58540
rect 12713 58531 12771 58537
rect 12713 58528 12725 58531
rect 12216 58500 12725 58528
rect 12216 58488 12222 58500
rect 12713 58497 12725 58500
rect 12759 58497 12771 58531
rect 12713 58491 12771 58497
rect 5721 58463 5779 58469
rect 5721 58429 5733 58463
rect 5767 58429 5779 58463
rect 5994 58460 6000 58472
rect 5955 58432 6000 58460
rect 5721 58423 5779 58429
rect 3881 58395 3939 58401
rect 3881 58361 3893 58395
rect 3927 58392 3939 58395
rect 5736 58392 5764 58423
rect 5994 58420 6000 58432
rect 6052 58420 6058 58472
rect 6362 58460 6368 58472
rect 6323 58432 6368 58460
rect 6362 58420 6368 58432
rect 6420 58420 6426 58472
rect 6641 58463 6699 58469
rect 6641 58429 6653 58463
rect 6687 58429 6699 58463
rect 6641 58423 6699 58429
rect 8205 58463 8263 58469
rect 8205 58429 8217 58463
rect 8251 58460 8263 58463
rect 8294 58460 8300 58472
rect 8251 58432 8300 58460
rect 8251 58429 8263 58432
rect 8205 58423 8263 58429
rect 3927 58364 5764 58392
rect 3927 58361 3939 58364
rect 3881 58355 3939 58361
rect 1762 58324 1768 58336
rect 1504 58296 1768 58324
rect 1762 58284 1768 58296
rect 1820 58284 1826 58336
rect 3050 58284 3056 58336
rect 3108 58324 3114 58336
rect 3418 58324 3424 58336
rect 3108 58296 3424 58324
rect 3108 58284 3114 58296
rect 3418 58284 3424 58296
rect 3476 58324 3482 58336
rect 4249 58327 4307 58333
rect 4249 58324 4261 58327
rect 3476 58296 4261 58324
rect 3476 58284 3482 58296
rect 4249 58293 4261 58296
rect 4295 58293 4307 58327
rect 4249 58287 4307 58293
rect 5074 58284 5080 58336
rect 5132 58324 5138 58336
rect 5353 58327 5411 58333
rect 5353 58324 5365 58327
rect 5132 58296 5365 58324
rect 5132 58284 5138 58296
rect 5353 58293 5365 58296
rect 5399 58324 5411 58327
rect 6656 58324 6684 58423
rect 8294 58420 8300 58432
rect 8352 58420 8358 58472
rect 8570 58460 8576 58472
rect 8531 58432 8576 58460
rect 8570 58420 8576 58432
rect 8628 58420 8634 58472
rect 9674 58460 9680 58472
rect 9635 58432 9680 58460
rect 9674 58420 9680 58432
rect 9732 58420 9738 58472
rect 10137 58463 10195 58469
rect 10137 58429 10149 58463
rect 10183 58429 10195 58463
rect 10137 58423 10195 58429
rect 10505 58463 10563 58469
rect 10505 58429 10517 58463
rect 10551 58460 10563 58463
rect 10594 58460 10600 58472
rect 10551 58432 10600 58460
rect 10551 58429 10563 58432
rect 10505 58423 10563 58429
rect 6914 58352 6920 58404
rect 6972 58392 6978 58404
rect 7745 58395 7803 58401
rect 7745 58392 7757 58395
rect 6972 58364 7757 58392
rect 6972 58352 6978 58364
rect 7745 58361 7757 58364
rect 7791 58361 7803 58395
rect 10152 58392 10180 58423
rect 10594 58420 10600 58432
rect 10652 58420 10658 58472
rect 12434 58460 12440 58472
rect 12084 58432 12440 58460
rect 7745 58355 7803 58361
rect 9508 58364 10180 58392
rect 9508 58336 9536 58364
rect 12084 58336 12112 58432
rect 12434 58420 12440 58432
rect 12492 58460 12498 58472
rect 12492 58432 12537 58460
rect 12492 58420 12498 58432
rect 12802 58420 12808 58472
rect 12860 58460 12866 58472
rect 12989 58463 13047 58469
rect 12989 58460 13001 58463
rect 12860 58432 13001 58460
rect 12860 58420 12866 58432
rect 12989 58429 13001 58432
rect 13035 58460 13047 58463
rect 13630 58460 13636 58472
rect 13035 58432 13636 58460
rect 13035 58429 13047 58432
rect 12989 58423 13047 58429
rect 13630 58420 13636 58432
rect 13688 58420 13694 58472
rect 5399 58296 6684 58324
rect 5399 58293 5411 58296
rect 5353 58287 5411 58293
rect 8018 58284 8024 58336
rect 8076 58324 8082 58336
rect 8202 58324 8208 58336
rect 8076 58296 8208 58324
rect 8076 58284 8082 58296
rect 8202 58284 8208 58296
rect 8260 58284 8266 58336
rect 9122 58324 9128 58336
rect 9083 58296 9128 58324
rect 9122 58284 9128 58296
rect 9180 58284 9186 58336
rect 9490 58324 9496 58336
rect 9451 58296 9496 58324
rect 9490 58284 9496 58296
rect 9548 58284 9554 58336
rect 11333 58327 11391 58333
rect 11333 58293 11345 58327
rect 11379 58324 11391 58327
rect 11422 58324 11428 58336
rect 11379 58296 11428 58324
rect 11379 58293 11391 58296
rect 11333 58287 11391 58293
rect 11422 58284 11428 58296
rect 11480 58324 11486 58336
rect 11606 58324 11612 58336
rect 11480 58296 11612 58324
rect 11480 58284 11486 58296
rect 11606 58284 11612 58296
rect 11664 58284 11670 58336
rect 12066 58324 12072 58336
rect 12027 58296 12072 58324
rect 12066 58284 12072 58296
rect 12124 58284 12130 58336
rect 12250 58324 12256 58336
rect 12211 58296 12256 58324
rect 12250 58284 12256 58296
rect 12308 58284 12314 58336
rect 14090 58324 14096 58336
rect 14051 58296 14096 58324
rect 14090 58284 14096 58296
rect 14148 58284 14154 58336
rect 1104 58234 18860 58256
rect 1104 58182 7648 58234
rect 7700 58182 7712 58234
rect 7764 58182 7776 58234
rect 7828 58182 7840 58234
rect 7892 58182 14315 58234
rect 14367 58182 14379 58234
rect 14431 58182 14443 58234
rect 14495 58182 14507 58234
rect 14559 58182 18860 58234
rect 1104 58160 18860 58182
rect 1302 58080 1308 58132
rect 1360 58120 1366 58132
rect 5537 58123 5595 58129
rect 1360 58092 4016 58120
rect 1360 58080 1366 58092
rect 1394 58012 1400 58064
rect 1452 58052 1458 58064
rect 3988 58061 4016 58092
rect 5537 58089 5549 58123
rect 5583 58120 5595 58123
rect 6270 58120 6276 58132
rect 5583 58092 6276 58120
rect 5583 58089 5595 58092
rect 5537 58083 5595 58089
rect 6270 58080 6276 58092
rect 6328 58080 6334 58132
rect 6454 58120 6460 58132
rect 6415 58092 6460 58120
rect 6454 58080 6460 58092
rect 6512 58080 6518 58132
rect 6730 58080 6736 58132
rect 6788 58120 6794 58132
rect 11146 58120 11152 58132
rect 6788 58092 7972 58120
rect 11107 58092 11152 58120
rect 6788 58080 6794 58092
rect 7944 58064 7972 58092
rect 11146 58080 11152 58092
rect 11204 58080 11210 58132
rect 12250 58080 12256 58132
rect 12308 58120 12314 58132
rect 15930 58120 15936 58132
rect 12308 58092 15936 58120
rect 12308 58080 12314 58092
rect 15930 58080 15936 58092
rect 15988 58080 15994 58132
rect 1581 58055 1639 58061
rect 1581 58052 1593 58055
rect 1452 58024 1593 58052
rect 1452 58012 1458 58024
rect 1581 58021 1593 58024
rect 1627 58021 1639 58055
rect 1581 58015 1639 58021
rect 3973 58055 4031 58061
rect 3973 58021 3985 58055
rect 4019 58021 4031 58055
rect 3973 58015 4031 58021
rect 4448 58024 5672 58052
rect 2317 57987 2375 57993
rect 2317 57953 2329 57987
rect 2363 57984 2375 57987
rect 2363 57956 2728 57984
rect 2363 57953 2375 57956
rect 2317 57947 2375 57953
rect 1486 57916 1492 57928
rect 1447 57888 1492 57916
rect 1486 57876 1492 57888
rect 1544 57876 1550 57928
rect 2222 57876 2228 57928
rect 2280 57916 2286 57928
rect 2409 57919 2467 57925
rect 2409 57916 2421 57919
rect 2280 57888 2421 57916
rect 2280 57876 2286 57888
rect 2409 57885 2421 57888
rect 2455 57885 2467 57919
rect 2409 57879 2467 57885
rect 1394 57808 1400 57860
rect 1452 57848 1458 57860
rect 1946 57848 1952 57860
rect 1452 57820 1952 57848
rect 1452 57808 1458 57820
rect 1946 57808 1952 57820
rect 2004 57808 2010 57860
rect 2700 57848 2728 57956
rect 2869 57919 2927 57925
rect 2869 57885 2881 57919
rect 2915 57916 2927 57919
rect 3694 57916 3700 57928
rect 2915 57888 3700 57916
rect 2915 57885 2927 57888
rect 2869 57879 2927 57885
rect 3694 57876 3700 57888
rect 3752 57876 3758 57928
rect 3881 57919 3939 57925
rect 3881 57885 3893 57919
rect 3927 57916 3939 57919
rect 4448 57916 4476 58024
rect 4798 57984 4804 57996
rect 4759 57956 4804 57984
rect 4798 57944 4804 57956
rect 4856 57944 4862 57996
rect 5644 57984 5672 58024
rect 5718 58012 5724 58064
rect 5776 58052 5782 58064
rect 6825 58055 6883 58061
rect 6825 58052 6837 58055
rect 5776 58024 6837 58052
rect 5776 58012 5782 58024
rect 6825 58021 6837 58024
rect 6871 58021 6883 58055
rect 6825 58015 6883 58021
rect 7926 58012 7932 58064
rect 7984 58012 7990 58064
rect 8570 58012 8576 58064
rect 8628 58052 8634 58064
rect 8849 58055 8907 58061
rect 8849 58052 8861 58055
rect 8628 58024 8861 58052
rect 8628 58012 8634 58024
rect 8849 58021 8861 58024
rect 8895 58021 8907 58055
rect 8849 58015 8907 58021
rect 6454 57984 6460 57996
rect 5644 57956 6460 57984
rect 6454 57944 6460 57956
rect 6512 57984 6518 57996
rect 6641 57987 6699 57993
rect 6641 57984 6653 57987
rect 6512 57956 6653 57984
rect 6512 57944 6518 57956
rect 6641 57953 6653 57956
rect 6687 57953 6699 57987
rect 6641 57947 6699 57953
rect 7469 57987 7527 57993
rect 7469 57953 7481 57987
rect 7515 57984 7527 57987
rect 7650 57984 7656 57996
rect 7515 57956 7656 57984
rect 7515 57953 7527 57956
rect 7469 57947 7527 57953
rect 7650 57944 7656 57956
rect 7708 57944 7714 57996
rect 7834 57984 7840 57996
rect 7795 57956 7840 57984
rect 7834 57944 7840 57956
rect 7892 57944 7898 57996
rect 9677 57987 9735 57993
rect 9677 57953 9689 57987
rect 9723 57984 9735 57987
rect 9766 57984 9772 57996
rect 9723 57956 9772 57984
rect 9723 57953 9735 57956
rect 9677 57947 9735 57953
rect 9766 57944 9772 57956
rect 9824 57944 9830 57996
rect 11057 57987 11115 57993
rect 11057 57953 11069 57987
rect 11103 57953 11115 57987
rect 12526 57984 12532 57996
rect 12487 57956 12532 57984
rect 11057 57947 11115 57953
rect 3927 57888 4476 57916
rect 4525 57919 4583 57925
rect 3927 57885 3939 57888
rect 3881 57879 3939 57885
rect 4525 57885 4537 57919
rect 4571 57916 4583 57919
rect 4614 57916 4620 57928
rect 4571 57888 4620 57916
rect 4571 57885 4583 57888
rect 4525 57879 4583 57885
rect 4614 57876 4620 57888
rect 4672 57876 4678 57928
rect 4985 57919 5043 57925
rect 4985 57885 4997 57919
rect 5031 57885 5043 57919
rect 4985 57879 5043 57885
rect 3510 57848 3516 57860
rect 2700 57820 3516 57848
rect 3510 57808 3516 57820
rect 3568 57808 3574 57860
rect 3712 57848 3740 57876
rect 5000 57848 5028 57879
rect 6178 57876 6184 57928
rect 6236 57916 6242 57928
rect 7285 57919 7343 57925
rect 7285 57916 7297 57919
rect 6236 57888 7297 57916
rect 6236 57876 6242 57888
rect 7285 57885 7297 57888
rect 7331 57885 7343 57919
rect 7285 57879 7343 57885
rect 7745 57919 7803 57925
rect 7745 57885 7757 57919
rect 7791 57916 7803 57919
rect 8386 57916 8392 57928
rect 7791 57888 8392 57916
rect 7791 57885 7803 57888
rect 7745 57879 7803 57885
rect 8386 57876 8392 57888
rect 8444 57876 8450 57928
rect 9306 57876 9312 57928
rect 9364 57916 9370 57928
rect 9401 57919 9459 57925
rect 9401 57916 9413 57919
rect 9364 57888 9413 57916
rect 9364 57876 9370 57888
rect 9401 57885 9413 57888
rect 9447 57885 9459 57919
rect 9401 57879 9459 57885
rect 9861 57919 9919 57925
rect 9861 57885 9873 57919
rect 9907 57885 9919 57919
rect 9861 57879 9919 57885
rect 3712 57820 5028 57848
rect 5905 57851 5963 57857
rect 5905 57817 5917 57851
rect 5951 57848 5963 57851
rect 6730 57848 6736 57860
rect 5951 57820 6736 57848
rect 5951 57817 5963 57820
rect 5905 57811 5963 57817
rect 6730 57808 6736 57820
rect 6788 57808 6794 57860
rect 8404 57848 8432 57876
rect 9876 57848 9904 57879
rect 10686 57876 10692 57928
rect 10744 57916 10750 57928
rect 10870 57916 10876 57928
rect 10744 57888 10876 57916
rect 10744 57876 10750 57888
rect 10870 57876 10876 57888
rect 10928 57916 10934 57928
rect 11072 57916 11100 57947
rect 12526 57944 12532 57956
rect 12584 57944 12590 57996
rect 12802 57984 12808 57996
rect 12763 57956 12808 57984
rect 12802 57944 12808 57956
rect 12860 57944 12866 57996
rect 13170 57984 13176 57996
rect 13131 57956 13176 57984
rect 13170 57944 13176 57956
rect 13228 57944 13234 57996
rect 11698 57916 11704 57928
rect 10928 57888 11100 57916
rect 11659 57888 11704 57916
rect 10928 57876 10934 57888
rect 11698 57876 11704 57888
rect 11756 57916 11762 57928
rect 12250 57916 12256 57928
rect 11756 57888 12256 57916
rect 11756 57876 11762 57888
rect 12250 57876 12256 57888
rect 12308 57876 12314 57928
rect 13538 57916 13544 57928
rect 13499 57888 13544 57916
rect 13538 57876 13544 57888
rect 13596 57876 13602 57928
rect 13814 57876 13820 57928
rect 13872 57916 13878 57928
rect 14277 57919 14335 57925
rect 14277 57916 14289 57919
rect 13872 57888 14289 57916
rect 13872 57876 13878 57888
rect 14277 57885 14289 57888
rect 14323 57885 14335 57919
rect 14277 57879 14335 57885
rect 8404 57820 9904 57848
rect 11238 57808 11244 57860
rect 11296 57848 11302 57860
rect 11606 57848 11612 57860
rect 11296 57820 11612 57848
rect 11296 57808 11302 57820
rect 11606 57808 11612 57820
rect 11664 57808 11670 57860
rect 3050 57740 3056 57792
rect 3108 57780 3114 57792
rect 3145 57783 3203 57789
rect 3145 57780 3157 57783
rect 3108 57752 3157 57780
rect 3108 57740 3114 57752
rect 3145 57749 3157 57752
rect 3191 57749 3203 57783
rect 6270 57780 6276 57792
rect 6231 57752 6276 57780
rect 3145 57743 3203 57749
rect 6270 57740 6276 57752
rect 6328 57780 6334 57792
rect 7834 57780 7840 57792
rect 6328 57752 7840 57780
rect 6328 57740 6334 57752
rect 7834 57740 7840 57752
rect 7892 57740 7898 57792
rect 8570 57780 8576 57792
rect 8531 57752 8576 57780
rect 8570 57740 8576 57752
rect 8628 57740 8634 57792
rect 9030 57740 9036 57792
rect 9088 57780 9094 57792
rect 9674 57780 9680 57792
rect 9088 57752 9680 57780
rect 9088 57740 9094 57752
rect 9674 57740 9680 57752
rect 9732 57780 9738 57792
rect 10137 57783 10195 57789
rect 10137 57780 10149 57783
rect 9732 57752 10149 57780
rect 9732 57740 9738 57752
rect 10137 57749 10149 57752
rect 10183 57749 10195 57783
rect 10137 57743 10195 57749
rect 10597 57783 10655 57789
rect 10597 57749 10609 57783
rect 10643 57780 10655 57783
rect 10686 57780 10692 57792
rect 10643 57752 10692 57780
rect 10643 57749 10655 57752
rect 10597 57743 10655 57749
rect 10686 57740 10692 57752
rect 10744 57740 10750 57792
rect 13906 57740 13912 57792
rect 13964 57780 13970 57792
rect 14001 57783 14059 57789
rect 14001 57780 14013 57783
rect 13964 57752 14013 57780
rect 13964 57740 13970 57752
rect 14001 57749 14013 57752
rect 14047 57780 14059 57783
rect 15562 57780 15568 57792
rect 14047 57752 15568 57780
rect 14047 57749 14059 57752
rect 14001 57743 14059 57749
rect 15562 57740 15568 57752
rect 15620 57740 15626 57792
rect 1104 57690 18860 57712
rect 1104 57638 4315 57690
rect 4367 57638 4379 57690
rect 4431 57638 4443 57690
rect 4495 57638 4507 57690
rect 4559 57638 10982 57690
rect 11034 57638 11046 57690
rect 11098 57638 11110 57690
rect 11162 57638 11174 57690
rect 11226 57638 17648 57690
rect 17700 57638 17712 57690
rect 17764 57638 17776 57690
rect 17828 57638 17840 57690
rect 17892 57638 18860 57690
rect 1104 57616 18860 57638
rect 4985 57579 5043 57585
rect 4985 57545 4997 57579
rect 5031 57576 5043 57579
rect 5442 57576 5448 57588
rect 5031 57548 5448 57576
rect 5031 57545 5043 57548
rect 4985 57539 5043 57545
rect 5442 57536 5448 57548
rect 5500 57536 5506 57588
rect 8941 57579 8999 57585
rect 8941 57545 8953 57579
rect 8987 57576 8999 57579
rect 9306 57576 9312 57588
rect 8987 57548 9312 57576
rect 8987 57545 8999 57548
rect 8941 57539 8999 57545
rect 9306 57536 9312 57548
rect 9364 57576 9370 57588
rect 9582 57576 9588 57588
rect 9364 57548 9588 57576
rect 9364 57536 9370 57548
rect 9582 57536 9588 57548
rect 9640 57536 9646 57588
rect 10318 57536 10324 57588
rect 10376 57576 10382 57588
rect 10597 57579 10655 57585
rect 10597 57576 10609 57579
rect 10376 57548 10609 57576
rect 10376 57536 10382 57548
rect 10597 57545 10609 57548
rect 10643 57545 10655 57579
rect 10597 57539 10655 57545
rect 12713 57579 12771 57585
rect 12713 57545 12725 57579
rect 12759 57576 12771 57579
rect 12802 57576 12808 57588
rect 12759 57548 12808 57576
rect 12759 57545 12771 57548
rect 12713 57539 12771 57545
rect 12802 57536 12808 57548
rect 12860 57536 12866 57588
rect 6362 57468 6368 57520
rect 6420 57508 6426 57520
rect 7558 57508 7564 57520
rect 6420 57480 7564 57508
rect 6420 57468 6426 57480
rect 7558 57468 7564 57480
rect 7616 57468 7622 57520
rect 14642 57508 14648 57520
rect 11532 57480 14648 57508
rect 2038 57400 2044 57452
rect 2096 57440 2102 57452
rect 2133 57443 2191 57449
rect 2133 57440 2145 57443
rect 2096 57412 2145 57440
rect 2096 57400 2102 57412
rect 2133 57409 2145 57412
rect 2179 57409 2191 57443
rect 2133 57403 2191 57409
rect 3145 57443 3203 57449
rect 3145 57409 3157 57443
rect 3191 57440 3203 57443
rect 3694 57440 3700 57452
rect 3191 57412 3700 57440
rect 3191 57409 3203 57412
rect 3145 57403 3203 57409
rect 3694 57400 3700 57412
rect 3752 57440 3758 57452
rect 4249 57443 4307 57449
rect 4249 57440 4261 57443
rect 3752 57412 4261 57440
rect 3752 57400 3758 57412
rect 4249 57409 4261 57412
rect 4295 57409 4307 57443
rect 4249 57403 4307 57409
rect 5353 57443 5411 57449
rect 5353 57409 5365 57443
rect 5399 57440 5411 57443
rect 6457 57443 6515 57449
rect 5399 57412 6408 57440
rect 5399 57409 5411 57412
rect 5353 57403 5411 57409
rect 2685 57375 2743 57381
rect 2685 57341 2697 57375
rect 2731 57341 2743 57375
rect 2685 57335 2743 57341
rect 2961 57375 3019 57381
rect 2961 57341 2973 57375
rect 3007 57372 3019 57375
rect 3050 57372 3056 57384
rect 3007 57344 3056 57372
rect 3007 57341 3019 57344
rect 2961 57335 3019 57341
rect 2700 57304 2728 57335
rect 3050 57332 3056 57344
rect 3108 57332 3114 57384
rect 6380 57381 6408 57412
rect 6457 57409 6469 57443
rect 6503 57440 6515 57443
rect 6730 57440 6736 57452
rect 6503 57412 6736 57440
rect 6503 57409 6515 57412
rect 6457 57403 6515 57409
rect 6730 57400 6736 57412
rect 6788 57400 6794 57452
rect 9858 57400 9864 57452
rect 9916 57440 9922 57452
rect 10870 57440 10876 57452
rect 9916 57412 10876 57440
rect 9916 57400 9922 57412
rect 10870 57400 10876 57412
rect 10928 57400 10934 57452
rect 6365 57375 6423 57381
rect 6365 57341 6377 57375
rect 6411 57372 6423 57375
rect 6822 57372 6828 57384
rect 6411 57344 6828 57372
rect 6411 57341 6423 57344
rect 6365 57335 6423 57341
rect 6822 57332 6828 57344
rect 6880 57332 6886 57384
rect 7193 57375 7251 57381
rect 7193 57341 7205 57375
rect 7239 57372 7251 57375
rect 7282 57372 7288 57384
rect 7239 57344 7288 57372
rect 7239 57341 7251 57344
rect 7193 57335 7251 57341
rect 7282 57332 7288 57344
rect 7340 57332 7346 57384
rect 7377 57375 7435 57381
rect 7377 57341 7389 57375
rect 7423 57341 7435 57375
rect 7377 57335 7435 57341
rect 10137 57375 10195 57381
rect 10137 57341 10149 57375
rect 10183 57372 10195 57375
rect 10318 57372 10324 57384
rect 10183 57344 10324 57372
rect 10183 57341 10195 57344
rect 10137 57335 10195 57341
rect 5629 57307 5687 57313
rect 2700 57276 3556 57304
rect 1673 57239 1731 57245
rect 1673 57205 1685 57239
rect 1719 57236 1731 57239
rect 2041 57239 2099 57245
rect 2041 57236 2053 57239
rect 1719 57208 2053 57236
rect 1719 57205 1731 57208
rect 1673 57199 1731 57205
rect 2041 57205 2053 57208
rect 2087 57236 2099 57239
rect 2222 57236 2228 57248
rect 2087 57208 2228 57236
rect 2087 57205 2099 57208
rect 2041 57199 2099 57205
rect 2222 57196 2228 57208
rect 2280 57196 2286 57248
rect 3528 57245 3556 57276
rect 5629 57273 5641 57307
rect 5675 57304 5687 57307
rect 6638 57304 6644 57316
rect 5675 57276 6644 57304
rect 5675 57273 5687 57276
rect 5629 57267 5687 57273
rect 6638 57264 6644 57276
rect 6696 57304 6702 57316
rect 7392 57304 7420 57335
rect 10318 57332 10324 57344
rect 10376 57332 10382 57384
rect 10962 57332 10968 57384
rect 11020 57372 11026 57384
rect 11057 57375 11115 57381
rect 11057 57372 11069 57375
rect 11020 57344 11069 57372
rect 11020 57332 11026 57344
rect 11057 57341 11069 57344
rect 11103 57372 11115 57375
rect 11425 57375 11483 57381
rect 11425 57372 11437 57375
rect 11103 57344 11437 57372
rect 11103 57341 11115 57344
rect 11057 57335 11115 57341
rect 11425 57341 11437 57344
rect 11471 57372 11483 57375
rect 11532 57372 11560 57480
rect 14642 57468 14648 57480
rect 14700 57468 14706 57520
rect 11790 57440 11796 57452
rect 11751 57412 11796 57440
rect 11790 57400 11796 57412
rect 11848 57400 11854 57452
rect 12250 57440 12256 57452
rect 11900 57412 12256 57440
rect 11471 57344 11560 57372
rect 11701 57375 11759 57381
rect 11471 57341 11483 57344
rect 11425 57335 11483 57341
rect 11701 57341 11713 57375
rect 11747 57372 11759 57375
rect 11900 57372 11928 57412
rect 12250 57400 12256 57412
rect 12308 57400 12314 57452
rect 15841 57443 15899 57449
rect 15841 57409 15853 57443
rect 15887 57440 15899 57443
rect 15887 57412 16252 57440
rect 15887 57409 15899 57412
rect 15841 57403 15899 57409
rect 16224 57384 16252 57412
rect 11747 57344 11928 57372
rect 12161 57375 12219 57381
rect 11747 57341 11759 57344
rect 11701 57335 11759 57341
rect 12161 57341 12173 57375
rect 12207 57341 12219 57375
rect 12161 57335 12219 57341
rect 6696 57276 7420 57304
rect 6696 57264 6702 57276
rect 7650 57264 7656 57316
rect 7708 57264 7714 57316
rect 9766 57264 9772 57316
rect 9824 57304 9830 57316
rect 9824 57276 10364 57304
rect 9824 57264 9830 57276
rect 3513 57239 3571 57245
rect 3513 57205 3525 57239
rect 3559 57236 3571 57239
rect 3694 57236 3700 57248
rect 3559 57208 3700 57236
rect 3559 57205 3571 57208
rect 3513 57199 3571 57205
rect 3694 57196 3700 57208
rect 3752 57196 3758 57248
rect 3881 57239 3939 57245
rect 3881 57205 3893 57239
rect 3927 57236 3939 57239
rect 4614 57236 4620 57248
rect 3927 57208 4620 57236
rect 3927 57205 3939 57208
rect 3881 57199 3939 57205
rect 4614 57196 4620 57208
rect 4672 57236 4678 57248
rect 5442 57236 5448 57248
rect 4672 57208 5448 57236
rect 4672 57196 4678 57208
rect 5442 57196 5448 57208
rect 5500 57196 5506 57248
rect 5718 57196 5724 57248
rect 5776 57236 5782 57248
rect 6733 57239 6791 57245
rect 6733 57236 6745 57239
rect 5776 57208 6745 57236
rect 5776 57196 5782 57208
rect 6733 57205 6745 57208
rect 6779 57205 6791 57239
rect 6733 57199 6791 57205
rect 7374 57196 7380 57248
rect 7432 57236 7438 57248
rect 7668 57236 7696 57264
rect 7929 57239 7987 57245
rect 7929 57236 7941 57239
rect 7432 57208 7941 57236
rect 7432 57196 7438 57208
rect 7929 57205 7941 57208
rect 7975 57205 7987 57239
rect 8386 57236 8392 57248
rect 8347 57208 8392 57236
rect 7929 57199 7987 57205
rect 8386 57196 8392 57208
rect 8444 57236 8450 57248
rect 9217 57239 9275 57245
rect 9217 57236 9229 57239
rect 8444 57208 9229 57236
rect 8444 57196 8450 57208
rect 9217 57205 9229 57208
rect 9263 57205 9275 57239
rect 9217 57199 9275 57205
rect 9858 57196 9864 57248
rect 9916 57236 9922 57248
rect 10336 57245 10364 57276
rect 9953 57239 10011 57245
rect 9953 57236 9965 57239
rect 9916 57208 9965 57236
rect 9916 57196 9922 57208
rect 9953 57205 9965 57208
rect 9999 57205 10011 57239
rect 9953 57199 10011 57205
rect 10321 57239 10379 57245
rect 10321 57205 10333 57239
rect 10367 57205 10379 57239
rect 12176 57236 12204 57335
rect 12526 57332 12532 57384
rect 12584 57372 12590 57384
rect 15930 57372 15936 57384
rect 12584 57344 13492 57372
rect 15891 57344 15936 57372
rect 12584 57332 12590 57344
rect 12710 57264 12716 57316
rect 12768 57304 12774 57316
rect 12989 57307 13047 57313
rect 12989 57304 13001 57307
rect 12768 57276 13001 57304
rect 12768 57264 12774 57276
rect 12989 57273 13001 57276
rect 13035 57304 13047 57307
rect 13170 57304 13176 57316
rect 13035 57276 13176 57304
rect 13035 57273 13047 57276
rect 12989 57267 13047 57273
rect 13170 57264 13176 57276
rect 13228 57264 13234 57316
rect 13464 57248 13492 57344
rect 15930 57332 15936 57344
rect 15988 57332 15994 57384
rect 16206 57372 16212 57384
rect 16167 57344 16212 57372
rect 16206 57332 16212 57344
rect 16264 57332 16270 57384
rect 12250 57236 12256 57248
rect 12176 57208 12256 57236
rect 10321 57199 10379 57205
rect 12250 57196 12256 57208
rect 12308 57236 12314 57248
rect 12802 57236 12808 57248
rect 12308 57208 12808 57236
rect 12308 57196 12314 57208
rect 12802 57196 12808 57208
rect 12860 57196 12866 57248
rect 13446 57236 13452 57248
rect 13407 57208 13452 57236
rect 13446 57196 13452 57208
rect 13504 57196 13510 57248
rect 17310 57236 17316 57248
rect 17271 57208 17316 57236
rect 17310 57196 17316 57208
rect 17368 57196 17374 57248
rect 1104 57146 18860 57168
rect 1104 57094 7648 57146
rect 7700 57094 7712 57146
rect 7764 57094 7776 57146
rect 7828 57094 7840 57146
rect 7892 57094 14315 57146
rect 14367 57094 14379 57146
rect 14431 57094 14443 57146
rect 14495 57094 14507 57146
rect 14559 57094 18860 57146
rect 1104 57072 18860 57094
rect 4065 57035 4123 57041
rect 4065 57001 4077 57035
rect 4111 57032 4123 57035
rect 4798 57032 4804 57044
rect 4111 57004 4804 57032
rect 4111 57001 4123 57004
rect 4065 56995 4123 57001
rect 4798 56992 4804 57004
rect 4856 57032 4862 57044
rect 5629 57035 5687 57041
rect 5629 57032 5641 57035
rect 4856 57004 5641 57032
rect 4856 56992 4862 57004
rect 5629 57001 5641 57004
rect 5675 57001 5687 57035
rect 6178 57032 6184 57044
rect 6139 57004 6184 57032
rect 5629 56995 5687 57001
rect 6178 56992 6184 57004
rect 6236 56992 6242 57044
rect 9033 57035 9091 57041
rect 9033 57001 9045 57035
rect 9079 57032 9091 57035
rect 9674 57032 9680 57044
rect 9079 57004 9680 57032
rect 9079 57001 9091 57004
rect 9033 56995 9091 57001
rect 9674 56992 9680 57004
rect 9732 56992 9738 57044
rect 11517 57035 11575 57041
rect 11517 57001 11529 57035
rect 11563 57032 11575 57035
rect 12066 57032 12072 57044
rect 11563 57004 12072 57032
rect 11563 57001 11575 57004
rect 11517 56995 11575 57001
rect 12066 56992 12072 57004
rect 12124 56992 12130 57044
rect 12161 57035 12219 57041
rect 12161 57001 12173 57035
rect 12207 57032 12219 57035
rect 12526 57032 12532 57044
rect 12207 57004 12532 57032
rect 12207 57001 12219 57004
rect 12161 56995 12219 57001
rect 12526 56992 12532 57004
rect 12584 56992 12590 57044
rect 3050 56924 3056 56976
rect 3108 56964 3114 56976
rect 3418 56964 3424 56976
rect 3108 56936 3424 56964
rect 3108 56924 3114 56936
rect 3418 56924 3424 56936
rect 3476 56924 3482 56976
rect 6822 56924 6828 56976
rect 6880 56964 6886 56976
rect 8205 56967 8263 56973
rect 8205 56964 8217 56967
rect 6880 56936 8217 56964
rect 6880 56924 6886 56936
rect 1670 56856 1676 56908
rect 1728 56896 1734 56908
rect 1857 56899 1915 56905
rect 1857 56896 1869 56899
rect 1728 56868 1869 56896
rect 1728 56856 1734 56868
rect 1857 56865 1869 56868
rect 1903 56896 1915 56899
rect 3510 56896 3516 56908
rect 1903 56868 3516 56896
rect 1903 56865 1915 56868
rect 1857 56859 1915 56865
rect 3510 56856 3516 56868
rect 3568 56856 3574 56908
rect 4525 56899 4583 56905
rect 4525 56865 4537 56899
rect 4571 56896 4583 56899
rect 4798 56896 4804 56908
rect 4571 56868 4804 56896
rect 4571 56865 4583 56868
rect 4525 56859 4583 56865
rect 4798 56856 4804 56868
rect 4856 56856 4862 56908
rect 6178 56856 6184 56908
rect 6236 56896 6242 56908
rect 7668 56905 7696 56936
rect 8205 56933 8217 56936
rect 8251 56933 8263 56967
rect 8205 56927 8263 56933
rect 8570 56924 8576 56976
rect 8628 56964 8634 56976
rect 9306 56964 9312 56976
rect 8628 56936 9312 56964
rect 8628 56924 8634 56936
rect 9306 56924 9312 56936
rect 9364 56924 9370 56976
rect 12434 56924 12440 56976
rect 12492 56964 12498 56976
rect 12492 56936 12537 56964
rect 12492 56924 12498 56936
rect 7193 56899 7251 56905
rect 7193 56896 7205 56899
rect 6236 56868 7205 56896
rect 6236 56856 6242 56868
rect 7193 56865 7205 56868
rect 7239 56865 7251 56899
rect 7193 56859 7251 56865
rect 7653 56899 7711 56905
rect 7653 56865 7665 56899
rect 7699 56865 7711 56899
rect 7653 56859 7711 56865
rect 8846 56856 8852 56908
rect 8904 56896 8910 56908
rect 9217 56899 9275 56905
rect 9217 56896 9229 56899
rect 8904 56868 9229 56896
rect 8904 56856 8910 56868
rect 9217 56865 9229 56868
rect 9263 56865 9275 56899
rect 9324 56896 9352 56924
rect 9490 56896 9496 56908
rect 9324 56868 9496 56896
rect 9217 56859 9275 56865
rect 9490 56856 9496 56868
rect 9548 56896 9554 56908
rect 9585 56899 9643 56905
rect 9585 56896 9597 56899
rect 9548 56868 9597 56896
rect 9548 56856 9554 56868
rect 9585 56865 9597 56868
rect 9631 56865 9643 56899
rect 9585 56859 9643 56865
rect 9674 56856 9680 56908
rect 9732 56896 9738 56908
rect 10229 56899 10287 56905
rect 10229 56896 10241 56899
rect 9732 56868 10241 56896
rect 9732 56856 9738 56868
rect 10229 56865 10241 56868
rect 10275 56896 10287 56899
rect 10594 56896 10600 56908
rect 10275 56868 10600 56896
rect 10275 56865 10287 56868
rect 10229 56859 10287 56865
rect 10594 56856 10600 56868
rect 10652 56856 10658 56908
rect 10689 56899 10747 56905
rect 10689 56865 10701 56899
rect 10735 56865 10747 56899
rect 11698 56896 11704 56908
rect 11659 56868 11704 56896
rect 10689 56859 10747 56865
rect 1581 56831 1639 56837
rect 1581 56797 1593 56831
rect 1627 56828 1639 56831
rect 1762 56828 1768 56840
rect 1627 56800 1768 56828
rect 1627 56797 1639 56800
rect 1581 56791 1639 56797
rect 1762 56788 1768 56800
rect 1820 56828 1826 56840
rect 4249 56831 4307 56837
rect 4249 56828 4261 56831
rect 1820 56800 4261 56828
rect 1820 56788 1826 56800
rect 4249 56797 4261 56800
rect 4295 56797 4307 56831
rect 4249 56791 4307 56797
rect 6270 56788 6276 56840
rect 6328 56828 6334 56840
rect 6917 56831 6975 56837
rect 6917 56828 6929 56831
rect 6328 56800 6929 56828
rect 6328 56788 6334 56800
rect 6917 56797 6929 56800
rect 6963 56828 6975 56831
rect 7834 56828 7840 56840
rect 6963 56800 7840 56828
rect 6963 56797 6975 56800
rect 6917 56791 6975 56797
rect 7834 56788 7840 56800
rect 7892 56788 7898 56840
rect 8202 56788 8208 56840
rect 8260 56828 8266 56840
rect 9309 56831 9367 56837
rect 9309 56828 9321 56831
rect 8260 56800 9321 56828
rect 8260 56788 8266 56800
rect 9309 56797 9321 56800
rect 9355 56797 9367 56831
rect 9309 56791 9367 56797
rect 10410 56788 10416 56840
rect 10468 56828 10474 56840
rect 10704 56828 10732 56859
rect 11698 56856 11704 56868
rect 11756 56856 11762 56908
rect 12618 56856 12624 56908
rect 12676 56896 12682 56908
rect 12986 56896 12992 56908
rect 12676 56868 12992 56896
rect 12676 56856 12682 56868
rect 12986 56856 12992 56868
rect 13044 56856 13050 56908
rect 15289 56831 15347 56837
rect 15289 56828 15301 56831
rect 10468 56800 10732 56828
rect 14200 56800 15301 56828
rect 10468 56788 10474 56800
rect 7466 56720 7472 56772
rect 7524 56760 7530 56772
rect 7653 56763 7711 56769
rect 7653 56760 7665 56763
rect 7524 56732 7665 56760
rect 7524 56720 7530 56732
rect 7653 56729 7665 56732
rect 7699 56729 7711 56763
rect 7653 56723 7711 56729
rect 14200 56704 14228 56800
rect 15289 56797 15301 56800
rect 15335 56797 15347 56831
rect 15289 56791 15347 56797
rect 15565 56831 15623 56837
rect 15565 56797 15577 56831
rect 15611 56828 15623 56831
rect 15654 56828 15660 56840
rect 15611 56800 15660 56828
rect 15611 56797 15623 56800
rect 15565 56791 15623 56797
rect 15654 56788 15660 56800
rect 15712 56788 15718 56840
rect 2682 56652 2688 56704
rect 2740 56692 2746 56704
rect 2961 56695 3019 56701
rect 2961 56692 2973 56695
rect 2740 56664 2973 56692
rect 2740 56652 2746 56664
rect 2961 56661 2973 56664
rect 3007 56661 3019 56695
rect 2961 56655 3019 56661
rect 3510 56652 3516 56704
rect 3568 56692 3574 56704
rect 3605 56695 3663 56701
rect 3605 56692 3617 56695
rect 3568 56664 3617 56692
rect 3568 56652 3574 56664
rect 3605 56661 3617 56664
rect 3651 56692 3663 56695
rect 5718 56692 5724 56704
rect 3651 56664 5724 56692
rect 3651 56661 3663 56664
rect 3605 56655 3663 56661
rect 5718 56652 5724 56664
rect 5776 56652 5782 56704
rect 6641 56695 6699 56701
rect 6641 56661 6653 56695
rect 6687 56692 6699 56695
rect 6730 56692 6736 56704
rect 6687 56664 6736 56692
rect 6687 56661 6699 56664
rect 6641 56655 6699 56661
rect 6730 56652 6736 56664
rect 6788 56652 6794 56704
rect 8570 56652 8576 56704
rect 8628 56692 8634 56704
rect 8849 56695 8907 56701
rect 8849 56692 8861 56695
rect 8628 56664 8861 56692
rect 8628 56652 8634 56664
rect 8849 56661 8861 56664
rect 8895 56692 8907 56695
rect 9033 56695 9091 56701
rect 9033 56692 9045 56695
rect 8895 56664 9045 56692
rect 8895 56661 8907 56664
rect 8849 56655 8907 56661
rect 9033 56661 9045 56664
rect 9079 56661 9091 56695
rect 9033 56655 9091 56661
rect 11241 56695 11299 56701
rect 11241 56661 11253 56695
rect 11287 56692 11299 56695
rect 12250 56692 12256 56704
rect 11287 56664 12256 56692
rect 11287 56661 11299 56664
rect 11241 56655 11299 56661
rect 12250 56652 12256 56664
rect 12308 56652 12314 56704
rect 12802 56652 12808 56704
rect 12860 56692 12866 56704
rect 13449 56695 13507 56701
rect 13449 56692 13461 56695
rect 12860 56664 13461 56692
rect 12860 56652 12866 56664
rect 13449 56661 13461 56664
rect 13495 56661 13507 56695
rect 13449 56655 13507 56661
rect 13909 56695 13967 56701
rect 13909 56661 13921 56695
rect 13955 56692 13967 56695
rect 14182 56692 14188 56704
rect 13955 56664 14188 56692
rect 13955 56661 13967 56664
rect 13909 56655 13967 56661
rect 14182 56652 14188 56664
rect 14240 56652 14246 56704
rect 16666 56692 16672 56704
rect 16627 56664 16672 56692
rect 16666 56652 16672 56664
rect 16724 56652 16730 56704
rect 1104 56602 18860 56624
rect 1104 56550 4315 56602
rect 4367 56550 4379 56602
rect 4431 56550 4443 56602
rect 4495 56550 4507 56602
rect 4559 56550 10982 56602
rect 11034 56550 11046 56602
rect 11098 56550 11110 56602
rect 11162 56550 11174 56602
rect 11226 56550 17648 56602
rect 17700 56550 17712 56602
rect 17764 56550 17776 56602
rect 17828 56550 17840 56602
rect 17892 56550 18860 56602
rect 1104 56528 18860 56550
rect 1486 56448 1492 56500
rect 1544 56488 1550 56500
rect 1581 56491 1639 56497
rect 1581 56488 1593 56491
rect 1544 56460 1593 56488
rect 1544 56448 1550 56460
rect 1581 56457 1593 56460
rect 1627 56488 1639 56491
rect 2317 56491 2375 56497
rect 2317 56488 2329 56491
rect 1627 56460 2329 56488
rect 1627 56457 1639 56460
rect 1581 56451 1639 56457
rect 2317 56457 2329 56460
rect 2363 56457 2375 56491
rect 2317 56451 2375 56457
rect 3881 56491 3939 56497
rect 3881 56457 3893 56491
rect 3927 56488 3939 56491
rect 4798 56488 4804 56500
rect 3927 56460 4804 56488
rect 3927 56457 3939 56460
rect 3881 56451 3939 56457
rect 4798 56448 4804 56460
rect 4856 56448 4862 56500
rect 4982 56448 4988 56500
rect 5040 56488 5046 56500
rect 5626 56488 5632 56500
rect 5040 56460 5120 56488
rect 5587 56460 5632 56488
rect 5040 56448 5046 56460
rect 3510 56380 3516 56432
rect 3568 56420 3574 56432
rect 4062 56420 4068 56432
rect 3568 56392 4068 56420
rect 3568 56380 3574 56392
rect 4062 56380 4068 56392
rect 4120 56380 4126 56432
rect 2682 56352 2688 56364
rect 2516 56324 2688 56352
rect 2516 56293 2544 56324
rect 2682 56312 2688 56324
rect 2740 56312 2746 56364
rect 3694 56312 3700 56364
rect 3752 56352 3758 56364
rect 4982 56352 4988 56364
rect 3752 56324 4988 56352
rect 3752 56312 3758 56324
rect 4982 56312 4988 56324
rect 5040 56312 5046 56364
rect 2501 56287 2559 56293
rect 2501 56253 2513 56287
rect 2547 56253 2559 56287
rect 2866 56284 2872 56296
rect 2827 56256 2872 56284
rect 2501 56247 2559 56253
rect 2866 56244 2872 56256
rect 2924 56244 2930 56296
rect 4065 56287 4123 56293
rect 4065 56253 4077 56287
rect 4111 56253 4123 56287
rect 4338 56284 4344 56296
rect 4299 56256 4344 56284
rect 4065 56247 4123 56253
rect 2133 56219 2191 56225
rect 2133 56185 2145 56219
rect 2179 56216 2191 56219
rect 2884 56216 2912 56244
rect 2179 56188 2912 56216
rect 2179 56185 2191 56188
rect 2133 56179 2191 56185
rect 4080 56160 4108 56247
rect 4338 56244 4344 56256
rect 4396 56244 4402 56296
rect 3513 56151 3571 56157
rect 3513 56117 3525 56151
rect 3559 56148 3571 56151
rect 4062 56148 4068 56160
rect 3559 56120 4068 56148
rect 3559 56117 3571 56120
rect 3513 56111 3571 56117
rect 4062 56108 4068 56120
rect 4120 56108 4126 56160
rect 4798 56108 4804 56160
rect 4856 56148 4862 56160
rect 5092 56148 5120 56460
rect 5626 56448 5632 56460
rect 5684 56448 5690 56500
rect 7098 56448 7104 56500
rect 7156 56488 7162 56500
rect 7282 56488 7288 56500
rect 7156 56460 7288 56488
rect 7156 56448 7162 56460
rect 7282 56448 7288 56460
rect 7340 56448 7346 56500
rect 7834 56448 7840 56500
rect 7892 56488 7898 56500
rect 7929 56491 7987 56497
rect 7929 56488 7941 56491
rect 7892 56460 7941 56488
rect 7892 56448 7898 56460
rect 7929 56457 7941 56460
rect 7975 56457 7987 56491
rect 7929 56451 7987 56457
rect 8481 56491 8539 56497
rect 8481 56457 8493 56491
rect 8527 56488 8539 56491
rect 8662 56488 8668 56500
rect 8527 56460 8668 56488
rect 8527 56457 8539 56460
rect 8481 56451 8539 56457
rect 7006 56380 7012 56432
rect 7064 56420 7070 56432
rect 7377 56423 7435 56429
rect 7377 56420 7389 56423
rect 7064 56392 7389 56420
rect 7064 56380 7070 56392
rect 7377 56389 7389 56392
rect 7423 56389 7435 56423
rect 7377 56383 7435 56389
rect 6362 56244 6368 56296
rect 6420 56284 6426 56296
rect 6549 56287 6607 56293
rect 6549 56284 6561 56287
rect 6420 56256 6561 56284
rect 6420 56244 6426 56256
rect 6549 56253 6561 56256
rect 6595 56253 6607 56287
rect 6549 56247 6607 56253
rect 6730 56244 6736 56296
rect 6788 56284 6794 56296
rect 7006 56284 7012 56296
rect 6788 56256 7012 56284
rect 6788 56244 6794 56256
rect 7006 56244 7012 56256
rect 7064 56244 7070 56296
rect 7377 56287 7435 56293
rect 7377 56253 7389 56287
rect 7423 56284 7435 56287
rect 8294 56284 8300 56296
rect 7423 56256 8300 56284
rect 7423 56253 7435 56256
rect 7377 56247 7435 56253
rect 7392 56216 7420 56247
rect 8294 56244 8300 56256
rect 8352 56244 8358 56296
rect 8588 56293 8616 56460
rect 8662 56448 8668 56460
rect 8720 56448 8726 56500
rect 11882 56488 11888 56500
rect 11843 56460 11888 56488
rect 11882 56448 11888 56460
rect 11940 56448 11946 56500
rect 9953 56423 10011 56429
rect 9953 56389 9965 56423
rect 9999 56420 10011 56423
rect 10410 56420 10416 56432
rect 9999 56392 10416 56420
rect 9999 56389 10011 56392
rect 9953 56383 10011 56389
rect 10410 56380 10416 56392
rect 10468 56380 10474 56432
rect 11609 56423 11667 56429
rect 11609 56389 11621 56423
rect 11655 56420 11667 56423
rect 12066 56420 12072 56432
rect 11655 56392 12072 56420
rect 11655 56389 11667 56392
rect 11609 56383 11667 56389
rect 10229 56355 10287 56361
rect 10229 56321 10241 56355
rect 10275 56352 10287 56355
rect 11624 56352 11652 56383
rect 12066 56380 12072 56392
rect 12124 56380 12130 56432
rect 10275 56324 11652 56352
rect 16025 56355 16083 56361
rect 10275 56321 10287 56324
rect 10229 56315 10287 56321
rect 16025 56321 16037 56355
rect 16071 56352 16083 56355
rect 16071 56324 16436 56352
rect 16071 56321 16083 56324
rect 16025 56315 16083 56321
rect 16408 56296 16436 56324
rect 8573 56287 8631 56293
rect 8573 56253 8585 56287
rect 8619 56284 8631 56287
rect 9858 56284 9864 56296
rect 8619 56256 9864 56284
rect 8619 56253 8631 56256
rect 8573 56247 8631 56253
rect 9858 56244 9864 56256
rect 9916 56244 9922 56296
rect 11057 56287 11115 56293
rect 11057 56253 11069 56287
rect 11103 56253 11115 56287
rect 11057 56247 11115 56253
rect 7466 56216 7472 56228
rect 6748 56188 7472 56216
rect 6748 56160 6776 56188
rect 7466 56176 7472 56188
rect 7524 56176 7530 56228
rect 10321 56219 10379 56225
rect 10321 56185 10333 56219
rect 10367 56216 10379 56219
rect 10410 56216 10416 56228
rect 10367 56188 10416 56216
rect 10367 56185 10379 56188
rect 10321 56179 10379 56185
rect 10410 56176 10416 56188
rect 10468 56176 10474 56228
rect 11072 56216 11100 56247
rect 11146 56244 11152 56296
rect 11204 56284 11210 56296
rect 12526 56284 12532 56296
rect 11204 56256 11249 56284
rect 12487 56256 12532 56284
rect 11204 56244 11210 56256
rect 12526 56244 12532 56256
rect 12584 56244 12590 56296
rect 16117 56287 16175 56293
rect 16117 56284 16129 56287
rect 15028 56256 16129 56284
rect 11882 56216 11888 56228
rect 11072 56188 11888 56216
rect 11882 56176 11888 56188
rect 11940 56176 11946 56228
rect 13541 56219 13599 56225
rect 13541 56185 13553 56219
rect 13587 56216 13599 56219
rect 13722 56216 13728 56228
rect 13587 56188 13728 56216
rect 13587 56185 13599 56188
rect 13541 56179 13599 56185
rect 13722 56176 13728 56188
rect 13780 56216 13786 56228
rect 13817 56219 13875 56225
rect 13817 56216 13829 56219
rect 13780 56188 13829 56216
rect 13780 56176 13786 56188
rect 13817 56185 13829 56188
rect 13863 56185 13875 56219
rect 13817 56179 13875 56185
rect 4856 56120 5120 56148
rect 6089 56151 6147 56157
rect 4856 56108 4862 56120
rect 6089 56117 6101 56151
rect 6135 56148 6147 56151
rect 6178 56148 6184 56160
rect 6135 56120 6184 56148
rect 6135 56117 6147 56120
rect 6089 56111 6147 56117
rect 6178 56108 6184 56120
rect 6236 56108 6242 56160
rect 6457 56151 6515 56157
rect 6457 56117 6469 56151
rect 6503 56148 6515 56151
rect 6730 56148 6736 56160
rect 6503 56120 6736 56148
rect 6503 56117 6515 56120
rect 6457 56111 6515 56117
rect 6730 56108 6736 56120
rect 6788 56108 6794 56160
rect 8757 56151 8815 56157
rect 8757 56117 8769 56151
rect 8803 56148 8815 56151
rect 8938 56148 8944 56160
rect 8803 56120 8944 56148
rect 8803 56117 8815 56120
rect 8757 56111 8815 56117
rect 8938 56108 8944 56120
rect 8996 56108 9002 56160
rect 9306 56148 9312 56160
rect 9267 56120 9312 56148
rect 9306 56108 9312 56120
rect 9364 56108 9370 56160
rect 12526 56148 12532 56160
rect 12487 56120 12532 56148
rect 12526 56108 12532 56120
rect 12584 56108 12590 56160
rect 12986 56108 12992 56160
rect 13044 56148 13050 56160
rect 13081 56151 13139 56157
rect 13081 56148 13093 56151
rect 13044 56120 13093 56148
rect 13044 56108 13050 56120
rect 13081 56117 13093 56120
rect 13127 56117 13139 56151
rect 14182 56148 14188 56160
rect 14143 56120 14188 56148
rect 13081 56111 13139 56117
rect 14182 56108 14188 56120
rect 14240 56148 14246 56160
rect 15028 56157 15056 56256
rect 16117 56253 16129 56256
rect 16163 56253 16175 56287
rect 16390 56284 16396 56296
rect 16351 56256 16396 56284
rect 16117 56247 16175 56253
rect 16390 56244 16396 56256
rect 16448 56244 16454 56296
rect 14645 56151 14703 56157
rect 14645 56148 14657 56151
rect 14240 56120 14657 56148
rect 14240 56108 14246 56120
rect 14645 56117 14657 56120
rect 14691 56148 14703 56151
rect 15013 56151 15071 56157
rect 15013 56148 15025 56151
rect 14691 56120 15025 56148
rect 14691 56117 14703 56120
rect 14645 56111 14703 56117
rect 15013 56117 15025 56120
rect 15059 56117 15071 56151
rect 15013 56111 15071 56117
rect 15565 56151 15623 56157
rect 15565 56117 15577 56151
rect 15611 56148 15623 56151
rect 15654 56148 15660 56160
rect 15611 56120 15660 56148
rect 15611 56117 15623 56120
rect 15565 56111 15623 56117
rect 15654 56108 15660 56120
rect 15712 56108 15718 56160
rect 17494 56148 17500 56160
rect 17455 56120 17500 56148
rect 17494 56108 17500 56120
rect 17552 56108 17558 56160
rect 1104 56058 18860 56080
rect 1104 56006 7648 56058
rect 7700 56006 7712 56058
rect 7764 56006 7776 56058
rect 7828 56006 7840 56058
rect 7892 56006 14315 56058
rect 14367 56006 14379 56058
rect 14431 56006 14443 56058
rect 14495 56006 14507 56058
rect 14559 56006 18860 56058
rect 1104 55984 18860 56006
rect 1670 55944 1676 55956
rect 1631 55916 1676 55944
rect 1670 55904 1676 55916
rect 1728 55904 1734 55956
rect 2317 55947 2375 55953
rect 2317 55913 2329 55947
rect 2363 55944 2375 55947
rect 2682 55944 2688 55956
rect 2363 55916 2688 55944
rect 2363 55913 2375 55916
rect 2317 55907 2375 55913
rect 2682 55904 2688 55916
rect 2740 55904 2746 55956
rect 4525 55947 4583 55953
rect 4525 55913 4537 55947
rect 4571 55944 4583 55947
rect 6270 55944 6276 55956
rect 4571 55916 6276 55944
rect 4571 55913 4583 55916
rect 4525 55907 4583 55913
rect 6270 55904 6276 55916
rect 6328 55904 6334 55956
rect 6454 55944 6460 55956
rect 6415 55916 6460 55944
rect 6454 55904 6460 55916
rect 6512 55904 6518 55956
rect 8294 55944 8300 55956
rect 8255 55916 8300 55944
rect 8294 55904 8300 55916
rect 8352 55904 8358 55956
rect 8846 55944 8852 55956
rect 8807 55916 8852 55944
rect 8846 55904 8852 55916
rect 8904 55904 8910 55956
rect 9401 55947 9459 55953
rect 9401 55913 9413 55947
rect 9447 55944 9459 55947
rect 9490 55944 9496 55956
rect 9447 55916 9496 55944
rect 9447 55913 9459 55916
rect 9401 55907 9459 55913
rect 9490 55904 9496 55916
rect 9548 55904 9554 55956
rect 9674 55944 9680 55956
rect 9600 55916 9680 55944
rect 1762 55836 1768 55888
rect 1820 55876 1826 55888
rect 3697 55879 3755 55885
rect 3697 55876 3709 55879
rect 1820 55848 3709 55876
rect 1820 55836 1826 55848
rect 3697 55845 3709 55848
rect 3743 55845 3755 55879
rect 4890 55876 4896 55888
rect 3697 55839 3755 55845
rect 4816 55848 4896 55876
rect 2406 55768 2412 55820
rect 2464 55808 2470 55820
rect 2682 55808 2688 55820
rect 2464 55780 2688 55808
rect 2464 55768 2470 55780
rect 2682 55768 2688 55780
rect 2740 55768 2746 55820
rect 4816 55817 4844 55848
rect 4890 55836 4896 55848
rect 4948 55836 4954 55888
rect 6914 55836 6920 55888
rect 6972 55876 6978 55888
rect 7929 55879 7987 55885
rect 7929 55876 7941 55879
rect 6972 55848 7941 55876
rect 6972 55836 6978 55848
rect 7929 55845 7941 55848
rect 7975 55845 7987 55879
rect 7929 55839 7987 55845
rect 9309 55879 9367 55885
rect 9309 55845 9321 55879
rect 9355 55876 9367 55879
rect 9600 55876 9628 55916
rect 9674 55904 9680 55916
rect 9732 55904 9738 55956
rect 10962 55904 10968 55956
rect 11020 55904 11026 55956
rect 11146 55904 11152 55956
rect 11204 55944 11210 55956
rect 11517 55947 11575 55953
rect 11517 55944 11529 55947
rect 11204 55916 11529 55944
rect 11204 55904 11210 55916
rect 11517 55913 11529 55916
rect 11563 55913 11575 55947
rect 11517 55907 11575 55913
rect 12069 55947 12127 55953
rect 12069 55913 12081 55947
rect 12115 55944 12127 55947
rect 12158 55944 12164 55956
rect 12115 55916 12164 55944
rect 12115 55913 12127 55916
rect 12069 55907 12127 55913
rect 12158 55904 12164 55916
rect 12216 55904 12222 55956
rect 12805 55947 12863 55953
rect 12805 55913 12817 55947
rect 12851 55944 12863 55947
rect 12989 55947 13047 55953
rect 12989 55944 13001 55947
rect 12851 55916 13001 55944
rect 12851 55913 12863 55916
rect 12805 55907 12863 55913
rect 12989 55913 13001 55916
rect 13035 55944 13047 55947
rect 17310 55944 17316 55956
rect 13035 55916 17316 55944
rect 13035 55913 13047 55916
rect 12989 55907 13047 55913
rect 17310 55904 17316 55916
rect 17368 55904 17374 55956
rect 10980 55876 11008 55904
rect 12526 55876 12532 55888
rect 9355 55848 9628 55876
rect 9692 55848 11008 55876
rect 12360 55848 12532 55876
rect 9355 55845 9367 55848
rect 9309 55839 9367 55845
rect 9692 55820 9720 55848
rect 4801 55811 4859 55817
rect 4801 55777 4813 55811
rect 4847 55777 4859 55811
rect 4982 55808 4988 55820
rect 4943 55780 4988 55808
rect 4801 55771 4859 55777
rect 4982 55768 4988 55780
rect 5040 55768 5046 55820
rect 5166 55808 5172 55820
rect 5127 55780 5172 55808
rect 5166 55768 5172 55780
rect 5224 55768 5230 55820
rect 6641 55811 6699 55817
rect 6641 55777 6653 55811
rect 6687 55777 6699 55811
rect 6641 55771 6699 55777
rect 4338 55632 4344 55684
rect 4396 55632 4402 55684
rect 6178 55632 6184 55684
rect 6236 55672 6242 55684
rect 6656 55672 6684 55771
rect 7006 55768 7012 55820
rect 7064 55808 7070 55820
rect 7193 55811 7251 55817
rect 7193 55808 7205 55811
rect 7064 55780 7205 55808
rect 7064 55768 7070 55780
rect 7193 55777 7205 55780
rect 7239 55777 7251 55811
rect 7193 55771 7251 55777
rect 7466 55768 7472 55820
rect 7524 55808 7530 55820
rect 7653 55811 7711 55817
rect 7653 55808 7665 55811
rect 7524 55780 7665 55808
rect 7524 55768 7530 55780
rect 7653 55777 7665 55780
rect 7699 55777 7711 55811
rect 7653 55771 7711 55777
rect 9585 55811 9643 55817
rect 9585 55777 9597 55811
rect 9631 55808 9643 55811
rect 9674 55808 9680 55820
rect 9631 55780 9680 55808
rect 9631 55777 9643 55780
rect 9585 55771 9643 55777
rect 6914 55740 6920 55752
rect 6875 55712 6920 55740
rect 6914 55700 6920 55712
rect 6972 55740 6978 55752
rect 7282 55740 7288 55752
rect 6972 55712 7288 55740
rect 6972 55700 6978 55712
rect 7282 55700 7288 55712
rect 7340 55700 7346 55752
rect 9600 55740 9628 55771
rect 9674 55768 9680 55780
rect 9732 55768 9738 55820
rect 9769 55811 9827 55817
rect 9769 55777 9781 55811
rect 9815 55777 9827 55811
rect 9769 55771 9827 55777
rect 8312 55712 9628 55740
rect 8312 55672 8340 55712
rect 6236 55644 8340 55672
rect 6236 55632 6242 55644
rect 8846 55632 8852 55684
rect 8904 55672 8910 55684
rect 9784 55672 9812 55771
rect 9858 55768 9864 55820
rect 9916 55808 9922 55820
rect 10045 55811 10103 55817
rect 10045 55808 10057 55811
rect 9916 55780 10057 55808
rect 9916 55768 9922 55780
rect 10045 55777 10057 55780
rect 10091 55777 10103 55811
rect 10045 55771 10103 55777
rect 10060 55740 10088 55771
rect 10318 55768 10324 55820
rect 10376 55808 10382 55820
rect 10413 55811 10471 55817
rect 10413 55808 10425 55811
rect 10376 55780 10425 55808
rect 10376 55768 10382 55780
rect 10413 55777 10425 55780
rect 10459 55777 10471 55811
rect 10413 55771 10471 55777
rect 12253 55811 12311 55817
rect 12253 55777 12265 55811
rect 12299 55808 12311 55811
rect 12360 55808 12388 55848
rect 12526 55836 12532 55848
rect 12584 55876 12590 55888
rect 12710 55876 12716 55888
rect 12584 55848 12716 55876
rect 12584 55836 12590 55848
rect 12710 55836 12716 55848
rect 12768 55836 12774 55888
rect 13078 55836 13084 55888
rect 13136 55836 13142 55888
rect 13449 55879 13507 55885
rect 13449 55845 13461 55879
rect 13495 55876 13507 55879
rect 13722 55876 13728 55888
rect 13495 55848 13728 55876
rect 13495 55845 13507 55848
rect 13449 55839 13507 55845
rect 13722 55836 13728 55848
rect 13780 55836 13786 55888
rect 12299 55780 12388 55808
rect 12437 55811 12495 55817
rect 12299 55777 12311 55780
rect 12253 55771 12311 55777
rect 12437 55777 12449 55811
rect 12483 55808 12495 55811
rect 12802 55808 12808 55820
rect 12483 55780 12808 55808
rect 12483 55777 12495 55780
rect 12437 55771 12495 55777
rect 12802 55768 12808 55780
rect 12860 55808 12866 55820
rect 13096 55808 13124 55836
rect 14182 55808 14188 55820
rect 12860 55780 13124 55808
rect 13648 55780 14188 55808
rect 12860 55768 12866 55780
rect 10502 55740 10508 55752
rect 10060 55712 10508 55740
rect 10502 55700 10508 55712
rect 10560 55700 10566 55752
rect 10594 55700 10600 55752
rect 10652 55740 10658 55752
rect 11241 55743 11299 55749
rect 10652 55712 10697 55740
rect 10652 55700 10658 55712
rect 11241 55709 11253 55743
rect 11287 55740 11299 55743
rect 12066 55740 12072 55752
rect 11287 55712 12072 55740
rect 11287 55709 11299 55712
rect 11241 55703 11299 55709
rect 12066 55700 12072 55712
rect 12124 55700 12130 55752
rect 12158 55700 12164 55752
rect 12216 55740 12222 55752
rect 13078 55740 13084 55752
rect 12216 55712 13084 55740
rect 12216 55700 12222 55712
rect 13078 55700 13084 55712
rect 13136 55740 13142 55752
rect 13648 55749 13676 55780
rect 14182 55768 14188 55780
rect 14240 55808 14246 55820
rect 15378 55808 15384 55820
rect 14240 55780 15384 55808
rect 14240 55768 14246 55780
rect 15378 55768 15384 55780
rect 15436 55808 15442 55820
rect 15565 55811 15623 55817
rect 15565 55808 15577 55811
rect 15436 55780 15577 55808
rect 15436 55768 15442 55780
rect 15565 55777 15577 55780
rect 15611 55777 15623 55811
rect 15565 55771 15623 55777
rect 16945 55811 17003 55817
rect 16945 55777 16957 55811
rect 16991 55808 17003 55811
rect 17402 55808 17408 55820
rect 16991 55780 17408 55808
rect 16991 55777 17003 55780
rect 16945 55771 17003 55777
rect 17402 55768 17408 55780
rect 17460 55768 17466 55820
rect 13633 55743 13691 55749
rect 13633 55740 13645 55743
rect 13136 55712 13645 55740
rect 13136 55700 13142 55712
rect 13633 55709 13645 55712
rect 13679 55709 13691 55743
rect 13906 55740 13912 55752
rect 13867 55712 13912 55740
rect 13633 55703 13691 55709
rect 13906 55700 13912 55712
rect 13964 55700 13970 55752
rect 15470 55700 15476 55752
rect 15528 55740 15534 55752
rect 16117 55743 16175 55749
rect 16117 55740 16129 55743
rect 15528 55712 16129 55740
rect 15528 55700 15534 55712
rect 16117 55709 16129 55712
rect 16163 55709 16175 55743
rect 16117 55703 16175 55709
rect 16298 55700 16304 55752
rect 16356 55740 16362 55752
rect 16669 55743 16727 55749
rect 16669 55740 16681 55743
rect 16356 55712 16681 55740
rect 16356 55700 16362 55712
rect 16669 55709 16681 55712
rect 16715 55709 16727 55743
rect 17126 55740 17132 55752
rect 17087 55712 17132 55740
rect 16669 55703 16727 55709
rect 17126 55700 17132 55712
rect 17184 55700 17190 55752
rect 10870 55672 10876 55684
rect 8904 55644 10876 55672
rect 8904 55632 8910 55644
rect 10870 55632 10876 55644
rect 10928 55672 10934 55684
rect 12805 55675 12863 55681
rect 12805 55672 12817 55675
rect 10928 55644 12817 55672
rect 10928 55632 10934 55644
rect 12805 55641 12817 55644
rect 12851 55641 12863 55675
rect 12805 55635 12863 55641
rect 16025 55675 16083 55681
rect 16025 55641 16037 55675
rect 16071 55672 16083 55675
rect 16316 55672 16344 55700
rect 16071 55644 16344 55672
rect 16071 55641 16083 55644
rect 16025 55635 16083 55641
rect 4157 55607 4215 55613
rect 4157 55573 4169 55607
rect 4203 55604 4215 55607
rect 4356 55604 4384 55632
rect 4706 55604 4712 55616
rect 4203 55576 4712 55604
rect 4203 55573 4215 55576
rect 4157 55567 4215 55573
rect 4706 55564 4712 55576
rect 4764 55564 4770 55616
rect 5718 55604 5724 55616
rect 5679 55576 5724 55604
rect 5718 55564 5724 55576
rect 5776 55564 5782 55616
rect 6089 55607 6147 55613
rect 6089 55573 6101 55607
rect 6135 55604 6147 55607
rect 6270 55604 6276 55616
rect 6135 55576 6276 55604
rect 6135 55573 6147 55576
rect 6089 55567 6147 55573
rect 6270 55564 6276 55576
rect 6328 55564 6334 55616
rect 11882 55604 11888 55616
rect 11843 55576 11888 55604
rect 11882 55564 11888 55576
rect 11940 55564 11946 55616
rect 12066 55564 12072 55616
rect 12124 55604 12130 55616
rect 12621 55607 12679 55613
rect 12621 55604 12633 55607
rect 12124 55576 12633 55604
rect 12124 55564 12130 55576
rect 12621 55573 12633 55576
rect 12667 55573 12679 55607
rect 12621 55567 12679 55573
rect 15197 55607 15255 55613
rect 15197 55573 15209 55607
rect 15243 55604 15255 55607
rect 15286 55604 15292 55616
rect 15243 55576 15292 55604
rect 15243 55573 15255 55576
rect 15197 55567 15255 55573
rect 15286 55564 15292 55576
rect 15344 55564 15350 55616
rect 1104 55514 18860 55536
rect 1104 55462 4315 55514
rect 4367 55462 4379 55514
rect 4431 55462 4443 55514
rect 4495 55462 4507 55514
rect 4559 55462 10982 55514
rect 11034 55462 11046 55514
rect 11098 55462 11110 55514
rect 11162 55462 11174 55514
rect 11226 55462 17648 55514
rect 17700 55462 17712 55514
rect 17764 55462 17776 55514
rect 17828 55462 17840 55514
rect 17892 55462 18860 55514
rect 1104 55440 18860 55462
rect 1673 55403 1731 55409
rect 1673 55369 1685 55403
rect 1719 55400 1731 55403
rect 1762 55400 1768 55412
rect 1719 55372 1768 55400
rect 1719 55369 1731 55372
rect 1673 55363 1731 55369
rect 1762 55360 1768 55372
rect 1820 55360 1826 55412
rect 3142 55360 3148 55412
rect 3200 55400 3206 55412
rect 3418 55400 3424 55412
rect 3200 55372 3424 55400
rect 3200 55360 3206 55372
rect 3418 55360 3424 55372
rect 3476 55360 3482 55412
rect 3510 55360 3516 55412
rect 3568 55400 3574 55412
rect 3789 55403 3847 55409
rect 3789 55400 3801 55403
rect 3568 55372 3801 55400
rect 3568 55360 3574 55372
rect 3789 55369 3801 55372
rect 3835 55369 3847 55403
rect 3789 55363 3847 55369
rect 5353 55403 5411 55409
rect 5353 55369 5365 55403
rect 5399 55400 5411 55403
rect 6086 55400 6092 55412
rect 5399 55372 6092 55400
rect 5399 55369 5411 55372
rect 5353 55363 5411 55369
rect 2961 55199 3019 55205
rect 2961 55165 2973 55199
rect 3007 55196 3019 55199
rect 3142 55196 3148 55208
rect 3007 55168 3148 55196
rect 3007 55165 3019 55168
rect 2961 55159 3019 55165
rect 3142 55156 3148 55168
rect 3200 55156 3206 55208
rect 3804 55196 3832 55363
rect 6086 55360 6092 55372
rect 6144 55360 6150 55412
rect 8846 55360 8852 55412
rect 8904 55400 8910 55412
rect 9033 55403 9091 55409
rect 9033 55400 9045 55403
rect 8904 55372 9045 55400
rect 8904 55360 8910 55372
rect 9033 55369 9045 55372
rect 9079 55369 9091 55403
rect 9033 55363 9091 55369
rect 9401 55403 9459 55409
rect 9401 55369 9413 55403
rect 9447 55400 9459 55403
rect 10318 55400 10324 55412
rect 9447 55372 10324 55400
rect 9447 55369 9459 55372
rect 9401 55363 9459 55369
rect 10318 55360 10324 55372
rect 10376 55360 10382 55412
rect 10502 55400 10508 55412
rect 10463 55372 10508 55400
rect 10502 55360 10508 55372
rect 10560 55360 10566 55412
rect 11514 55360 11520 55412
rect 11572 55400 11578 55412
rect 12158 55400 12164 55412
rect 11572 55372 12164 55400
rect 11572 55360 11578 55372
rect 12158 55360 12164 55372
rect 12216 55360 12222 55412
rect 13906 55360 13912 55412
rect 13964 55360 13970 55412
rect 16298 55400 16304 55412
rect 14936 55372 16304 55400
rect 5534 55292 5540 55344
rect 5592 55332 5598 55344
rect 6273 55335 6331 55341
rect 6273 55332 6285 55335
rect 5592 55304 6285 55332
rect 5592 55292 5598 55304
rect 6273 55301 6285 55304
rect 6319 55301 6331 55335
rect 8757 55335 8815 55341
rect 8757 55332 8769 55335
rect 6273 55295 6331 55301
rect 7944 55304 8769 55332
rect 4801 55267 4859 55273
rect 4801 55233 4813 55267
rect 4847 55264 4859 55267
rect 5166 55264 5172 55276
rect 4847 55236 5172 55264
rect 4847 55233 4859 55236
rect 4801 55227 4859 55233
rect 5166 55224 5172 55236
rect 5224 55264 5230 55276
rect 5629 55267 5687 55273
rect 5224 55236 5488 55264
rect 5224 55224 5230 55236
rect 4249 55199 4307 55205
rect 4249 55196 4261 55199
rect 3804 55168 4261 55196
rect 4249 55165 4261 55168
rect 4295 55165 4307 55199
rect 5460 55196 5488 55236
rect 5629 55233 5641 55267
rect 5675 55264 5687 55267
rect 5718 55264 5724 55276
rect 5675 55236 5724 55264
rect 5675 55233 5687 55236
rect 5629 55227 5687 55233
rect 5718 55224 5724 55236
rect 5776 55264 5782 55276
rect 6917 55267 6975 55273
rect 5776 55236 6408 55264
rect 5776 55224 5782 55236
rect 5997 55199 6055 55205
rect 5460 55168 5764 55196
rect 4249 55159 4307 55165
rect 5736 55140 5764 55168
rect 5997 55165 6009 55199
rect 6043 55196 6055 55199
rect 6086 55196 6092 55208
rect 6043 55168 6092 55196
rect 6043 55165 6055 55168
rect 5997 55159 6055 55165
rect 6086 55156 6092 55168
rect 6144 55156 6150 55208
rect 6270 55196 6276 55208
rect 6231 55168 6276 55196
rect 6270 55156 6276 55168
rect 6328 55156 6334 55208
rect 6380 55196 6408 55236
rect 6917 55233 6929 55267
rect 6963 55264 6975 55267
rect 7006 55264 7012 55276
rect 6963 55236 7012 55264
rect 6963 55233 6975 55236
rect 6917 55227 6975 55233
rect 7006 55224 7012 55236
rect 7064 55224 7070 55276
rect 7944 55273 7972 55304
rect 8757 55301 8769 55304
rect 8803 55332 8815 55335
rect 9490 55332 9496 55344
rect 8803 55304 9496 55332
rect 8803 55301 8815 55304
rect 8757 55295 8815 55301
rect 9490 55292 9496 55304
rect 9548 55292 9554 55344
rect 13265 55335 13323 55341
rect 13265 55301 13277 55335
rect 13311 55332 13323 55335
rect 13924 55332 13952 55360
rect 14182 55332 14188 55344
rect 13311 55304 14188 55332
rect 13311 55301 13323 55304
rect 13265 55295 13323 55301
rect 14182 55292 14188 55304
rect 14240 55292 14246 55344
rect 7929 55267 7987 55273
rect 7929 55233 7941 55267
rect 7975 55233 7987 55267
rect 8294 55264 8300 55276
rect 7929 55227 7987 55233
rect 8220 55236 8300 55264
rect 8220 55205 8248 55236
rect 8294 55224 8300 55236
rect 8352 55224 8358 55276
rect 8662 55224 8668 55276
rect 8720 55264 8726 55276
rect 8846 55264 8852 55276
rect 8720 55236 8852 55264
rect 8720 55224 8726 55236
rect 8846 55224 8852 55236
rect 8904 55224 8910 55276
rect 9306 55224 9312 55276
rect 9364 55264 9370 55276
rect 11514 55264 11520 55276
rect 9364 55236 9720 55264
rect 11475 55236 11520 55264
rect 9364 55224 9370 55236
rect 8205 55199 8263 55205
rect 6380 55168 7512 55196
rect 4706 55088 4712 55140
rect 4764 55128 4770 55140
rect 5534 55128 5540 55140
rect 4764 55100 5540 55128
rect 4764 55088 4770 55100
rect 5534 55088 5540 55100
rect 5592 55088 5598 55140
rect 5718 55088 5724 55140
rect 5776 55088 5782 55140
rect 7374 55128 7380 55140
rect 7335 55100 7380 55128
rect 7374 55088 7380 55100
rect 7432 55088 7438 55140
rect 7484 55128 7512 55168
rect 8205 55165 8217 55199
rect 8251 55165 8263 55199
rect 8386 55196 8392 55208
rect 8299 55168 8392 55196
rect 8205 55159 8263 55165
rect 8220 55128 8248 55159
rect 8386 55156 8392 55168
rect 8444 55156 8450 55208
rect 9692 55205 9720 55236
rect 11514 55224 11520 55236
rect 11572 55224 11578 55276
rect 12066 55264 12072 55276
rect 11808 55236 12072 55264
rect 9677 55199 9735 55205
rect 9677 55165 9689 55199
rect 9723 55196 9735 55199
rect 9950 55196 9956 55208
rect 9723 55168 9956 55196
rect 9723 55165 9735 55168
rect 9677 55159 9735 55165
rect 9950 55156 9956 55168
rect 10008 55196 10014 55208
rect 10137 55199 10195 55205
rect 10137 55196 10149 55199
rect 10008 55168 10149 55196
rect 10008 55156 10014 55168
rect 10137 55165 10149 55168
rect 10183 55165 10195 55199
rect 10137 55159 10195 55165
rect 10870 55156 10876 55208
rect 10928 55196 10934 55208
rect 11808 55205 11836 55236
rect 12066 55224 12072 55236
rect 12124 55224 12130 55276
rect 13814 55224 13820 55276
rect 13872 55264 13878 55276
rect 13909 55267 13967 55273
rect 13909 55264 13921 55267
rect 13872 55236 13921 55264
rect 13872 55224 13878 55236
rect 13909 55233 13921 55236
rect 13955 55264 13967 55267
rect 14936 55264 14964 55372
rect 16298 55360 16304 55372
rect 16356 55360 16362 55412
rect 17126 55360 17132 55412
rect 17184 55400 17190 55412
rect 17221 55403 17279 55409
rect 17221 55400 17233 55403
rect 17184 55372 17233 55400
rect 17184 55360 17190 55372
rect 17221 55369 17233 55372
rect 17267 55369 17279 55403
rect 17221 55363 17279 55369
rect 13955 55236 14964 55264
rect 15105 55267 15163 55273
rect 13955 55233 13967 55236
rect 13909 55227 13967 55233
rect 15105 55233 15117 55267
rect 15151 55264 15163 55267
rect 15151 55236 15608 55264
rect 15151 55233 15163 55236
rect 15105 55227 15163 55233
rect 11057 55199 11115 55205
rect 11057 55196 11069 55199
rect 10928 55168 11069 55196
rect 10928 55156 10934 55168
rect 11057 55165 11069 55168
rect 11103 55165 11115 55199
rect 11057 55159 11115 55165
rect 11793 55199 11851 55205
rect 11793 55165 11805 55199
rect 11839 55165 11851 55199
rect 11793 55159 11851 55165
rect 11885 55199 11943 55205
rect 11885 55165 11897 55199
rect 11931 55196 11943 55199
rect 11974 55196 11980 55208
rect 11931 55168 11980 55196
rect 11931 55165 11943 55168
rect 11885 55159 11943 55165
rect 7484 55100 8248 55128
rect 2222 55020 2228 55072
rect 2280 55060 2286 55072
rect 3145 55063 3203 55069
rect 3145 55060 3157 55063
rect 2280 55032 3157 55060
rect 2280 55020 2286 55032
rect 3145 55029 3157 55032
rect 3191 55029 3203 55063
rect 4430 55060 4436 55072
rect 4391 55032 4436 55060
rect 3145 55023 3203 55029
rect 4430 55020 4436 55032
rect 4488 55060 4494 55072
rect 4798 55060 4804 55072
rect 4488 55032 4804 55060
rect 4488 55020 4494 55032
rect 4798 55020 4804 55032
rect 4856 55020 4862 55072
rect 7282 55060 7288 55072
rect 7243 55032 7288 55060
rect 7282 55020 7288 55032
rect 7340 55060 7346 55072
rect 8404 55060 8432 55156
rect 10965 55131 11023 55137
rect 10965 55097 10977 55131
rect 11011 55128 11023 55131
rect 11900 55128 11928 55159
rect 11974 55156 11980 55168
rect 12032 55156 12038 55208
rect 12253 55199 12311 55205
rect 12253 55165 12265 55199
rect 12299 55165 12311 55199
rect 12253 55159 12311 55165
rect 14185 55199 14243 55205
rect 14185 55165 14197 55199
rect 14231 55165 14243 55199
rect 14366 55196 14372 55208
rect 14327 55168 14372 55196
rect 14185 55159 14243 55165
rect 11011 55100 11928 55128
rect 11011 55097 11023 55100
rect 10965 55091 11023 55097
rect 7340 55032 8432 55060
rect 7340 55020 7346 55032
rect 9582 55020 9588 55072
rect 9640 55060 9646 55072
rect 9861 55063 9919 55069
rect 9861 55060 9873 55063
rect 9640 55032 9873 55060
rect 9640 55020 9646 55032
rect 9861 55029 9873 55032
rect 9907 55029 9919 55063
rect 9861 55023 9919 55029
rect 11422 55020 11428 55072
rect 11480 55060 11486 55072
rect 11606 55060 11612 55072
rect 11480 55032 11612 55060
rect 11480 55020 11486 55032
rect 11606 55020 11612 55032
rect 11664 55020 11670 55072
rect 11882 55020 11888 55072
rect 11940 55060 11946 55072
rect 12268 55060 12296 55159
rect 13262 55088 13268 55140
rect 13320 55128 13326 55140
rect 13357 55131 13415 55137
rect 13357 55128 13369 55131
rect 13320 55100 13369 55128
rect 13320 55088 13326 55100
rect 13357 55097 13369 55100
rect 13403 55097 13415 55131
rect 14200 55128 14228 55159
rect 14366 55156 14372 55168
rect 14424 55156 14430 55208
rect 15289 55199 15347 55205
rect 15289 55165 15301 55199
rect 15335 55196 15347 55199
rect 15378 55196 15384 55208
rect 15335 55168 15384 55196
rect 15335 55165 15347 55168
rect 15289 55159 15347 55165
rect 15378 55156 15384 55168
rect 15436 55156 15442 55208
rect 15580 55205 15608 55236
rect 17402 55224 17408 55276
rect 17460 55264 17466 55276
rect 17589 55267 17647 55273
rect 17589 55264 17601 55267
rect 17460 55236 17601 55264
rect 17460 55224 17466 55236
rect 17589 55233 17601 55236
rect 17635 55233 17647 55267
rect 17589 55227 17647 55233
rect 15565 55199 15623 55205
rect 15565 55165 15577 55199
rect 15611 55196 15623 55199
rect 18138 55196 18144 55208
rect 15611 55168 18144 55196
rect 15611 55165 15623 55168
rect 15565 55159 15623 55165
rect 18138 55156 18144 55168
rect 18196 55156 18202 55208
rect 14200 55100 14780 55128
rect 13357 55091 13415 55097
rect 14752 55072 14780 55100
rect 12802 55060 12808 55072
rect 11940 55032 12296 55060
rect 12763 55032 12808 55060
rect 11940 55020 11946 55032
rect 12802 55020 12808 55032
rect 12860 55020 12866 55072
rect 14734 55060 14740 55072
rect 14695 55032 14740 55060
rect 14734 55020 14740 55032
rect 14792 55020 14798 55072
rect 16669 55063 16727 55069
rect 16669 55029 16681 55063
rect 16715 55060 16727 55063
rect 16758 55060 16764 55072
rect 16715 55032 16764 55060
rect 16715 55029 16727 55032
rect 16669 55023 16727 55029
rect 16758 55020 16764 55032
rect 16816 55020 16822 55072
rect 1104 54970 18860 54992
rect 1104 54918 7648 54970
rect 7700 54918 7712 54970
rect 7764 54918 7776 54970
rect 7828 54918 7840 54970
rect 7892 54918 14315 54970
rect 14367 54918 14379 54970
rect 14431 54918 14443 54970
rect 14495 54918 14507 54970
rect 14559 54918 18860 54970
rect 1104 54896 18860 54918
rect 4709 54859 4767 54865
rect 4709 54825 4721 54859
rect 4755 54856 4767 54859
rect 4890 54856 4896 54868
rect 4755 54828 4896 54856
rect 4755 54825 4767 54828
rect 4709 54819 4767 54825
rect 4890 54816 4896 54828
rect 4948 54816 4954 54868
rect 11790 54856 11796 54868
rect 11751 54828 11796 54856
rect 11790 54816 11796 54828
rect 11848 54816 11854 54868
rect 12710 54816 12716 54868
rect 12768 54856 12774 54868
rect 12894 54856 12900 54868
rect 12768 54828 12900 54856
rect 12768 54816 12774 54828
rect 12894 54816 12900 54828
rect 12952 54816 12958 54868
rect 13173 54859 13231 54865
rect 13173 54825 13185 54859
rect 13219 54856 13231 54859
rect 13814 54856 13820 54868
rect 13219 54828 13820 54856
rect 13219 54825 13231 54828
rect 13173 54819 13231 54825
rect 13814 54816 13820 54828
rect 13872 54816 13878 54868
rect 9766 54748 9772 54800
rect 9824 54788 9830 54800
rect 9824 54760 9904 54788
rect 9824 54748 9830 54760
rect 2406 54720 2412 54732
rect 2367 54692 2412 54720
rect 2406 54680 2412 54692
rect 2464 54680 2470 54732
rect 2866 54720 2872 54732
rect 2827 54692 2872 54720
rect 2866 54680 2872 54692
rect 2924 54680 2930 54732
rect 5534 54720 5540 54732
rect 5495 54692 5540 54720
rect 5534 54680 5540 54692
rect 5592 54680 5598 54732
rect 7193 54723 7251 54729
rect 7193 54689 7205 54723
rect 7239 54720 7251 54723
rect 7929 54723 7987 54729
rect 7929 54720 7941 54723
rect 7239 54692 7941 54720
rect 7239 54689 7251 54692
rect 7193 54683 7251 54689
rect 7929 54689 7941 54692
rect 7975 54720 7987 54723
rect 8202 54720 8208 54732
rect 7975 54692 8208 54720
rect 7975 54689 7987 54692
rect 7929 54683 7987 54689
rect 8202 54680 8208 54692
rect 8260 54680 8266 54732
rect 8386 54680 8392 54732
rect 8444 54720 8450 54732
rect 8846 54720 8852 54732
rect 8444 54692 8852 54720
rect 8444 54680 8450 54692
rect 8846 54680 8852 54692
rect 8904 54680 8910 54732
rect 9030 54680 9036 54732
rect 9088 54720 9094 54732
rect 9876 54729 9904 54760
rect 16500 54760 16896 54788
rect 9217 54723 9275 54729
rect 9217 54720 9229 54723
rect 9088 54692 9229 54720
rect 9088 54680 9094 54692
rect 9217 54689 9229 54692
rect 9263 54689 9275 54723
rect 9217 54683 9275 54689
rect 9861 54723 9919 54729
rect 9861 54689 9873 54723
rect 9907 54689 9919 54723
rect 9861 54683 9919 54689
rect 10778 54680 10784 54732
rect 10836 54720 10842 54732
rect 10965 54723 11023 54729
rect 10965 54720 10977 54723
rect 10836 54692 10977 54720
rect 10836 54680 10842 54692
rect 10965 54689 10977 54692
rect 11011 54689 11023 54723
rect 10965 54683 11023 54689
rect 13078 54680 13084 54732
rect 13136 54720 13142 54732
rect 13265 54723 13323 54729
rect 13265 54720 13277 54723
rect 13136 54692 13277 54720
rect 13136 54680 13142 54692
rect 13265 54689 13277 54692
rect 13311 54689 13323 54723
rect 16500 54720 16528 54760
rect 16868 54732 16896 54760
rect 13265 54683 13323 54689
rect 13464 54692 16528 54720
rect 16577 54723 16635 54729
rect 7282 54652 7288 54664
rect 7243 54624 7288 54652
rect 7282 54612 7288 54624
rect 7340 54612 7346 54664
rect 9490 54652 9496 54664
rect 9451 54624 9496 54652
rect 9490 54612 9496 54624
rect 9548 54612 9554 54664
rect 10594 54612 10600 54664
rect 10652 54652 10658 54664
rect 10873 54655 10931 54661
rect 10873 54652 10885 54655
rect 10652 54624 10885 54652
rect 10652 54612 10658 54624
rect 10873 54621 10885 54624
rect 10919 54621 10931 54655
rect 11422 54652 11428 54664
rect 11383 54624 11428 54652
rect 10873 54615 10931 54621
rect 11422 54612 11428 54624
rect 11480 54612 11486 54664
rect 13464 54652 13492 54692
rect 16577 54689 16589 54723
rect 16623 54689 16635 54723
rect 16850 54720 16856 54732
rect 16763 54692 16856 54720
rect 16577 54683 16635 54689
rect 13280 54624 13492 54652
rect 13541 54655 13599 54661
rect 13280 54596 13308 54624
rect 13541 54621 13553 54655
rect 13587 54652 13599 54655
rect 13722 54652 13728 54664
rect 13587 54624 13728 54652
rect 13587 54621 13599 54624
rect 13541 54615 13599 54621
rect 13722 54612 13728 54624
rect 13780 54612 13786 54664
rect 16114 54652 16120 54664
rect 16075 54624 16120 54652
rect 16114 54612 16120 54624
rect 16172 54612 16178 54664
rect 16592 54652 16620 54683
rect 16850 54680 16856 54692
rect 16908 54680 16914 54732
rect 17126 54652 17132 54664
rect 16592 54624 17132 54652
rect 17126 54612 17132 54624
rect 17184 54612 17190 54664
rect 1486 54544 1492 54596
rect 1544 54584 1550 54596
rect 1673 54587 1731 54593
rect 1673 54584 1685 54587
rect 1544 54556 1685 54584
rect 1544 54544 1550 54556
rect 1673 54553 1685 54556
rect 1719 54584 1731 54587
rect 2317 54587 2375 54593
rect 2317 54584 2329 54587
rect 1719 54556 2329 54584
rect 1719 54553 1731 54556
rect 1673 54547 1731 54553
rect 2317 54553 2329 54556
rect 2363 54553 2375 54587
rect 2317 54547 2375 54553
rect 5077 54587 5135 54593
rect 5077 54553 5089 54587
rect 5123 54584 5135 54587
rect 5810 54584 5816 54596
rect 5123 54556 5816 54584
rect 5123 54553 5135 54556
rect 5077 54547 5135 54553
rect 5810 54544 5816 54556
rect 5868 54544 5874 54596
rect 6914 54584 6920 54596
rect 6380 54556 6920 54584
rect 6380 54528 6408 54556
rect 6914 54544 6920 54556
rect 6972 54544 6978 54596
rect 12161 54587 12219 54593
rect 12161 54553 12173 54587
rect 12207 54584 12219 54587
rect 12894 54584 12900 54596
rect 12207 54556 12900 54584
rect 12207 54553 12219 54556
rect 12161 54547 12219 54553
rect 12894 54544 12900 54556
rect 12952 54544 12958 54596
rect 13262 54544 13268 54596
rect 13320 54544 13326 54596
rect 15381 54587 15439 54593
rect 15381 54553 15393 54587
rect 15427 54584 15439 54587
rect 16390 54584 16396 54596
rect 15427 54556 16396 54584
rect 15427 54553 15439 54556
rect 15381 54547 15439 54553
rect 16390 54544 16396 54556
rect 16448 54544 16454 54596
rect 16942 54584 16948 54596
rect 16903 54556 16948 54584
rect 16942 54544 16948 54556
rect 17000 54544 17006 54596
rect 1762 54476 1768 54528
rect 1820 54516 1826 54528
rect 1949 54519 2007 54525
rect 1949 54516 1961 54519
rect 1820 54488 1961 54516
rect 1820 54476 1826 54488
rect 1949 54485 1961 54488
rect 1995 54485 2007 54519
rect 1949 54479 2007 54485
rect 4062 54476 4068 54528
rect 4120 54516 4126 54528
rect 4249 54519 4307 54525
rect 4249 54516 4261 54519
rect 4120 54488 4261 54516
rect 4120 54476 4126 54488
rect 4249 54485 4261 54488
rect 4295 54485 4307 54519
rect 4249 54479 4307 54485
rect 5629 54519 5687 54525
rect 5629 54485 5641 54519
rect 5675 54516 5687 54519
rect 5718 54516 5724 54528
rect 5675 54488 5724 54516
rect 5675 54485 5687 54488
rect 5629 54479 5687 54485
rect 5718 54476 5724 54488
rect 5776 54476 5782 54528
rect 6273 54519 6331 54525
rect 6273 54485 6285 54519
rect 6319 54516 6331 54519
rect 6362 54516 6368 54528
rect 6319 54488 6368 54516
rect 6319 54485 6331 54488
rect 6273 54479 6331 54485
rect 6362 54476 6368 54488
rect 6420 54476 6426 54528
rect 6641 54519 6699 54525
rect 6641 54485 6653 54519
rect 6687 54516 6699 54519
rect 6730 54516 6736 54528
rect 6687 54488 6736 54516
rect 6687 54485 6699 54488
rect 6641 54479 6699 54485
rect 6730 54476 6736 54488
rect 6788 54476 6794 54528
rect 8294 54516 8300 54528
rect 8255 54488 8300 54516
rect 8294 54476 8300 54488
rect 8352 54516 8358 54528
rect 8570 54516 8576 54528
rect 8352 54488 8576 54516
rect 8352 54476 8358 54488
rect 8570 54476 8576 54488
rect 8628 54476 8634 54528
rect 8757 54519 8815 54525
rect 8757 54485 8769 54519
rect 8803 54516 8815 54519
rect 9030 54516 9036 54528
rect 8803 54488 9036 54516
rect 8803 54485 8815 54488
rect 8757 54479 8815 54485
rect 9030 54476 9036 54488
rect 9088 54476 9094 54528
rect 9490 54476 9496 54528
rect 9548 54516 9554 54528
rect 9766 54516 9772 54528
rect 9548 54488 9772 54516
rect 9548 54476 9554 54488
rect 9766 54476 9772 54488
rect 9824 54476 9830 54528
rect 10505 54519 10563 54525
rect 10505 54485 10517 54519
rect 10551 54516 10563 54519
rect 10870 54516 10876 54528
rect 10551 54488 10876 54516
rect 10551 54485 10563 54488
rect 10505 54479 10563 54485
rect 10870 54476 10876 54488
rect 10928 54476 10934 54528
rect 12618 54516 12624 54528
rect 12579 54488 12624 54516
rect 12618 54476 12624 54488
rect 12676 54476 12682 54528
rect 13446 54476 13452 54528
rect 13504 54516 13510 54528
rect 14645 54519 14703 54525
rect 14645 54516 14657 54519
rect 13504 54488 14657 54516
rect 13504 54476 13510 54488
rect 14645 54485 14657 54488
rect 14691 54485 14703 54519
rect 14645 54479 14703 54485
rect 15749 54519 15807 54525
rect 15749 54485 15761 54519
rect 15795 54516 15807 54519
rect 15930 54516 15936 54528
rect 15795 54488 15936 54516
rect 15795 54485 15807 54488
rect 15749 54479 15807 54485
rect 15930 54476 15936 54488
rect 15988 54476 15994 54528
rect 1104 54426 18860 54448
rect 1104 54374 4315 54426
rect 4367 54374 4379 54426
rect 4431 54374 4443 54426
rect 4495 54374 4507 54426
rect 4559 54374 10982 54426
rect 11034 54374 11046 54426
rect 11098 54374 11110 54426
rect 11162 54374 11174 54426
rect 11226 54374 17648 54426
rect 17700 54374 17712 54426
rect 17764 54374 17776 54426
rect 17828 54374 17840 54426
rect 17892 54374 18860 54426
rect 1104 54352 18860 54374
rect 2866 54312 2872 54324
rect 2827 54284 2872 54312
rect 2866 54272 2872 54284
rect 2924 54272 2930 54324
rect 5353 54315 5411 54321
rect 5353 54281 5365 54315
rect 5399 54312 5411 54315
rect 5534 54312 5540 54324
rect 5399 54284 5540 54312
rect 5399 54281 5411 54284
rect 5353 54275 5411 54281
rect 5534 54272 5540 54284
rect 5592 54272 5598 54324
rect 5721 54315 5779 54321
rect 5721 54281 5733 54315
rect 5767 54312 5779 54315
rect 6178 54312 6184 54324
rect 5767 54284 6184 54312
rect 5767 54281 5779 54284
rect 5721 54275 5779 54281
rect 6178 54272 6184 54284
rect 6236 54272 6242 54324
rect 9214 54272 9220 54324
rect 9272 54312 9278 54324
rect 9401 54315 9459 54321
rect 9401 54312 9413 54315
rect 9272 54284 9413 54312
rect 9272 54272 9278 54284
rect 9401 54281 9413 54284
rect 9447 54281 9459 54315
rect 9401 54275 9459 54281
rect 6730 54204 6736 54256
rect 6788 54244 6794 54256
rect 6825 54247 6883 54253
rect 6825 54244 6837 54247
rect 6788 54216 6837 54244
rect 6788 54204 6794 54216
rect 6825 54213 6837 54216
rect 6871 54213 6883 54247
rect 6825 54207 6883 54213
rect 1578 54176 1584 54188
rect 1539 54148 1584 54176
rect 1578 54136 1584 54148
rect 1636 54136 1642 54188
rect 1670 54136 1676 54188
rect 1728 54176 1734 54188
rect 2222 54176 2228 54188
rect 1728 54148 2228 54176
rect 1728 54136 1734 54148
rect 2222 54136 2228 54148
rect 2280 54176 2286 54188
rect 2409 54179 2467 54185
rect 2409 54176 2421 54179
rect 2280 54148 2421 54176
rect 2280 54136 2286 54148
rect 2409 54145 2421 54148
rect 2455 54145 2467 54179
rect 2409 54139 2467 54145
rect 6914 54136 6920 54188
rect 6972 54176 6978 54188
rect 8294 54176 8300 54188
rect 6972 54148 8300 54176
rect 6972 54136 6978 54148
rect 1486 54108 1492 54120
rect 1447 54080 1492 54108
rect 1486 54068 1492 54080
rect 1544 54068 1550 54120
rect 1762 54068 1768 54120
rect 1820 54108 1826 54120
rect 2317 54111 2375 54117
rect 2317 54108 2329 54111
rect 1820 54080 2329 54108
rect 1820 54068 1826 54080
rect 2317 54077 2329 54080
rect 2363 54077 2375 54111
rect 2317 54071 2375 54077
rect 3510 54068 3516 54120
rect 3568 54068 3574 54120
rect 3881 54111 3939 54117
rect 3881 54077 3893 54111
rect 3927 54108 3939 54111
rect 4249 54111 4307 54117
rect 4249 54108 4261 54111
rect 3927 54080 4261 54108
rect 3927 54077 3939 54080
rect 3881 54071 3939 54077
rect 4249 54077 4261 54080
rect 4295 54108 4307 54111
rect 4706 54108 4712 54120
rect 4295 54080 4712 54108
rect 4295 54077 4307 54080
rect 4249 54071 4307 54077
rect 4706 54068 4712 54080
rect 4764 54068 4770 54120
rect 6089 54111 6147 54117
rect 6089 54077 6101 54111
rect 6135 54108 6147 54111
rect 6178 54108 6184 54120
rect 6135 54080 6184 54108
rect 6135 54077 6147 54080
rect 6089 54071 6147 54077
rect 6178 54068 6184 54080
rect 6236 54068 6242 54120
rect 6365 54111 6423 54117
rect 6365 54077 6377 54111
rect 6411 54108 6423 54111
rect 6454 54108 6460 54120
rect 6411 54080 6460 54108
rect 6411 54077 6423 54080
rect 6365 54071 6423 54077
rect 6454 54068 6460 54080
rect 6512 54068 6518 54120
rect 6641 54111 6699 54117
rect 6641 54077 6653 54111
rect 6687 54108 6699 54111
rect 7101 54111 7159 54117
rect 7101 54108 7113 54111
rect 6687 54080 7113 54108
rect 6687 54077 6699 54080
rect 6641 54071 6699 54077
rect 7101 54077 7113 54080
rect 7147 54108 7159 54111
rect 7834 54108 7840 54120
rect 7147 54080 7840 54108
rect 7147 54077 7159 54080
rect 7101 54071 7159 54077
rect 7834 54068 7840 54080
rect 7892 54068 7898 54120
rect 8128 54117 8156 54148
rect 8294 54136 8300 54148
rect 8352 54136 8358 54188
rect 9416 54176 9444 54275
rect 10778 54272 10784 54324
rect 10836 54312 10842 54324
rect 11425 54315 11483 54321
rect 11425 54312 11437 54315
rect 10836 54284 11437 54312
rect 10836 54272 10842 54284
rect 11425 54281 11437 54284
rect 11471 54281 11483 54315
rect 11425 54275 11483 54281
rect 11974 54272 11980 54324
rect 12032 54312 12038 54324
rect 12526 54312 12532 54324
rect 12032 54284 12532 54312
rect 12032 54272 12038 54284
rect 12526 54272 12532 54284
rect 12584 54272 12590 54324
rect 16850 54272 16856 54324
rect 16908 54312 16914 54324
rect 17773 54315 17831 54321
rect 17773 54312 17785 54315
rect 16908 54284 17785 54312
rect 16908 54272 16914 54284
rect 17773 54281 17785 54284
rect 17819 54281 17831 54315
rect 17773 54275 17831 54281
rect 9766 54204 9772 54256
rect 9824 54244 9830 54256
rect 10134 54244 10140 54256
rect 9824 54216 10140 54244
rect 9824 54204 9830 54216
rect 10134 54204 10140 54216
rect 10192 54204 10198 54256
rect 10318 54204 10324 54256
rect 10376 54244 10382 54256
rect 10505 54247 10563 54253
rect 10505 54244 10517 54247
rect 10376 54216 10517 54244
rect 10376 54204 10382 54216
rect 10505 54213 10517 54216
rect 10551 54213 10563 54247
rect 10505 54207 10563 54213
rect 9861 54179 9919 54185
rect 9861 54176 9873 54179
rect 9416 54148 9873 54176
rect 9861 54145 9873 54148
rect 9907 54145 9919 54179
rect 12526 54176 12532 54188
rect 12487 54148 12532 54176
rect 9861 54139 9919 54145
rect 12526 54136 12532 54148
rect 12584 54136 12590 54188
rect 14001 54179 14059 54185
rect 14001 54145 14013 54179
rect 14047 54176 14059 54179
rect 15838 54176 15844 54188
rect 14047 54148 15332 54176
rect 15799 54148 15844 54176
rect 14047 54145 14059 54148
rect 14001 54139 14059 54145
rect 15304 54120 15332 54148
rect 15838 54136 15844 54148
rect 15896 54136 15902 54188
rect 7929 54111 7987 54117
rect 7929 54077 7941 54111
rect 7975 54077 7987 54111
rect 7929 54071 7987 54077
rect 8113 54111 8171 54117
rect 8113 54077 8125 54111
rect 8159 54077 8171 54111
rect 8113 54071 8171 54077
rect 3528 54040 3556 54068
rect 4065 54043 4123 54049
rect 4065 54040 4077 54043
rect 3528 54012 4077 54040
rect 4065 54009 4077 54012
rect 4111 54040 4123 54043
rect 4522 54040 4528 54052
rect 4111 54012 4528 54040
rect 4111 54009 4123 54012
rect 4065 54003 4123 54009
rect 4522 54000 4528 54012
rect 4580 54040 4586 54052
rect 4893 54043 4951 54049
rect 4893 54040 4905 54043
rect 4580 54012 4905 54040
rect 4580 54000 4586 54012
rect 4893 54009 4905 54012
rect 4939 54009 4951 54043
rect 4893 54003 4951 54009
rect 7561 54043 7619 54049
rect 7561 54009 7573 54043
rect 7607 54040 7619 54043
rect 7944 54040 7972 54071
rect 8386 54068 8392 54120
rect 8444 54108 8450 54120
rect 8481 54111 8539 54117
rect 8481 54108 8493 54111
rect 8444 54080 8493 54108
rect 8444 54068 8450 54080
rect 8481 54077 8493 54080
rect 8527 54077 8539 54111
rect 8481 54071 8539 54077
rect 9125 54111 9183 54117
rect 9125 54077 9137 54111
rect 9171 54108 9183 54111
rect 9490 54108 9496 54120
rect 9171 54080 9496 54108
rect 9171 54077 9183 54080
rect 9125 54071 9183 54077
rect 9490 54068 9496 54080
rect 9548 54068 9554 54120
rect 9674 54068 9680 54120
rect 9732 54108 9738 54120
rect 10045 54111 10103 54117
rect 10045 54108 10057 54111
rect 9732 54080 10057 54108
rect 9732 54068 9738 54080
rect 10045 54077 10057 54080
rect 10091 54077 10103 54111
rect 10045 54071 10103 54077
rect 10134 54068 10140 54120
rect 10192 54108 10198 54120
rect 10505 54111 10563 54117
rect 10505 54108 10517 54111
rect 10192 54080 10517 54108
rect 10192 54068 10198 54080
rect 10505 54077 10517 54080
rect 10551 54077 10563 54111
rect 10505 54071 10563 54077
rect 11698 54068 11704 54120
rect 11756 54108 11762 54120
rect 11793 54111 11851 54117
rect 11793 54108 11805 54111
rect 11756 54080 11805 54108
rect 11756 54068 11762 54080
rect 11793 54077 11805 54080
rect 11839 54077 11851 54111
rect 11793 54071 11851 54077
rect 11882 54068 11888 54120
rect 11940 54108 11946 54120
rect 12069 54111 12127 54117
rect 12069 54108 12081 54111
rect 11940 54080 12081 54108
rect 11940 54068 11946 54080
rect 12069 54077 12081 54080
rect 12115 54077 12127 54111
rect 12069 54071 12127 54077
rect 12158 54068 12164 54120
rect 12216 54108 12222 54120
rect 12342 54108 12348 54120
rect 12216 54080 12348 54108
rect 12216 54068 12222 54080
rect 12342 54068 12348 54080
rect 12400 54068 12406 54120
rect 12618 54108 12624 54120
rect 12579 54080 12624 54108
rect 12618 54068 12624 54080
rect 12676 54068 12682 54120
rect 12894 54108 12900 54120
rect 12855 54080 12900 54108
rect 12894 54068 12900 54080
rect 12952 54068 12958 54120
rect 14090 54108 14096 54120
rect 14051 54080 14096 54108
rect 14090 54068 14096 54080
rect 14148 54108 14154 54120
rect 14553 54111 14611 54117
rect 14553 54108 14565 54111
rect 14148 54080 14565 54108
rect 14148 54068 14154 54080
rect 14553 54077 14565 54080
rect 14599 54077 14611 54111
rect 15286 54108 15292 54120
rect 15247 54080 15292 54108
rect 14553 54071 14611 54077
rect 15286 54068 15292 54080
rect 15344 54068 15350 54120
rect 15930 54108 15936 54120
rect 15891 54080 15936 54108
rect 15930 54068 15936 54080
rect 15988 54068 15994 54120
rect 16301 54111 16359 54117
rect 16301 54077 16313 54111
rect 16347 54108 16359 54111
rect 16390 54108 16396 54120
rect 16347 54080 16396 54108
rect 16347 54077 16359 54080
rect 16301 54071 16359 54077
rect 16390 54068 16396 54080
rect 16448 54068 16454 54120
rect 16666 54108 16672 54120
rect 16627 54080 16672 54108
rect 16666 54068 16672 54080
rect 16724 54068 16730 54120
rect 8294 54040 8300 54052
rect 7607 54012 8300 54040
rect 7607 54009 7619 54012
rect 7561 54003 7619 54009
rect 8294 54000 8300 54012
rect 8352 54000 8358 54052
rect 4246 53932 4252 53984
rect 4304 53972 4310 53984
rect 4341 53975 4399 53981
rect 4341 53972 4353 53975
rect 4304 53944 4353 53972
rect 4304 53932 4310 53944
rect 4341 53941 4353 53944
rect 4387 53941 4399 53975
rect 6178 53972 6184 53984
rect 6139 53944 6184 53972
rect 4341 53935 4399 53941
rect 6178 53932 6184 53944
rect 6236 53932 6242 53984
rect 8570 53972 8576 53984
rect 8531 53944 8576 53972
rect 8570 53932 8576 53944
rect 8628 53932 8634 53984
rect 10594 53932 10600 53984
rect 10652 53972 10658 53984
rect 11146 53972 11152 53984
rect 10652 53944 11152 53972
rect 10652 53932 10658 53944
rect 11146 53932 11152 53944
rect 11204 53932 11210 53984
rect 11609 53975 11667 53981
rect 11609 53941 11621 53975
rect 11655 53972 11667 53975
rect 12434 53972 12440 53984
rect 11655 53944 12440 53972
rect 11655 53941 11667 53944
rect 11609 53935 11667 53941
rect 12434 53932 12440 53944
rect 12492 53932 12498 53984
rect 13633 53975 13691 53981
rect 13633 53941 13645 53975
rect 13679 53972 13691 53975
rect 13722 53972 13728 53984
rect 13679 53944 13728 53972
rect 13679 53941 13691 53944
rect 13633 53935 13691 53941
rect 13722 53932 13728 53944
rect 13780 53932 13786 53984
rect 13998 53932 14004 53984
rect 14056 53972 14062 53984
rect 14277 53975 14335 53981
rect 14277 53972 14289 53975
rect 14056 53944 14289 53972
rect 14056 53932 14062 53944
rect 14277 53941 14289 53944
rect 14323 53941 14335 53975
rect 15102 53972 15108 53984
rect 15063 53944 15108 53972
rect 14277 53935 14335 53941
rect 15102 53932 15108 53944
rect 15160 53932 15166 53984
rect 16114 53932 16120 53984
rect 16172 53972 16178 53984
rect 17037 53975 17095 53981
rect 17037 53972 17049 53975
rect 16172 53944 17049 53972
rect 16172 53932 16178 53944
rect 17037 53941 17049 53944
rect 17083 53941 17095 53975
rect 17037 53935 17095 53941
rect 17126 53932 17132 53984
rect 17184 53972 17190 53984
rect 17405 53975 17463 53981
rect 17405 53972 17417 53975
rect 17184 53944 17417 53972
rect 17184 53932 17190 53944
rect 17405 53941 17417 53944
rect 17451 53941 17463 53975
rect 17405 53935 17463 53941
rect 1104 53882 18860 53904
rect 1104 53830 7648 53882
rect 7700 53830 7712 53882
rect 7764 53830 7776 53882
rect 7828 53830 7840 53882
rect 7892 53830 14315 53882
rect 14367 53830 14379 53882
rect 14431 53830 14443 53882
rect 14495 53830 14507 53882
rect 14559 53830 18860 53882
rect 1104 53808 18860 53830
rect 1670 53768 1676 53780
rect 1631 53740 1676 53768
rect 1670 53728 1676 53740
rect 1728 53728 1734 53780
rect 5629 53771 5687 53777
rect 5629 53737 5641 53771
rect 5675 53768 5687 53771
rect 6454 53768 6460 53780
rect 5675 53740 6460 53768
rect 5675 53737 5687 53740
rect 5629 53731 5687 53737
rect 6454 53728 6460 53740
rect 6512 53728 6518 53780
rect 8662 53768 8668 53780
rect 8496 53740 8668 53768
rect 2222 53660 2228 53712
rect 2280 53700 2286 53712
rect 2866 53700 2872 53712
rect 2280 53672 2872 53700
rect 2280 53660 2286 53672
rect 2866 53660 2872 53672
rect 2924 53660 2930 53712
rect 4246 53700 4252 53712
rect 3436 53672 4252 53700
rect 3050 53592 3056 53644
rect 3108 53632 3114 53644
rect 3436 53641 3464 53672
rect 4246 53660 4252 53672
rect 4304 53660 4310 53712
rect 4522 53660 4528 53712
rect 4580 53700 4586 53712
rect 4709 53703 4767 53709
rect 4709 53700 4721 53703
rect 4580 53672 4721 53700
rect 4580 53660 4586 53672
rect 4709 53669 4721 53672
rect 4755 53700 4767 53703
rect 5166 53700 5172 53712
rect 4755 53672 5172 53700
rect 4755 53669 4767 53672
rect 4709 53663 4767 53669
rect 5166 53660 5172 53672
rect 5224 53660 5230 53712
rect 5534 53660 5540 53712
rect 5592 53700 5598 53712
rect 5997 53703 6055 53709
rect 5997 53700 6009 53703
rect 5592 53672 6009 53700
rect 5592 53660 5598 53672
rect 5997 53669 6009 53672
rect 6043 53700 6055 53703
rect 8496 53700 8524 53740
rect 8662 53728 8668 53740
rect 8720 53728 8726 53780
rect 9674 53728 9680 53780
rect 9732 53768 9738 53780
rect 9769 53771 9827 53777
rect 9769 53768 9781 53771
rect 9732 53740 9781 53768
rect 9732 53728 9738 53740
rect 9769 53737 9781 53740
rect 9815 53737 9827 53771
rect 9769 53731 9827 53737
rect 11146 53728 11152 53780
rect 11204 53768 11210 53780
rect 11422 53768 11428 53780
rect 11204 53740 11428 53768
rect 11204 53728 11210 53740
rect 11422 53728 11428 53740
rect 11480 53728 11486 53780
rect 12069 53771 12127 53777
rect 12069 53737 12081 53771
rect 12115 53768 12127 53771
rect 12250 53768 12256 53780
rect 12115 53740 12256 53768
rect 12115 53737 12127 53740
rect 12069 53731 12127 53737
rect 12250 53728 12256 53740
rect 12308 53768 12314 53780
rect 12526 53768 12532 53780
rect 12308 53740 12532 53768
rect 12308 53728 12314 53740
rect 12526 53728 12532 53740
rect 12584 53728 12590 53780
rect 14001 53771 14059 53777
rect 14001 53737 14013 53771
rect 14047 53768 14059 53771
rect 14182 53768 14188 53780
rect 14047 53740 14188 53768
rect 14047 53737 14059 53740
rect 14001 53731 14059 53737
rect 14182 53728 14188 53740
rect 14240 53728 14246 53780
rect 9582 53700 9588 53712
rect 6043 53672 8524 53700
rect 8680 53672 9588 53700
rect 6043 53669 6055 53672
rect 5997 53663 6055 53669
rect 3421 53635 3479 53641
rect 3421 53632 3433 53635
rect 3108 53604 3433 53632
rect 3108 53592 3114 53604
rect 3421 53601 3433 53604
rect 3467 53601 3479 53635
rect 3421 53595 3479 53601
rect 3697 53635 3755 53641
rect 3697 53601 3709 53635
rect 3743 53601 3755 53635
rect 4890 53632 4896 53644
rect 4851 53604 4896 53632
rect 3697 53595 3755 53601
rect 2869 53567 2927 53573
rect 2869 53533 2881 53567
rect 2915 53564 2927 53567
rect 3602 53564 3608 53576
rect 2915 53536 3608 53564
rect 2915 53533 2927 53536
rect 2869 53527 2927 53533
rect 3602 53524 3608 53536
rect 3660 53524 3666 53576
rect 3712 53496 3740 53595
rect 4890 53592 4896 53604
rect 4948 53592 4954 53644
rect 5810 53592 5816 53644
rect 5868 53632 5874 53644
rect 6178 53632 6184 53644
rect 5868 53604 6184 53632
rect 5868 53592 5874 53604
rect 6178 53592 6184 53604
rect 6236 53632 6242 53644
rect 8220 53641 8248 53672
rect 8680 53644 8708 53672
rect 9582 53660 9588 53672
rect 9640 53660 9646 53712
rect 10870 53660 10876 53712
rect 10928 53700 10934 53712
rect 10928 53672 11376 53700
rect 10928 53660 10934 53672
rect 6273 53635 6331 53641
rect 6273 53632 6285 53635
rect 6236 53604 6285 53632
rect 6236 53592 6242 53604
rect 6273 53601 6285 53604
rect 6319 53601 6331 53635
rect 6273 53595 6331 53601
rect 7009 53635 7067 53641
rect 7009 53601 7021 53635
rect 7055 53601 7067 53635
rect 7009 53595 7067 53601
rect 8205 53635 8263 53641
rect 8205 53601 8217 53635
rect 8251 53601 8263 53635
rect 8662 53632 8668 53644
rect 8575 53604 8668 53632
rect 8205 53595 8263 53601
rect 3881 53567 3939 53573
rect 3881 53533 3893 53567
rect 3927 53533 3939 53567
rect 3881 53527 3939 53533
rect 2792 53468 3740 53496
rect 2792 53440 2820 53468
rect 2317 53431 2375 53437
rect 2317 53397 2329 53431
rect 2363 53428 2375 53431
rect 2406 53428 2412 53440
rect 2363 53400 2412 53428
rect 2363 53397 2375 53400
rect 2317 53391 2375 53397
rect 2406 53388 2412 53400
rect 2464 53388 2470 53440
rect 2774 53428 2780 53440
rect 2735 53400 2780 53428
rect 2774 53388 2780 53400
rect 2832 53388 2838 53440
rect 3142 53388 3148 53440
rect 3200 53428 3206 53440
rect 3896 53428 3924 53527
rect 5534 53524 5540 53576
rect 5592 53564 5598 53576
rect 6914 53564 6920 53576
rect 5592 53536 6920 53564
rect 5592 53524 5598 53536
rect 6914 53524 6920 53536
rect 6972 53524 6978 53576
rect 7024 53564 7052 53595
rect 8662 53592 8668 53604
rect 8720 53592 8726 53644
rect 8846 53632 8852 53644
rect 8807 53604 8852 53632
rect 8846 53592 8852 53604
rect 8904 53592 8910 53644
rect 9490 53632 9496 53644
rect 9451 53604 9496 53632
rect 9490 53592 9496 53604
rect 9548 53592 9554 53644
rect 10594 53632 10600 53644
rect 10555 53604 10600 53632
rect 10594 53592 10600 53604
rect 10652 53592 10658 53644
rect 10778 53632 10784 53644
rect 10739 53604 10784 53632
rect 10778 53592 10784 53604
rect 10836 53592 10842 53644
rect 11348 53641 11376 53672
rect 12544 53672 13032 53700
rect 11333 53635 11391 53641
rect 11333 53601 11345 53635
rect 11379 53632 11391 53635
rect 11606 53632 11612 53644
rect 11379 53604 11612 53632
rect 11379 53601 11391 53604
rect 11333 53595 11391 53601
rect 11606 53592 11612 53604
rect 11664 53592 11670 53644
rect 12544 53641 12572 53672
rect 12529 53635 12587 53641
rect 12529 53601 12541 53635
rect 12575 53601 12587 53635
rect 12802 53632 12808 53644
rect 12529 53595 12587 53601
rect 12636 53604 12808 53632
rect 8110 53564 8116 53576
rect 7024 53536 8116 53564
rect 8110 53524 8116 53536
rect 8168 53524 8174 53576
rect 9401 53567 9459 53573
rect 9401 53533 9413 53567
rect 9447 53564 9459 53567
rect 10134 53564 10140 53576
rect 9447 53536 10140 53564
rect 9447 53533 9459 53536
rect 9401 53527 9459 53533
rect 10134 53524 10140 53536
rect 10192 53524 10198 53576
rect 11517 53567 11575 53573
rect 11517 53533 11529 53567
rect 11563 53564 11575 53567
rect 11882 53564 11888 53576
rect 11563 53536 11888 53564
rect 11563 53533 11575 53536
rect 11517 53527 11575 53533
rect 11882 53524 11888 53536
rect 11940 53524 11946 53576
rect 12066 53524 12072 53576
rect 12124 53564 12130 53576
rect 12636 53564 12664 53604
rect 12802 53592 12808 53604
rect 12860 53592 12866 53644
rect 12894 53564 12900 53576
rect 12124 53536 12664 53564
rect 12855 53536 12900 53564
rect 12124 53524 12130 53536
rect 12894 53524 12900 53536
rect 12952 53524 12958 53576
rect 4338 53496 4344 53508
rect 4299 53468 4344 53496
rect 4338 53456 4344 53468
rect 4396 53456 4402 53508
rect 7466 53456 7472 53508
rect 7524 53496 7530 53508
rect 7524 53468 7788 53496
rect 7524 53456 7530 53468
rect 4982 53428 4988 53440
rect 3200 53400 3924 53428
rect 4943 53400 4988 53428
rect 3200 53388 3206 53400
rect 4982 53388 4988 53400
rect 5040 53388 5046 53440
rect 6086 53428 6092 53440
rect 6047 53400 6092 53428
rect 6086 53388 6092 53400
rect 6144 53388 6150 53440
rect 6638 53428 6644 53440
rect 6599 53400 6644 53428
rect 6638 53388 6644 53400
rect 6696 53388 6702 53440
rect 7193 53431 7251 53437
rect 7193 53397 7205 53431
rect 7239 53428 7251 53431
rect 7374 53428 7380 53440
rect 7239 53400 7380 53428
rect 7239 53397 7251 53400
rect 7193 53391 7251 53397
rect 7374 53388 7380 53400
rect 7432 53388 7438 53440
rect 7760 53437 7788 53468
rect 9214 53456 9220 53508
rect 9272 53496 9278 53508
rect 9582 53496 9588 53508
rect 9272 53468 9588 53496
rect 9272 53456 9278 53468
rect 9582 53456 9588 53468
rect 9640 53456 9646 53508
rect 12434 53456 12440 53508
rect 12492 53496 12498 53508
rect 12802 53496 12808 53508
rect 12492 53468 12808 53496
rect 12492 53456 12498 53468
rect 12802 53456 12808 53468
rect 12860 53456 12866 53508
rect 7745 53431 7803 53437
rect 7745 53397 7757 53431
rect 7791 53428 7803 53431
rect 8386 53428 8392 53440
rect 7791 53400 8392 53428
rect 7791 53397 7803 53400
rect 7745 53391 7803 53397
rect 8386 53388 8392 53400
rect 8444 53388 8450 53440
rect 10134 53388 10140 53440
rect 10192 53428 10198 53440
rect 10318 53428 10324 53440
rect 10192 53400 10324 53428
rect 10192 53388 10198 53400
rect 10318 53388 10324 53400
rect 10376 53388 10382 53440
rect 12894 53388 12900 53440
rect 12952 53428 12958 53440
rect 13004 53428 13032 53672
rect 13078 53592 13084 53644
rect 13136 53632 13142 53644
rect 13173 53635 13231 53641
rect 13173 53632 13185 53635
rect 13136 53604 13185 53632
rect 13136 53592 13142 53604
rect 13173 53601 13185 53604
rect 13219 53601 13231 53635
rect 13173 53595 13231 53601
rect 14642 53592 14648 53644
rect 14700 53632 14706 53644
rect 15286 53632 15292 53644
rect 14700 53604 15292 53632
rect 14700 53592 14706 53604
rect 15286 53592 15292 53604
rect 15344 53592 15350 53644
rect 15930 53632 15936 53644
rect 15891 53604 15936 53632
rect 15930 53592 15936 53604
rect 15988 53592 15994 53644
rect 16206 53632 16212 53644
rect 16167 53604 16212 53632
rect 16206 53592 16212 53604
rect 16264 53592 16270 53644
rect 16577 53635 16635 53641
rect 16577 53601 16589 53635
rect 16623 53601 16635 53635
rect 16577 53595 16635 53601
rect 16592 53564 16620 53595
rect 16666 53564 16672 53576
rect 15120 53536 16672 53564
rect 15120 53508 15148 53536
rect 16666 53524 16672 53536
rect 16724 53524 16730 53576
rect 14090 53456 14096 53508
rect 14148 53496 14154 53508
rect 14737 53499 14795 53505
rect 14737 53496 14749 53499
rect 14148 53468 14749 53496
rect 14148 53456 14154 53468
rect 14737 53465 14749 53468
rect 14783 53496 14795 53499
rect 15102 53496 15108 53508
rect 14783 53468 15108 53496
rect 14783 53465 14795 53468
rect 14737 53459 14795 53465
rect 15102 53456 15108 53468
rect 15160 53456 15166 53508
rect 12952 53400 13032 53428
rect 14461 53431 14519 53437
rect 12952 53388 12958 53400
rect 14461 53397 14473 53431
rect 14507 53428 14519 53431
rect 14642 53428 14648 53440
rect 14507 53400 14648 53428
rect 14507 53397 14519 53400
rect 14461 53391 14519 53397
rect 14642 53388 14648 53400
rect 14700 53388 14706 53440
rect 16485 53431 16543 53437
rect 16485 53397 16497 53431
rect 16531 53428 16543 53431
rect 16574 53428 16580 53440
rect 16531 53400 16580 53428
rect 16531 53397 16543 53400
rect 16485 53391 16543 53397
rect 16574 53388 16580 53400
rect 16632 53388 16638 53440
rect 17034 53428 17040 53440
rect 16995 53400 17040 53428
rect 17034 53388 17040 53400
rect 17092 53388 17098 53440
rect 1104 53338 18860 53360
rect 1104 53286 4315 53338
rect 4367 53286 4379 53338
rect 4431 53286 4443 53338
rect 4495 53286 4507 53338
rect 4559 53286 10982 53338
rect 11034 53286 11046 53338
rect 11098 53286 11110 53338
rect 11162 53286 11174 53338
rect 11226 53286 17648 53338
rect 17700 53286 17712 53338
rect 17764 53286 17776 53338
rect 17828 53286 17840 53338
rect 17892 53286 18860 53338
rect 1104 53264 18860 53286
rect 2406 53184 2412 53236
rect 2464 53224 2470 53236
rect 2869 53227 2927 53233
rect 2869 53224 2881 53227
rect 2464 53196 2881 53224
rect 2464 53184 2470 53196
rect 2869 53193 2881 53196
rect 2915 53193 2927 53227
rect 2869 53187 2927 53193
rect 3881 53227 3939 53233
rect 3881 53193 3893 53227
rect 3927 53224 3939 53227
rect 4890 53224 4896 53236
rect 3927 53196 4896 53224
rect 3927 53193 3939 53196
rect 3881 53187 3939 53193
rect 4890 53184 4896 53196
rect 4948 53224 4954 53236
rect 5629 53227 5687 53233
rect 5629 53224 5641 53227
rect 4948 53196 5641 53224
rect 4948 53184 4954 53196
rect 5629 53193 5641 53196
rect 5675 53193 5687 53227
rect 5629 53187 5687 53193
rect 6641 53227 6699 53233
rect 6641 53193 6653 53227
rect 6687 53224 6699 53227
rect 8110 53224 8116 53236
rect 6687 53196 8116 53224
rect 6687 53193 6699 53196
rect 6641 53187 6699 53193
rect 8110 53184 8116 53196
rect 8168 53184 8174 53236
rect 8573 53227 8631 53233
rect 8573 53193 8585 53227
rect 8619 53224 8631 53227
rect 8662 53224 8668 53236
rect 8619 53196 8668 53224
rect 8619 53193 8631 53196
rect 8573 53187 8631 53193
rect 8662 53184 8668 53196
rect 8720 53184 8726 53236
rect 8846 53224 8852 53236
rect 8807 53196 8852 53224
rect 8846 53184 8852 53196
rect 8904 53184 8910 53236
rect 9490 53184 9496 53236
rect 9548 53184 9554 53236
rect 9953 53227 10011 53233
rect 9953 53193 9965 53227
rect 9999 53224 10011 53227
rect 10594 53224 10600 53236
rect 9999 53196 10600 53224
rect 9999 53193 10011 53196
rect 9953 53187 10011 53193
rect 10594 53184 10600 53196
rect 10652 53184 10658 53236
rect 11422 53224 11428 53236
rect 11256 53196 11428 53224
rect 6914 53156 6920 53168
rect 6875 53128 6920 53156
rect 6914 53116 6920 53128
rect 6972 53116 6978 53168
rect 7374 53116 7380 53168
rect 7432 53156 7438 53168
rect 8205 53159 8263 53165
rect 8205 53156 8217 53159
rect 7432 53128 8217 53156
rect 7432 53116 7438 53128
rect 8205 53125 8217 53128
rect 8251 53156 8263 53159
rect 9508 53156 9536 53184
rect 11256 53168 11284 53196
rect 11422 53184 11428 53196
rect 11480 53184 11486 53236
rect 17034 53224 17040 53236
rect 12728 53196 17040 53224
rect 8251 53128 9536 53156
rect 8251 53125 8263 53128
rect 8205 53119 8263 53125
rect 11238 53116 11244 53168
rect 11296 53116 11302 53168
rect 11517 53159 11575 53165
rect 11517 53125 11529 53159
rect 11563 53156 11575 53159
rect 11790 53156 11796 53168
rect 11563 53128 11796 53156
rect 11563 53125 11575 53128
rect 11517 53119 11575 53125
rect 1670 53048 1676 53100
rect 1728 53088 1734 53100
rect 1765 53091 1823 53097
rect 1765 53088 1777 53091
rect 1728 53060 1777 53088
rect 1728 53048 1734 53060
rect 1765 53057 1777 53060
rect 1811 53057 1823 53091
rect 1765 53051 1823 53057
rect 6638 53048 6644 53100
rect 6696 53088 6702 53100
rect 7466 53088 7472 53100
rect 6696 53060 7472 53088
rect 6696 53048 6702 53060
rect 7466 53048 7472 53060
rect 7524 53088 7530 53100
rect 7561 53091 7619 53097
rect 7561 53088 7573 53091
rect 7524 53060 7573 53088
rect 7524 53048 7530 53060
rect 7561 53057 7573 53060
rect 7607 53057 7619 53091
rect 7561 53051 7619 53057
rect 9493 53091 9551 53097
rect 9493 53057 9505 53091
rect 9539 53088 9551 53091
rect 10226 53088 10232 53100
rect 9539 53060 10232 53088
rect 9539 53057 9551 53060
rect 9493 53051 9551 53057
rect 10226 53048 10232 53060
rect 10284 53048 10290 53100
rect 11532 53088 11560 53119
rect 11790 53116 11796 53128
rect 11848 53116 11854 53168
rect 12728 53088 12756 53196
rect 17034 53184 17040 53196
rect 17092 53184 17098 53236
rect 13909 53159 13967 53165
rect 13909 53125 13921 53159
rect 13955 53156 13967 53159
rect 14642 53156 14648 53168
rect 13955 53128 14648 53156
rect 13955 53125 13967 53128
rect 13909 53119 13967 53125
rect 14642 53116 14648 53128
rect 14700 53116 14706 53168
rect 13170 53088 13176 53100
rect 10612 53060 11560 53088
rect 12636 53060 12756 53088
rect 13131 53060 13176 53088
rect 1489 53023 1547 53029
rect 1489 52989 1501 53023
rect 1535 53020 1547 53023
rect 2406 53020 2412 53032
rect 1535 52992 2412 53020
rect 1535 52989 1547 52992
rect 1489 52983 1547 52989
rect 2406 52980 2412 52992
rect 2464 53020 2470 53032
rect 4062 53020 4068 53032
rect 2464 52992 4068 53020
rect 2464 52980 2470 52992
rect 4062 52980 4068 52992
rect 4120 53020 4126 53032
rect 4249 53023 4307 53029
rect 4249 53020 4261 53023
rect 4120 52992 4261 53020
rect 4120 52980 4126 52992
rect 4249 52989 4261 52992
rect 4295 52989 4307 53023
rect 4522 53020 4528 53032
rect 4483 52992 4528 53020
rect 4249 52983 4307 52989
rect 4522 52980 4528 52992
rect 4580 52980 4586 53032
rect 6733 53023 6791 53029
rect 6733 53020 6745 53023
rect 6196 52992 6745 53020
rect 3142 52844 3148 52896
rect 3200 52884 3206 52896
rect 3510 52884 3516 52896
rect 3200 52856 3516 52884
rect 3200 52844 3206 52856
rect 3510 52844 3516 52856
rect 3568 52844 3574 52896
rect 4062 52844 4068 52896
rect 4120 52884 4126 52896
rect 5534 52884 5540 52896
rect 4120 52856 5540 52884
rect 4120 52844 4126 52856
rect 5534 52844 5540 52856
rect 5592 52844 5598 52896
rect 5626 52844 5632 52896
rect 5684 52884 5690 52896
rect 6196 52893 6224 52992
rect 6733 52989 6745 52992
rect 6779 53020 6791 53023
rect 7006 53020 7012 53032
rect 6779 52992 7012 53020
rect 6779 52989 6791 52992
rect 6733 52983 6791 52989
rect 7006 52980 7012 52992
rect 7064 52980 7070 53032
rect 7098 52980 7104 53032
rect 7156 53020 7162 53032
rect 10612 53029 10640 53060
rect 7285 53023 7343 53029
rect 7285 53020 7297 53023
rect 7156 52992 7297 53020
rect 7156 52980 7162 52992
rect 7285 52989 7297 52992
rect 7331 52989 7343 53023
rect 7285 52983 7343 52989
rect 10597 53023 10655 53029
rect 10597 52989 10609 53023
rect 10643 52989 10655 53023
rect 10597 52983 10655 52989
rect 10873 53023 10931 53029
rect 10873 52989 10885 53023
rect 10919 53020 10931 53023
rect 11606 53020 11612 53032
rect 10919 52992 11612 53020
rect 10919 52989 10931 52992
rect 10873 52983 10931 52989
rect 6638 52912 6644 52964
rect 6696 52952 6702 52964
rect 6822 52952 6828 52964
rect 6696 52924 6828 52952
rect 6696 52912 6702 52924
rect 6822 52912 6828 52924
rect 6880 52912 6886 52964
rect 9214 52912 9220 52964
rect 9272 52952 9278 52964
rect 10888 52952 10916 52983
rect 11606 52980 11612 52992
rect 11664 52980 11670 53032
rect 11790 52980 11796 53032
rect 11848 53020 11854 53032
rect 12636 53029 12664 53060
rect 13170 53048 13176 53060
rect 13228 53048 13234 53100
rect 14182 53088 14188 53100
rect 13280 53060 14188 53088
rect 11977 53023 12035 53029
rect 11977 53020 11989 53023
rect 11848 52992 11989 53020
rect 11848 52980 11854 52992
rect 11977 52989 11989 52992
rect 12023 52989 12035 53023
rect 11977 52983 12035 52989
rect 12621 53023 12679 53029
rect 12621 52989 12633 53023
rect 12667 52989 12679 53023
rect 12621 52983 12679 52989
rect 12713 53023 12771 53029
rect 12713 52989 12725 53023
rect 12759 52989 12771 53023
rect 12713 52983 12771 52989
rect 11149 52955 11207 52961
rect 11149 52952 11161 52955
rect 9272 52924 10916 52952
rect 10980 52924 11161 52952
rect 9272 52912 9278 52924
rect 6181 52887 6239 52893
rect 6181 52884 6193 52887
rect 5684 52856 6193 52884
rect 5684 52844 5690 52856
rect 6181 52853 6193 52856
rect 6227 52853 6239 52887
rect 6181 52847 6239 52853
rect 6362 52844 6368 52896
rect 6420 52884 6426 52896
rect 6546 52884 6552 52896
rect 6420 52856 6552 52884
rect 6420 52844 6426 52856
rect 6546 52844 6552 52856
rect 6604 52844 6610 52896
rect 7374 52844 7380 52896
rect 7432 52884 7438 52896
rect 8202 52884 8208 52896
rect 7432 52856 8208 52884
rect 7432 52844 7438 52856
rect 8202 52844 8208 52856
rect 8260 52844 8266 52896
rect 10594 52844 10600 52896
rect 10652 52884 10658 52896
rect 10980 52884 11008 52924
rect 11149 52921 11161 52924
rect 11195 52921 11207 52955
rect 11149 52915 11207 52921
rect 11330 52912 11336 52964
rect 11388 52952 11394 52964
rect 11514 52952 11520 52964
rect 11388 52924 11520 52952
rect 11388 52912 11394 52924
rect 11514 52912 11520 52924
rect 11572 52912 11578 52964
rect 10652 52856 11008 52884
rect 11885 52887 11943 52893
rect 10652 52844 10658 52856
rect 11885 52853 11897 52887
rect 11931 52884 11943 52887
rect 12066 52884 12072 52896
rect 11931 52856 12072 52884
rect 11931 52853 11943 52856
rect 11885 52847 11943 52853
rect 12066 52844 12072 52856
rect 12124 52844 12130 52896
rect 12526 52844 12532 52896
rect 12584 52884 12590 52896
rect 12728 52884 12756 52983
rect 13170 52912 13176 52964
rect 13228 52952 13234 52964
rect 13280 52952 13308 53060
rect 14182 53048 14188 53060
rect 14240 53048 14246 53100
rect 14734 53048 14740 53100
rect 14792 53088 14798 53100
rect 15286 53088 15292 53100
rect 14792 53060 15292 53088
rect 14792 53048 14798 53060
rect 15286 53048 15292 53060
rect 15344 53088 15350 53100
rect 15473 53091 15531 53097
rect 15473 53088 15485 53091
rect 15344 53060 15485 53088
rect 15344 53048 15350 53060
rect 15473 53057 15485 53060
rect 15519 53057 15531 53091
rect 17129 53091 17187 53097
rect 17129 53088 17141 53091
rect 15473 53051 15531 53057
rect 15580 53060 17141 53088
rect 15580 53032 15608 53060
rect 17129 53057 17141 53060
rect 17175 53057 17187 53091
rect 17129 53051 17187 53057
rect 14001 53023 14059 53029
rect 14001 52989 14013 53023
rect 14047 53020 14059 53023
rect 14461 53023 14519 53029
rect 14461 53020 14473 53023
rect 14047 52992 14473 53020
rect 14047 52989 14059 52992
rect 14001 52983 14059 52989
rect 14461 52989 14473 52992
rect 14507 53020 14519 53023
rect 14550 53020 14556 53032
rect 14507 52992 14556 53020
rect 14507 52989 14519 52992
rect 14461 52983 14519 52989
rect 14550 52980 14556 52992
rect 14608 52980 14614 53032
rect 15562 53020 15568 53032
rect 15523 52992 15568 53020
rect 15562 52980 15568 52992
rect 15620 52980 15626 53032
rect 15930 53020 15936 53032
rect 15891 52992 15936 53020
rect 15930 52980 15936 52992
rect 15988 52980 15994 53032
rect 16117 53023 16175 53029
rect 16117 52989 16129 53023
rect 16163 52989 16175 53023
rect 16666 53020 16672 53032
rect 16627 52992 16672 53020
rect 16117 52983 16175 52989
rect 13228 52924 13308 52952
rect 13228 52912 13234 52924
rect 15010 52912 15016 52964
rect 15068 52952 15074 52964
rect 15105 52955 15163 52961
rect 15105 52952 15117 52955
rect 15068 52924 15117 52952
rect 15068 52912 15074 52924
rect 15105 52921 15117 52924
rect 15151 52952 15163 52955
rect 16132 52952 16160 52983
rect 16666 52980 16672 52992
rect 16724 52980 16730 53032
rect 17954 53020 17960 53032
rect 17915 52992 17960 53020
rect 17954 52980 17960 52992
rect 18012 52980 18018 53032
rect 15151 52924 16160 52952
rect 15151 52921 15163 52924
rect 15105 52915 15163 52921
rect 12584 52856 12756 52884
rect 12584 52844 12590 52856
rect 13078 52844 13084 52896
rect 13136 52884 13142 52896
rect 13449 52887 13507 52893
rect 13449 52884 13461 52887
rect 13136 52856 13461 52884
rect 13136 52844 13142 52856
rect 13449 52853 13461 52856
rect 13495 52853 13507 52887
rect 14182 52884 14188 52896
rect 14143 52856 14188 52884
rect 13449 52847 13507 52853
rect 14182 52844 14188 52856
rect 14240 52844 14246 52896
rect 15930 52844 15936 52896
rect 15988 52884 15994 52896
rect 17497 52887 17555 52893
rect 17497 52884 17509 52887
rect 15988 52856 17509 52884
rect 15988 52844 15994 52856
rect 17497 52853 17509 52856
rect 17543 52884 17555 52887
rect 17954 52884 17960 52896
rect 17543 52856 17960 52884
rect 17543 52853 17555 52856
rect 17497 52847 17555 52853
rect 17954 52844 17960 52856
rect 18012 52844 18018 52896
rect 1104 52794 18860 52816
rect 1104 52742 7648 52794
rect 7700 52742 7712 52794
rect 7764 52742 7776 52794
rect 7828 52742 7840 52794
rect 7892 52742 14315 52794
rect 14367 52742 14379 52794
rect 14431 52742 14443 52794
rect 14495 52742 14507 52794
rect 14559 52742 18860 52794
rect 1104 52720 18860 52742
rect 2961 52683 3019 52689
rect 2961 52649 2973 52683
rect 3007 52680 3019 52683
rect 3050 52680 3056 52692
rect 3007 52652 3056 52680
rect 3007 52649 3019 52652
rect 2961 52643 3019 52649
rect 3050 52640 3056 52652
rect 3108 52640 3114 52692
rect 3510 52680 3516 52692
rect 3252 52652 3516 52680
rect 1670 52612 1676 52624
rect 1631 52584 1676 52612
rect 1670 52572 1676 52584
rect 1728 52572 1734 52624
rect 3142 52544 3148 52556
rect 3103 52516 3148 52544
rect 3142 52504 3148 52516
rect 3200 52504 3206 52556
rect 3050 52436 3056 52488
rect 3108 52476 3114 52488
rect 3252 52476 3280 52652
rect 3510 52640 3516 52652
rect 3568 52640 3574 52692
rect 4706 52680 4712 52692
rect 4667 52652 4712 52680
rect 4706 52640 4712 52652
rect 4764 52640 4770 52692
rect 5166 52680 5172 52692
rect 5127 52652 5172 52680
rect 5166 52640 5172 52652
rect 5224 52640 5230 52692
rect 5534 52640 5540 52692
rect 5592 52680 5598 52692
rect 5813 52683 5871 52689
rect 5813 52680 5825 52683
rect 5592 52652 5825 52680
rect 5592 52640 5598 52652
rect 5813 52649 5825 52652
rect 5859 52680 5871 52683
rect 6362 52680 6368 52692
rect 5859 52652 6368 52680
rect 5859 52649 5871 52652
rect 5813 52643 5871 52649
rect 6362 52640 6368 52652
rect 6420 52640 6426 52692
rect 7466 52640 7472 52692
rect 7524 52680 7530 52692
rect 7745 52683 7803 52689
rect 7745 52680 7757 52683
rect 7524 52652 7757 52680
rect 7524 52640 7530 52652
rect 7745 52649 7757 52652
rect 7791 52649 7803 52683
rect 7745 52643 7803 52649
rect 9125 52683 9183 52689
rect 9125 52649 9137 52683
rect 9171 52680 9183 52683
rect 9214 52680 9220 52692
rect 9171 52652 9220 52680
rect 9171 52649 9183 52652
rect 9125 52643 9183 52649
rect 9214 52640 9220 52652
rect 9272 52640 9278 52692
rect 9493 52683 9551 52689
rect 9493 52649 9505 52683
rect 9539 52680 9551 52683
rect 10778 52680 10784 52692
rect 9539 52652 10784 52680
rect 9539 52649 9551 52652
rect 9493 52643 9551 52649
rect 10778 52640 10784 52652
rect 10836 52680 10842 52692
rect 12158 52680 12164 52692
rect 10836 52652 12164 52680
rect 10836 52640 10842 52652
rect 12158 52640 12164 52652
rect 12216 52680 12222 52692
rect 16206 52680 16212 52692
rect 12216 52652 16068 52680
rect 16167 52652 16212 52680
rect 12216 52640 12222 52652
rect 4522 52572 4528 52624
rect 4580 52612 4586 52624
rect 5445 52615 5503 52621
rect 5445 52612 5457 52615
rect 4580 52584 5457 52612
rect 4580 52572 4586 52584
rect 5445 52581 5457 52584
rect 5491 52612 5503 52615
rect 8202 52612 8208 52624
rect 5491 52584 8208 52612
rect 5491 52581 5503 52584
rect 5445 52575 5503 52581
rect 5644 52553 5672 52584
rect 8202 52572 8208 52584
rect 8260 52572 8266 52624
rect 11238 52572 11244 52624
rect 11296 52612 11302 52624
rect 11698 52612 11704 52624
rect 11296 52584 11704 52612
rect 11296 52572 11302 52584
rect 11698 52572 11704 52584
rect 11756 52572 11762 52624
rect 5629 52547 5687 52553
rect 5629 52513 5641 52547
rect 5675 52544 5687 52547
rect 7377 52547 7435 52553
rect 5675 52516 5709 52544
rect 5675 52513 5687 52516
rect 5629 52507 5687 52513
rect 7377 52513 7389 52547
rect 7423 52544 7435 52547
rect 8113 52547 8171 52553
rect 7423 52516 7788 52544
rect 7423 52513 7435 52516
rect 7377 52507 7435 52513
rect 3108 52448 3280 52476
rect 3421 52479 3479 52485
rect 3108 52436 3114 52448
rect 3421 52445 3433 52479
rect 3467 52476 3479 52479
rect 3510 52476 3516 52488
rect 3467 52448 3516 52476
rect 3467 52445 3479 52448
rect 3421 52439 3479 52445
rect 3510 52436 3516 52448
rect 3568 52436 3574 52488
rect 6641 52479 6699 52485
rect 6641 52445 6653 52479
rect 6687 52476 6699 52479
rect 7098 52476 7104 52488
rect 6687 52448 7104 52476
rect 6687 52445 6699 52448
rect 6641 52439 6699 52445
rect 7098 52436 7104 52448
rect 7156 52436 7162 52488
rect 7466 52476 7472 52488
rect 7427 52448 7472 52476
rect 7466 52436 7472 52448
rect 7524 52436 7530 52488
rect 7760 52476 7788 52516
rect 8113 52513 8125 52547
rect 8159 52544 8171 52547
rect 8159 52516 8340 52544
rect 8159 52513 8171 52516
rect 8113 52507 8171 52513
rect 8202 52476 8208 52488
rect 7760 52448 8208 52476
rect 8202 52436 8208 52448
rect 8260 52436 8266 52488
rect 8312 52408 8340 52516
rect 8386 52504 8392 52556
rect 8444 52544 8450 52556
rect 8481 52547 8539 52553
rect 8481 52544 8493 52547
rect 8444 52516 8493 52544
rect 8444 52504 8450 52516
rect 8481 52513 8493 52516
rect 8527 52544 8539 52547
rect 8846 52544 8852 52556
rect 8527 52516 8852 52544
rect 8527 52513 8539 52516
rect 8481 52507 8539 52513
rect 8846 52504 8852 52516
rect 8904 52504 8910 52556
rect 9950 52504 9956 52556
rect 10008 52544 10014 52556
rect 10321 52547 10379 52553
rect 10321 52544 10333 52547
rect 10008 52516 10333 52544
rect 10008 52504 10014 52516
rect 10321 52513 10333 52516
rect 10367 52513 10379 52547
rect 10778 52544 10784 52556
rect 10739 52516 10784 52544
rect 10321 52507 10379 52513
rect 10778 52504 10784 52516
rect 10836 52504 10842 52556
rect 10870 52504 10876 52556
rect 10928 52544 10934 52556
rect 11057 52547 11115 52553
rect 11057 52544 11069 52547
rect 10928 52516 11069 52544
rect 10928 52504 10934 52516
rect 11057 52513 11069 52516
rect 11103 52513 11115 52547
rect 11057 52507 11115 52513
rect 11422 52504 11428 52556
rect 11480 52504 11486 52556
rect 13004 52553 13032 52652
rect 13262 52572 13268 52624
rect 13320 52612 13326 52624
rect 13906 52612 13912 52624
rect 13320 52584 13912 52612
rect 13320 52572 13326 52584
rect 13372 52553 13400 52584
rect 13906 52572 13912 52584
rect 13964 52572 13970 52624
rect 12989 52547 13047 52553
rect 12989 52513 13001 52547
rect 13035 52513 13047 52547
rect 12989 52507 13047 52513
rect 13357 52547 13415 52553
rect 13357 52513 13369 52547
rect 13403 52513 13415 52547
rect 13357 52507 13415 52513
rect 13446 52504 13452 52556
rect 13504 52504 13510 52556
rect 14642 52544 14648 52556
rect 14555 52516 14648 52544
rect 14642 52504 14648 52516
rect 14700 52504 14706 52556
rect 15010 52544 15016 52556
rect 14971 52516 15016 52544
rect 15010 52504 15016 52516
rect 15068 52504 15074 52556
rect 15102 52504 15108 52556
rect 15160 52544 15166 52556
rect 15197 52547 15255 52553
rect 15197 52544 15209 52547
rect 15160 52516 15209 52544
rect 15160 52504 15166 52516
rect 15197 52513 15209 52516
rect 15243 52513 15255 52547
rect 15657 52547 15715 52553
rect 15657 52544 15669 52547
rect 15197 52507 15255 52513
rect 15580 52516 15669 52544
rect 10134 52476 10140 52488
rect 10095 52448 10140 52476
rect 10134 52436 10140 52448
rect 10192 52436 10198 52488
rect 8386 52408 8392 52420
rect 8299 52380 8392 52408
rect 8386 52368 8392 52380
rect 8444 52408 8450 52420
rect 8754 52408 8760 52420
rect 8444 52380 8760 52408
rect 8444 52368 8450 52380
rect 8754 52368 8760 52380
rect 8812 52368 8818 52420
rect 10413 52411 10471 52417
rect 10413 52377 10425 52411
rect 10459 52408 10471 52411
rect 10502 52408 10508 52420
rect 10459 52380 10508 52408
rect 10459 52377 10471 52380
rect 10413 52371 10471 52377
rect 10502 52368 10508 52380
rect 10560 52368 10566 52420
rect 2041 52343 2099 52349
rect 2041 52309 2053 52343
rect 2087 52340 2099 52343
rect 2406 52340 2412 52352
rect 2087 52312 2412 52340
rect 2087 52309 2099 52312
rect 2041 52303 2099 52309
rect 2406 52300 2412 52312
rect 2464 52300 2470 52352
rect 6086 52340 6092 52352
rect 6047 52312 6092 52340
rect 6086 52300 6092 52312
rect 6144 52300 6150 52352
rect 9861 52343 9919 52349
rect 9861 52309 9873 52343
rect 9907 52340 9919 52343
rect 9950 52340 9956 52352
rect 9907 52312 9956 52340
rect 9907 52309 9919 52312
rect 9861 52303 9919 52309
rect 9950 52300 9956 52312
rect 10008 52300 10014 52352
rect 11440 52340 11468 52504
rect 11882 52436 11888 52488
rect 11940 52476 11946 52488
rect 12250 52476 12256 52488
rect 11940 52448 12256 52476
rect 11940 52436 11946 52448
rect 12250 52436 12256 52448
rect 12308 52436 12314 52488
rect 12621 52479 12679 52485
rect 12621 52445 12633 52479
rect 12667 52476 12679 52479
rect 12894 52476 12900 52488
rect 12667 52448 12900 52476
rect 12667 52445 12679 52448
rect 12621 52439 12679 52445
rect 12894 52436 12900 52448
rect 12952 52436 12958 52488
rect 13464 52476 13492 52504
rect 13280 52448 13492 52476
rect 14660 52476 14688 52504
rect 15470 52476 15476 52488
rect 14660 52448 15476 52476
rect 13280 52420 13308 52448
rect 15470 52436 15476 52448
rect 15528 52436 15534 52488
rect 11790 52368 11796 52420
rect 11848 52408 11854 52420
rect 11977 52411 12035 52417
rect 11977 52408 11989 52411
rect 11848 52380 11989 52408
rect 11848 52368 11854 52380
rect 11977 52377 11989 52380
rect 12023 52377 12035 52411
rect 11977 52371 12035 52377
rect 13262 52368 13268 52420
rect 13320 52368 13326 52420
rect 13357 52411 13415 52417
rect 13357 52377 13369 52411
rect 13403 52408 13415 52411
rect 13446 52408 13452 52420
rect 13403 52380 13452 52408
rect 13403 52377 13415 52380
rect 13357 52371 13415 52377
rect 13446 52368 13452 52380
rect 13504 52368 13510 52420
rect 14090 52368 14096 52420
rect 14148 52408 14154 52420
rect 14185 52411 14243 52417
rect 14185 52408 14197 52411
rect 14148 52380 14197 52408
rect 14148 52368 14154 52380
rect 14185 52377 14197 52380
rect 14231 52408 14243 52411
rect 15580 52408 15608 52516
rect 15657 52513 15669 52516
rect 15703 52513 15715 52547
rect 15657 52507 15715 52513
rect 14231 52380 15608 52408
rect 16040 52408 16068 52652
rect 16206 52640 16212 52652
rect 16264 52640 16270 52692
rect 16850 52504 16856 52556
rect 16908 52544 16914 52556
rect 16945 52547 17003 52553
rect 16945 52544 16957 52547
rect 16908 52516 16957 52544
rect 16908 52504 16914 52516
rect 16945 52513 16957 52516
rect 16991 52513 17003 52547
rect 16945 52507 17003 52513
rect 17126 52408 17132 52420
rect 16040 52380 17132 52408
rect 14231 52377 14243 52380
rect 14185 52371 14243 52377
rect 17126 52368 17132 52380
rect 17184 52368 17190 52420
rect 12250 52340 12256 52352
rect 11440 52312 12256 52340
rect 12250 52300 12256 52312
rect 12308 52300 12314 52352
rect 13909 52343 13967 52349
rect 13909 52309 13921 52343
rect 13955 52340 13967 52343
rect 14274 52340 14280 52352
rect 13955 52312 14280 52340
rect 13955 52309 13967 52312
rect 13909 52303 13967 52309
rect 14274 52300 14280 52312
rect 14332 52300 14338 52352
rect 14461 52343 14519 52349
rect 14461 52309 14473 52343
rect 14507 52340 14519 52343
rect 14734 52340 14740 52352
rect 14507 52312 14740 52340
rect 14507 52309 14519 52312
rect 14461 52303 14519 52309
rect 14734 52300 14740 52312
rect 14792 52300 14798 52352
rect 15930 52300 15936 52352
rect 15988 52340 15994 52352
rect 16485 52343 16543 52349
rect 16485 52340 16497 52343
rect 15988 52312 16497 52340
rect 15988 52300 15994 52312
rect 16485 52309 16497 52312
rect 16531 52309 16543 52343
rect 16485 52303 16543 52309
rect 1104 52250 18860 52272
rect 1104 52198 4315 52250
rect 4367 52198 4379 52250
rect 4431 52198 4443 52250
rect 4495 52198 4507 52250
rect 4559 52198 10982 52250
rect 11034 52198 11046 52250
rect 11098 52198 11110 52250
rect 11162 52198 11174 52250
rect 11226 52198 17648 52250
rect 17700 52198 17712 52250
rect 17764 52198 17776 52250
rect 17828 52198 17840 52250
rect 17892 52198 18860 52250
rect 1104 52176 18860 52198
rect 3881 52139 3939 52145
rect 3881 52105 3893 52139
rect 3927 52136 3939 52139
rect 5445 52139 5503 52145
rect 3927 52108 5120 52136
rect 3927 52105 3939 52108
rect 3881 52099 3939 52105
rect 3513 52071 3571 52077
rect 3513 52037 3525 52071
rect 3559 52068 3571 52071
rect 3559 52040 4660 52068
rect 3559 52037 3571 52040
rect 3513 52031 3571 52037
rect 4065 52003 4123 52009
rect 4065 51969 4077 52003
rect 4111 52000 4123 52003
rect 4154 52000 4160 52012
rect 4111 51972 4160 52000
rect 4111 51969 4123 51972
rect 4065 51963 4123 51969
rect 4154 51960 4160 51972
rect 4212 51960 4218 52012
rect 4632 52009 4660 52040
rect 4617 52003 4675 52009
rect 4617 51969 4629 52003
rect 4663 52000 4675 52003
rect 4982 52000 4988 52012
rect 4663 51972 4988 52000
rect 4663 51969 4675 51972
rect 4617 51963 4675 51969
rect 4982 51960 4988 51972
rect 5040 51960 5046 52012
rect 5092 52009 5120 52108
rect 5445 52105 5457 52139
rect 5491 52136 5503 52139
rect 6546 52136 6552 52148
rect 5491 52108 6552 52136
rect 5491 52105 5503 52108
rect 5445 52099 5503 52105
rect 6546 52096 6552 52108
rect 6604 52096 6610 52148
rect 8386 52136 8392 52148
rect 8347 52108 8392 52136
rect 8386 52096 8392 52108
rect 8444 52096 8450 52148
rect 8846 52096 8852 52148
rect 8904 52136 8910 52148
rect 9030 52136 9036 52148
rect 8904 52108 9036 52136
rect 8904 52096 8910 52108
rect 9030 52096 9036 52108
rect 9088 52096 9094 52148
rect 10045 52139 10103 52145
rect 10045 52105 10057 52139
rect 10091 52136 10103 52139
rect 10870 52136 10876 52148
rect 10091 52108 10876 52136
rect 10091 52105 10103 52108
rect 10045 52099 10103 52105
rect 10870 52096 10876 52108
rect 10928 52096 10934 52148
rect 11330 52096 11336 52148
rect 11388 52136 11394 52148
rect 13906 52136 13912 52148
rect 11388 52108 13912 52136
rect 11388 52096 11394 52108
rect 13906 52096 13912 52108
rect 13964 52096 13970 52148
rect 13998 52096 14004 52148
rect 14056 52136 14062 52148
rect 14737 52139 14795 52145
rect 14737 52136 14749 52139
rect 14056 52108 14749 52136
rect 14056 52096 14062 52108
rect 14737 52105 14749 52108
rect 14783 52136 14795 52139
rect 15102 52136 15108 52148
rect 14783 52108 15108 52136
rect 14783 52105 14795 52108
rect 14737 52099 14795 52105
rect 15102 52096 15108 52108
rect 15160 52096 15166 52148
rect 16850 52096 16856 52148
rect 16908 52136 16914 52148
rect 17589 52139 17647 52145
rect 17589 52136 17601 52139
rect 16908 52108 17601 52136
rect 16908 52096 16914 52108
rect 17589 52105 17601 52108
rect 17635 52105 17647 52139
rect 17954 52136 17960 52148
rect 17915 52108 17960 52136
rect 17589 52099 17647 52105
rect 17954 52096 17960 52108
rect 18012 52096 18018 52148
rect 6178 52068 6184 52080
rect 6012 52040 6184 52068
rect 5077 52003 5135 52009
rect 5077 51969 5089 52003
rect 5123 52000 5135 52003
rect 5534 52000 5540 52012
rect 5123 51972 5540 52000
rect 5123 51969 5135 51972
rect 5077 51963 5135 51969
rect 5534 51960 5540 51972
rect 5592 51960 5598 52012
rect 6012 52009 6040 52040
rect 6178 52028 6184 52040
rect 6236 52068 6242 52080
rect 6822 52068 6828 52080
rect 6236 52040 6828 52068
rect 6236 52028 6242 52040
rect 6822 52028 6828 52040
rect 6880 52028 6886 52080
rect 7006 52068 7012 52080
rect 6967 52040 7012 52068
rect 7006 52028 7012 52040
rect 7064 52028 7070 52080
rect 7653 52071 7711 52077
rect 7653 52037 7665 52071
rect 7699 52068 7711 52071
rect 8754 52068 8760 52080
rect 7699 52040 8760 52068
rect 7699 52037 7711 52040
rect 7653 52031 7711 52037
rect 8754 52028 8760 52040
rect 8812 52028 8818 52080
rect 11238 52028 11244 52080
rect 11296 52068 11302 52080
rect 11606 52068 11612 52080
rect 11296 52040 11612 52068
rect 11296 52028 11302 52040
rect 11606 52028 11612 52040
rect 11664 52028 11670 52080
rect 13265 52071 13323 52077
rect 13265 52037 13277 52071
rect 13311 52068 13323 52071
rect 13814 52068 13820 52080
rect 13311 52040 13820 52068
rect 13311 52037 13323 52040
rect 13265 52031 13323 52037
rect 13814 52028 13820 52040
rect 13872 52068 13878 52080
rect 13872 52040 14412 52068
rect 13872 52028 13878 52040
rect 5997 52003 6055 52009
rect 5997 51969 6009 52003
rect 6043 51969 6055 52003
rect 5997 51963 6055 51969
rect 9493 52003 9551 52009
rect 9493 51969 9505 52003
rect 9539 52000 9551 52003
rect 12250 52000 12256 52012
rect 9539 51972 10916 52000
rect 9539 51969 9551 51972
rect 9493 51963 9551 51969
rect 10888 51944 10916 51972
rect 12084 51972 12256 52000
rect 4522 51892 4528 51944
rect 4580 51932 4586 51944
rect 4893 51935 4951 51941
rect 4893 51932 4905 51935
rect 4580 51904 4905 51932
rect 4580 51892 4586 51904
rect 4893 51901 4905 51904
rect 4939 51901 4951 51935
rect 6086 51932 6092 51944
rect 5999 51904 6092 51932
rect 4893 51895 4951 51901
rect 6086 51892 6092 51904
rect 6144 51892 6150 51944
rect 6546 51932 6552 51944
rect 6507 51904 6552 51932
rect 6546 51892 6552 51904
rect 6604 51892 6610 51944
rect 6641 51935 6699 51941
rect 6641 51901 6653 51935
rect 6687 51932 6699 51935
rect 8573 51935 8631 51941
rect 6687 51904 6960 51932
rect 6687 51901 6699 51904
rect 6641 51895 6699 51901
rect 4154 51824 4160 51876
rect 4212 51864 4218 51876
rect 5074 51864 5080 51876
rect 4212 51836 5080 51864
rect 4212 51824 4218 51836
rect 5074 51824 5080 51836
rect 5132 51824 5138 51876
rect 6104 51864 6132 51892
rect 6822 51864 6828 51876
rect 6104 51836 6828 51864
rect 6822 51824 6828 51836
rect 6880 51824 6886 51876
rect 2774 51796 2780 51808
rect 2735 51768 2780 51796
rect 2774 51756 2780 51768
rect 2832 51756 2838 51808
rect 3145 51799 3203 51805
rect 3145 51765 3157 51799
rect 3191 51796 3203 51799
rect 4706 51796 4712 51808
rect 3191 51768 4712 51796
rect 3191 51765 3203 51768
rect 3145 51759 3203 51765
rect 4706 51756 4712 51768
rect 4764 51756 4770 51808
rect 4798 51756 4804 51808
rect 4856 51796 4862 51808
rect 5258 51796 5264 51808
rect 4856 51768 5264 51796
rect 4856 51756 4862 51768
rect 5258 51756 5264 51768
rect 5316 51756 5322 51808
rect 5813 51799 5871 51805
rect 5813 51765 5825 51799
rect 5859 51796 5871 51799
rect 6454 51796 6460 51808
rect 5859 51768 6460 51796
rect 5859 51765 5871 51768
rect 5813 51759 5871 51765
rect 6454 51756 6460 51768
rect 6512 51796 6518 51808
rect 6932 51796 6960 51904
rect 8573 51901 8585 51935
rect 8619 51932 8631 51935
rect 9033 51935 9091 51941
rect 9033 51932 9045 51935
rect 8619 51904 9045 51932
rect 8619 51901 8631 51904
rect 8573 51895 8631 51901
rect 9033 51901 9045 51904
rect 9079 51932 9091 51935
rect 9582 51932 9588 51944
rect 9079 51904 9588 51932
rect 9079 51901 9091 51904
rect 9033 51895 9091 51901
rect 9582 51892 9588 51904
rect 9640 51892 9646 51944
rect 9950 51892 9956 51944
rect 10008 51932 10014 51944
rect 10226 51932 10232 51944
rect 10008 51904 10232 51932
rect 10008 51892 10014 51904
rect 10226 51892 10232 51904
rect 10284 51932 10290 51944
rect 10689 51935 10747 51941
rect 10689 51932 10701 51935
rect 10284 51904 10701 51932
rect 10284 51892 10290 51904
rect 10689 51901 10701 51904
rect 10735 51901 10747 51935
rect 10689 51895 10747 51901
rect 10870 51892 10876 51944
rect 10928 51932 10934 51944
rect 11057 51935 11115 51941
rect 11057 51932 11069 51935
rect 10928 51904 11069 51932
rect 10928 51892 10934 51904
rect 11057 51901 11069 51904
rect 11103 51901 11115 51935
rect 11422 51932 11428 51944
rect 11383 51904 11428 51932
rect 11057 51895 11115 51901
rect 11422 51892 11428 51904
rect 11480 51892 11486 51944
rect 12084 51941 12112 51972
rect 12250 51960 12256 51972
rect 12308 51960 12314 52012
rect 12894 52000 12900 52012
rect 12807 51972 12900 52000
rect 12894 51960 12900 51972
rect 12952 52000 12958 52012
rect 14384 52009 14412 52040
rect 16298 52028 16304 52080
rect 16356 52068 16362 52080
rect 16666 52068 16672 52080
rect 16356 52040 16672 52068
rect 16356 52028 16362 52040
rect 16666 52028 16672 52040
rect 16724 52028 16730 52080
rect 14369 52003 14427 52009
rect 12952 51972 14228 52000
rect 12952 51960 12958 51972
rect 12069 51935 12127 51941
rect 12069 51901 12081 51935
rect 12115 51901 12127 51935
rect 12069 51895 12127 51901
rect 12529 51935 12587 51941
rect 12529 51901 12541 51935
rect 12575 51932 12587 51935
rect 13170 51932 13176 51944
rect 12575 51904 13176 51932
rect 12575 51901 12587 51904
rect 12529 51895 12587 51901
rect 10594 51864 10600 51876
rect 10555 51836 10600 51864
rect 10594 51824 10600 51836
rect 10652 51824 10658 51876
rect 10962 51824 10968 51876
rect 11020 51864 11026 51876
rect 12084 51864 12112 51895
rect 12544 51864 12572 51895
rect 13170 51892 13176 51904
rect 13228 51892 13234 51944
rect 13906 51932 13912 51944
rect 13867 51904 13912 51932
rect 13906 51892 13912 51904
rect 13964 51892 13970 51944
rect 14200 51941 14228 51972
rect 14369 51969 14381 52003
rect 14415 51969 14427 52003
rect 14369 51963 14427 51969
rect 14642 51960 14648 52012
rect 14700 52000 14706 52012
rect 15930 52000 15936 52012
rect 14700 51972 15936 52000
rect 14700 51960 14706 51972
rect 14185 51935 14243 51941
rect 14185 51901 14197 51935
rect 14231 51932 14243 51935
rect 14274 51932 14280 51944
rect 14231 51904 14280 51932
rect 14231 51901 14243 51904
rect 14185 51895 14243 51901
rect 14274 51892 14280 51904
rect 14332 51892 14338 51944
rect 15378 51892 15384 51944
rect 15436 51932 15442 51944
rect 15473 51935 15531 51941
rect 15473 51932 15485 51935
rect 15436 51904 15485 51932
rect 15436 51892 15442 51904
rect 15473 51901 15485 51904
rect 15519 51932 15531 51935
rect 15562 51932 15568 51944
rect 15519 51904 15568 51932
rect 15519 51901 15531 51904
rect 15473 51895 15531 51901
rect 15562 51892 15568 51904
rect 15620 51892 15626 51944
rect 15856 51941 15884 51972
rect 15930 51960 15936 51972
rect 15988 51960 15994 52012
rect 17221 52003 17279 52009
rect 17221 52000 17233 52003
rect 16224 51972 17233 52000
rect 16224 51944 16252 51972
rect 17221 51969 17233 51972
rect 17267 51969 17279 52003
rect 17221 51963 17279 51969
rect 15841 51935 15899 51941
rect 15841 51901 15853 51935
rect 15887 51901 15899 51935
rect 16206 51932 16212 51944
rect 16167 51904 16212 51932
rect 15841 51895 15899 51901
rect 16206 51892 16212 51904
rect 16264 51892 16270 51944
rect 16758 51932 16764 51944
rect 16592 51904 16764 51932
rect 11020 51836 12112 51864
rect 12176 51836 12572 51864
rect 13357 51867 13415 51873
rect 11020 51824 11026 51836
rect 6512 51768 6960 51796
rect 8021 51799 8079 51805
rect 6512 51756 6518 51768
rect 8021 51765 8033 51799
rect 8067 51796 8079 51799
rect 8202 51796 8208 51808
rect 8067 51768 8208 51796
rect 8067 51765 8079 51768
rect 8021 51759 8079 51765
rect 8202 51756 8208 51768
rect 8260 51756 8266 51808
rect 8386 51756 8392 51808
rect 8444 51796 8450 51808
rect 8757 51799 8815 51805
rect 8757 51796 8769 51799
rect 8444 51768 8769 51796
rect 8444 51756 8450 51768
rect 8757 51765 8769 51768
rect 8803 51765 8815 51799
rect 8757 51759 8815 51765
rect 10413 51799 10471 51805
rect 10413 51765 10425 51799
rect 10459 51796 10471 51799
rect 10778 51796 10784 51808
rect 10459 51768 10784 51796
rect 10459 51765 10471 51768
rect 10413 51759 10471 51765
rect 10778 51756 10784 51768
rect 10836 51796 10842 51808
rect 11422 51796 11428 51808
rect 10836 51768 11428 51796
rect 10836 51756 10842 51768
rect 11422 51756 11428 51768
rect 11480 51756 11486 51808
rect 11606 51756 11612 51808
rect 11664 51796 11670 51808
rect 12176 51796 12204 51836
rect 13357 51833 13369 51867
rect 13403 51864 13415 51867
rect 13722 51864 13728 51876
rect 13403 51836 13728 51864
rect 13403 51833 13415 51836
rect 13357 51827 13415 51833
rect 13722 51824 13728 51836
rect 13780 51824 13786 51876
rect 11664 51768 12204 51796
rect 14292 51796 14320 51892
rect 15105 51867 15163 51873
rect 15105 51833 15117 51867
rect 15151 51864 15163 51867
rect 16592 51864 16620 51904
rect 16758 51892 16764 51904
rect 16816 51892 16822 51944
rect 15151 51836 16620 51864
rect 16669 51867 16727 51873
rect 15151 51833 15163 51836
rect 15105 51827 15163 51833
rect 16669 51833 16681 51867
rect 16715 51864 16727 51867
rect 17402 51864 17408 51876
rect 16715 51836 17408 51864
rect 16715 51833 16727 51836
rect 16669 51827 16727 51833
rect 16684 51796 16712 51827
rect 17402 51824 17408 51836
rect 17460 51824 17466 51876
rect 14292 51768 16712 51796
rect 11664 51756 11670 51768
rect 1104 51706 18860 51728
rect 1104 51654 7648 51706
rect 7700 51654 7712 51706
rect 7764 51654 7776 51706
rect 7828 51654 7840 51706
rect 7892 51654 14315 51706
rect 14367 51654 14379 51706
rect 14431 51654 14443 51706
rect 14495 51654 14507 51706
rect 14559 51654 18860 51706
rect 1104 51632 18860 51654
rect 1578 51552 1584 51604
rect 1636 51592 1642 51604
rect 1673 51595 1731 51601
rect 1673 51592 1685 51595
rect 1636 51564 1685 51592
rect 1636 51552 1642 51564
rect 1673 51561 1685 51564
rect 1719 51592 1731 51595
rect 3142 51592 3148 51604
rect 1719 51564 3148 51592
rect 1719 51561 1731 51564
rect 1673 51555 1731 51561
rect 3142 51552 3148 51564
rect 3200 51552 3206 51604
rect 4617 51595 4675 51601
rect 4617 51561 4629 51595
rect 4663 51592 4675 51595
rect 5905 51595 5963 51601
rect 5905 51592 5917 51595
rect 4663 51564 5917 51592
rect 4663 51561 4675 51564
rect 4617 51555 4675 51561
rect 5905 51561 5917 51564
rect 5951 51561 5963 51595
rect 6178 51592 6184 51604
rect 6139 51564 6184 51592
rect 5905 51555 5963 51561
rect 6178 51552 6184 51564
rect 6236 51552 6242 51604
rect 7101 51595 7159 51601
rect 7101 51561 7113 51595
rect 7147 51592 7159 51595
rect 8938 51592 8944 51604
rect 7147 51564 8944 51592
rect 7147 51561 7159 51564
rect 7101 51555 7159 51561
rect 7576 51536 7604 51564
rect 8938 51552 8944 51564
rect 8996 51552 9002 51604
rect 9950 51552 9956 51604
rect 10008 51592 10014 51604
rect 10318 51592 10324 51604
rect 10008 51564 10324 51592
rect 10008 51552 10014 51564
rect 10318 51552 10324 51564
rect 10376 51552 10382 51604
rect 10689 51595 10747 51601
rect 10689 51561 10701 51595
rect 10735 51592 10747 51595
rect 10962 51592 10968 51604
rect 10735 51564 10968 51592
rect 10735 51561 10747 51564
rect 10689 51555 10747 51561
rect 10962 51552 10968 51564
rect 11020 51552 11026 51604
rect 11057 51595 11115 51601
rect 11057 51561 11069 51595
rect 11103 51592 11115 51595
rect 11330 51592 11336 51604
rect 11103 51564 11336 51592
rect 11103 51561 11115 51564
rect 11057 51555 11115 51561
rect 7006 51484 7012 51536
rect 7064 51524 7070 51536
rect 7285 51527 7343 51533
rect 7285 51524 7297 51527
rect 7064 51496 7297 51524
rect 7064 51484 7070 51496
rect 7285 51493 7297 51496
rect 7331 51493 7343 51527
rect 7285 51487 7343 51493
rect 7558 51484 7564 51536
rect 7616 51484 7622 51536
rect 7653 51527 7711 51533
rect 7653 51493 7665 51527
rect 7699 51524 7711 51527
rect 8110 51524 8116 51536
rect 7699 51496 8116 51524
rect 7699 51493 7711 51496
rect 7653 51487 7711 51493
rect 8110 51484 8116 51496
rect 8168 51484 8174 51536
rect 8389 51527 8447 51533
rect 8389 51493 8401 51527
rect 8435 51524 8447 51527
rect 8662 51524 8668 51536
rect 8435 51496 8668 51524
rect 8435 51493 8447 51496
rect 8389 51487 8447 51493
rect 8662 51484 8668 51496
rect 8720 51524 8726 51536
rect 9030 51524 9036 51536
rect 8720 51496 9036 51524
rect 8720 51484 8726 51496
rect 9030 51484 9036 51496
rect 9088 51524 9094 51536
rect 9582 51524 9588 51536
rect 9088 51496 9352 51524
rect 9088 51484 9094 51496
rect 3142 51416 3148 51468
rect 3200 51456 3206 51468
rect 3786 51456 3792 51468
rect 3200 51428 3792 51456
rect 3200 51416 3206 51428
rect 3786 51416 3792 51428
rect 3844 51416 3850 51468
rect 5166 51456 5172 51468
rect 5127 51428 5172 51456
rect 5166 51416 5172 51428
rect 5224 51416 5230 51468
rect 5442 51456 5448 51468
rect 5276 51428 5448 51456
rect 4062 51348 4068 51400
rect 4120 51388 4126 51400
rect 4801 51391 4859 51397
rect 4801 51388 4813 51391
rect 4120 51360 4813 51388
rect 4120 51348 4126 51360
rect 4801 51357 4813 51360
rect 4847 51357 4859 51391
rect 4801 51351 4859 51357
rect 3050 51280 3056 51332
rect 3108 51320 3114 51332
rect 3786 51320 3792 51332
rect 3108 51292 3792 51320
rect 3108 51280 3114 51292
rect 3786 51280 3792 51292
rect 3844 51280 3850 51332
rect 4522 51320 4528 51332
rect 4080 51292 4528 51320
rect 3510 51212 3516 51264
rect 3568 51252 3574 51264
rect 4080 51261 4108 51292
rect 4522 51280 4528 51292
rect 4580 51280 4586 51332
rect 5074 51280 5080 51332
rect 5132 51320 5138 51332
rect 5276 51320 5304 51428
rect 5442 51416 5448 51428
rect 5500 51416 5506 51468
rect 5537 51459 5595 51465
rect 5537 51425 5549 51459
rect 5583 51456 5595 51459
rect 6086 51456 6092 51468
rect 5583 51428 6092 51456
rect 5583 51425 5595 51428
rect 5537 51419 5595 51425
rect 6086 51416 6092 51428
rect 6144 51416 6150 51468
rect 7193 51459 7251 51465
rect 7193 51425 7205 51459
rect 7239 51456 7251 51459
rect 7742 51456 7748 51468
rect 7239 51428 7748 51456
rect 7239 51425 7251 51428
rect 7193 51419 7251 51425
rect 7742 51416 7748 51428
rect 7800 51416 7806 51468
rect 7926 51456 7932 51468
rect 7887 51428 7932 51456
rect 7926 51416 7932 51428
rect 7984 51416 7990 51468
rect 8941 51459 8999 51465
rect 8941 51425 8953 51459
rect 8987 51425 8999 51459
rect 9214 51456 9220 51468
rect 9175 51428 9220 51456
rect 8941 51419 8999 51425
rect 6822 51348 6828 51400
rect 6880 51348 6886 51400
rect 6917 51391 6975 51397
rect 6917 51357 6929 51391
rect 6963 51388 6975 51391
rect 7006 51388 7012 51400
rect 6963 51360 7012 51388
rect 6963 51357 6975 51360
rect 6917 51351 6975 51357
rect 7006 51348 7012 51360
rect 7064 51348 7070 51400
rect 8110 51348 8116 51400
rect 8168 51388 8174 51400
rect 8481 51391 8539 51397
rect 8481 51388 8493 51391
rect 8168 51360 8493 51388
rect 8168 51348 8174 51360
rect 8481 51357 8493 51360
rect 8527 51357 8539 51391
rect 8481 51351 8539 51357
rect 8956 51388 8984 51419
rect 9214 51416 9220 51428
rect 9272 51416 9278 51468
rect 9324 51465 9352 51496
rect 9416 51496 9588 51524
rect 9309 51459 9367 51465
rect 9309 51425 9321 51459
rect 9355 51425 9367 51459
rect 9309 51419 9367 51425
rect 9416 51388 9444 51496
rect 9582 51484 9588 51496
rect 9640 51484 9646 51536
rect 9766 51484 9772 51536
rect 9824 51524 9830 51536
rect 10229 51527 10287 51533
rect 10229 51524 10241 51527
rect 9824 51496 10241 51524
rect 9824 51484 9830 51496
rect 10229 51493 10241 51496
rect 10275 51524 10287 51527
rect 10502 51524 10508 51536
rect 10275 51496 10508 51524
rect 10275 51493 10287 51496
rect 10229 51487 10287 51493
rect 10502 51484 10508 51496
rect 10560 51484 10566 51536
rect 9953 51459 10011 51465
rect 9953 51425 9965 51459
rect 9999 51456 10011 51459
rect 10318 51456 10324 51468
rect 9999 51428 10324 51456
rect 9999 51425 10011 51428
rect 9953 51419 10011 51425
rect 10318 51416 10324 51428
rect 10376 51416 10382 51468
rect 10962 51456 10968 51468
rect 10923 51428 10968 51456
rect 10962 51416 10968 51428
rect 11020 51416 11026 51468
rect 8956 51360 9444 51388
rect 9585 51391 9643 51397
rect 5132 51292 5304 51320
rect 5132 51280 5138 51292
rect 5442 51280 5448 51332
rect 5500 51320 5506 51332
rect 5629 51323 5687 51329
rect 5629 51320 5641 51323
rect 5500 51292 5641 51320
rect 5500 51280 5506 51292
rect 5629 51289 5641 51292
rect 5675 51289 5687 51323
rect 6840 51320 6868 51348
rect 5629 51283 5687 51289
rect 6380 51292 6868 51320
rect 6380 51264 6408 51292
rect 7466 51280 7472 51332
rect 7524 51320 7530 51332
rect 8956 51320 8984 51360
rect 9585 51357 9597 51391
rect 9631 51357 9643 51391
rect 9585 51351 9643 51357
rect 7524 51292 8984 51320
rect 7524 51280 7530 51292
rect 4065 51255 4123 51261
rect 4065 51252 4077 51255
rect 3568 51224 4077 51252
rect 3568 51212 3574 51224
rect 4065 51221 4077 51224
rect 4111 51221 4123 51255
rect 4065 51215 4123 51221
rect 5534 51212 5540 51264
rect 5592 51252 5598 51264
rect 5905 51255 5963 51261
rect 5905 51252 5917 51255
rect 5592 51224 5917 51252
rect 5592 51212 5598 51224
rect 5905 51221 5917 51224
rect 5951 51221 5963 51255
rect 5905 51215 5963 51221
rect 6362 51212 6368 51264
rect 6420 51212 6426 51264
rect 6641 51255 6699 51261
rect 6641 51221 6653 51255
rect 6687 51252 6699 51255
rect 7742 51252 7748 51264
rect 6687 51224 7748 51252
rect 6687 51221 6699 51224
rect 6641 51215 6699 51221
rect 7742 51212 7748 51224
rect 7800 51212 7806 51264
rect 8754 51212 8760 51264
rect 8812 51252 8818 51264
rect 9600 51252 9628 51351
rect 10134 51348 10140 51400
rect 10192 51388 10198 51400
rect 10781 51391 10839 51397
rect 10781 51388 10793 51391
rect 10192 51360 10793 51388
rect 10192 51348 10198 51360
rect 10781 51357 10793 51360
rect 10827 51357 10839 51391
rect 10781 51351 10839 51357
rect 9766 51280 9772 51332
rect 9824 51320 9830 51332
rect 11072 51320 11100 51555
rect 11330 51552 11336 51564
rect 11388 51552 11394 51604
rect 12805 51595 12863 51601
rect 12805 51592 12817 51595
rect 12544 51564 12817 51592
rect 11149 51527 11207 51533
rect 11149 51493 11161 51527
rect 11195 51524 11207 51527
rect 12158 51524 12164 51536
rect 11195 51496 11652 51524
rect 12119 51496 12164 51524
rect 11195 51493 11207 51496
rect 11149 51487 11207 51493
rect 11330 51416 11336 51468
rect 11388 51416 11394 51468
rect 11624 51456 11652 51496
rect 12158 51484 12164 51496
rect 12216 51484 12222 51536
rect 12434 51484 12440 51536
rect 12492 51524 12498 51536
rect 12544 51524 12572 51564
rect 12805 51561 12817 51564
rect 12851 51592 12863 51595
rect 13906 51592 13912 51604
rect 12851 51564 13912 51592
rect 12851 51561 12863 51564
rect 12805 51555 12863 51561
rect 13906 51552 13912 51564
rect 13964 51552 13970 51604
rect 14921 51595 14979 51601
rect 14921 51561 14933 51595
rect 14967 51592 14979 51595
rect 15010 51592 15016 51604
rect 14967 51564 15016 51592
rect 14967 51561 14979 51564
rect 14921 51555 14979 51561
rect 15010 51552 15016 51564
rect 15068 51552 15074 51604
rect 17126 51592 17132 51604
rect 17087 51564 17132 51592
rect 17126 51552 17132 51564
rect 17184 51552 17190 51604
rect 17494 51592 17500 51604
rect 17455 51564 17500 51592
rect 17494 51552 17500 51564
rect 17552 51552 17558 51604
rect 12492 51496 12572 51524
rect 12492 51484 12498 51496
rect 12894 51484 12900 51536
rect 12952 51484 12958 51536
rect 14553 51527 14611 51533
rect 14553 51493 14565 51527
rect 14599 51524 14611 51527
rect 17034 51524 17040 51536
rect 14599 51496 17040 51524
rect 14599 51493 14611 51496
rect 14553 51487 14611 51493
rect 11624 51428 12204 51456
rect 9824 51292 11100 51320
rect 11348 51320 11376 51416
rect 11517 51391 11575 51397
rect 11517 51357 11529 51391
rect 11563 51388 11575 51391
rect 11606 51388 11612 51400
rect 11563 51360 11612 51388
rect 11563 51357 11575 51360
rect 11517 51351 11575 51357
rect 11606 51348 11612 51360
rect 11664 51388 11670 51400
rect 11793 51391 11851 51397
rect 11793 51388 11805 51391
rect 11664 51360 11805 51388
rect 11664 51348 11670 51360
rect 11793 51357 11805 51360
rect 11839 51357 11851 51391
rect 12176 51388 12204 51428
rect 12250 51416 12256 51468
rect 12308 51456 12314 51468
rect 12526 51456 12532 51468
rect 12308 51428 12532 51456
rect 12308 51416 12314 51428
rect 12526 51416 12532 51428
rect 12584 51416 12590 51468
rect 12912 51456 12940 51484
rect 14568 51456 14596 51487
rect 17034 51484 17040 51496
rect 17092 51484 17098 51536
rect 15562 51456 15568 51468
rect 12636 51428 14596 51456
rect 15523 51428 15568 51456
rect 12636 51388 12664 51428
rect 15562 51416 15568 51428
rect 15620 51416 15626 51468
rect 16022 51456 16028 51468
rect 15983 51428 16028 51456
rect 16022 51416 16028 51428
rect 16080 51416 16086 51468
rect 16206 51456 16212 51468
rect 16167 51428 16212 51456
rect 16206 51416 16212 51428
rect 16264 51456 16270 51468
rect 16390 51456 16396 51468
rect 16264 51428 16396 51456
rect 16264 51416 16270 51428
rect 16390 51416 16396 51428
rect 16448 51416 16454 51468
rect 16758 51456 16764 51468
rect 16719 51428 16764 51456
rect 16758 51416 16764 51428
rect 16816 51456 16822 51468
rect 17310 51456 17316 51468
rect 16816 51428 17316 51456
rect 16816 51416 16822 51428
rect 17310 51416 17316 51428
rect 17368 51416 17374 51468
rect 12894 51388 12900 51400
rect 12176 51360 12664 51388
rect 12855 51360 12900 51388
rect 11793 51351 11851 51357
rect 12894 51348 12900 51360
rect 12952 51348 12958 51400
rect 13170 51388 13176 51400
rect 13131 51360 13176 51388
rect 13170 51348 13176 51360
rect 13228 51348 13234 51400
rect 15289 51391 15347 51397
rect 15289 51357 15301 51391
rect 15335 51388 15347 51391
rect 15378 51388 15384 51400
rect 15335 51360 15384 51388
rect 15335 51357 15347 51360
rect 15289 51351 15347 51357
rect 15378 51348 15384 51360
rect 15436 51348 15442 51400
rect 11348 51292 12112 51320
rect 9824 51280 9830 51292
rect 12084 51264 12112 51292
rect 8812 51224 9628 51252
rect 8812 51212 8818 51224
rect 12066 51212 12072 51264
rect 12124 51212 12130 51264
rect 12618 51212 12624 51264
rect 12676 51252 12682 51264
rect 13262 51252 13268 51264
rect 12676 51224 13268 51252
rect 12676 51212 12682 51224
rect 13262 51212 13268 51224
rect 13320 51212 13326 51264
rect 15378 51212 15384 51264
rect 15436 51252 15442 51264
rect 15473 51255 15531 51261
rect 15473 51252 15485 51255
rect 15436 51224 15485 51252
rect 15436 51212 15442 51224
rect 15473 51221 15485 51224
rect 15519 51221 15531 51255
rect 15473 51215 15531 51221
rect 1104 51162 18860 51184
rect 1104 51110 4315 51162
rect 4367 51110 4379 51162
rect 4431 51110 4443 51162
rect 4495 51110 4507 51162
rect 4559 51110 10982 51162
rect 11034 51110 11046 51162
rect 11098 51110 11110 51162
rect 11162 51110 11174 51162
rect 11226 51110 17648 51162
rect 17700 51110 17712 51162
rect 17764 51110 17776 51162
rect 17828 51110 17840 51162
rect 17892 51110 18860 51162
rect 1104 51088 18860 51110
rect 3053 51051 3111 51057
rect 3053 51017 3065 51051
rect 3099 51048 3111 51051
rect 3234 51048 3240 51060
rect 3099 51020 3240 51048
rect 3099 51017 3111 51020
rect 3053 51011 3111 51017
rect 3234 51008 3240 51020
rect 3292 51008 3298 51060
rect 3881 51051 3939 51057
rect 3881 51017 3893 51051
rect 3927 51048 3939 51051
rect 4062 51048 4068 51060
rect 3927 51020 4068 51048
rect 3927 51017 3939 51020
rect 3881 51011 3939 51017
rect 4062 51008 4068 51020
rect 4120 51008 4126 51060
rect 4985 51051 5043 51057
rect 4985 51017 4997 51051
rect 5031 51048 5043 51051
rect 5166 51048 5172 51060
rect 5031 51020 5172 51048
rect 5031 51017 5043 51020
rect 4985 51011 5043 51017
rect 4522 50940 4528 50992
rect 4580 50980 4586 50992
rect 5000 50980 5028 51011
rect 5166 51008 5172 51020
rect 5224 51008 5230 51060
rect 5445 51051 5503 51057
rect 5445 51017 5457 51051
rect 5491 51048 5503 51051
rect 5718 51048 5724 51060
rect 5491 51020 5724 51048
rect 5491 51017 5503 51020
rect 5445 51011 5503 51017
rect 5718 51008 5724 51020
rect 5776 51008 5782 51060
rect 6086 51008 6092 51060
rect 6144 51048 6150 51060
rect 6181 51051 6239 51057
rect 6181 51048 6193 51051
rect 6144 51020 6193 51048
rect 6144 51008 6150 51020
rect 6181 51017 6193 51020
rect 6227 51017 6239 51051
rect 6181 51011 6239 51017
rect 6733 51051 6791 51057
rect 6733 51017 6745 51051
rect 6779 51048 6791 51051
rect 7558 51048 7564 51060
rect 6779 51020 7564 51048
rect 6779 51017 6791 51020
rect 6733 51011 6791 51017
rect 7558 51008 7564 51020
rect 7616 51008 7622 51060
rect 7834 51008 7840 51060
rect 7892 51048 7898 51060
rect 7892 51020 8156 51048
rect 7892 51008 7898 51020
rect 4580 50952 5028 50980
rect 4580 50940 4586 50952
rect 5534 50940 5540 50992
rect 5592 50980 5598 50992
rect 7466 50980 7472 50992
rect 5592 50952 7472 50980
rect 5592 50940 5598 50952
rect 7466 50940 7472 50952
rect 7524 50940 7530 50992
rect 7926 50940 7932 50992
rect 7984 50940 7990 50992
rect 8128 50980 8156 51020
rect 8202 51008 8208 51060
rect 8260 51048 8266 51060
rect 8757 51051 8815 51057
rect 8757 51048 8769 51051
rect 8260 51020 8769 51048
rect 8260 51008 8266 51020
rect 8757 51017 8769 51020
rect 8803 51017 8815 51051
rect 8757 51011 8815 51017
rect 9214 51008 9220 51060
rect 9272 51048 9278 51060
rect 9309 51051 9367 51057
rect 9309 51048 9321 51051
rect 9272 51020 9321 51048
rect 9272 51008 9278 51020
rect 9309 51017 9321 51020
rect 9355 51048 9367 51051
rect 9674 51048 9680 51060
rect 9355 51020 9680 51048
rect 9355 51017 9367 51020
rect 9309 51011 9367 51017
rect 9674 51008 9680 51020
rect 9732 51008 9738 51060
rect 9766 51008 9772 51060
rect 9824 51048 9830 51060
rect 10045 51051 10103 51057
rect 10045 51048 10057 51051
rect 9824 51020 10057 51048
rect 9824 51008 9830 51020
rect 10045 51017 10057 51020
rect 10091 51017 10103 51051
rect 10045 51011 10103 51017
rect 10318 51008 10324 51060
rect 10376 51048 10382 51060
rect 11974 51048 11980 51060
rect 10376 51020 11980 51048
rect 10376 51008 10382 51020
rect 11974 51008 11980 51020
rect 12032 51008 12038 51060
rect 12434 51008 12440 51060
rect 12492 51048 12498 51060
rect 12492 51020 12537 51048
rect 12492 51008 12498 51020
rect 12802 51008 12808 51060
rect 12860 51008 12866 51060
rect 13170 51048 13176 51060
rect 13131 51020 13176 51048
rect 13170 51008 13176 51020
rect 13228 51008 13234 51060
rect 13446 51008 13452 51060
rect 13504 51048 13510 51060
rect 13722 51048 13728 51060
rect 13504 51020 13728 51048
rect 13504 51008 13510 51020
rect 13722 51008 13728 51020
rect 13780 51008 13786 51060
rect 14461 51051 14519 51057
rect 14461 51017 14473 51051
rect 14507 51048 14519 51051
rect 14737 51051 14795 51057
rect 14737 51048 14749 51051
rect 14507 51020 14749 51048
rect 14507 51017 14519 51020
rect 14461 51011 14519 51017
rect 14737 51017 14749 51020
rect 14783 51048 14795 51051
rect 15286 51048 15292 51060
rect 14783 51020 15292 51048
rect 14783 51017 14795 51020
rect 14737 51011 14795 51017
rect 15286 51008 15292 51020
rect 15344 51008 15350 51060
rect 8128 50952 8708 50980
rect 3513 50915 3571 50921
rect 3513 50881 3525 50915
rect 3559 50912 3571 50915
rect 5810 50912 5816 50924
rect 3559 50884 5816 50912
rect 3559 50881 3571 50884
rect 3513 50875 3571 50881
rect 1489 50847 1547 50853
rect 1489 50813 1501 50847
rect 1535 50844 1547 50847
rect 1578 50844 1584 50856
rect 1535 50816 1584 50844
rect 1535 50813 1547 50816
rect 1489 50807 1547 50813
rect 1578 50804 1584 50816
rect 1636 50804 1642 50856
rect 1762 50844 1768 50856
rect 1723 50816 1768 50844
rect 1762 50804 1768 50816
rect 1820 50804 1826 50856
rect 2222 50804 2228 50856
rect 2280 50844 2286 50856
rect 4065 50847 4123 50853
rect 4065 50844 4077 50847
rect 2280 50816 4077 50844
rect 2280 50804 2286 50816
rect 4065 50813 4077 50816
rect 4111 50844 4123 50847
rect 4525 50847 4583 50853
rect 4525 50844 4537 50847
rect 4111 50816 4537 50844
rect 4111 50813 4123 50816
rect 4065 50807 4123 50813
rect 4525 50813 4537 50816
rect 4571 50813 4583 50847
rect 4525 50807 4583 50813
rect 5166 50804 5172 50856
rect 5224 50844 5230 50856
rect 5368 50853 5396 50884
rect 5810 50872 5816 50884
rect 5868 50872 5874 50924
rect 7190 50912 7196 50924
rect 6472 50884 7196 50912
rect 6472 50856 6500 50884
rect 7190 50872 7196 50884
rect 7248 50872 7254 50924
rect 7944 50912 7972 50940
rect 8570 50912 8576 50924
rect 7944 50884 8156 50912
rect 5353 50847 5411 50853
rect 5224 50816 5304 50844
rect 5224 50804 5230 50816
rect 5276 50776 5304 50816
rect 5353 50813 5365 50847
rect 5399 50813 5411 50847
rect 5353 50807 5411 50813
rect 5626 50804 5632 50856
rect 5684 50804 5690 50856
rect 6454 50804 6460 50856
rect 6512 50804 6518 50856
rect 7006 50804 7012 50856
rect 7064 50804 7070 50856
rect 7466 50804 7472 50856
rect 7524 50844 7530 50856
rect 7742 50844 7748 50856
rect 7524 50816 7748 50844
rect 7524 50804 7530 50816
rect 7742 50804 7748 50816
rect 7800 50804 7806 50856
rect 8128 50853 8156 50884
rect 8312 50884 8576 50912
rect 8312 50853 8340 50884
rect 8570 50872 8576 50884
rect 8628 50872 8634 50924
rect 8680 50912 8708 50952
rect 9784 50912 9812 51008
rect 8680 50884 9812 50912
rect 11606 50872 11612 50924
rect 11664 50872 11670 50924
rect 7837 50847 7895 50853
rect 7837 50813 7849 50847
rect 7883 50813 7895 50847
rect 7837 50807 7895 50813
rect 8113 50847 8171 50853
rect 8113 50813 8125 50847
rect 8159 50813 8171 50847
rect 8113 50807 8171 50813
rect 8297 50847 8355 50853
rect 8297 50813 8309 50847
rect 8343 50813 8355 50847
rect 8297 50807 8355 50813
rect 8481 50847 8539 50853
rect 8481 50813 8493 50847
rect 8527 50813 8539 50847
rect 8754 50844 8760 50856
rect 8715 50816 8760 50844
rect 8481 50807 8539 50813
rect 5445 50779 5503 50785
rect 5445 50776 5457 50779
rect 2424 50748 5212 50776
rect 5276 50748 5457 50776
rect 2424 50720 2452 50748
rect 2406 50668 2412 50720
rect 2464 50668 2470 50720
rect 4246 50708 4252 50720
rect 4207 50680 4252 50708
rect 4246 50668 4252 50680
rect 4304 50668 4310 50720
rect 5184 50717 5212 50748
rect 5445 50745 5457 50748
rect 5491 50745 5503 50779
rect 5644 50776 5672 50804
rect 6730 50776 6736 50788
rect 5644 50748 6736 50776
rect 5445 50739 5503 50745
rect 6730 50736 6736 50748
rect 6788 50736 6794 50788
rect 7024 50776 7052 50804
rect 6840 50748 7052 50776
rect 5169 50711 5227 50717
rect 5169 50677 5181 50711
rect 5215 50677 5227 50711
rect 5626 50708 5632 50720
rect 5587 50680 5632 50708
rect 5169 50671 5227 50677
rect 5626 50668 5632 50680
rect 5684 50708 5690 50720
rect 6181 50711 6239 50717
rect 6181 50708 6193 50711
rect 5684 50680 6193 50708
rect 5684 50668 5690 50680
rect 6181 50677 6193 50680
rect 6227 50677 6239 50711
rect 6181 50671 6239 50677
rect 6365 50711 6423 50717
rect 6365 50677 6377 50711
rect 6411 50708 6423 50711
rect 6840 50708 6868 50748
rect 7374 50736 7380 50788
rect 7432 50776 7438 50788
rect 7852 50776 7880 50807
rect 7432 50748 7880 50776
rect 7432 50736 7438 50748
rect 8202 50736 8208 50788
rect 8260 50776 8266 50788
rect 8312 50776 8340 50807
rect 8260 50748 8340 50776
rect 8260 50736 8266 50748
rect 8496 50720 8524 50807
rect 8754 50804 8760 50816
rect 8812 50804 8818 50856
rect 10318 50844 10324 50856
rect 10152 50816 10324 50844
rect 7006 50708 7012 50720
rect 6411 50680 6868 50708
rect 6967 50680 7012 50708
rect 6411 50677 6423 50680
rect 6365 50671 6423 50677
rect 7006 50668 7012 50680
rect 7064 50668 7070 50720
rect 7282 50708 7288 50720
rect 7243 50680 7288 50708
rect 7282 50668 7288 50680
rect 7340 50668 7346 50720
rect 8478 50668 8484 50720
rect 8536 50668 8542 50720
rect 8938 50708 8944 50720
rect 8899 50680 8944 50708
rect 8938 50668 8944 50680
rect 8996 50668 9002 50720
rect 9766 50668 9772 50720
rect 9824 50708 9830 50720
rect 10152 50708 10180 50816
rect 10318 50804 10324 50816
rect 10376 50804 10382 50856
rect 10502 50844 10508 50856
rect 10463 50816 10508 50844
rect 10502 50804 10508 50816
rect 10560 50804 10566 50856
rect 10965 50847 11023 50853
rect 10965 50813 10977 50847
rect 11011 50813 11023 50847
rect 11238 50844 11244 50856
rect 11199 50816 11244 50844
rect 10965 50807 11023 50813
rect 10686 50736 10692 50788
rect 10744 50776 10750 50788
rect 10980 50776 11008 50807
rect 11238 50804 11244 50816
rect 11296 50804 11302 50856
rect 11517 50847 11575 50853
rect 11517 50813 11529 50847
rect 11563 50844 11575 50847
rect 11624 50844 11652 50872
rect 11563 50816 11652 50844
rect 12713 50847 12771 50853
rect 11563 50813 11575 50816
rect 11517 50807 11575 50813
rect 12713 50813 12725 50847
rect 12759 50844 12771 50847
rect 12820 50844 12848 51008
rect 17034 50940 17040 50992
rect 17092 50980 17098 50992
rect 17497 50983 17555 50989
rect 17497 50980 17509 50983
rect 17092 50952 17509 50980
rect 17092 50940 17098 50952
rect 17497 50949 17509 50952
rect 17543 50949 17555 50983
rect 17497 50943 17555 50949
rect 13170 50872 13176 50924
rect 13228 50912 13234 50924
rect 14369 50915 14427 50921
rect 14369 50912 14381 50915
rect 13228 50884 14381 50912
rect 13228 50872 13234 50884
rect 14369 50881 14381 50884
rect 14415 50912 14427 50915
rect 15010 50912 15016 50924
rect 14415 50884 15016 50912
rect 14415 50881 14427 50884
rect 14369 50875 14427 50881
rect 15010 50872 15016 50884
rect 15068 50872 15074 50924
rect 15102 50872 15108 50924
rect 15160 50912 15166 50924
rect 15746 50912 15752 50924
rect 15160 50884 15752 50912
rect 15160 50872 15166 50884
rect 15746 50872 15752 50884
rect 15804 50872 15810 50924
rect 15841 50915 15899 50921
rect 15841 50881 15853 50915
rect 15887 50912 15899 50915
rect 17310 50912 17316 50924
rect 15887 50884 17316 50912
rect 15887 50881 15899 50884
rect 15841 50875 15899 50881
rect 17310 50872 17316 50884
rect 17368 50872 17374 50924
rect 13722 50844 13728 50856
rect 12759 50816 13728 50844
rect 12759 50813 12771 50816
rect 12713 50807 12771 50813
rect 13722 50804 13728 50816
rect 13780 50804 13786 50856
rect 13906 50844 13912 50856
rect 13819 50816 13912 50844
rect 13906 50804 13912 50816
rect 13964 50804 13970 50856
rect 14185 50847 14243 50853
rect 14185 50813 14197 50847
rect 14231 50844 14243 50847
rect 14461 50847 14519 50853
rect 14461 50844 14473 50847
rect 14231 50816 14473 50844
rect 14231 50813 14243 50816
rect 14185 50807 14243 50813
rect 14461 50813 14473 50816
rect 14507 50813 14519 50847
rect 14461 50807 14519 50813
rect 15289 50847 15347 50853
rect 15289 50813 15301 50847
rect 15335 50844 15347 50847
rect 16117 50847 16175 50853
rect 16117 50844 16129 50847
rect 15335 50816 16129 50844
rect 15335 50813 15347 50816
rect 15289 50807 15347 50813
rect 16117 50813 16129 50816
rect 16163 50844 16175 50847
rect 16574 50844 16580 50856
rect 16163 50816 16580 50844
rect 16163 50813 16175 50816
rect 16117 50807 16175 50813
rect 16574 50804 16580 50816
rect 16632 50804 16638 50856
rect 16669 50847 16727 50853
rect 16669 50813 16681 50847
rect 16715 50813 16727 50847
rect 17126 50844 17132 50856
rect 17087 50816 17132 50844
rect 16669 50807 16727 50813
rect 11977 50779 12035 50785
rect 11977 50776 11989 50779
rect 10744 50748 11989 50776
rect 10744 50736 10750 50748
rect 11977 50745 11989 50748
rect 12023 50745 12035 50779
rect 11977 50739 12035 50745
rect 13262 50736 13268 50788
rect 13320 50776 13326 50788
rect 13357 50779 13415 50785
rect 13357 50776 13369 50779
rect 13320 50748 13369 50776
rect 13320 50736 13326 50748
rect 13357 50745 13369 50748
rect 13403 50745 13415 50779
rect 13924 50776 13952 50804
rect 13924 50748 15148 50776
rect 13357 50739 13415 50745
rect 10318 50708 10324 50720
rect 9824 50680 10180 50708
rect 10279 50680 10324 50708
rect 9824 50668 9830 50680
rect 10318 50668 10324 50680
rect 10376 50668 10382 50720
rect 12529 50711 12587 50717
rect 12529 50677 12541 50711
rect 12575 50708 12587 50711
rect 12802 50708 12808 50720
rect 12575 50680 12808 50708
rect 12575 50677 12587 50680
rect 12529 50671 12587 50677
rect 12802 50668 12808 50680
rect 12860 50668 12866 50720
rect 12894 50668 12900 50720
rect 12952 50708 12958 50720
rect 13081 50711 13139 50717
rect 13081 50708 13093 50711
rect 12952 50680 13093 50708
rect 12952 50668 12958 50680
rect 13081 50677 13093 50680
rect 13127 50708 13139 50711
rect 13173 50711 13231 50717
rect 13173 50708 13185 50711
rect 13127 50680 13185 50708
rect 13127 50677 13139 50680
rect 13081 50671 13139 50677
rect 13173 50677 13185 50680
rect 13219 50677 13231 50711
rect 13173 50671 13231 50677
rect 14826 50668 14832 50720
rect 14884 50708 14890 50720
rect 15013 50711 15071 50717
rect 15013 50708 15025 50711
rect 14884 50680 15025 50708
rect 14884 50668 14890 50680
rect 15013 50677 15025 50680
rect 15059 50677 15071 50711
rect 15120 50708 15148 50748
rect 15286 50708 15292 50720
rect 15120 50680 15292 50708
rect 15013 50671 15071 50677
rect 15286 50668 15292 50680
rect 15344 50668 15350 50720
rect 15470 50708 15476 50720
rect 15431 50680 15476 50708
rect 15470 50668 15476 50680
rect 15528 50668 15534 50720
rect 16574 50708 16580 50720
rect 16535 50680 16580 50708
rect 16574 50668 16580 50680
rect 16632 50708 16638 50720
rect 16684 50708 16712 50807
rect 17126 50804 17132 50816
rect 17184 50804 17190 50856
rect 17494 50844 17500 50856
rect 17455 50816 17500 50844
rect 17494 50804 17500 50816
rect 17552 50804 17558 50856
rect 18046 50708 18052 50720
rect 16632 50680 16712 50708
rect 18007 50680 18052 50708
rect 16632 50668 16638 50680
rect 18046 50668 18052 50680
rect 18104 50668 18110 50720
rect 1104 50618 18860 50640
rect 1104 50566 7648 50618
rect 7700 50566 7712 50618
rect 7764 50566 7776 50618
rect 7828 50566 7840 50618
rect 7892 50566 14315 50618
rect 14367 50566 14379 50618
rect 14431 50566 14443 50618
rect 14495 50566 14507 50618
rect 14559 50566 18860 50618
rect 1104 50544 18860 50566
rect 4709 50507 4767 50513
rect 4709 50473 4721 50507
rect 4755 50504 4767 50507
rect 4890 50504 4896 50516
rect 4755 50476 4896 50504
rect 4755 50473 4767 50476
rect 4709 50467 4767 50473
rect 4890 50464 4896 50476
rect 4948 50464 4954 50516
rect 5077 50507 5135 50513
rect 5077 50473 5089 50507
rect 5123 50504 5135 50507
rect 5166 50504 5172 50516
rect 5123 50476 5172 50504
rect 5123 50473 5135 50476
rect 5077 50467 5135 50473
rect 5166 50464 5172 50476
rect 5224 50464 5230 50516
rect 5534 50504 5540 50516
rect 5495 50476 5540 50504
rect 5534 50464 5540 50476
rect 5592 50464 5598 50516
rect 6641 50507 6699 50513
rect 6641 50473 6653 50507
rect 6687 50504 6699 50507
rect 7374 50504 7380 50516
rect 6687 50476 7380 50504
rect 6687 50473 6699 50476
rect 6641 50467 6699 50473
rect 7374 50464 7380 50476
rect 7432 50464 7438 50516
rect 7469 50507 7527 50513
rect 7469 50473 7481 50507
rect 7515 50504 7527 50507
rect 8202 50504 8208 50516
rect 7515 50476 8208 50504
rect 7515 50473 7527 50476
rect 7469 50467 7527 50473
rect 8202 50464 8208 50476
rect 8260 50464 8266 50516
rect 8294 50464 8300 50516
rect 8352 50504 8358 50516
rect 8389 50507 8447 50513
rect 8389 50504 8401 50507
rect 8352 50476 8401 50504
rect 8352 50464 8358 50476
rect 8389 50473 8401 50476
rect 8435 50473 8447 50507
rect 9398 50504 9404 50516
rect 8389 50467 8447 50473
rect 9048 50476 9404 50504
rect 3329 50439 3387 50445
rect 3329 50405 3341 50439
rect 3375 50436 3387 50439
rect 3694 50436 3700 50448
rect 3375 50408 3700 50436
rect 3375 50405 3387 50408
rect 3329 50399 3387 50405
rect 3694 50396 3700 50408
rect 3752 50396 3758 50448
rect 5905 50439 5963 50445
rect 5905 50405 5917 50439
rect 5951 50436 5963 50439
rect 6822 50436 6828 50448
rect 5951 50408 6828 50436
rect 5951 50405 5963 50408
rect 5905 50399 5963 50405
rect 6822 50396 6828 50408
rect 6880 50396 6886 50448
rect 7190 50396 7196 50448
rect 7248 50436 7254 50448
rect 7837 50439 7895 50445
rect 7837 50436 7849 50439
rect 7248 50408 7849 50436
rect 7248 50396 7254 50408
rect 7837 50405 7849 50408
rect 7883 50405 7895 50439
rect 9048 50436 9076 50476
rect 9398 50464 9404 50476
rect 9456 50464 9462 50516
rect 10778 50504 10784 50516
rect 10739 50476 10784 50504
rect 10778 50464 10784 50476
rect 10836 50464 10842 50516
rect 11238 50464 11244 50516
rect 11296 50504 11302 50516
rect 11793 50507 11851 50513
rect 11793 50504 11805 50507
rect 11296 50476 11805 50504
rect 11296 50464 11302 50476
rect 11793 50473 11805 50476
rect 11839 50473 11851 50507
rect 11793 50467 11851 50473
rect 12989 50507 13047 50513
rect 12989 50473 13001 50507
rect 13035 50504 13047 50507
rect 13170 50504 13176 50516
rect 13035 50476 13176 50504
rect 13035 50473 13047 50476
rect 12989 50467 13047 50473
rect 7837 50399 7895 50405
rect 8312 50408 9076 50436
rect 4062 50368 4068 50380
rect 4023 50340 4068 50368
rect 4062 50328 4068 50340
rect 4120 50328 4126 50380
rect 4154 50328 4160 50380
rect 4212 50368 4218 50380
rect 4212 50340 4257 50368
rect 4212 50328 4218 50340
rect 3234 50300 3240 50312
rect 3195 50272 3240 50300
rect 3234 50260 3240 50272
rect 3292 50260 3298 50312
rect 3510 50260 3516 50312
rect 3568 50300 3574 50312
rect 3694 50300 3700 50312
rect 3568 50272 3700 50300
rect 3568 50260 3574 50272
rect 3694 50260 3700 50272
rect 3752 50300 3758 50312
rect 4246 50300 4252 50312
rect 3752 50272 4252 50300
rect 3752 50260 3758 50272
rect 4246 50260 4252 50272
rect 4304 50260 4310 50312
rect 6362 50260 6368 50312
rect 6420 50300 6426 50312
rect 7190 50300 7196 50312
rect 6420 50272 7196 50300
rect 6420 50260 6426 50272
rect 7190 50260 7196 50272
rect 7248 50260 7254 50312
rect 7852 50300 7880 50399
rect 8312 50377 8340 50408
rect 9048 50377 9076 50408
rect 10134 50396 10140 50448
rect 10192 50436 10198 50448
rect 11149 50439 11207 50445
rect 11149 50436 11161 50439
rect 10192 50408 11161 50436
rect 10192 50396 10198 50408
rect 11149 50405 11161 50408
rect 11195 50405 11207 50439
rect 11149 50399 11207 50405
rect 8297 50371 8355 50377
rect 8297 50337 8309 50371
rect 8343 50337 8355 50371
rect 8297 50331 8355 50337
rect 8573 50371 8631 50377
rect 8573 50337 8585 50371
rect 8619 50368 8631 50371
rect 9033 50371 9091 50377
rect 8619 50340 8800 50368
rect 8619 50337 8631 50340
rect 8573 50331 8631 50337
rect 8665 50303 8723 50309
rect 8665 50300 8677 50303
rect 7852 50272 8677 50300
rect 8665 50269 8677 50272
rect 8711 50269 8723 50303
rect 8665 50263 8723 50269
rect 7101 50235 7159 50241
rect 7101 50201 7113 50235
rect 7147 50232 7159 50235
rect 7466 50232 7472 50244
rect 7147 50204 7472 50232
rect 7147 50201 7159 50204
rect 7101 50195 7159 50201
rect 7466 50192 7472 50204
rect 7524 50192 7530 50244
rect 8294 50192 8300 50244
rect 8352 50232 8358 50244
rect 8772 50232 8800 50340
rect 9033 50337 9045 50371
rect 9079 50337 9091 50371
rect 9214 50368 9220 50380
rect 9175 50340 9220 50368
rect 9033 50331 9091 50337
rect 9214 50328 9220 50340
rect 9272 50328 9278 50380
rect 9398 50368 9404 50380
rect 9359 50340 9404 50368
rect 9398 50328 9404 50340
rect 9456 50328 9462 50380
rect 9677 50371 9735 50377
rect 9677 50337 9689 50371
rect 9723 50368 9735 50371
rect 10962 50368 10968 50380
rect 9723 50340 10968 50368
rect 9723 50337 9735 50340
rect 9677 50331 9735 50337
rect 10962 50328 10968 50340
rect 11020 50328 11026 50380
rect 11333 50371 11391 50377
rect 11333 50337 11345 50371
rect 11379 50368 11391 50371
rect 11514 50368 11520 50380
rect 11379 50340 11520 50368
rect 11379 50337 11391 50340
rect 11333 50331 11391 50337
rect 11514 50328 11520 50340
rect 11572 50328 11578 50380
rect 8938 50260 8944 50312
rect 8996 50300 9002 50312
rect 9416 50300 9444 50328
rect 8996 50272 9444 50300
rect 11808 50300 11836 50467
rect 13170 50464 13176 50476
rect 13228 50464 13234 50516
rect 15473 50507 15531 50513
rect 15473 50473 15485 50507
rect 15519 50504 15531 50507
rect 16022 50504 16028 50516
rect 15519 50476 16028 50504
rect 15519 50473 15531 50476
rect 15473 50467 15531 50473
rect 16022 50464 16028 50476
rect 16080 50464 16086 50516
rect 17126 50464 17132 50516
rect 17184 50504 17190 50516
rect 17313 50507 17371 50513
rect 17313 50504 17325 50507
rect 17184 50476 17325 50504
rect 17184 50464 17190 50476
rect 17313 50473 17325 50476
rect 17359 50473 17371 50507
rect 17313 50467 17371 50473
rect 14826 50396 14832 50448
rect 14884 50436 14890 50448
rect 16206 50436 16212 50448
rect 14884 50408 16212 50436
rect 14884 50396 14890 50408
rect 16206 50396 16212 50408
rect 16264 50436 16270 50448
rect 16264 50408 16344 50436
rect 16264 50396 16270 50408
rect 12253 50371 12311 50377
rect 12253 50337 12265 50371
rect 12299 50368 12311 50371
rect 13170 50368 13176 50380
rect 12299 50340 13176 50368
rect 12299 50337 12311 50340
rect 12253 50331 12311 50337
rect 13170 50328 13176 50340
rect 13228 50328 13234 50380
rect 13354 50368 13360 50380
rect 13315 50340 13360 50368
rect 13354 50328 13360 50340
rect 13412 50328 13418 50380
rect 15105 50371 15163 50377
rect 15105 50337 15117 50371
rect 15151 50368 15163 50371
rect 15562 50368 15568 50380
rect 15151 50340 15568 50368
rect 15151 50337 15163 50340
rect 15105 50331 15163 50337
rect 15562 50328 15568 50340
rect 15620 50328 15626 50380
rect 15746 50328 15752 50380
rect 15804 50368 15810 50380
rect 16316 50377 16344 50408
rect 15933 50371 15991 50377
rect 15933 50368 15945 50371
rect 15804 50340 15945 50368
rect 15804 50328 15810 50340
rect 15933 50337 15945 50340
rect 15979 50337 15991 50371
rect 15933 50331 15991 50337
rect 16301 50371 16359 50377
rect 16301 50337 16313 50371
rect 16347 50337 16359 50371
rect 16301 50331 16359 50337
rect 16853 50371 16911 50377
rect 16853 50337 16865 50371
rect 16899 50368 16911 50371
rect 17126 50368 17132 50380
rect 16899 50340 17132 50368
rect 16899 50337 16911 50340
rect 16853 50331 16911 50337
rect 12434 50300 12440 50312
rect 11808 50272 12440 50300
rect 8996 50260 9002 50272
rect 12434 50260 12440 50272
rect 12492 50260 12498 50312
rect 12802 50260 12808 50312
rect 12860 50300 12866 50312
rect 13081 50303 13139 50309
rect 13081 50300 13093 50303
rect 12860 50272 13093 50300
rect 12860 50260 12866 50272
rect 13081 50269 13093 50272
rect 13127 50300 13139 50303
rect 15838 50300 15844 50312
rect 13127 50272 14044 50300
rect 15799 50272 15844 50300
rect 13127 50269 13139 50272
rect 13081 50263 13139 50269
rect 8352 50204 8800 50232
rect 11517 50235 11575 50241
rect 8352 50192 8358 50204
rect 11517 50201 11529 50235
rect 11563 50232 11575 50235
rect 11882 50232 11888 50244
rect 11563 50204 11888 50232
rect 11563 50201 11575 50204
rect 11517 50195 11575 50201
rect 11882 50192 11888 50204
rect 11940 50232 11946 50244
rect 12250 50232 12256 50244
rect 11940 50204 12256 50232
rect 11940 50192 11946 50204
rect 12250 50192 12256 50204
rect 12308 50192 12314 50244
rect 14016 50232 14044 50272
rect 15838 50260 15844 50272
rect 15896 50260 15902 50312
rect 16206 50260 16212 50312
rect 16264 50300 16270 50312
rect 16868 50300 16896 50331
rect 17126 50328 17132 50340
rect 17184 50368 17190 50380
rect 17310 50368 17316 50380
rect 17184 50340 17316 50368
rect 17184 50328 17190 50340
rect 17310 50328 17316 50340
rect 17368 50328 17374 50380
rect 16264 50272 16896 50300
rect 16264 50260 16270 50272
rect 18046 50232 18052 50244
rect 14016 50204 18052 50232
rect 18046 50192 18052 50204
rect 18104 50192 18110 50244
rect 1673 50167 1731 50173
rect 1673 50133 1685 50167
rect 1719 50164 1731 50167
rect 1762 50164 1768 50176
rect 1719 50136 1768 50164
rect 1719 50133 1731 50136
rect 1673 50127 1731 50133
rect 1762 50124 1768 50136
rect 1820 50124 1826 50176
rect 6273 50167 6331 50173
rect 6273 50133 6285 50167
rect 6319 50164 6331 50167
rect 7742 50164 7748 50176
rect 6319 50136 7748 50164
rect 6319 50133 6331 50136
rect 6273 50127 6331 50133
rect 7742 50124 7748 50136
rect 7800 50124 7806 50176
rect 8938 50124 8944 50176
rect 8996 50164 9002 50176
rect 10045 50167 10103 50173
rect 10045 50164 10057 50167
rect 8996 50136 10057 50164
rect 8996 50124 9002 50136
rect 10045 50133 10057 50136
rect 10091 50133 10103 50167
rect 10045 50127 10103 50133
rect 10505 50167 10563 50173
rect 10505 50133 10517 50167
rect 10551 50164 10563 50167
rect 10778 50164 10784 50176
rect 10551 50136 10784 50164
rect 10551 50133 10563 50136
rect 10505 50127 10563 50133
rect 10778 50124 10784 50136
rect 10836 50124 10842 50176
rect 13998 50124 14004 50176
rect 14056 50164 14062 50176
rect 14461 50167 14519 50173
rect 14461 50164 14473 50167
rect 14056 50136 14473 50164
rect 14056 50124 14062 50136
rect 14461 50133 14473 50136
rect 14507 50133 14519 50167
rect 14461 50127 14519 50133
rect 1104 50074 18860 50096
rect 1104 50022 4315 50074
rect 4367 50022 4379 50074
rect 4431 50022 4443 50074
rect 4495 50022 4507 50074
rect 4559 50022 10982 50074
rect 11034 50022 11046 50074
rect 11098 50022 11110 50074
rect 11162 50022 11174 50074
rect 11226 50022 17648 50074
rect 17700 50022 17712 50074
rect 17764 50022 17776 50074
rect 17828 50022 17840 50074
rect 17892 50022 18860 50074
rect 1104 50000 18860 50022
rect 2222 49960 2228 49972
rect 2183 49932 2228 49960
rect 2222 49920 2228 49932
rect 2280 49920 2286 49972
rect 3513 49963 3571 49969
rect 3513 49929 3525 49963
rect 3559 49960 3571 49963
rect 4154 49960 4160 49972
rect 3559 49932 4160 49960
rect 3559 49929 3571 49932
rect 3513 49923 3571 49929
rect 4154 49920 4160 49932
rect 4212 49920 4218 49972
rect 4893 49963 4951 49969
rect 4893 49929 4905 49963
rect 4939 49960 4951 49963
rect 5810 49960 5816 49972
rect 4939 49932 5816 49960
rect 4939 49929 4951 49932
rect 4893 49923 4951 49929
rect 5810 49920 5816 49932
rect 5868 49920 5874 49972
rect 6454 49920 6460 49972
rect 6512 49960 6518 49972
rect 7926 49960 7932 49972
rect 6512 49932 7932 49960
rect 6512 49920 6518 49932
rect 7926 49920 7932 49932
rect 7984 49920 7990 49972
rect 9214 49960 9220 49972
rect 9175 49932 9220 49960
rect 9214 49920 9220 49932
rect 9272 49920 9278 49972
rect 9493 49963 9551 49969
rect 9493 49929 9505 49963
rect 9539 49960 9551 49963
rect 9582 49960 9588 49972
rect 9539 49932 9588 49960
rect 9539 49929 9551 49932
rect 9493 49923 9551 49929
rect 9582 49920 9588 49932
rect 9640 49920 9646 49972
rect 10134 49920 10140 49972
rect 10192 49960 10198 49972
rect 11882 49960 11888 49972
rect 10192 49932 10456 49960
rect 11843 49932 11888 49960
rect 10192 49920 10198 49932
rect 2240 49824 2268 49920
rect 5166 49852 5172 49904
rect 5224 49852 5230 49904
rect 6086 49892 6092 49904
rect 6047 49864 6092 49892
rect 6086 49852 6092 49864
rect 6144 49852 6150 49904
rect 7006 49852 7012 49904
rect 7064 49892 7070 49904
rect 7101 49895 7159 49901
rect 7101 49892 7113 49895
rect 7064 49864 7113 49892
rect 7064 49852 7070 49864
rect 7101 49861 7113 49864
rect 7147 49892 7159 49895
rect 8478 49892 8484 49904
rect 7147 49864 8484 49892
rect 7147 49861 7159 49864
rect 7101 49855 7159 49861
rect 2777 49827 2835 49833
rect 2240 49796 2728 49824
rect 2498 49756 2504 49768
rect 2459 49728 2504 49756
rect 2498 49716 2504 49728
rect 2556 49716 2562 49768
rect 2700 49756 2728 49796
rect 2777 49793 2789 49827
rect 2823 49824 2835 49827
rect 3234 49824 3240 49836
rect 2823 49796 3240 49824
rect 2823 49793 2835 49796
rect 2777 49787 2835 49793
rect 3234 49784 3240 49796
rect 3292 49824 3298 49836
rect 3789 49827 3847 49833
rect 3789 49824 3801 49827
rect 3292 49796 3801 49824
rect 3292 49784 3298 49796
rect 3789 49793 3801 49796
rect 3835 49793 3847 49827
rect 5184 49824 5212 49852
rect 8110 49824 8116 49836
rect 5184 49796 5396 49824
rect 3789 49787 3847 49793
rect 2961 49759 3019 49765
rect 2961 49756 2973 49759
rect 2700 49728 2973 49756
rect 2961 49725 2973 49728
rect 3007 49725 3019 49759
rect 2961 49719 3019 49725
rect 4525 49759 4583 49765
rect 4525 49725 4537 49759
rect 4571 49756 4583 49759
rect 4982 49756 4988 49768
rect 4571 49728 4988 49756
rect 4571 49725 4583 49728
rect 4525 49719 4583 49725
rect 4982 49716 4988 49728
rect 5040 49716 5046 49768
rect 5166 49756 5172 49768
rect 5127 49728 5172 49756
rect 5166 49716 5172 49728
rect 5224 49716 5230 49768
rect 5368 49756 5396 49796
rect 6932 49796 8116 49824
rect 5629 49759 5687 49765
rect 5629 49756 5641 49759
rect 5368 49728 5641 49756
rect 5629 49725 5641 49728
rect 5675 49725 5687 49759
rect 5629 49719 5687 49725
rect 5721 49759 5779 49765
rect 5721 49725 5733 49759
rect 5767 49756 5779 49759
rect 5810 49756 5816 49768
rect 5767 49728 5816 49756
rect 5767 49725 5779 49728
rect 5721 49719 5779 49725
rect 5810 49716 5816 49728
rect 5868 49756 5874 49768
rect 6362 49756 6368 49768
rect 5868 49728 6368 49756
rect 5868 49716 5874 49728
rect 6362 49716 6368 49728
rect 6420 49716 6426 49768
rect 6086 49648 6092 49700
rect 6144 49688 6150 49700
rect 6270 49688 6276 49700
rect 6144 49660 6276 49688
rect 6144 49648 6150 49660
rect 6270 49648 6276 49660
rect 6328 49648 6334 49700
rect 6822 49648 6828 49700
rect 6880 49688 6886 49700
rect 6932 49688 6960 49796
rect 7006 49716 7012 49768
rect 7064 49756 7070 49768
rect 7193 49759 7251 49765
rect 7193 49756 7205 49759
rect 7064 49728 7205 49756
rect 7064 49716 7070 49728
rect 7193 49725 7205 49728
rect 7239 49725 7251 49759
rect 7193 49719 7251 49725
rect 7466 49716 7472 49768
rect 7524 49756 7530 49768
rect 7742 49756 7748 49768
rect 7524 49728 7748 49756
rect 7524 49716 7530 49728
rect 7742 49716 7748 49728
rect 7800 49716 7806 49768
rect 7834 49716 7840 49768
rect 7892 49756 7898 49768
rect 8036 49765 8064 49796
rect 8110 49784 8116 49796
rect 8168 49784 8174 49836
rect 8220 49768 8248 49864
rect 8478 49852 8484 49864
rect 8536 49852 8542 49904
rect 8570 49852 8576 49904
rect 8628 49892 8634 49904
rect 8846 49892 8852 49904
rect 8628 49864 8852 49892
rect 8628 49852 8634 49864
rect 8846 49852 8852 49864
rect 8904 49852 8910 49904
rect 10134 49824 10140 49836
rect 10095 49796 10140 49824
rect 10134 49784 10140 49796
rect 10192 49784 10198 49836
rect 8021 49759 8079 49765
rect 7892 49728 7937 49756
rect 7892 49716 7898 49728
rect 8021 49725 8033 49759
rect 8067 49725 8079 49759
rect 8202 49756 8208 49768
rect 8163 49728 8208 49756
rect 8021 49719 8079 49725
rect 8202 49716 8208 49728
rect 8260 49716 8266 49768
rect 8478 49756 8484 49768
rect 8312 49728 8484 49756
rect 6880 49660 6960 49688
rect 6880 49648 6886 49660
rect 2314 49580 2320 49632
rect 2372 49620 2378 49632
rect 2866 49620 2872 49632
rect 2372 49592 2872 49620
rect 2372 49580 2378 49592
rect 2866 49580 2872 49592
rect 2924 49580 2930 49632
rect 6733 49623 6791 49629
rect 6733 49589 6745 49623
rect 6779 49620 6791 49623
rect 8312 49620 8340 49728
rect 8478 49716 8484 49728
rect 8536 49716 8542 49768
rect 9033 49759 9091 49765
rect 9033 49725 9045 49759
rect 9079 49756 9091 49759
rect 9398 49756 9404 49768
rect 9079 49728 9404 49756
rect 9079 49725 9091 49728
rect 9033 49719 9091 49725
rect 9398 49716 9404 49728
rect 9456 49716 9462 49768
rect 9674 49756 9680 49768
rect 9635 49728 9680 49756
rect 9674 49716 9680 49728
rect 9732 49716 9738 49768
rect 10318 49756 10324 49768
rect 9784 49728 10324 49756
rect 8754 49648 8760 49700
rect 8812 49688 8818 49700
rect 9784 49688 9812 49728
rect 10318 49716 10324 49728
rect 10376 49716 10382 49768
rect 8812 49660 9812 49688
rect 8812 49648 8818 49660
rect 6779 49592 8340 49620
rect 6779 49589 6791 49592
rect 6733 49583 6791 49589
rect 8846 49580 8852 49632
rect 8904 49620 8910 49632
rect 9217 49623 9275 49629
rect 9217 49620 9229 49623
rect 8904 49592 9229 49620
rect 8904 49580 8910 49592
rect 9217 49589 9229 49592
rect 9263 49620 9275 49623
rect 9309 49623 9367 49629
rect 9309 49620 9321 49623
rect 9263 49592 9321 49620
rect 9263 49589 9275 49592
rect 9217 49583 9275 49589
rect 9309 49589 9321 49592
rect 9355 49589 9367 49623
rect 9309 49583 9367 49589
rect 9493 49623 9551 49629
rect 9493 49589 9505 49623
rect 9539 49620 9551 49623
rect 9674 49620 9680 49632
rect 9539 49592 9680 49620
rect 9539 49589 9551 49592
rect 9493 49583 9551 49589
rect 9674 49580 9680 49592
rect 9732 49580 9738 49632
rect 10428 49620 10456 49932
rect 11882 49920 11888 49932
rect 11940 49920 11946 49972
rect 12434 49960 12440 49972
rect 12395 49932 12440 49960
rect 12434 49920 12440 49932
rect 12492 49920 12498 49972
rect 13173 49963 13231 49969
rect 13173 49929 13185 49963
rect 13219 49960 13231 49963
rect 13354 49960 13360 49972
rect 13219 49932 13360 49960
rect 13219 49929 13231 49932
rect 13173 49923 13231 49929
rect 13354 49920 13360 49932
rect 13412 49920 13418 49972
rect 13541 49963 13599 49969
rect 13541 49929 13553 49963
rect 13587 49960 13599 49963
rect 13633 49963 13691 49969
rect 13633 49960 13645 49963
rect 13587 49932 13645 49960
rect 13587 49929 13599 49932
rect 13541 49923 13599 49929
rect 13633 49929 13645 49932
rect 13679 49960 13691 49963
rect 13906 49960 13912 49972
rect 13679 49932 13912 49960
rect 13679 49929 13691 49932
rect 13633 49923 13691 49929
rect 13906 49920 13912 49932
rect 13964 49920 13970 49972
rect 14826 49920 14832 49972
rect 14884 49960 14890 49972
rect 14921 49963 14979 49969
rect 14921 49960 14933 49963
rect 14884 49932 14933 49960
rect 14884 49920 14890 49932
rect 14921 49929 14933 49932
rect 14967 49929 14979 49963
rect 14921 49923 14979 49929
rect 16022 49920 16028 49972
rect 16080 49960 16086 49972
rect 16390 49960 16396 49972
rect 16080 49932 16396 49960
rect 16080 49920 16086 49932
rect 16390 49920 16396 49932
rect 16448 49920 16454 49972
rect 11054 49824 11060 49836
rect 10612 49796 11060 49824
rect 10612 49768 10640 49796
rect 11054 49784 11060 49796
rect 11112 49784 11118 49836
rect 11900 49824 11928 49920
rect 11974 49852 11980 49904
rect 12032 49892 12038 49904
rect 14645 49895 14703 49901
rect 14645 49892 14657 49895
rect 12032 49864 14657 49892
rect 12032 49852 12038 49864
rect 11900 49796 12204 49824
rect 10594 49756 10600 49768
rect 10555 49728 10600 49756
rect 10594 49716 10600 49728
rect 10652 49716 10658 49768
rect 10778 49716 10784 49768
rect 10836 49756 10842 49768
rect 10965 49759 11023 49765
rect 10965 49756 10977 49759
rect 10836 49728 10977 49756
rect 10836 49716 10842 49728
rect 10965 49725 10977 49728
rect 11011 49725 11023 49759
rect 11514 49756 11520 49768
rect 11475 49728 11520 49756
rect 10965 49719 11023 49725
rect 11514 49716 11520 49728
rect 11572 49716 11578 49768
rect 12066 49756 12072 49768
rect 12027 49728 12072 49756
rect 12066 49716 12072 49728
rect 12124 49716 12130 49768
rect 12176 49765 12204 49796
rect 12268 49765 12296 49864
rect 14645 49861 14657 49864
rect 14691 49861 14703 49895
rect 16206 49892 16212 49904
rect 16167 49864 16212 49892
rect 14645 49855 14703 49861
rect 16206 49852 16212 49864
rect 16264 49852 16270 49904
rect 16666 49892 16672 49904
rect 16500 49864 16672 49892
rect 12434 49784 12440 49836
rect 12492 49824 12498 49836
rect 12802 49824 12808 49836
rect 12492 49796 12808 49824
rect 12492 49784 12498 49796
rect 12802 49784 12808 49796
rect 12860 49784 12866 49836
rect 12894 49784 12900 49836
rect 12952 49824 12958 49836
rect 13170 49824 13176 49836
rect 12952 49796 13176 49824
rect 12952 49784 12958 49796
rect 13170 49784 13176 49796
rect 13228 49784 13234 49836
rect 14090 49824 14096 49836
rect 13924 49796 14096 49824
rect 13924 49765 13952 49796
rect 14090 49784 14096 49796
rect 14148 49824 14154 49836
rect 15378 49824 15384 49836
rect 14148 49796 15384 49824
rect 14148 49784 14154 49796
rect 15378 49784 15384 49796
rect 15436 49784 15442 49836
rect 12161 49759 12219 49765
rect 12161 49725 12173 49759
rect 12207 49725 12219 49759
rect 12161 49719 12219 49725
rect 12253 49759 12311 49765
rect 12253 49725 12265 49759
rect 12299 49725 12311 49759
rect 13817 49759 13875 49765
rect 13817 49756 13829 49759
rect 12253 49719 12311 49725
rect 13740 49728 13829 49756
rect 13740 49688 13768 49728
rect 13817 49725 13829 49728
rect 13863 49725 13875 49759
rect 13817 49719 13875 49725
rect 13909 49759 13967 49765
rect 13909 49725 13921 49759
rect 13955 49725 13967 49759
rect 13909 49719 13967 49725
rect 15102 49716 15108 49768
rect 15160 49756 15166 49768
rect 15289 49759 15347 49765
rect 15289 49756 15301 49759
rect 15160 49728 15301 49756
rect 15160 49716 15166 49728
rect 15289 49725 15301 49728
rect 15335 49756 15347 49759
rect 15749 49759 15807 49765
rect 15749 49756 15761 49759
rect 15335 49728 15761 49756
rect 15335 49725 15347 49728
rect 15289 49719 15347 49725
rect 15749 49725 15761 49728
rect 15795 49725 15807 49759
rect 15749 49719 15807 49725
rect 16298 49716 16304 49768
rect 16356 49756 16362 49768
rect 16500 49756 16528 49864
rect 16666 49852 16672 49864
rect 16724 49852 16730 49904
rect 17589 49827 17647 49833
rect 17589 49824 17601 49827
rect 16356 49728 16528 49756
rect 16592 49796 17601 49824
rect 16356 49716 16362 49728
rect 13648 49660 13768 49688
rect 14369 49691 14427 49697
rect 13648 49632 13676 49660
rect 14369 49657 14381 49691
rect 14415 49688 14427 49691
rect 14826 49688 14832 49700
rect 14415 49660 14832 49688
rect 14415 49657 14427 49660
rect 14369 49651 14427 49657
rect 14826 49648 14832 49660
rect 14884 49648 14890 49700
rect 16206 49648 16212 49700
rect 16264 49688 16270 49700
rect 16592 49688 16620 49796
rect 17589 49793 17601 49796
rect 17635 49793 17647 49827
rect 17589 49787 17647 49793
rect 16669 49759 16727 49765
rect 16669 49725 16681 49759
rect 16715 49725 16727 49759
rect 17218 49756 17224 49768
rect 17179 49728 17224 49756
rect 16669 49719 16727 49725
rect 16264 49660 16620 49688
rect 16264 49648 16270 49660
rect 10502 49620 10508 49632
rect 10428 49592 10508 49620
rect 10502 49580 10508 49592
rect 10560 49580 10566 49632
rect 13630 49580 13636 49632
rect 13688 49580 13694 49632
rect 14921 49623 14979 49629
rect 14921 49589 14933 49623
rect 14967 49620 14979 49623
rect 15010 49620 15016 49632
rect 14967 49592 15016 49620
rect 14967 49589 14979 49592
rect 14921 49583 14979 49589
rect 15010 49580 15016 49592
rect 15068 49620 15074 49632
rect 15473 49623 15531 49629
rect 15473 49620 15485 49623
rect 15068 49592 15485 49620
rect 15068 49580 15074 49592
rect 15473 49589 15485 49592
rect 15519 49589 15531 49623
rect 15473 49583 15531 49589
rect 16577 49623 16635 49629
rect 16577 49589 16589 49623
rect 16623 49620 16635 49623
rect 16684 49620 16712 49719
rect 17218 49716 17224 49728
rect 17276 49716 17282 49768
rect 17494 49756 17500 49768
rect 17455 49728 17500 49756
rect 17494 49716 17500 49728
rect 17552 49716 17558 49768
rect 16758 49620 16764 49632
rect 16623 49592 16764 49620
rect 16623 49589 16635 49592
rect 16577 49583 16635 49589
rect 16758 49580 16764 49592
rect 16816 49580 16822 49632
rect 1104 49530 18860 49552
rect 1104 49478 7648 49530
rect 7700 49478 7712 49530
rect 7764 49478 7776 49530
rect 7828 49478 7840 49530
rect 7892 49478 14315 49530
rect 14367 49478 14379 49530
rect 14431 49478 14443 49530
rect 14495 49478 14507 49530
rect 14559 49478 18860 49530
rect 1104 49456 18860 49478
rect 2498 49416 2504 49428
rect 2459 49388 2504 49416
rect 2498 49376 2504 49388
rect 2556 49416 2562 49428
rect 4525 49419 4583 49425
rect 4525 49416 4537 49419
rect 2556 49388 4537 49416
rect 2556 49376 2562 49388
rect 4525 49385 4537 49388
rect 4571 49385 4583 49419
rect 6270 49416 6276 49428
rect 6231 49388 6276 49416
rect 4525 49379 4583 49385
rect 6270 49376 6276 49388
rect 6328 49376 6334 49428
rect 6641 49419 6699 49425
rect 6641 49385 6653 49419
rect 6687 49416 6699 49419
rect 6822 49416 6828 49428
rect 6687 49388 6828 49416
rect 6687 49385 6699 49388
rect 6641 49379 6699 49385
rect 6822 49376 6828 49388
rect 6880 49376 6886 49428
rect 8754 49416 8760 49428
rect 8715 49388 8760 49416
rect 8754 49376 8760 49388
rect 8812 49376 8818 49428
rect 9493 49419 9551 49425
rect 9493 49385 9505 49419
rect 9539 49416 9551 49419
rect 9950 49416 9956 49428
rect 9539 49388 9956 49416
rect 9539 49385 9551 49388
rect 9493 49379 9551 49385
rect 9950 49376 9956 49388
rect 10008 49416 10014 49428
rect 10134 49416 10140 49428
rect 10008 49388 10140 49416
rect 10008 49376 10014 49388
rect 10134 49376 10140 49388
rect 10192 49416 10198 49428
rect 10413 49419 10471 49425
rect 10413 49416 10425 49419
rect 10192 49388 10425 49416
rect 10192 49376 10198 49388
rect 10413 49385 10425 49388
rect 10459 49385 10471 49419
rect 10413 49379 10471 49385
rect 11054 49376 11060 49428
rect 11112 49416 11118 49428
rect 11149 49419 11207 49425
rect 11149 49416 11161 49419
rect 11112 49388 11161 49416
rect 11112 49376 11118 49388
rect 11149 49385 11161 49388
rect 11195 49385 11207 49419
rect 12066 49416 12072 49428
rect 12027 49388 12072 49416
rect 11149 49379 11207 49385
rect 12066 49376 12072 49388
rect 12124 49416 12130 49428
rect 14090 49416 14096 49428
rect 12124 49388 12664 49416
rect 14051 49388 14096 49416
rect 12124 49376 12130 49388
rect 5905 49351 5963 49357
rect 5905 49317 5917 49351
rect 5951 49348 5963 49351
rect 8389 49351 8447 49357
rect 5951 49320 7880 49348
rect 5951 49317 5963 49320
rect 5905 49311 5963 49317
rect 3053 49283 3111 49289
rect 3053 49249 3065 49283
rect 3099 49280 3111 49283
rect 3421 49283 3479 49289
rect 3421 49280 3433 49283
rect 3099 49252 3433 49280
rect 3099 49249 3111 49252
rect 3053 49243 3111 49249
rect 3421 49249 3433 49252
rect 3467 49280 3479 49283
rect 3510 49280 3516 49292
rect 3467 49252 3516 49280
rect 3467 49249 3479 49252
rect 3421 49243 3479 49249
rect 3510 49240 3516 49252
rect 3568 49280 3574 49292
rect 4062 49280 4068 49292
rect 3568 49252 4068 49280
rect 3568 49240 3574 49252
rect 4062 49240 4068 49252
rect 4120 49240 4126 49292
rect 6825 49283 6883 49289
rect 6825 49249 6837 49283
rect 6871 49280 6883 49283
rect 6914 49280 6920 49292
rect 6871 49252 6920 49280
rect 6871 49249 6883 49252
rect 6825 49243 6883 49249
rect 6914 49240 6920 49252
rect 6972 49240 6978 49292
rect 7006 49240 7012 49292
rect 7064 49280 7070 49292
rect 7852 49289 7880 49320
rect 8389 49317 8401 49351
rect 8435 49348 8447 49351
rect 9582 49348 9588 49360
rect 8435 49320 9588 49348
rect 8435 49317 8447 49320
rect 8389 49311 8447 49317
rect 9582 49308 9588 49320
rect 9640 49308 9646 49360
rect 10505 49351 10563 49357
rect 10505 49317 10517 49351
rect 10551 49348 10563 49351
rect 10594 49348 10600 49360
rect 10551 49320 10600 49348
rect 10551 49317 10563 49320
rect 10505 49311 10563 49317
rect 10594 49308 10600 49320
rect 10652 49308 10658 49360
rect 10686 49308 10692 49360
rect 10744 49348 10750 49360
rect 12636 49357 12664 49388
rect 14090 49376 14096 49388
rect 14148 49376 14154 49428
rect 15562 49376 15568 49428
rect 15620 49416 15626 49428
rect 15933 49419 15991 49425
rect 15933 49416 15945 49419
rect 15620 49388 15945 49416
rect 15620 49376 15626 49388
rect 15933 49385 15945 49388
rect 15979 49385 15991 49419
rect 17494 49416 17500 49428
rect 17455 49388 17500 49416
rect 15933 49379 15991 49385
rect 17494 49376 17500 49388
rect 17552 49376 17558 49428
rect 10873 49351 10931 49357
rect 10873 49348 10885 49351
rect 10744 49320 10885 49348
rect 10744 49308 10750 49320
rect 10873 49317 10885 49320
rect 10919 49317 10931 49351
rect 10873 49311 10931 49317
rect 12621 49351 12679 49357
rect 12621 49317 12633 49351
rect 12667 49317 12679 49351
rect 12621 49311 12679 49317
rect 13722 49308 13728 49360
rect 13780 49348 13786 49360
rect 14369 49351 14427 49357
rect 14369 49348 14381 49351
rect 13780 49320 14381 49348
rect 13780 49308 13786 49320
rect 14369 49317 14381 49320
rect 14415 49317 14427 49351
rect 14734 49348 14740 49360
rect 14695 49320 14740 49348
rect 14369 49311 14427 49317
rect 14734 49308 14740 49320
rect 14792 49308 14798 49360
rect 15010 49348 15016 49360
rect 14936 49320 15016 49348
rect 7469 49283 7527 49289
rect 7469 49280 7481 49283
rect 7064 49252 7481 49280
rect 7064 49240 7070 49252
rect 7469 49249 7481 49252
rect 7515 49249 7527 49283
rect 7469 49243 7527 49249
rect 7837 49283 7895 49289
rect 7837 49249 7849 49283
rect 7883 49280 7895 49283
rect 8110 49280 8116 49292
rect 7883 49252 8116 49280
rect 7883 49249 7895 49252
rect 7837 49243 7895 49249
rect 8110 49240 8116 49252
rect 8168 49240 8174 49292
rect 8846 49280 8852 49292
rect 8807 49252 8852 49280
rect 8846 49240 8852 49252
rect 8904 49240 8910 49292
rect 10042 49240 10048 49292
rect 10100 49280 10106 49292
rect 10321 49283 10379 49289
rect 10321 49280 10333 49283
rect 10100 49252 10333 49280
rect 10100 49240 10106 49252
rect 10321 49249 10333 49252
rect 10367 49249 10379 49283
rect 10321 49243 10379 49249
rect 11974 49240 11980 49292
rect 12032 49280 12038 49292
rect 12250 49280 12256 49292
rect 12032 49252 12256 49280
rect 12032 49240 12038 49252
rect 12250 49240 12256 49252
rect 12308 49280 12314 49292
rect 12437 49283 12495 49289
rect 12437 49280 12449 49283
rect 12308 49252 12449 49280
rect 12308 49240 12314 49252
rect 12437 49249 12449 49252
rect 12483 49249 12495 49283
rect 12710 49280 12716 49292
rect 12671 49252 12716 49280
rect 12437 49243 12495 49249
rect 12710 49240 12716 49252
rect 12768 49240 12774 49292
rect 14090 49240 14096 49292
rect 14148 49280 14154 49292
rect 14829 49283 14887 49289
rect 14829 49280 14841 49283
rect 14148 49252 14841 49280
rect 14148 49240 14154 49252
rect 14829 49249 14841 49252
rect 14875 49249 14887 49283
rect 14829 49243 14887 49249
rect 2406 49172 2412 49224
rect 2464 49212 2470 49224
rect 3145 49215 3203 49221
rect 3145 49212 3157 49215
rect 2464 49184 3157 49212
rect 2464 49172 2470 49184
rect 3145 49181 3157 49184
rect 3191 49181 3203 49215
rect 7558 49212 7564 49224
rect 7519 49184 7564 49212
rect 3145 49175 3203 49181
rect 7558 49172 7564 49184
rect 7616 49172 7622 49224
rect 7926 49212 7932 49224
rect 7887 49184 7932 49212
rect 7926 49172 7932 49184
rect 7984 49172 7990 49224
rect 9674 49172 9680 49224
rect 9732 49212 9738 49224
rect 10137 49215 10195 49221
rect 10137 49212 10149 49215
rect 9732 49184 10149 49212
rect 9732 49172 9738 49184
rect 10137 49181 10149 49184
rect 10183 49212 10195 49215
rect 11422 49212 11428 49224
rect 10183 49184 11428 49212
rect 10183 49181 10195 49184
rect 10137 49175 10195 49181
rect 11422 49172 11428 49184
rect 11480 49172 11486 49224
rect 12526 49172 12532 49224
rect 12584 49212 12590 49224
rect 12802 49212 12808 49224
rect 12584 49184 12808 49212
rect 12584 49172 12590 49184
rect 12802 49172 12808 49184
rect 12860 49172 12866 49224
rect 14274 49172 14280 49224
rect 14332 49212 14338 49224
rect 14936 49212 14964 49320
rect 15010 49308 15016 49320
rect 15068 49308 15074 49360
rect 15286 49348 15292 49360
rect 15247 49320 15292 49348
rect 15286 49308 15292 49320
rect 15344 49308 15350 49360
rect 15378 49308 15384 49360
rect 15436 49348 15442 49360
rect 15657 49351 15715 49357
rect 15657 49348 15669 49351
rect 15436 49320 15669 49348
rect 15436 49308 15442 49320
rect 15657 49317 15669 49320
rect 15703 49348 15715 49351
rect 15746 49348 15752 49360
rect 15703 49320 15752 49348
rect 15703 49317 15715 49320
rect 15657 49311 15715 49317
rect 15746 49308 15752 49320
rect 15804 49308 15810 49360
rect 16666 49308 16672 49360
rect 16724 49348 16730 49360
rect 16724 49320 17172 49348
rect 16724 49308 16730 49320
rect 16758 49240 16764 49292
rect 16816 49280 16822 49292
rect 17144 49289 17172 49320
rect 16945 49283 17003 49289
rect 16945 49280 16957 49283
rect 16816 49252 16957 49280
rect 16816 49240 16822 49252
rect 16945 49249 16957 49252
rect 16991 49249 17003 49283
rect 16945 49243 17003 49249
rect 17129 49283 17187 49289
rect 17129 49249 17141 49283
rect 17175 49280 17187 49283
rect 17494 49280 17500 49292
rect 17175 49252 17500 49280
rect 17175 49249 17187 49252
rect 17129 49243 17187 49249
rect 17494 49240 17500 49252
rect 17552 49240 17558 49292
rect 14332 49184 14964 49212
rect 14332 49172 14338 49184
rect 15010 49172 15016 49224
rect 15068 49212 15074 49224
rect 16117 49215 16175 49221
rect 16117 49212 16129 49215
rect 15068 49184 16129 49212
rect 15068 49172 15074 49184
rect 16117 49181 16129 49184
rect 16163 49181 16175 49215
rect 16666 49212 16672 49224
rect 16627 49184 16672 49212
rect 16117 49175 16175 49181
rect 16666 49172 16672 49184
rect 16724 49172 16730 49224
rect 5534 49144 5540 49156
rect 5495 49116 5540 49144
rect 5534 49104 5540 49116
rect 5592 49104 5598 49156
rect 10686 49104 10692 49156
rect 10744 49144 10750 49156
rect 10962 49144 10968 49156
rect 10744 49116 10968 49144
rect 10744 49104 10750 49116
rect 10962 49104 10968 49116
rect 11020 49104 11026 49156
rect 1578 49076 1584 49088
rect 1539 49048 1584 49076
rect 1578 49036 1584 49048
rect 1636 49036 1642 49088
rect 5166 49076 5172 49088
rect 5127 49048 5172 49076
rect 5166 49036 5172 49048
rect 5224 49036 5230 49088
rect 8294 49036 8300 49088
rect 8352 49076 8358 49088
rect 9033 49079 9091 49085
rect 9033 49076 9045 49079
rect 8352 49048 9045 49076
rect 8352 49036 8358 49048
rect 9033 49045 9045 49048
rect 9079 49045 9091 49079
rect 9033 49039 9091 49045
rect 9861 49079 9919 49085
rect 9861 49045 9873 49079
rect 9907 49076 9919 49079
rect 10318 49076 10324 49088
rect 9907 49048 10324 49076
rect 9907 49045 9919 49048
rect 9861 49039 9919 49045
rect 10318 49036 10324 49048
rect 10376 49036 10382 49088
rect 11606 49076 11612 49088
rect 11567 49048 11612 49076
rect 11606 49036 11612 49048
rect 11664 49036 11670 49088
rect 12894 49076 12900 49088
rect 12855 49048 12900 49076
rect 12894 49036 12900 49048
rect 12952 49036 12958 49088
rect 13630 49076 13636 49088
rect 13591 49048 13636 49076
rect 13630 49036 13636 49048
rect 13688 49036 13694 49088
rect 13906 49036 13912 49088
rect 13964 49076 13970 49088
rect 14550 49076 14556 49088
rect 13964 49048 14556 49076
rect 13964 49036 13970 49048
rect 14550 49036 14556 49048
rect 14608 49036 14614 49088
rect 1104 48986 18860 49008
rect 1104 48934 4315 48986
rect 4367 48934 4379 48986
rect 4431 48934 4443 48986
rect 4495 48934 4507 48986
rect 4559 48934 10982 48986
rect 11034 48934 11046 48986
rect 11098 48934 11110 48986
rect 11162 48934 11174 48986
rect 11226 48934 17648 48986
rect 17700 48934 17712 48986
rect 17764 48934 17776 48986
rect 17828 48934 17840 48986
rect 17892 48934 18860 48986
rect 1104 48912 18860 48934
rect 3053 48875 3111 48881
rect 3053 48841 3065 48875
rect 3099 48872 3111 48875
rect 3234 48872 3240 48884
rect 3099 48844 3240 48872
rect 3099 48841 3111 48844
rect 3053 48835 3111 48841
rect 3234 48832 3240 48844
rect 3292 48832 3298 48884
rect 3510 48872 3516 48884
rect 3471 48844 3516 48872
rect 3510 48832 3516 48844
rect 3568 48832 3574 48884
rect 4893 48875 4951 48881
rect 4893 48841 4905 48875
rect 4939 48872 4951 48875
rect 5074 48872 5080 48884
rect 4939 48844 5080 48872
rect 4939 48841 4951 48844
rect 4893 48835 4951 48841
rect 5074 48832 5080 48844
rect 5132 48832 5138 48884
rect 7282 48832 7288 48884
rect 7340 48872 7346 48884
rect 8205 48875 8263 48881
rect 8205 48872 8217 48875
rect 7340 48844 8217 48872
rect 7340 48832 7346 48844
rect 8205 48841 8217 48844
rect 8251 48841 8263 48875
rect 8205 48835 8263 48841
rect 10502 48832 10508 48884
rect 10560 48832 10566 48884
rect 10594 48832 10600 48884
rect 10652 48872 10658 48884
rect 10652 48844 11376 48872
rect 10652 48832 10658 48844
rect 5994 48764 6000 48816
rect 6052 48804 6058 48816
rect 6270 48804 6276 48816
rect 6052 48776 6276 48804
rect 6052 48764 6058 48776
rect 6270 48764 6276 48776
rect 6328 48764 6334 48816
rect 7558 48804 7564 48816
rect 7484 48776 7564 48804
rect 1489 48739 1547 48745
rect 1489 48705 1501 48739
rect 1535 48736 1547 48739
rect 1670 48736 1676 48748
rect 1535 48708 1676 48736
rect 1535 48705 1547 48708
rect 1489 48699 1547 48705
rect 1670 48696 1676 48708
rect 1728 48736 1734 48748
rect 1728 48708 2084 48736
rect 1728 48696 1734 48708
rect 2056 48680 2084 48708
rect 3694 48696 3700 48748
rect 3752 48736 3758 48748
rect 5074 48736 5080 48748
rect 3752 48708 5080 48736
rect 3752 48696 3758 48708
rect 5074 48696 5080 48708
rect 5132 48696 5138 48748
rect 5166 48696 5172 48748
rect 5224 48736 5230 48748
rect 6733 48739 6791 48745
rect 6733 48736 6745 48739
rect 5224 48708 6745 48736
rect 5224 48696 5230 48708
rect 6733 48705 6745 48708
rect 6779 48705 6791 48739
rect 6733 48699 6791 48705
rect 6914 48696 6920 48748
rect 6972 48736 6978 48748
rect 7484 48745 7512 48776
rect 7558 48764 7564 48776
rect 7616 48764 7622 48816
rect 10520 48804 10548 48832
rect 11054 48804 11060 48816
rect 10520 48776 11060 48804
rect 11054 48764 11060 48776
rect 11112 48764 11118 48816
rect 7469 48739 7527 48745
rect 7469 48736 7481 48739
rect 6972 48708 7481 48736
rect 6972 48696 6978 48708
rect 7469 48705 7481 48708
rect 7515 48705 7527 48739
rect 10594 48736 10600 48748
rect 10555 48708 10600 48736
rect 7469 48699 7527 48705
rect 10594 48696 10600 48708
rect 10652 48696 10658 48748
rect 1578 48628 1584 48680
rect 1636 48668 1642 48680
rect 1765 48671 1823 48677
rect 1765 48668 1777 48671
rect 1636 48640 1777 48668
rect 1636 48628 1642 48640
rect 1765 48637 1777 48640
rect 1811 48637 1823 48671
rect 1765 48631 1823 48637
rect 2038 48628 2044 48680
rect 2096 48628 2102 48680
rect 4890 48668 4896 48680
rect 4851 48640 4896 48668
rect 4890 48628 4896 48640
rect 4948 48628 4954 48680
rect 5350 48668 5356 48680
rect 5311 48640 5356 48668
rect 5350 48628 5356 48640
rect 5408 48628 5414 48680
rect 6273 48671 6331 48677
rect 6273 48637 6285 48671
rect 6319 48668 6331 48671
rect 6641 48671 6699 48677
rect 6641 48668 6653 48671
rect 6319 48640 6653 48668
rect 6319 48637 6331 48640
rect 6273 48631 6331 48637
rect 6641 48637 6653 48640
rect 6687 48668 6699 48671
rect 6822 48668 6828 48680
rect 6687 48640 6828 48668
rect 6687 48637 6699 48640
rect 6641 48631 6699 48637
rect 6822 48628 6828 48640
rect 6880 48628 6886 48680
rect 7282 48628 7288 48680
rect 7340 48668 7346 48680
rect 7377 48671 7435 48677
rect 7377 48668 7389 48671
rect 7340 48640 7389 48668
rect 7340 48628 7346 48640
rect 7377 48637 7389 48640
rect 7423 48637 7435 48671
rect 7742 48668 7748 48680
rect 7703 48640 7748 48668
rect 7377 48631 7435 48637
rect 7742 48628 7748 48640
rect 7800 48628 7806 48680
rect 7837 48671 7895 48677
rect 7837 48637 7849 48671
rect 7883 48668 7895 48671
rect 7926 48668 7932 48680
rect 7883 48640 7932 48668
rect 7883 48637 7895 48640
rect 7837 48631 7895 48637
rect 4709 48603 4767 48609
rect 4709 48569 4721 48603
rect 4755 48600 4767 48603
rect 5368 48600 5396 48628
rect 4755 48572 5396 48600
rect 6840 48600 6868 48628
rect 7852 48600 7880 48631
rect 7926 48628 7932 48640
rect 7984 48628 7990 48680
rect 9493 48671 9551 48677
rect 9493 48637 9505 48671
rect 9539 48668 9551 48671
rect 9582 48668 9588 48680
rect 9539 48640 9588 48668
rect 9539 48637 9551 48640
rect 9493 48631 9551 48637
rect 9582 48628 9588 48640
rect 9640 48628 9646 48680
rect 9858 48668 9864 48680
rect 9819 48640 9864 48668
rect 9858 48628 9864 48640
rect 9916 48628 9922 48680
rect 10134 48668 10140 48680
rect 10095 48640 10140 48668
rect 10134 48628 10140 48640
rect 10192 48628 10198 48680
rect 10318 48628 10324 48680
rect 10376 48668 10382 48680
rect 10781 48671 10839 48677
rect 10781 48668 10793 48671
rect 10376 48640 10793 48668
rect 10376 48628 10382 48640
rect 10781 48637 10793 48640
rect 10827 48668 10839 48671
rect 10962 48668 10968 48680
rect 10827 48640 10968 48668
rect 10827 48637 10839 48640
rect 10781 48631 10839 48637
rect 10962 48628 10968 48640
rect 11020 48628 11026 48680
rect 11238 48668 11244 48680
rect 11199 48640 11244 48668
rect 11238 48628 11244 48640
rect 11296 48628 11302 48680
rect 11348 48668 11376 48844
rect 11422 48832 11428 48884
rect 11480 48872 11486 48884
rect 11517 48875 11575 48881
rect 11517 48872 11529 48875
rect 11480 48844 11529 48872
rect 11480 48832 11486 48844
rect 11517 48841 11529 48844
rect 11563 48841 11575 48875
rect 11517 48835 11575 48841
rect 11532 48736 11560 48835
rect 12066 48832 12072 48884
rect 12124 48872 12130 48884
rect 12253 48875 12311 48881
rect 12253 48872 12265 48875
rect 12124 48844 12265 48872
rect 12124 48832 12130 48844
rect 12253 48841 12265 48844
rect 12299 48841 12311 48875
rect 12253 48835 12311 48841
rect 12268 48804 12296 48835
rect 12434 48832 12440 48884
rect 12492 48872 12498 48884
rect 12894 48872 12900 48884
rect 12492 48844 12900 48872
rect 12492 48832 12498 48844
rect 12894 48832 12900 48844
rect 12952 48832 12958 48884
rect 14277 48875 14335 48881
rect 14277 48841 14289 48875
rect 14323 48872 14335 48875
rect 14734 48872 14740 48884
rect 14323 48844 14740 48872
rect 14323 48841 14335 48844
rect 14277 48835 14335 48841
rect 14734 48832 14740 48844
rect 14792 48832 14798 48884
rect 14826 48832 14832 48884
rect 14884 48872 14890 48884
rect 15013 48875 15071 48881
rect 15013 48872 15025 48875
rect 14884 48844 15025 48872
rect 14884 48832 14890 48844
rect 15013 48841 15025 48844
rect 15059 48841 15071 48875
rect 15013 48835 15071 48841
rect 15473 48875 15531 48881
rect 15473 48841 15485 48875
rect 15519 48872 15531 48875
rect 15562 48872 15568 48884
rect 15519 48844 15568 48872
rect 15519 48841 15531 48844
rect 15473 48835 15531 48841
rect 15562 48832 15568 48844
rect 15620 48832 15626 48884
rect 13265 48807 13323 48813
rect 13265 48804 13277 48807
rect 12268 48776 13277 48804
rect 13265 48773 13277 48776
rect 13311 48773 13323 48807
rect 13265 48767 13323 48773
rect 12434 48736 12440 48748
rect 11532 48708 12440 48736
rect 12434 48696 12440 48708
rect 12492 48696 12498 48748
rect 13354 48696 13360 48748
rect 13412 48736 13418 48748
rect 14826 48736 14832 48748
rect 13412 48708 14832 48736
rect 13412 48696 13418 48708
rect 14826 48696 14832 48708
rect 14884 48696 14890 48748
rect 16666 48696 16672 48748
rect 16724 48736 16730 48748
rect 17310 48736 17316 48748
rect 16724 48708 17316 48736
rect 16724 48696 16730 48708
rect 17310 48696 17316 48708
rect 17368 48696 17374 48748
rect 17494 48696 17500 48748
rect 17552 48736 17558 48748
rect 17773 48739 17831 48745
rect 17773 48736 17785 48739
rect 17552 48708 17785 48736
rect 17552 48696 17558 48708
rect 17773 48705 17785 48708
rect 17819 48705 17831 48739
rect 17773 48699 17831 48705
rect 11885 48671 11943 48677
rect 11885 48668 11897 48671
rect 11348 48640 11897 48668
rect 11885 48637 11897 48640
rect 11931 48637 11943 48671
rect 11885 48631 11943 48637
rect 12069 48671 12127 48677
rect 12069 48637 12081 48671
rect 12115 48668 12127 48671
rect 12250 48668 12256 48680
rect 12115 48640 12256 48668
rect 12115 48637 12127 48640
rect 12069 48631 12127 48637
rect 12250 48628 12256 48640
rect 12308 48668 12314 48680
rect 12897 48671 12955 48677
rect 12897 48668 12909 48671
rect 12308 48640 12909 48668
rect 12308 48628 12314 48640
rect 12897 48637 12909 48640
rect 12943 48637 12955 48671
rect 15286 48668 15292 48680
rect 15247 48640 15292 48668
rect 12897 48631 12955 48637
rect 15286 48628 15292 48640
rect 15344 48668 15350 48680
rect 15749 48671 15807 48677
rect 15749 48668 15761 48671
rect 15344 48640 15761 48668
rect 15344 48628 15350 48640
rect 15749 48637 15761 48640
rect 15795 48668 15807 48671
rect 16298 48668 16304 48680
rect 15795 48640 16304 48668
rect 15795 48637 15807 48640
rect 15749 48631 15807 48637
rect 16298 48628 16304 48640
rect 16356 48628 16362 48680
rect 17589 48671 17647 48677
rect 17589 48637 17601 48671
rect 17635 48637 17647 48671
rect 17589 48631 17647 48637
rect 6840 48572 7880 48600
rect 4755 48569 4767 48572
rect 4709 48563 4767 48569
rect 11974 48560 11980 48612
rect 12032 48600 12038 48612
rect 12529 48603 12587 48609
rect 12529 48600 12541 48603
rect 12032 48572 12541 48600
rect 12032 48560 12038 48572
rect 12529 48569 12541 48572
rect 12575 48569 12587 48603
rect 12529 48563 12587 48569
rect 14550 48560 14556 48612
rect 14608 48560 14614 48612
rect 16209 48603 16267 48609
rect 16209 48569 16221 48603
rect 16255 48600 16267 48603
rect 16666 48600 16672 48612
rect 16255 48572 16672 48600
rect 16255 48569 16267 48572
rect 16209 48563 16267 48569
rect 16666 48560 16672 48572
rect 16724 48560 16730 48612
rect 16761 48603 16819 48609
rect 16761 48569 16773 48603
rect 16807 48600 16819 48603
rect 17494 48600 17500 48612
rect 16807 48572 17500 48600
rect 16807 48569 16819 48572
rect 16761 48563 16819 48569
rect 17494 48560 17500 48572
rect 17552 48560 17558 48612
rect 2406 48492 2412 48544
rect 2464 48532 2470 48544
rect 3789 48535 3847 48541
rect 3789 48532 3801 48535
rect 2464 48504 3801 48532
rect 2464 48492 2470 48504
rect 3789 48501 3801 48504
rect 3835 48501 3847 48535
rect 3789 48495 3847 48501
rect 5905 48535 5963 48541
rect 5905 48501 5917 48535
rect 5951 48532 5963 48535
rect 6914 48532 6920 48544
rect 5951 48504 6920 48532
rect 5951 48501 5963 48504
rect 5905 48495 5963 48501
rect 6914 48492 6920 48504
rect 6972 48492 6978 48544
rect 8846 48492 8852 48544
rect 8904 48532 8910 48544
rect 8941 48535 8999 48541
rect 8941 48532 8953 48535
rect 8904 48504 8953 48532
rect 8904 48492 8910 48504
rect 8941 48501 8953 48504
rect 8987 48532 8999 48535
rect 9582 48532 9588 48544
rect 8987 48504 9588 48532
rect 8987 48501 8999 48504
rect 8941 48495 8999 48501
rect 9582 48492 9588 48504
rect 9640 48492 9646 48544
rect 13538 48492 13544 48544
rect 13596 48532 13602 48544
rect 13817 48535 13875 48541
rect 13817 48532 13829 48535
rect 13596 48504 13829 48532
rect 13596 48492 13602 48504
rect 13817 48501 13829 48504
rect 13863 48532 13875 48535
rect 14090 48532 14096 48544
rect 13863 48504 14096 48532
rect 13863 48501 13875 48504
rect 13817 48495 13875 48501
rect 14090 48492 14096 48504
rect 14148 48492 14154 48544
rect 14568 48532 14596 48560
rect 14645 48535 14703 48541
rect 14645 48532 14657 48535
rect 14568 48504 14657 48532
rect 14645 48501 14657 48504
rect 14691 48532 14703 48535
rect 14734 48532 14740 48544
rect 14691 48504 14740 48532
rect 14691 48501 14703 48504
rect 14645 48495 14703 48501
rect 14734 48492 14740 48504
rect 14792 48492 14798 48544
rect 16574 48532 16580 48544
rect 16535 48504 16580 48532
rect 16574 48492 16580 48504
rect 16632 48532 16638 48544
rect 17604 48532 17632 48631
rect 16632 48504 17632 48532
rect 16632 48492 16638 48504
rect 1104 48442 18860 48464
rect 1104 48390 7648 48442
rect 7700 48390 7712 48442
rect 7764 48390 7776 48442
rect 7828 48390 7840 48442
rect 7892 48390 14315 48442
rect 14367 48390 14379 48442
rect 14431 48390 14443 48442
rect 14495 48390 14507 48442
rect 14559 48390 18860 48442
rect 1104 48368 18860 48390
rect 3418 48288 3424 48340
rect 3476 48328 3482 48340
rect 3694 48328 3700 48340
rect 3476 48300 3700 48328
rect 3476 48288 3482 48300
rect 3694 48288 3700 48300
rect 3752 48288 3758 48340
rect 6273 48331 6331 48337
rect 6273 48297 6285 48331
rect 6319 48328 6331 48331
rect 7374 48328 7380 48340
rect 6319 48300 7380 48328
rect 6319 48297 6331 48300
rect 6273 48291 6331 48297
rect 7374 48288 7380 48300
rect 7432 48328 7438 48340
rect 8110 48328 8116 48340
rect 7432 48300 8116 48328
rect 7432 48288 7438 48300
rect 8110 48288 8116 48300
rect 8168 48288 8174 48340
rect 8386 48288 8392 48340
rect 8444 48328 8450 48340
rect 8846 48328 8852 48340
rect 8444 48300 8852 48328
rect 8444 48288 8450 48300
rect 8846 48288 8852 48300
rect 8904 48288 8910 48340
rect 9125 48331 9183 48337
rect 9125 48297 9137 48331
rect 9171 48328 9183 48331
rect 10134 48328 10140 48340
rect 9171 48300 10140 48328
rect 9171 48297 9183 48300
rect 9125 48291 9183 48297
rect 10134 48288 10140 48300
rect 10192 48288 10198 48340
rect 10318 48288 10324 48340
rect 10376 48328 10382 48340
rect 10686 48328 10692 48340
rect 10376 48300 10692 48328
rect 10376 48288 10382 48300
rect 10686 48288 10692 48300
rect 10744 48288 10750 48340
rect 11238 48328 11244 48340
rect 11072 48300 11244 48328
rect 6641 48263 6699 48269
rect 6641 48229 6653 48263
rect 6687 48260 6699 48263
rect 7006 48260 7012 48272
rect 6687 48232 7012 48260
rect 6687 48229 6699 48232
rect 6641 48223 6699 48229
rect 7006 48220 7012 48232
rect 7064 48220 7070 48272
rect 7190 48260 7196 48272
rect 7151 48232 7196 48260
rect 7190 48220 7196 48232
rect 7248 48220 7254 48272
rect 9398 48220 9404 48272
rect 9456 48260 9462 48272
rect 9582 48260 9588 48272
rect 9456 48232 9588 48260
rect 9456 48220 9462 48232
rect 9582 48220 9588 48232
rect 9640 48220 9646 48272
rect 9769 48263 9827 48269
rect 9769 48229 9781 48263
rect 9815 48260 9827 48263
rect 11072 48260 11100 48300
rect 11238 48288 11244 48300
rect 11296 48288 11302 48340
rect 12710 48328 12716 48340
rect 12671 48300 12716 48328
rect 12710 48288 12716 48300
rect 12768 48288 12774 48340
rect 14090 48288 14096 48340
rect 14148 48328 14154 48340
rect 14148 48300 15148 48328
rect 14148 48288 14154 48300
rect 9815 48232 11100 48260
rect 11701 48263 11759 48269
rect 9815 48229 9827 48232
rect 9769 48223 9827 48229
rect 5166 48152 5172 48204
rect 5224 48192 5230 48204
rect 5810 48192 5816 48204
rect 5224 48164 5816 48192
rect 5224 48152 5230 48164
rect 5810 48152 5816 48164
rect 5868 48152 5874 48204
rect 7374 48192 7380 48204
rect 7335 48164 7380 48192
rect 7374 48152 7380 48164
rect 7432 48152 7438 48204
rect 8021 48195 8079 48201
rect 8021 48161 8033 48195
rect 8067 48192 8079 48195
rect 8386 48192 8392 48204
rect 8067 48164 8392 48192
rect 8067 48161 8079 48164
rect 8021 48155 8079 48161
rect 8386 48152 8392 48164
rect 8444 48152 8450 48204
rect 9122 48152 9128 48204
rect 9180 48192 9186 48204
rect 9217 48195 9275 48201
rect 9217 48192 9229 48195
rect 9180 48164 9229 48192
rect 9180 48152 9186 48164
rect 9217 48161 9229 48164
rect 9263 48161 9275 48195
rect 9217 48155 9275 48161
rect 5350 48084 5356 48136
rect 5408 48124 5414 48136
rect 5905 48127 5963 48133
rect 5905 48124 5917 48127
rect 5408 48096 5917 48124
rect 5408 48084 5414 48096
rect 5905 48093 5917 48096
rect 5951 48124 5963 48127
rect 6086 48124 6092 48136
rect 5951 48096 6092 48124
rect 5951 48093 5963 48096
rect 5905 48087 5963 48093
rect 6086 48084 6092 48096
rect 6144 48084 6150 48136
rect 6914 48084 6920 48136
rect 6972 48124 6978 48136
rect 7009 48127 7067 48133
rect 7009 48124 7021 48127
rect 6972 48096 7021 48124
rect 6972 48084 6978 48096
rect 7009 48093 7021 48096
rect 7055 48093 7067 48127
rect 7009 48087 7067 48093
rect 7190 48084 7196 48136
rect 7248 48124 7254 48136
rect 8113 48127 8171 48133
rect 8113 48124 8125 48127
rect 7248 48096 8125 48124
rect 7248 48084 7254 48096
rect 8113 48093 8125 48096
rect 8159 48124 8171 48127
rect 8202 48124 8208 48136
rect 8159 48096 8208 48124
rect 8159 48093 8171 48096
rect 8113 48087 8171 48093
rect 8202 48084 8208 48096
rect 8260 48084 8266 48136
rect 7466 48056 7472 48068
rect 7427 48028 7472 48056
rect 7466 48016 7472 48028
rect 7524 48016 7530 48068
rect 10060 48056 10088 48232
rect 11701 48229 11713 48263
rect 11747 48260 11759 48263
rect 11790 48260 11796 48272
rect 11747 48232 11796 48260
rect 11747 48229 11759 48232
rect 11701 48223 11759 48229
rect 11790 48220 11796 48232
rect 11848 48220 11854 48272
rect 12069 48263 12127 48269
rect 12069 48229 12081 48263
rect 12115 48260 12127 48263
rect 12618 48260 12624 48272
rect 12115 48232 12624 48260
rect 12115 48229 12127 48232
rect 12069 48223 12127 48229
rect 12618 48220 12624 48232
rect 12676 48220 12682 48272
rect 15120 48260 15148 48300
rect 17310 48288 17316 48340
rect 17368 48328 17374 48340
rect 17405 48331 17463 48337
rect 17405 48328 17417 48331
rect 17368 48300 17417 48328
rect 17368 48288 17374 48300
rect 17405 48297 17417 48300
rect 17451 48297 17463 48331
rect 17405 48291 17463 48297
rect 15841 48263 15899 48269
rect 15841 48260 15853 48263
rect 15120 48232 15853 48260
rect 15841 48229 15853 48232
rect 15887 48260 15899 48263
rect 16298 48260 16304 48272
rect 15887 48232 16304 48260
rect 15887 48229 15899 48232
rect 15841 48223 15899 48229
rect 16298 48220 16304 48232
rect 16356 48220 16362 48272
rect 16393 48263 16451 48269
rect 16393 48229 16405 48263
rect 16439 48260 16451 48263
rect 16482 48260 16488 48272
rect 16439 48232 16488 48260
rect 16439 48229 16451 48232
rect 16393 48223 16451 48229
rect 16482 48220 16488 48232
rect 16540 48220 16546 48272
rect 16761 48263 16819 48269
rect 16761 48229 16773 48263
rect 16807 48260 16819 48263
rect 17129 48263 17187 48269
rect 17129 48260 17141 48263
rect 16807 48232 17141 48260
rect 16807 48229 16819 48232
rect 16761 48223 16819 48229
rect 17129 48229 17141 48232
rect 17175 48260 17187 48263
rect 17586 48260 17592 48272
rect 17175 48232 17592 48260
rect 17175 48229 17187 48232
rect 17129 48223 17187 48229
rect 17328 48204 17356 48232
rect 17586 48220 17592 48232
rect 17644 48220 17650 48272
rect 10410 48192 10416 48204
rect 10371 48164 10416 48192
rect 10410 48152 10416 48164
rect 10468 48152 10474 48204
rect 10502 48152 10508 48204
rect 10560 48192 10566 48204
rect 10686 48201 10692 48204
rect 10638 48195 10692 48201
rect 10560 48164 10605 48192
rect 10560 48152 10566 48164
rect 10638 48161 10650 48195
rect 10684 48161 10692 48195
rect 10638 48155 10692 48161
rect 10686 48152 10692 48155
rect 10744 48152 10750 48204
rect 15930 48192 15936 48204
rect 15891 48164 15936 48192
rect 15930 48152 15936 48164
rect 15988 48152 15994 48204
rect 17310 48152 17316 48204
rect 17368 48152 17374 48204
rect 10134 48084 10140 48136
rect 10192 48124 10198 48136
rect 11054 48124 11060 48136
rect 10192 48096 11060 48124
rect 10192 48084 10198 48096
rect 11054 48084 11060 48096
rect 11112 48084 11118 48136
rect 12894 48084 12900 48136
rect 12952 48124 12958 48136
rect 12989 48127 13047 48133
rect 12989 48124 13001 48127
rect 12952 48096 13001 48124
rect 12952 48084 12958 48096
rect 12989 48093 13001 48096
rect 13035 48093 13047 48127
rect 13262 48124 13268 48136
rect 13223 48096 13268 48124
rect 12989 48087 13047 48093
rect 13262 48084 13268 48096
rect 13320 48084 13326 48136
rect 15470 48084 15476 48136
rect 15528 48124 15534 48136
rect 15746 48124 15752 48136
rect 15528 48096 15752 48124
rect 15528 48084 15534 48096
rect 15746 48084 15752 48096
rect 15804 48084 15810 48136
rect 10594 48056 10600 48068
rect 10060 48028 10600 48056
rect 10594 48016 10600 48028
rect 10652 48016 10658 48068
rect 1578 47988 1584 48000
rect 1539 47960 1584 47988
rect 1578 47948 1584 47960
rect 1636 47948 1642 48000
rect 4890 47988 4896 48000
rect 4803 47960 4896 47988
rect 4890 47948 4896 47960
rect 4948 47988 4954 48000
rect 5350 47988 5356 48000
rect 4948 47960 5356 47988
rect 4948 47948 4954 47960
rect 5350 47948 5356 47960
rect 5408 47948 5414 48000
rect 6914 47948 6920 48000
rect 6972 47988 6978 48000
rect 7193 47991 7251 47997
rect 7193 47988 7205 47991
rect 6972 47960 7205 47988
rect 6972 47948 6978 47960
rect 7193 47957 7205 47960
rect 7239 47957 7251 47991
rect 7193 47951 7251 47957
rect 7558 47948 7564 48000
rect 7616 47988 7622 48000
rect 8018 47988 8024 48000
rect 7616 47960 8024 47988
rect 7616 47948 7622 47960
rect 8018 47948 8024 47960
rect 8076 47948 8082 48000
rect 8294 47948 8300 48000
rect 8352 47988 8358 48000
rect 8665 47991 8723 47997
rect 8665 47988 8677 47991
rect 8352 47960 8677 47988
rect 8352 47948 8358 47960
rect 8665 47957 8677 47960
rect 8711 47957 8723 47991
rect 8665 47951 8723 47957
rect 8754 47948 8760 48000
rect 8812 47988 8818 48000
rect 9401 47991 9459 47997
rect 9401 47988 9413 47991
rect 8812 47960 9413 47988
rect 8812 47948 8818 47960
rect 9401 47957 9413 47960
rect 9447 47957 9459 47991
rect 9401 47951 9459 47957
rect 10042 47948 10048 48000
rect 10100 47988 10106 48000
rect 10137 47991 10195 47997
rect 10137 47988 10149 47991
rect 10100 47960 10149 47988
rect 10100 47948 10106 47960
rect 10137 47957 10149 47960
rect 10183 47957 10195 47991
rect 10778 47988 10784 48000
rect 10739 47960 10784 47988
rect 10137 47951 10195 47957
rect 10778 47948 10784 47960
rect 10836 47948 10842 48000
rect 13906 47948 13912 48000
rect 13964 47988 13970 48000
rect 14369 47991 14427 47997
rect 14369 47988 14381 47991
rect 13964 47960 14381 47988
rect 13964 47948 13970 47960
rect 14369 47957 14381 47960
rect 14415 47957 14427 47991
rect 14369 47951 14427 47957
rect 15470 47948 15476 48000
rect 15528 47988 15534 48000
rect 15657 47991 15715 47997
rect 15657 47988 15669 47991
rect 15528 47960 15669 47988
rect 15528 47948 15534 47960
rect 15657 47957 15669 47960
rect 15703 47957 15715 47991
rect 15657 47951 15715 47957
rect 1104 47898 18860 47920
rect 1104 47846 4315 47898
rect 4367 47846 4379 47898
rect 4431 47846 4443 47898
rect 4495 47846 4507 47898
rect 4559 47846 10982 47898
rect 11034 47846 11046 47898
rect 11098 47846 11110 47898
rect 11162 47846 11174 47898
rect 11226 47846 17648 47898
rect 17700 47846 17712 47898
rect 17764 47846 17776 47898
rect 17828 47846 17840 47898
rect 17892 47846 18860 47898
rect 1104 47824 18860 47846
rect 2869 47787 2927 47793
rect 2869 47753 2881 47787
rect 2915 47784 2927 47787
rect 2958 47784 2964 47796
rect 2915 47756 2964 47784
rect 2915 47753 2927 47756
rect 2869 47747 2927 47753
rect 2958 47744 2964 47756
rect 3016 47744 3022 47796
rect 4341 47787 4399 47793
rect 4341 47753 4353 47787
rect 4387 47784 4399 47787
rect 5166 47784 5172 47796
rect 4387 47756 5172 47784
rect 4387 47753 4399 47756
rect 4341 47747 4399 47753
rect 5166 47744 5172 47756
rect 5224 47744 5230 47796
rect 5460 47756 6132 47784
rect 4709 47719 4767 47725
rect 4709 47685 4721 47719
rect 4755 47716 4767 47719
rect 5460 47716 5488 47756
rect 5810 47716 5816 47728
rect 4755 47688 5488 47716
rect 5736 47688 5816 47716
rect 4755 47685 4767 47688
rect 4709 47679 4767 47685
rect 1670 47608 1676 47660
rect 1728 47648 1734 47660
rect 1765 47651 1823 47657
rect 1765 47648 1777 47651
rect 1728 47620 1777 47648
rect 1728 47608 1734 47620
rect 1765 47617 1777 47620
rect 1811 47617 1823 47651
rect 1765 47611 1823 47617
rect 1489 47583 1547 47589
rect 1489 47549 1501 47583
rect 1535 47580 1547 47583
rect 2038 47580 2044 47592
rect 1535 47552 2044 47580
rect 1535 47549 1547 47552
rect 1489 47543 1547 47549
rect 2038 47540 2044 47552
rect 2096 47540 2102 47592
rect 5736 47589 5764 47688
rect 5810 47676 5816 47688
rect 5868 47676 5874 47728
rect 6104 47716 6132 47756
rect 6638 47744 6644 47796
rect 6696 47784 6702 47796
rect 6733 47787 6791 47793
rect 6733 47784 6745 47787
rect 6696 47756 6745 47784
rect 6696 47744 6702 47756
rect 6733 47753 6745 47756
rect 6779 47753 6791 47787
rect 8478 47784 8484 47796
rect 8439 47756 8484 47784
rect 6733 47747 6791 47753
rect 8478 47744 8484 47756
rect 8536 47744 8542 47796
rect 9122 47784 9128 47796
rect 9083 47756 9128 47784
rect 9122 47744 9128 47756
rect 9180 47784 9186 47796
rect 9401 47787 9459 47793
rect 9401 47784 9413 47787
rect 9180 47756 9413 47784
rect 9180 47744 9186 47756
rect 9401 47753 9413 47756
rect 9447 47753 9459 47787
rect 9401 47747 9459 47753
rect 6104 47688 6960 47716
rect 6932 47592 6960 47688
rect 5721 47583 5779 47589
rect 5721 47549 5733 47583
rect 5767 47549 5779 47583
rect 5905 47583 5963 47589
rect 5905 47580 5917 47583
rect 5721 47543 5779 47549
rect 5828 47552 5917 47580
rect 5828 47456 5856 47552
rect 5905 47549 5917 47552
rect 5951 47549 5963 47583
rect 5905 47543 5963 47549
rect 6086 47540 6092 47592
rect 6144 47580 6150 47592
rect 6273 47583 6331 47589
rect 6273 47580 6285 47583
rect 6144 47552 6285 47580
rect 6144 47540 6150 47552
rect 6273 47549 6285 47552
rect 6319 47549 6331 47583
rect 6914 47580 6920 47592
rect 6875 47552 6920 47580
rect 6273 47543 6331 47549
rect 6914 47540 6920 47552
rect 6972 47540 6978 47592
rect 8294 47580 8300 47592
rect 8255 47552 8300 47580
rect 8294 47540 8300 47552
rect 8352 47540 8358 47592
rect 9416 47580 9444 47747
rect 10410 47744 10416 47796
rect 10468 47784 10474 47796
rect 11057 47787 11115 47793
rect 11057 47784 11069 47787
rect 10468 47756 11069 47784
rect 10468 47744 10474 47756
rect 11057 47753 11069 47756
rect 11103 47753 11115 47787
rect 11057 47747 11115 47753
rect 13173 47787 13231 47793
rect 13173 47753 13185 47787
rect 13219 47784 13231 47787
rect 13262 47784 13268 47796
rect 13219 47756 13268 47784
rect 13219 47753 13231 47756
rect 13173 47747 13231 47753
rect 13262 47744 13268 47756
rect 13320 47744 13326 47796
rect 16298 47744 16304 47796
rect 16356 47784 16362 47796
rect 16669 47787 16727 47793
rect 16669 47784 16681 47787
rect 16356 47756 16681 47784
rect 16356 47744 16362 47756
rect 16669 47753 16681 47756
rect 16715 47753 16727 47787
rect 16669 47747 16727 47753
rect 15105 47651 15163 47657
rect 15105 47617 15117 47651
rect 15151 47648 15163 47651
rect 15151 47620 15884 47648
rect 15151 47617 15163 47620
rect 15105 47611 15163 47617
rect 15856 47592 15884 47620
rect 16390 47608 16396 47660
rect 16448 47648 16454 47660
rect 17954 47648 17960 47660
rect 16448 47620 17960 47648
rect 16448 47608 16454 47620
rect 17954 47608 17960 47620
rect 18012 47608 18018 47660
rect 9677 47583 9735 47589
rect 9677 47580 9689 47583
rect 9416 47552 9689 47580
rect 9677 47549 9689 47552
rect 9723 47549 9735 47583
rect 9677 47543 9735 47549
rect 10229 47583 10287 47589
rect 10229 47549 10241 47583
rect 10275 47580 10287 47583
rect 10594 47580 10600 47592
rect 10275 47552 10600 47580
rect 10275 47549 10287 47552
rect 10229 47543 10287 47549
rect 9122 47472 9128 47524
rect 9180 47512 9186 47524
rect 10244 47512 10272 47543
rect 10594 47540 10600 47552
rect 10652 47540 10658 47592
rect 11790 47580 11796 47592
rect 11751 47552 11796 47580
rect 11790 47540 11796 47552
rect 11848 47540 11854 47592
rect 11882 47540 11888 47592
rect 11940 47580 11946 47592
rect 11977 47583 12035 47589
rect 11977 47580 11989 47583
rect 11940 47552 11989 47580
rect 11940 47540 11946 47552
rect 11977 47549 11989 47552
rect 12023 47549 12035 47583
rect 11977 47543 12035 47549
rect 12250 47540 12256 47592
rect 12308 47580 12314 47592
rect 12345 47583 12403 47589
rect 12345 47580 12357 47583
rect 12308 47552 12357 47580
rect 12308 47540 12314 47552
rect 12345 47549 12357 47552
rect 12391 47549 12403 47583
rect 15657 47583 15715 47589
rect 15657 47580 15669 47583
rect 12345 47543 12403 47549
rect 15488 47552 15669 47580
rect 11514 47512 11520 47524
rect 9180 47484 10272 47512
rect 11427 47484 11520 47512
rect 9180 47472 9186 47484
rect 11514 47472 11520 47484
rect 11572 47512 11578 47524
rect 11900 47512 11928 47540
rect 12710 47512 12716 47524
rect 11572 47484 11928 47512
rect 12671 47484 12716 47512
rect 11572 47472 11578 47484
rect 12710 47472 12716 47484
rect 12768 47472 12774 47524
rect 15488 47456 15516 47552
rect 15657 47549 15669 47552
rect 15703 47549 15715 47583
rect 15838 47580 15844 47592
rect 15799 47552 15844 47580
rect 15657 47543 15715 47549
rect 15838 47540 15844 47552
rect 15896 47540 15902 47592
rect 15933 47583 15991 47589
rect 15933 47549 15945 47583
rect 15979 47549 15991 47583
rect 15933 47543 15991 47549
rect 15562 47472 15568 47524
rect 15620 47512 15626 47524
rect 15948 47512 15976 47543
rect 15620 47484 15976 47512
rect 16393 47515 16451 47521
rect 15620 47472 15626 47484
rect 16393 47481 16405 47515
rect 16439 47512 16451 47515
rect 16482 47512 16488 47524
rect 16439 47484 16488 47512
rect 16439 47481 16451 47484
rect 16393 47475 16451 47481
rect 16482 47472 16488 47484
rect 16540 47472 16546 47524
rect 4706 47404 4712 47456
rect 4764 47444 4770 47456
rect 4890 47444 4896 47456
rect 4764 47416 4896 47444
rect 4764 47404 4770 47416
rect 4890 47404 4896 47416
rect 4948 47404 4954 47456
rect 5077 47447 5135 47453
rect 5077 47413 5089 47447
rect 5123 47444 5135 47447
rect 5166 47444 5172 47456
rect 5123 47416 5172 47444
rect 5123 47413 5135 47416
rect 5077 47407 5135 47413
rect 5166 47404 5172 47416
rect 5224 47404 5230 47456
rect 5445 47447 5503 47453
rect 5445 47413 5457 47447
rect 5491 47444 5503 47447
rect 5810 47444 5816 47456
rect 5491 47416 5816 47444
rect 5491 47413 5503 47416
rect 5445 47407 5503 47413
rect 5810 47404 5816 47416
rect 5868 47404 5874 47456
rect 7190 47404 7196 47456
rect 7248 47444 7254 47456
rect 7285 47447 7343 47453
rect 7285 47444 7297 47447
rect 7248 47416 7297 47444
rect 7248 47404 7254 47416
rect 7285 47413 7297 47416
rect 7331 47413 7343 47447
rect 7285 47407 7343 47413
rect 7374 47404 7380 47456
rect 7432 47444 7438 47456
rect 7745 47447 7803 47453
rect 7745 47444 7757 47447
rect 7432 47416 7757 47444
rect 7432 47404 7438 47416
rect 7745 47413 7757 47416
rect 7791 47444 7803 47447
rect 8202 47444 8208 47456
rect 7791 47416 8208 47444
rect 7791 47413 7803 47416
rect 7745 47407 7803 47413
rect 8202 47404 8208 47416
rect 8260 47404 8266 47456
rect 9674 47404 9680 47456
rect 9732 47444 9738 47456
rect 9769 47447 9827 47453
rect 9769 47444 9781 47447
rect 9732 47416 9781 47444
rect 9732 47404 9738 47416
rect 9769 47413 9781 47416
rect 9815 47413 9827 47447
rect 9769 47407 9827 47413
rect 10502 47404 10508 47456
rect 10560 47444 10566 47456
rect 10689 47447 10747 47453
rect 10689 47444 10701 47447
rect 10560 47416 10701 47444
rect 10560 47404 10566 47416
rect 10689 47413 10701 47416
rect 10735 47413 10747 47447
rect 10689 47407 10747 47413
rect 12894 47404 12900 47456
rect 12952 47444 12958 47456
rect 13449 47447 13507 47453
rect 13449 47444 13461 47447
rect 12952 47416 13461 47444
rect 12952 47404 12958 47416
rect 13449 47413 13461 47416
rect 13495 47444 13507 47447
rect 13817 47447 13875 47453
rect 13817 47444 13829 47447
rect 13495 47416 13829 47444
rect 13495 47413 13507 47416
rect 13449 47407 13507 47413
rect 13817 47413 13829 47416
rect 13863 47413 13875 47447
rect 15470 47444 15476 47456
rect 15431 47416 15476 47444
rect 13817 47407 13875 47413
rect 15470 47404 15476 47416
rect 15528 47404 15534 47456
rect 15838 47404 15844 47456
rect 15896 47444 15902 47456
rect 16114 47444 16120 47456
rect 15896 47416 16120 47444
rect 15896 47404 15902 47416
rect 16114 47404 16120 47416
rect 16172 47404 16178 47456
rect 1104 47354 18860 47376
rect 1104 47302 7648 47354
rect 7700 47302 7712 47354
rect 7764 47302 7776 47354
rect 7828 47302 7840 47354
rect 7892 47302 14315 47354
rect 14367 47302 14379 47354
rect 14431 47302 14443 47354
rect 14495 47302 14507 47354
rect 14559 47302 18860 47354
rect 1104 47280 18860 47302
rect 6273 47243 6331 47249
rect 6273 47209 6285 47243
rect 6319 47240 6331 47243
rect 6638 47240 6644 47252
rect 6319 47212 6644 47240
rect 6319 47209 6331 47212
rect 6273 47203 6331 47209
rect 6638 47200 6644 47212
rect 6696 47200 6702 47252
rect 7377 47243 7435 47249
rect 7377 47209 7389 47243
rect 7423 47240 7435 47243
rect 8386 47240 8392 47252
rect 7423 47212 8392 47240
rect 7423 47209 7435 47212
rect 7377 47203 7435 47209
rect 4709 47175 4767 47181
rect 4709 47141 4721 47175
rect 4755 47172 4767 47175
rect 4755 47144 5672 47172
rect 4755 47141 4767 47144
rect 4709 47135 4767 47141
rect 5644 47116 5672 47144
rect 3510 47104 3516 47116
rect 3471 47076 3516 47104
rect 3510 47064 3516 47076
rect 3568 47064 3574 47116
rect 3602 47064 3608 47116
rect 3660 47104 3666 47116
rect 3697 47107 3755 47113
rect 3697 47104 3709 47107
rect 3660 47076 3709 47104
rect 3660 47064 3666 47076
rect 3697 47073 3709 47076
rect 3743 47073 3755 47107
rect 5169 47107 5227 47113
rect 5169 47104 5181 47107
rect 3697 47067 3755 47073
rect 3804 47076 5181 47104
rect 1670 47036 1676 47048
rect 1583 47008 1676 47036
rect 1670 46996 1676 47008
rect 1728 47036 1734 47048
rect 2406 47036 2412 47048
rect 1728 47008 2412 47036
rect 1728 46996 1734 47008
rect 2406 46996 2412 47008
rect 2464 46996 2470 47048
rect 3234 46996 3240 47048
rect 3292 47036 3298 47048
rect 3804 47036 3832 47076
rect 5169 47073 5181 47076
rect 5215 47073 5227 47107
rect 5626 47104 5632 47116
rect 5587 47076 5632 47104
rect 5169 47067 5227 47073
rect 5626 47064 5632 47076
rect 5684 47064 5690 47116
rect 3970 47036 3976 47048
rect 3292 47008 3832 47036
rect 3931 47008 3976 47036
rect 3292 46996 3298 47008
rect 3970 46996 3976 47008
rect 4028 46996 4034 47048
rect 4062 46996 4068 47048
rect 4120 47036 4126 47048
rect 4985 47039 5043 47045
rect 4985 47036 4997 47039
rect 4120 47008 4997 47036
rect 4120 46996 4126 47008
rect 4985 47005 4997 47008
rect 5031 47036 5043 47039
rect 7392 47036 7420 47203
rect 8386 47200 8392 47212
rect 8444 47240 8450 47252
rect 12802 47240 12808 47252
rect 8444 47212 10364 47240
rect 12763 47212 12808 47240
rect 8444 47200 8450 47212
rect 9030 47172 9036 47184
rect 8588 47144 9036 47172
rect 8588 47116 8616 47144
rect 9030 47132 9036 47144
rect 9088 47132 9094 47184
rect 10336 47181 10364 47212
rect 12802 47200 12808 47212
rect 12860 47200 12866 47252
rect 14090 47200 14096 47252
rect 14148 47240 14154 47252
rect 14369 47243 14427 47249
rect 14369 47240 14381 47243
rect 14148 47212 14381 47240
rect 14148 47200 14154 47212
rect 14369 47209 14381 47212
rect 14415 47209 14427 47243
rect 14369 47203 14427 47209
rect 15930 47200 15936 47252
rect 15988 47240 15994 47252
rect 16393 47243 16451 47249
rect 16393 47240 16405 47243
rect 15988 47212 16405 47240
rect 15988 47200 15994 47212
rect 16393 47209 16405 47212
rect 16439 47209 16451 47243
rect 16393 47203 16451 47209
rect 10321 47175 10379 47181
rect 10321 47141 10333 47175
rect 10367 47141 10379 47175
rect 10321 47135 10379 47141
rect 15562 47132 15568 47184
rect 15620 47172 15626 47184
rect 16025 47175 16083 47181
rect 16025 47172 16037 47175
rect 15620 47144 16037 47172
rect 15620 47132 15626 47144
rect 16025 47141 16037 47144
rect 16071 47141 16083 47175
rect 16025 47135 16083 47141
rect 8021 47107 8079 47113
rect 8021 47104 8033 47107
rect 5031 47008 7420 47036
rect 7668 47076 8033 47104
rect 5031 47005 5043 47008
rect 4985 46999 5043 47005
rect 2038 46968 2044 46980
rect 1951 46940 2044 46968
rect 2038 46928 2044 46940
rect 2096 46968 2102 46980
rect 2498 46968 2504 46980
rect 2096 46940 2504 46968
rect 2096 46928 2102 46940
rect 2498 46928 2504 46940
rect 2556 46928 2562 46980
rect 5534 46928 5540 46980
rect 5592 46968 5598 46980
rect 5629 46971 5687 46977
rect 5629 46968 5641 46971
rect 5592 46940 5641 46968
rect 5592 46928 5598 46940
rect 5629 46937 5641 46940
rect 5675 46937 5687 46971
rect 5629 46931 5687 46937
rect 6638 46928 6644 46980
rect 6696 46968 6702 46980
rect 7668 46968 7696 47076
rect 8021 47073 8033 47076
rect 8067 47104 8079 47107
rect 8570 47104 8576 47116
rect 8067 47076 8432 47104
rect 8531 47076 8576 47104
rect 8067 47073 8079 47076
rect 8021 47067 8079 47073
rect 8294 47036 8300 47048
rect 8255 47008 8300 47036
rect 8294 46996 8300 47008
rect 8352 46996 8358 47048
rect 8404 47036 8432 47076
rect 8570 47064 8576 47076
rect 8628 47064 8634 47116
rect 8754 47104 8760 47116
rect 8715 47076 8760 47104
rect 8754 47064 8760 47076
rect 8812 47064 8818 47116
rect 9214 47064 9220 47116
rect 9272 47104 9278 47116
rect 9309 47107 9367 47113
rect 9309 47104 9321 47107
rect 9272 47076 9321 47104
rect 9272 47064 9278 47076
rect 9309 47073 9321 47076
rect 9355 47073 9367 47107
rect 9309 47067 9367 47073
rect 10594 47064 10600 47116
rect 10652 47104 10658 47116
rect 10962 47104 10968 47116
rect 10652 47076 10968 47104
rect 10652 47064 10658 47076
rect 10962 47064 10968 47076
rect 11020 47064 11026 47116
rect 16850 47064 16856 47116
rect 16908 47104 16914 47116
rect 16945 47107 17003 47113
rect 16945 47104 16957 47107
rect 16908 47076 16957 47104
rect 16908 47064 16914 47076
rect 16945 47073 16957 47076
rect 16991 47104 17003 47107
rect 17126 47104 17132 47116
rect 16991 47076 17132 47104
rect 16991 47073 17003 47076
rect 16945 47067 17003 47073
rect 17126 47064 17132 47076
rect 17184 47064 17190 47116
rect 9769 47039 9827 47045
rect 9769 47036 9781 47039
rect 8404 47008 9781 47036
rect 9769 47005 9781 47008
rect 9815 47036 9827 47039
rect 9858 47036 9864 47048
rect 9815 47008 9864 47036
rect 9815 47005 9827 47008
rect 9769 46999 9827 47005
rect 9858 46996 9864 47008
rect 9916 46996 9922 47048
rect 12161 47039 12219 47045
rect 12161 47005 12173 47039
rect 12207 47036 12219 47039
rect 12894 47036 12900 47048
rect 12207 47008 12900 47036
rect 12207 47005 12219 47008
rect 12161 46999 12219 47005
rect 12894 46996 12900 47008
rect 12952 47036 12958 47048
rect 12989 47039 13047 47045
rect 12989 47036 13001 47039
rect 12952 47008 13001 47036
rect 12952 46996 12958 47008
rect 12989 47005 13001 47008
rect 13035 47005 13047 47039
rect 13262 47036 13268 47048
rect 13223 47008 13268 47036
rect 12989 46999 13047 47005
rect 13262 46996 13268 47008
rect 13320 46996 13326 47048
rect 7742 46968 7748 46980
rect 6696 46940 7748 46968
rect 6696 46928 6702 46940
rect 7742 46928 7748 46940
rect 7800 46928 7806 46980
rect 8386 46928 8392 46980
rect 8444 46928 8450 46980
rect 10229 46971 10287 46977
rect 10229 46937 10241 46971
rect 10275 46968 10287 46971
rect 10686 46968 10692 46980
rect 10275 46940 10692 46968
rect 10275 46937 10287 46940
rect 10229 46931 10287 46937
rect 10686 46928 10692 46940
rect 10744 46928 10750 46980
rect 11514 46928 11520 46980
rect 11572 46968 11578 46980
rect 11609 46971 11667 46977
rect 11609 46968 11621 46971
rect 11572 46940 11621 46968
rect 11572 46928 11578 46940
rect 11609 46937 11621 46940
rect 11655 46968 11667 46971
rect 12250 46968 12256 46980
rect 11655 46940 12256 46968
rect 11655 46937 11667 46940
rect 11609 46931 11667 46937
rect 12250 46928 12256 46940
rect 12308 46928 12314 46980
rect 14734 46928 14740 46980
rect 14792 46968 14798 46980
rect 15470 46968 15476 46980
rect 14792 46940 15476 46968
rect 14792 46928 14798 46940
rect 15470 46928 15476 46940
rect 15528 46968 15534 46980
rect 15657 46971 15715 46977
rect 15657 46968 15669 46971
rect 15528 46940 15669 46968
rect 15528 46928 15534 46940
rect 15657 46937 15669 46940
rect 15703 46937 15715 46971
rect 15657 46931 15715 46937
rect 16850 46928 16856 46980
rect 16908 46968 16914 46980
rect 17129 46971 17187 46977
rect 17129 46968 17141 46971
rect 16908 46940 17141 46968
rect 16908 46928 16914 46940
rect 17129 46937 17141 46940
rect 17175 46937 17187 46971
rect 17129 46931 17187 46937
rect 8294 46860 8300 46912
rect 8352 46900 8358 46912
rect 8404 46900 8432 46928
rect 8352 46872 8432 46900
rect 8352 46860 8358 46872
rect 9858 46860 9864 46912
rect 9916 46900 9922 46912
rect 10134 46900 10140 46912
rect 9916 46872 10140 46900
rect 9916 46860 9922 46872
rect 10134 46860 10140 46872
rect 10192 46860 10198 46912
rect 1104 46810 18860 46832
rect 1104 46758 4315 46810
rect 4367 46758 4379 46810
rect 4431 46758 4443 46810
rect 4495 46758 4507 46810
rect 4559 46758 10982 46810
rect 11034 46758 11046 46810
rect 11098 46758 11110 46810
rect 11162 46758 11174 46810
rect 11226 46758 17648 46810
rect 17700 46758 17712 46810
rect 17764 46758 17776 46810
rect 17828 46758 17840 46810
rect 17892 46758 18860 46810
rect 1104 46736 18860 46758
rect 3513 46699 3571 46705
rect 3513 46665 3525 46699
rect 3559 46696 3571 46699
rect 3602 46696 3608 46708
rect 3559 46668 3608 46696
rect 3559 46665 3571 46668
rect 3513 46659 3571 46665
rect 3602 46656 3608 46668
rect 3660 46656 3666 46708
rect 4062 46656 4068 46708
rect 4120 46696 4126 46708
rect 4249 46699 4307 46705
rect 4249 46696 4261 46699
rect 4120 46668 4261 46696
rect 4120 46656 4126 46668
rect 4249 46665 4261 46668
rect 4295 46665 4307 46699
rect 5626 46696 5632 46708
rect 5587 46668 5632 46696
rect 4249 46659 4307 46665
rect 5626 46656 5632 46668
rect 5684 46656 5690 46708
rect 7742 46696 7748 46708
rect 7703 46668 7748 46696
rect 7742 46656 7748 46668
rect 7800 46656 7806 46708
rect 8481 46699 8539 46705
rect 8481 46665 8493 46699
rect 8527 46696 8539 46699
rect 9214 46696 9220 46708
rect 8527 46668 9220 46696
rect 8527 46665 8539 46668
rect 8481 46659 8539 46665
rect 9214 46656 9220 46668
rect 9272 46696 9278 46708
rect 9674 46696 9680 46708
rect 9272 46668 9680 46696
rect 9272 46656 9278 46668
rect 9674 46656 9680 46668
rect 9732 46656 9738 46708
rect 9766 46656 9772 46708
rect 9824 46696 9830 46708
rect 9861 46699 9919 46705
rect 9861 46696 9873 46699
rect 9824 46668 9873 46696
rect 9824 46656 9830 46668
rect 9861 46665 9873 46668
rect 9907 46696 9919 46699
rect 10134 46696 10140 46708
rect 9907 46668 10140 46696
rect 9907 46665 9919 46668
rect 9861 46659 9919 46665
rect 10134 46656 10140 46668
rect 10192 46656 10198 46708
rect 10594 46696 10600 46708
rect 10555 46668 10600 46696
rect 10594 46656 10600 46668
rect 10652 46656 10658 46708
rect 11422 46696 11428 46708
rect 10980 46668 11428 46696
rect 10980 46640 11008 46668
rect 11422 46656 11428 46668
rect 11480 46696 11486 46708
rect 11609 46699 11667 46705
rect 11609 46696 11621 46699
rect 11480 46668 11621 46696
rect 11480 46656 11486 46668
rect 11609 46665 11621 46668
rect 11655 46665 11667 46699
rect 11609 46659 11667 46665
rect 12621 46699 12679 46705
rect 12621 46665 12633 46699
rect 12667 46696 12679 46699
rect 13170 46696 13176 46708
rect 12667 46668 13176 46696
rect 12667 46665 12679 46668
rect 12621 46659 12679 46665
rect 13170 46656 13176 46668
rect 13228 46656 13234 46708
rect 17221 46699 17279 46705
rect 17221 46665 17233 46699
rect 17267 46696 17279 46699
rect 17310 46696 17316 46708
rect 17267 46668 17316 46696
rect 17267 46665 17279 46668
rect 17221 46659 17279 46665
rect 17310 46656 17316 46668
rect 17368 46656 17374 46708
rect 3234 46588 3240 46640
rect 3292 46628 3298 46640
rect 4617 46631 4675 46637
rect 4617 46628 4629 46631
rect 3292 46600 4629 46628
rect 3292 46588 3298 46600
rect 4617 46597 4629 46600
rect 4663 46628 4675 46631
rect 5534 46628 5540 46640
rect 4663 46600 5540 46628
rect 4663 46597 4675 46600
rect 4617 46591 4675 46597
rect 5534 46588 5540 46600
rect 5592 46588 5598 46640
rect 10962 46588 10968 46640
rect 11020 46588 11026 46640
rect 1489 46563 1547 46569
rect 1489 46529 1501 46563
rect 1535 46560 1547 46563
rect 1670 46560 1676 46572
rect 1535 46532 1676 46560
rect 1535 46529 1547 46532
rect 1489 46523 1547 46529
rect 1670 46520 1676 46532
rect 1728 46520 1734 46572
rect 3145 46563 3203 46569
rect 3145 46529 3157 46563
rect 3191 46560 3203 46563
rect 4522 46560 4528 46572
rect 3191 46532 4528 46560
rect 3191 46529 3203 46532
rect 3145 46523 3203 46529
rect 4522 46520 4528 46532
rect 4580 46520 4586 46572
rect 4706 46520 4712 46572
rect 4764 46520 4770 46572
rect 5077 46563 5135 46569
rect 5077 46529 5089 46563
rect 5123 46560 5135 46563
rect 5166 46560 5172 46572
rect 5123 46532 5172 46560
rect 5123 46529 5135 46532
rect 5077 46523 5135 46529
rect 5166 46520 5172 46532
rect 5224 46560 5230 46572
rect 12713 46563 12771 46569
rect 5224 46532 6132 46560
rect 5224 46520 5230 46532
rect 1765 46495 1823 46501
rect 1765 46492 1777 46495
rect 1504 46464 1777 46492
rect 1504 46436 1532 46464
rect 1765 46461 1777 46464
rect 1811 46461 1823 46495
rect 4724 46492 4752 46520
rect 6104 46504 6132 46532
rect 12713 46529 12725 46563
rect 12759 46560 12771 46563
rect 12894 46560 12900 46572
rect 12759 46532 12900 46560
rect 12759 46529 12771 46532
rect 12713 46523 12771 46529
rect 12894 46520 12900 46532
rect 12952 46560 12958 46572
rect 13170 46560 13176 46572
rect 12952 46532 13176 46560
rect 12952 46520 12958 46532
rect 13170 46520 13176 46532
rect 13228 46520 13234 46572
rect 14093 46563 14151 46569
rect 14093 46529 14105 46563
rect 14139 46529 14151 46563
rect 14093 46523 14151 46529
rect 5626 46492 5632 46504
rect 1765 46455 1823 46461
rect 4632 46464 4752 46492
rect 5587 46464 5632 46492
rect 1486 46384 1492 46436
rect 1544 46384 1550 46436
rect 3510 46316 3516 46368
rect 3568 46356 3574 46368
rect 3881 46359 3939 46365
rect 3881 46356 3893 46359
rect 3568 46328 3893 46356
rect 3568 46316 3574 46328
rect 3881 46325 3893 46328
rect 3927 46356 3939 46359
rect 4062 46356 4068 46368
rect 3927 46328 4068 46356
rect 3927 46325 3939 46328
rect 3881 46319 3939 46325
rect 4062 46316 4068 46328
rect 4120 46316 4126 46368
rect 4632 46356 4660 46464
rect 5626 46452 5632 46464
rect 5684 46452 5690 46504
rect 5905 46495 5963 46501
rect 5905 46492 5917 46495
rect 5828 46464 5917 46492
rect 4706 46384 4712 46436
rect 4764 46424 4770 46436
rect 5258 46424 5264 46436
rect 4764 46396 5264 46424
rect 4764 46384 4770 46396
rect 5258 46384 5264 46396
rect 5316 46384 5322 46436
rect 5828 46368 5856 46464
rect 5905 46461 5917 46464
rect 5951 46461 5963 46495
rect 5905 46455 5963 46461
rect 6086 46452 6092 46504
rect 6144 46492 6150 46504
rect 6273 46495 6331 46501
rect 6273 46492 6285 46495
rect 6144 46464 6285 46492
rect 6144 46452 6150 46464
rect 6273 46461 6285 46464
rect 6319 46461 6331 46495
rect 6914 46492 6920 46504
rect 6875 46464 6920 46492
rect 6273 46455 6331 46461
rect 6914 46452 6920 46464
rect 6972 46452 6978 46504
rect 9677 46495 9735 46501
rect 9677 46461 9689 46495
rect 9723 46492 9735 46495
rect 9950 46492 9956 46504
rect 9723 46464 9956 46492
rect 9723 46461 9735 46464
rect 9677 46455 9735 46461
rect 9950 46452 9956 46464
rect 10008 46492 10014 46504
rect 10137 46495 10195 46501
rect 10137 46492 10149 46495
rect 10008 46464 10149 46492
rect 10008 46452 10014 46464
rect 10137 46461 10149 46464
rect 10183 46461 10195 46495
rect 11422 46492 11428 46504
rect 11383 46464 11428 46492
rect 10137 46455 10195 46461
rect 11422 46452 11428 46464
rect 11480 46492 11486 46504
rect 11885 46495 11943 46501
rect 11885 46492 11897 46495
rect 11480 46464 11897 46492
rect 11480 46452 11486 46464
rect 11885 46461 11897 46464
rect 11931 46461 11943 46495
rect 11885 46455 11943 46461
rect 12802 46452 12808 46504
rect 12860 46492 12866 46504
rect 12989 46495 13047 46501
rect 12989 46492 13001 46495
rect 12860 46464 13001 46492
rect 12860 46452 12866 46464
rect 12989 46461 13001 46464
rect 13035 46461 13047 46495
rect 12989 46455 13047 46461
rect 13262 46452 13268 46504
rect 13320 46492 13326 46504
rect 14108 46492 14136 46523
rect 13320 46464 14136 46492
rect 16025 46495 16083 46501
rect 13320 46452 13326 46464
rect 16025 46461 16037 46495
rect 16071 46461 16083 46495
rect 17034 46492 17040 46504
rect 16995 46464 17040 46492
rect 16025 46455 16083 46461
rect 8113 46427 8171 46433
rect 8113 46393 8125 46427
rect 8159 46424 8171 46427
rect 8754 46424 8760 46436
rect 8159 46396 8760 46424
rect 8159 46393 8171 46396
rect 8113 46387 8171 46393
rect 8754 46384 8760 46396
rect 8812 46384 8818 46436
rect 16040 46424 16068 46455
rect 17034 46452 17040 46464
rect 17092 46492 17098 46504
rect 17497 46495 17555 46501
rect 17497 46492 17509 46495
rect 17092 46464 17509 46492
rect 17092 46452 17098 46464
rect 17497 46461 17509 46464
rect 17543 46461 17555 46495
rect 17497 46455 17555 46461
rect 16577 46427 16635 46433
rect 16577 46424 16589 46427
rect 16040 46396 16589 46424
rect 16577 46393 16589 46396
rect 16623 46424 16635 46427
rect 18138 46424 18144 46436
rect 16623 46396 18144 46424
rect 16623 46393 16635 46396
rect 16577 46387 16635 46393
rect 18138 46384 18144 46396
rect 18196 46384 18202 46436
rect 5166 46356 5172 46368
rect 4632 46328 5172 46356
rect 5166 46316 5172 46328
rect 5224 46316 5230 46368
rect 5445 46359 5503 46365
rect 5445 46325 5457 46359
rect 5491 46356 5503 46359
rect 5810 46356 5816 46368
rect 5491 46328 5816 46356
rect 5491 46325 5503 46328
rect 5445 46319 5503 46325
rect 5810 46316 5816 46328
rect 5868 46316 5874 46368
rect 8570 46316 8576 46368
rect 8628 46356 8634 46368
rect 8849 46359 8907 46365
rect 8849 46356 8861 46359
rect 8628 46328 8861 46356
rect 8628 46316 8634 46328
rect 8849 46325 8861 46328
rect 8895 46356 8907 46359
rect 9398 46356 9404 46368
rect 8895 46328 9404 46356
rect 8895 46325 8907 46328
rect 8849 46319 8907 46325
rect 9398 46316 9404 46328
rect 9456 46316 9462 46368
rect 12250 46316 12256 46368
rect 12308 46356 12314 46368
rect 13906 46356 13912 46368
rect 12308 46328 13912 46356
rect 12308 46316 12314 46328
rect 13906 46316 13912 46328
rect 13964 46316 13970 46368
rect 16206 46356 16212 46368
rect 16167 46328 16212 46356
rect 16206 46316 16212 46328
rect 16264 46316 16270 46368
rect 16945 46359 17003 46365
rect 16945 46325 16957 46359
rect 16991 46356 17003 46359
rect 17126 46356 17132 46368
rect 16991 46328 17132 46356
rect 16991 46325 17003 46328
rect 16945 46319 17003 46325
rect 17126 46316 17132 46328
rect 17184 46316 17190 46368
rect 1104 46266 18860 46288
rect 1104 46214 7648 46266
rect 7700 46214 7712 46266
rect 7764 46214 7776 46266
rect 7828 46214 7840 46266
rect 7892 46214 14315 46266
rect 14367 46214 14379 46266
rect 14431 46214 14443 46266
rect 14495 46214 14507 46266
rect 14559 46214 18860 46266
rect 1104 46192 18860 46214
rect 1670 46112 1676 46164
rect 1728 46152 1734 46164
rect 2041 46155 2099 46161
rect 2041 46152 2053 46155
rect 1728 46124 2053 46152
rect 1728 46112 1734 46124
rect 2041 46121 2053 46124
rect 2087 46152 2099 46155
rect 2314 46152 2320 46164
rect 2087 46124 2320 46152
rect 2087 46121 2099 46124
rect 2041 46115 2099 46121
rect 2314 46112 2320 46124
rect 2372 46112 2378 46164
rect 4062 46112 4068 46164
rect 4120 46152 4126 46164
rect 5169 46155 5227 46161
rect 5169 46152 5181 46155
rect 4120 46124 5181 46152
rect 4120 46112 4126 46124
rect 5169 46121 5181 46124
rect 5215 46121 5227 46155
rect 5169 46115 5227 46121
rect 5626 46112 5632 46164
rect 5684 46152 5690 46164
rect 6089 46155 6147 46161
rect 6089 46152 6101 46155
rect 5684 46124 6101 46152
rect 5684 46112 5690 46124
rect 6089 46121 6101 46124
rect 6135 46121 6147 46155
rect 6089 46115 6147 46121
rect 6730 46112 6736 46164
rect 6788 46112 6794 46164
rect 7006 46152 7012 46164
rect 6967 46124 7012 46152
rect 7006 46112 7012 46124
rect 7064 46112 7070 46164
rect 9122 46112 9128 46164
rect 9180 46152 9186 46164
rect 9306 46152 9312 46164
rect 9180 46124 9312 46152
rect 9180 46112 9186 46124
rect 9306 46112 9312 46124
rect 9364 46112 9370 46164
rect 9950 46112 9956 46164
rect 10008 46152 10014 46164
rect 10597 46155 10655 46161
rect 10597 46152 10609 46155
rect 10008 46124 10609 46152
rect 10008 46112 10014 46124
rect 10597 46121 10609 46124
rect 10643 46152 10655 46155
rect 10778 46152 10784 46164
rect 10643 46124 10784 46152
rect 10643 46121 10655 46124
rect 10597 46115 10655 46121
rect 10778 46112 10784 46124
rect 10836 46112 10842 46164
rect 11606 46112 11612 46164
rect 11664 46152 11670 46164
rect 12250 46152 12256 46164
rect 11664 46124 12256 46152
rect 11664 46112 11670 46124
rect 12250 46112 12256 46124
rect 12308 46112 12314 46164
rect 12621 46155 12679 46161
rect 12621 46121 12633 46155
rect 12667 46152 12679 46155
rect 12710 46152 12716 46164
rect 12667 46124 12716 46152
rect 12667 46121 12679 46124
rect 12621 46115 12679 46121
rect 12710 46112 12716 46124
rect 12768 46112 12774 46164
rect 13078 46112 13084 46164
rect 13136 46152 13142 46164
rect 13630 46152 13636 46164
rect 13136 46124 13636 46152
rect 13136 46112 13142 46124
rect 13630 46112 13636 46124
rect 13688 46112 13694 46164
rect 16574 46112 16580 46164
rect 16632 46152 16638 46164
rect 17126 46152 17132 46164
rect 16632 46124 17132 46152
rect 16632 46112 16638 46124
rect 17126 46112 17132 46124
rect 17184 46112 17190 46164
rect 17310 46112 17316 46164
rect 17368 46152 17374 46164
rect 17405 46155 17463 46161
rect 17405 46152 17417 46155
rect 17368 46124 17417 46152
rect 17368 46112 17374 46124
rect 17405 46121 17417 46124
rect 17451 46121 17463 46155
rect 17405 46115 17463 46121
rect 2498 45976 2504 46028
rect 2556 46016 2562 46028
rect 2556 45988 3556 46016
rect 2556 45976 2562 45988
rect 3528 45960 3556 45988
rect 3510 45908 3516 45960
rect 3568 45948 3574 45960
rect 3789 45951 3847 45957
rect 3789 45948 3801 45951
rect 3568 45920 3801 45948
rect 3568 45908 3574 45920
rect 3789 45917 3801 45920
rect 3835 45917 3847 45951
rect 4062 45948 4068 45960
rect 4023 45920 4068 45948
rect 3789 45911 3847 45917
rect 4062 45908 4068 45920
rect 4120 45908 4126 45960
rect 6546 45908 6552 45960
rect 6604 45948 6610 45960
rect 6748 45948 6776 46112
rect 8478 46084 8484 46096
rect 8036 46056 8484 46084
rect 8036 46028 8064 46056
rect 8478 46044 8484 46056
rect 8536 46044 8542 46096
rect 10229 46087 10287 46093
rect 10229 46053 10241 46087
rect 10275 46084 10287 46087
rect 10686 46084 10692 46096
rect 10275 46056 10692 46084
rect 10275 46053 10287 46056
rect 10229 46047 10287 46053
rect 10686 46044 10692 46056
rect 10744 46044 10750 46096
rect 10870 46044 10876 46096
rect 10928 46084 10934 46096
rect 11057 46087 11115 46093
rect 11057 46084 11069 46087
rect 10928 46056 11069 46084
rect 10928 46044 10934 46056
rect 11057 46053 11069 46056
rect 11103 46053 11115 46087
rect 11057 46047 11115 46053
rect 12805 46087 12863 46093
rect 12805 46053 12817 46087
rect 12851 46084 12863 46087
rect 12851 46056 13032 46084
rect 12851 46053 12863 46056
rect 12805 46047 12863 46053
rect 6825 46019 6883 46025
rect 6825 45985 6837 46019
rect 6871 46016 6883 46019
rect 7282 46016 7288 46028
rect 6871 45988 7288 46016
rect 6871 45985 6883 45988
rect 6825 45979 6883 45985
rect 7282 45976 7288 45988
rect 7340 45976 7346 46028
rect 8018 46016 8024 46028
rect 7931 45988 8024 46016
rect 8018 45976 8024 45988
rect 8076 45976 8082 46028
rect 8110 45976 8116 46028
rect 8168 46016 8174 46028
rect 8665 46019 8723 46025
rect 8665 46016 8677 46019
rect 8168 45988 8677 46016
rect 8168 45976 8174 45988
rect 8665 45985 8677 45988
rect 8711 45985 8723 46019
rect 8665 45979 8723 45985
rect 9674 45976 9680 46028
rect 9732 46016 9738 46028
rect 10410 46016 10416 46028
rect 9732 45988 10416 46016
rect 9732 45976 9738 45988
rect 10410 45976 10416 45988
rect 10468 46016 10474 46028
rect 10505 46019 10563 46025
rect 10505 46016 10517 46019
rect 10468 45988 10517 46016
rect 10468 45976 10474 45988
rect 10505 45985 10517 45988
rect 10551 45985 10563 46019
rect 10505 45979 10563 45985
rect 12710 45976 12716 46028
rect 12768 46016 12774 46028
rect 12768 45988 12813 46016
rect 12768 45976 12774 45988
rect 13004 45960 13032 46056
rect 13170 46044 13176 46096
rect 13228 46084 13234 46096
rect 13228 46056 13308 46084
rect 13228 46044 13234 46056
rect 6604 45920 6776 45948
rect 6604 45908 6610 45920
rect 8386 45908 8392 45960
rect 8444 45948 8450 45960
rect 8573 45951 8631 45957
rect 8573 45948 8585 45951
rect 8444 45920 8585 45948
rect 8444 45908 8450 45920
rect 8573 45917 8585 45920
rect 8619 45917 8631 45951
rect 8573 45911 8631 45917
rect 8846 45908 8852 45960
rect 8904 45948 8910 45960
rect 9030 45948 9036 45960
rect 8904 45920 9036 45948
rect 8904 45908 8910 45920
rect 9030 45908 9036 45920
rect 9088 45908 9094 45960
rect 9858 45908 9864 45960
rect 9916 45948 9922 45960
rect 10321 45951 10379 45957
rect 10321 45948 10333 45951
rect 9916 45920 10333 45948
rect 9916 45908 9922 45920
rect 10321 45917 10333 45920
rect 10367 45917 10379 45951
rect 10321 45911 10379 45917
rect 12437 45951 12495 45957
rect 12437 45917 12449 45951
rect 12483 45948 12495 45951
rect 12894 45948 12900 45960
rect 12483 45920 12900 45948
rect 12483 45917 12495 45920
rect 12437 45911 12495 45917
rect 12894 45908 12900 45920
rect 12952 45908 12958 45960
rect 12986 45908 12992 45960
rect 13044 45908 13050 45960
rect 13170 45948 13176 45960
rect 13131 45920 13176 45948
rect 13170 45908 13176 45920
rect 13228 45908 13234 45960
rect 11885 45883 11943 45889
rect 11885 45849 11897 45883
rect 11931 45880 11943 45883
rect 12342 45880 12348 45892
rect 11931 45852 12348 45880
rect 11931 45849 11943 45852
rect 11885 45843 11943 45849
rect 12342 45840 12348 45852
rect 12400 45840 12406 45892
rect 1486 45772 1492 45824
rect 1544 45812 1550 45824
rect 1581 45815 1639 45821
rect 1581 45812 1593 45815
rect 1544 45784 1593 45812
rect 1544 45772 1550 45784
rect 1581 45781 1593 45784
rect 1627 45781 1639 45815
rect 1581 45775 1639 45781
rect 5626 45772 5632 45824
rect 5684 45812 5690 45824
rect 5813 45815 5871 45821
rect 5813 45812 5825 45815
rect 5684 45784 5825 45812
rect 5684 45772 5690 45784
rect 5813 45781 5825 45784
rect 5859 45812 5871 45815
rect 6638 45812 6644 45824
rect 5859 45784 6644 45812
rect 5859 45781 5871 45784
rect 5813 45775 5871 45781
rect 6638 45772 6644 45784
rect 6696 45812 6702 45824
rect 6914 45812 6920 45824
rect 6696 45784 6920 45812
rect 6696 45772 6702 45784
rect 6914 45772 6920 45784
rect 6972 45772 6978 45824
rect 7282 45812 7288 45824
rect 7243 45784 7288 45812
rect 7282 45772 7288 45784
rect 7340 45772 7346 45824
rect 8941 45815 8999 45821
rect 8941 45781 8953 45815
rect 8987 45812 8999 45815
rect 9674 45812 9680 45824
rect 8987 45784 9680 45812
rect 8987 45781 8999 45784
rect 8941 45775 8999 45781
rect 9674 45772 9680 45784
rect 9732 45772 9738 45824
rect 9858 45812 9864 45824
rect 9819 45784 9864 45812
rect 9858 45772 9864 45784
rect 9916 45812 9922 45824
rect 10226 45812 10232 45824
rect 9916 45784 10232 45812
rect 9916 45772 9922 45784
rect 10226 45772 10232 45784
rect 10284 45772 10290 45824
rect 11422 45812 11428 45824
rect 11383 45784 11428 45812
rect 11422 45772 11428 45784
rect 11480 45772 11486 45824
rect 12434 45772 12440 45824
rect 12492 45812 12498 45824
rect 13280 45812 13308 46056
rect 14550 46044 14556 46096
rect 14608 46084 14614 46096
rect 15102 46084 15108 46096
rect 14608 46056 15108 46084
rect 14608 46044 14614 46056
rect 15102 46044 15108 46056
rect 15160 46044 15166 46096
rect 15657 46087 15715 46093
rect 15657 46053 15669 46087
rect 15703 46084 15715 46087
rect 17328 46084 17356 46112
rect 15703 46056 17356 46084
rect 15703 46053 15715 46056
rect 15657 46047 15715 46053
rect 14642 46016 14648 46028
rect 14603 45988 14648 46016
rect 14642 45976 14648 45988
rect 14700 45976 14706 46028
rect 16574 45976 16580 46028
rect 16632 46016 16638 46028
rect 16669 46019 16727 46025
rect 16669 46016 16681 46019
rect 16632 45988 16681 46016
rect 16632 45976 16638 45988
rect 16669 45985 16681 45988
rect 16715 45985 16727 46019
rect 16669 45979 16727 45985
rect 16945 46019 17003 46025
rect 16945 45985 16957 46019
rect 16991 45985 17003 46019
rect 16945 45979 17003 45985
rect 17129 46019 17187 46025
rect 17129 45985 17141 46019
rect 17175 46016 17187 46019
rect 17328 46016 17356 46056
rect 17175 45988 17356 46016
rect 17175 45985 17187 45988
rect 17129 45979 17187 45985
rect 15289 45951 15347 45957
rect 15289 45917 15301 45951
rect 15335 45948 15347 45951
rect 15470 45948 15476 45960
rect 15335 45920 15476 45948
rect 15335 45917 15347 45920
rect 15289 45911 15347 45917
rect 15470 45908 15476 45920
rect 15528 45908 15534 45960
rect 15930 45908 15936 45960
rect 15988 45948 15994 45960
rect 16117 45951 16175 45957
rect 16117 45948 16129 45951
rect 15988 45920 16129 45948
rect 15988 45908 15994 45920
rect 16117 45917 16129 45920
rect 16163 45917 16175 45951
rect 16117 45911 16175 45917
rect 16960 45948 16988 45979
rect 18414 45948 18420 45960
rect 16960 45920 18420 45948
rect 16025 45883 16083 45889
rect 16025 45849 16037 45883
rect 16071 45880 16083 45883
rect 16960 45880 16988 45920
rect 18414 45908 18420 45920
rect 18472 45908 18478 45960
rect 16071 45852 16988 45880
rect 16071 45849 16083 45852
rect 16025 45843 16083 45849
rect 13449 45815 13507 45821
rect 13449 45812 13461 45815
rect 12492 45784 13461 45812
rect 12492 45772 12498 45784
rect 13449 45781 13461 45784
rect 13495 45812 13507 45815
rect 13817 45815 13875 45821
rect 13817 45812 13829 45815
rect 13495 45784 13829 45812
rect 13495 45781 13507 45784
rect 13449 45775 13507 45781
rect 13817 45781 13829 45784
rect 13863 45781 13875 45815
rect 13817 45775 13875 45781
rect 1104 45722 18860 45744
rect 1104 45670 4315 45722
rect 4367 45670 4379 45722
rect 4431 45670 4443 45722
rect 4495 45670 4507 45722
rect 4559 45670 10982 45722
rect 11034 45670 11046 45722
rect 11098 45670 11110 45722
rect 11162 45670 11174 45722
rect 11226 45670 17648 45722
rect 17700 45670 17712 45722
rect 17764 45670 17776 45722
rect 17828 45670 17840 45722
rect 17892 45670 18860 45722
rect 1104 45648 18860 45670
rect 3510 45568 3516 45620
rect 3568 45608 3574 45620
rect 5626 45608 5632 45620
rect 3568 45580 4200 45608
rect 3568 45568 3574 45580
rect 4172 45540 4200 45580
rect 5552 45580 5632 45608
rect 4249 45543 4307 45549
rect 4249 45540 4261 45543
rect 4172 45512 4261 45540
rect 4249 45509 4261 45512
rect 4295 45509 4307 45543
rect 4249 45503 4307 45509
rect 5077 45543 5135 45549
rect 5077 45509 5089 45543
rect 5123 45540 5135 45543
rect 5552 45540 5580 45580
rect 5626 45568 5632 45580
rect 5684 45568 5690 45620
rect 6178 45568 6184 45620
rect 6236 45608 6242 45620
rect 6733 45611 6791 45617
rect 6733 45608 6745 45611
rect 6236 45580 6745 45608
rect 6236 45568 6242 45580
rect 6733 45577 6745 45580
rect 6779 45577 6791 45611
rect 6733 45571 6791 45577
rect 7377 45611 7435 45617
rect 7377 45577 7389 45611
rect 7423 45608 7435 45611
rect 8018 45608 8024 45620
rect 7423 45580 8024 45608
rect 7423 45577 7435 45580
rect 7377 45571 7435 45577
rect 8018 45568 8024 45580
rect 8076 45568 8082 45620
rect 8386 45608 8392 45620
rect 8312 45580 8392 45608
rect 5123 45512 5580 45540
rect 7745 45543 7803 45549
rect 5123 45509 5135 45512
rect 5077 45503 5135 45509
rect 7745 45509 7757 45543
rect 7791 45540 7803 45543
rect 8312 45540 8340 45580
rect 8386 45568 8392 45580
rect 8444 45568 8450 45620
rect 10778 45568 10784 45620
rect 10836 45608 10842 45620
rect 10836 45580 11100 45608
rect 10836 45568 10842 45580
rect 7791 45512 8340 45540
rect 7791 45509 7803 45512
rect 7745 45503 7803 45509
rect 9858 45500 9864 45552
rect 9916 45540 9922 45552
rect 9916 45512 10364 45540
rect 9916 45500 9922 45512
rect 1489 45475 1547 45481
rect 1489 45441 1501 45475
rect 1535 45472 1547 45475
rect 2222 45472 2228 45484
rect 1535 45444 2228 45472
rect 1535 45441 1547 45444
rect 1489 45435 1547 45441
rect 2222 45432 2228 45444
rect 2280 45432 2286 45484
rect 3145 45475 3203 45481
rect 3145 45441 3157 45475
rect 3191 45472 3203 45475
rect 3418 45472 3424 45484
rect 3191 45444 3424 45472
rect 3191 45441 3203 45444
rect 3145 45435 3203 45441
rect 3418 45432 3424 45444
rect 3476 45432 3482 45484
rect 9398 45432 9404 45484
rect 9456 45472 9462 45484
rect 9493 45475 9551 45481
rect 9493 45472 9505 45475
rect 9456 45444 9505 45472
rect 9456 45432 9462 45444
rect 9493 45441 9505 45444
rect 9539 45472 9551 45475
rect 9539 45444 10180 45472
rect 9539 45441 9551 45444
rect 9493 45435 9551 45441
rect 1578 45364 1584 45416
rect 1636 45404 1642 45416
rect 1765 45407 1823 45413
rect 1765 45404 1777 45407
rect 1636 45376 1777 45404
rect 1636 45364 1642 45376
rect 1765 45373 1777 45376
rect 1811 45373 1823 45407
rect 1765 45367 1823 45373
rect 4709 45407 4767 45413
rect 4709 45373 4721 45407
rect 4755 45404 4767 45407
rect 5626 45404 5632 45416
rect 4755 45376 5632 45404
rect 4755 45373 4767 45376
rect 4709 45367 4767 45373
rect 5626 45364 5632 45376
rect 5684 45364 5690 45416
rect 5905 45407 5963 45413
rect 5905 45404 5917 45407
rect 5828 45376 5917 45404
rect 5828 45280 5856 45376
rect 5905 45373 5917 45376
rect 5951 45373 5963 45407
rect 5905 45367 5963 45373
rect 6086 45364 6092 45416
rect 6144 45404 6150 45416
rect 6273 45407 6331 45413
rect 6273 45404 6285 45407
rect 6144 45376 6285 45404
rect 6144 45364 6150 45376
rect 6273 45373 6285 45376
rect 6319 45373 6331 45407
rect 6273 45367 6331 45373
rect 6638 45364 6644 45416
rect 6696 45404 6702 45416
rect 6917 45407 6975 45413
rect 6917 45404 6929 45407
rect 6696 45376 6929 45404
rect 6696 45364 6702 45376
rect 6917 45373 6929 45376
rect 6963 45373 6975 45407
rect 6917 45367 6975 45373
rect 8481 45407 8539 45413
rect 8481 45373 8493 45407
rect 8527 45404 8539 45407
rect 8849 45407 8907 45413
rect 8849 45404 8861 45407
rect 8527 45376 8861 45404
rect 8527 45373 8539 45376
rect 8481 45367 8539 45373
rect 8849 45373 8861 45376
rect 8895 45404 8907 45407
rect 9766 45404 9772 45416
rect 8895 45376 9772 45404
rect 8895 45373 8907 45376
rect 8849 45367 8907 45373
rect 9766 45364 9772 45376
rect 9824 45364 9830 45416
rect 10152 45413 10180 45444
rect 10137 45407 10195 45413
rect 10137 45373 10149 45407
rect 10183 45404 10195 45407
rect 10226 45404 10232 45416
rect 10183 45376 10232 45404
rect 10183 45373 10195 45376
rect 10137 45367 10195 45373
rect 10226 45364 10232 45376
rect 10284 45364 10290 45416
rect 10336 45413 10364 45512
rect 10410 45500 10416 45552
rect 10468 45540 10474 45552
rect 10686 45540 10692 45552
rect 10468 45512 10692 45540
rect 10468 45500 10474 45512
rect 10686 45500 10692 45512
rect 10744 45540 10750 45552
rect 10873 45543 10931 45549
rect 10873 45540 10885 45543
rect 10744 45512 10885 45540
rect 10744 45500 10750 45512
rect 10873 45509 10885 45512
rect 10919 45509 10931 45543
rect 11072 45540 11100 45580
rect 12250 45568 12256 45620
rect 12308 45608 12314 45620
rect 12526 45608 12532 45620
rect 12308 45580 12532 45608
rect 12308 45568 12314 45580
rect 12526 45568 12532 45580
rect 12584 45568 12590 45620
rect 12894 45608 12900 45620
rect 12855 45580 12900 45608
rect 12894 45568 12900 45580
rect 12952 45568 12958 45620
rect 15286 45568 15292 45620
rect 15344 45608 15350 45620
rect 15654 45608 15660 45620
rect 15344 45580 15660 45608
rect 15344 45568 15350 45580
rect 15654 45568 15660 45580
rect 15712 45568 15718 45620
rect 11241 45543 11299 45549
rect 11241 45540 11253 45543
rect 11072 45512 11253 45540
rect 10873 45503 10931 45509
rect 11241 45509 11253 45512
rect 11287 45509 11299 45543
rect 11241 45503 11299 45509
rect 12802 45500 12808 45552
rect 12860 45540 12866 45552
rect 13265 45543 13323 45549
rect 13265 45540 13277 45543
rect 12860 45512 13277 45540
rect 12860 45500 12866 45512
rect 13265 45509 13277 45512
rect 13311 45509 13323 45543
rect 13265 45503 13323 45509
rect 15746 45500 15752 45552
rect 15804 45540 15810 45552
rect 16301 45543 16359 45549
rect 16301 45540 16313 45543
rect 15804 45512 16313 45540
rect 15804 45500 15810 45512
rect 16301 45509 16313 45512
rect 16347 45509 16359 45543
rect 16301 45503 16359 45509
rect 13538 45472 13544 45484
rect 12820 45444 13544 45472
rect 12820 45416 12848 45444
rect 13538 45432 13544 45444
rect 13596 45432 13602 45484
rect 15105 45475 15163 45481
rect 15105 45441 15117 45475
rect 15151 45472 15163 45475
rect 16574 45472 16580 45484
rect 15151 45444 16580 45472
rect 15151 45441 15163 45444
rect 15105 45435 15163 45441
rect 16574 45432 16580 45444
rect 16632 45472 16638 45484
rect 17313 45475 17371 45481
rect 17313 45472 17325 45475
rect 16632 45444 17325 45472
rect 16632 45432 16638 45444
rect 17313 45441 17325 45444
rect 17359 45472 17371 45475
rect 18049 45475 18107 45481
rect 18049 45472 18061 45475
rect 17359 45444 18061 45472
rect 17359 45441 17371 45444
rect 17313 45435 17371 45441
rect 18049 45441 18061 45444
rect 18095 45441 18107 45475
rect 18049 45435 18107 45441
rect 10321 45407 10379 45413
rect 10321 45373 10333 45407
rect 10367 45373 10379 45407
rect 10321 45367 10379 45373
rect 10597 45407 10655 45413
rect 10597 45373 10609 45407
rect 10643 45404 10655 45407
rect 11422 45404 11428 45416
rect 10643 45376 11428 45404
rect 10643 45373 10655 45376
rect 10597 45367 10655 45373
rect 11422 45364 11428 45376
rect 11480 45364 11486 45416
rect 11606 45364 11612 45416
rect 11664 45404 11670 45416
rect 11793 45407 11851 45413
rect 11793 45404 11805 45407
rect 11664 45376 11805 45404
rect 11664 45364 11670 45376
rect 11793 45373 11805 45376
rect 11839 45373 11851 45407
rect 11793 45367 11851 45373
rect 11882 45364 11888 45416
rect 11940 45404 11946 45416
rect 12161 45407 12219 45413
rect 12161 45404 12173 45407
rect 11940 45376 12173 45404
rect 11940 45364 11946 45376
rect 12161 45373 12173 45376
rect 12207 45373 12219 45407
rect 12161 45367 12219 45373
rect 12802 45364 12808 45416
rect 12860 45364 12866 45416
rect 14185 45407 14243 45413
rect 14185 45404 14197 45407
rect 14016 45376 14197 45404
rect 12621 45339 12679 45345
rect 12621 45305 12633 45339
rect 12667 45336 12679 45339
rect 12986 45336 12992 45348
rect 12667 45308 12992 45336
rect 12667 45305 12679 45308
rect 12621 45299 12679 45305
rect 12986 45296 12992 45308
rect 13044 45296 13050 45348
rect 14016 45280 14044 45376
rect 14185 45373 14197 45376
rect 14231 45404 14243 45407
rect 14642 45404 14648 45416
rect 14231 45376 14648 45404
rect 14231 45373 14243 45376
rect 14185 45367 14243 45373
rect 14642 45364 14648 45376
rect 14700 45364 14706 45416
rect 15470 45404 15476 45416
rect 15431 45376 15476 45404
rect 15470 45364 15476 45376
rect 15528 45404 15534 45416
rect 15933 45407 15991 45413
rect 15933 45404 15945 45407
rect 15528 45376 15945 45404
rect 15528 45364 15534 45376
rect 15933 45373 15945 45376
rect 15979 45373 15991 45407
rect 17586 45404 17592 45416
rect 17547 45376 17592 45404
rect 15933 45367 15991 45373
rect 17586 45364 17592 45376
rect 17644 45364 17650 45416
rect 17773 45407 17831 45413
rect 17773 45373 17785 45407
rect 17819 45373 17831 45407
rect 17773 45367 17831 45373
rect 15562 45296 15568 45348
rect 15620 45336 15626 45348
rect 16761 45339 16819 45345
rect 15620 45308 15792 45336
rect 15620 45296 15626 45308
rect 2958 45228 2964 45280
rect 3016 45268 3022 45280
rect 3789 45271 3847 45277
rect 3789 45268 3801 45271
rect 3016 45240 3801 45268
rect 3016 45228 3022 45240
rect 3789 45237 3801 45240
rect 3835 45268 3847 45271
rect 4062 45268 4068 45280
rect 3835 45240 4068 45268
rect 3835 45237 3847 45240
rect 3789 45231 3847 45237
rect 4062 45228 4068 45240
rect 4120 45228 4126 45280
rect 5445 45271 5503 45277
rect 5445 45237 5457 45271
rect 5491 45268 5503 45271
rect 5810 45268 5816 45280
rect 5491 45240 5816 45268
rect 5491 45237 5503 45240
rect 5445 45231 5503 45237
rect 5810 45228 5816 45240
rect 5868 45228 5874 45280
rect 8018 45228 8024 45280
rect 8076 45268 8082 45280
rect 8113 45271 8171 45277
rect 8113 45268 8125 45271
rect 8076 45240 8125 45268
rect 8076 45228 8082 45240
rect 8113 45237 8125 45240
rect 8159 45237 8171 45271
rect 8113 45231 8171 45237
rect 12526 45228 12532 45280
rect 12584 45268 12590 45280
rect 13633 45271 13691 45277
rect 13633 45268 13645 45271
rect 12584 45240 13645 45268
rect 12584 45228 12590 45240
rect 13633 45237 13645 45240
rect 13679 45237 13691 45271
rect 13998 45268 14004 45280
rect 13959 45240 14004 45268
rect 13633 45231 13691 45237
rect 13998 45228 14004 45240
rect 14056 45228 14062 45280
rect 14369 45271 14427 45277
rect 14369 45237 14381 45271
rect 14415 45268 14427 45271
rect 14826 45268 14832 45280
rect 14415 45240 14832 45268
rect 14415 45237 14427 45240
rect 14369 45231 14427 45237
rect 14826 45228 14832 45240
rect 14884 45228 14890 45280
rect 15378 45228 15384 45280
rect 15436 45268 15442 45280
rect 15657 45271 15715 45277
rect 15657 45268 15669 45271
rect 15436 45240 15669 45268
rect 15436 45228 15442 45240
rect 15657 45237 15669 45240
rect 15703 45237 15715 45271
rect 15764 45268 15792 45308
rect 16761 45305 16773 45339
rect 16807 45336 16819 45339
rect 16850 45336 16856 45348
rect 16807 45308 16856 45336
rect 16807 45305 16819 45308
rect 16761 45299 16819 45305
rect 16850 45296 16856 45308
rect 16908 45296 16914 45348
rect 17310 45296 17316 45348
rect 17368 45336 17374 45348
rect 17788 45336 17816 45367
rect 17368 45308 17816 45336
rect 17368 45296 17374 45308
rect 18230 45268 18236 45280
rect 15764 45240 18236 45268
rect 15657 45231 15715 45237
rect 18230 45228 18236 45240
rect 18288 45228 18294 45280
rect 1104 45178 18860 45200
rect 1104 45126 7648 45178
rect 7700 45126 7712 45178
rect 7764 45126 7776 45178
rect 7828 45126 7840 45178
rect 7892 45126 14315 45178
rect 14367 45126 14379 45178
rect 14431 45126 14443 45178
rect 14495 45126 14507 45178
rect 14559 45126 18860 45178
rect 1104 45104 18860 45126
rect 2041 45067 2099 45073
rect 2041 45033 2053 45067
rect 2087 45064 2099 45067
rect 2314 45064 2320 45076
rect 2087 45036 2320 45064
rect 2087 45033 2099 45036
rect 2041 45027 2099 45033
rect 2314 45024 2320 45036
rect 2372 45024 2378 45076
rect 4246 45064 4252 45076
rect 4207 45036 4252 45064
rect 4246 45024 4252 45036
rect 4304 45024 4310 45076
rect 8110 45064 8116 45076
rect 8071 45036 8116 45064
rect 8110 45024 8116 45036
rect 8168 45024 8174 45076
rect 9674 45024 9680 45076
rect 9732 45064 9738 45076
rect 9769 45067 9827 45073
rect 9769 45064 9781 45067
rect 9732 45036 9781 45064
rect 9732 45024 9738 45036
rect 9769 45033 9781 45036
rect 9815 45033 9827 45067
rect 9769 45027 9827 45033
rect 9858 45024 9864 45076
rect 9916 45064 9922 45076
rect 10137 45067 10195 45073
rect 10137 45064 10149 45067
rect 9916 45036 10149 45064
rect 9916 45024 9922 45036
rect 10137 45033 10149 45036
rect 10183 45064 10195 45067
rect 11422 45064 11428 45076
rect 10183 45036 11428 45064
rect 10183 45033 10195 45036
rect 10137 45027 10195 45033
rect 11422 45024 11428 45036
rect 11480 45024 11486 45076
rect 12066 45024 12072 45076
rect 12124 45064 12130 45076
rect 12161 45067 12219 45073
rect 12161 45064 12173 45067
rect 12124 45036 12173 45064
rect 12124 45024 12130 45036
rect 12161 45033 12173 45036
rect 12207 45033 12219 45067
rect 12710 45064 12716 45076
rect 12671 45036 12716 45064
rect 12161 45027 12219 45033
rect 12710 45024 12716 45036
rect 12768 45024 12774 45076
rect 12986 45064 12992 45076
rect 12947 45036 12992 45064
rect 12986 45024 12992 45036
rect 13044 45024 13050 45076
rect 15562 45064 15568 45076
rect 15475 45036 15568 45064
rect 15562 45024 15568 45036
rect 15620 45064 15626 45076
rect 16206 45064 16212 45076
rect 15620 45036 16212 45064
rect 15620 45024 15626 45036
rect 16206 45024 16212 45036
rect 16264 45024 16270 45076
rect 17497 45067 17555 45073
rect 17497 45033 17509 45067
rect 17543 45064 17555 45067
rect 17586 45064 17592 45076
rect 17543 45036 17592 45064
rect 17543 45033 17555 45036
rect 17497 45027 17555 45033
rect 17586 45024 17592 45036
rect 17644 45064 17650 45076
rect 18322 45064 18328 45076
rect 17644 45036 18328 45064
rect 17644 45024 17650 45036
rect 18322 45024 18328 45036
rect 18380 45024 18386 45076
rect 1946 44956 1952 45008
rect 2004 44996 2010 45008
rect 2222 44996 2228 45008
rect 2004 44968 2228 44996
rect 2004 44956 2010 44968
rect 2222 44956 2228 44968
rect 2280 44956 2286 45008
rect 6825 44999 6883 45005
rect 6825 44965 6837 44999
rect 6871 44996 6883 44999
rect 7098 44996 7104 45008
rect 6871 44968 7104 44996
rect 6871 44965 6883 44968
rect 6825 44959 6883 44965
rect 7098 44956 7104 44968
rect 7156 44956 7162 45008
rect 8662 44956 8668 45008
rect 8720 44996 8726 45008
rect 11517 44999 11575 45005
rect 8720 44968 9260 44996
rect 8720 44956 8726 44968
rect 1302 44888 1308 44940
rect 1360 44928 1366 44940
rect 2406 44928 2412 44940
rect 1360 44900 2412 44928
rect 1360 44888 1366 44900
rect 2406 44888 2412 44900
rect 2464 44888 2470 44940
rect 3970 44888 3976 44940
rect 4028 44928 4034 44940
rect 4157 44931 4215 44937
rect 4157 44928 4169 44931
rect 4028 44900 4169 44928
rect 4028 44888 4034 44900
rect 4157 44897 4169 44900
rect 4203 44897 4215 44931
rect 4157 44891 4215 44897
rect 4709 44931 4767 44937
rect 4709 44897 4721 44931
rect 4755 44897 4767 44931
rect 4709 44891 4767 44897
rect 4062 44820 4068 44872
rect 4120 44860 4126 44872
rect 4724 44860 4752 44891
rect 6178 44888 6184 44940
rect 6236 44928 6242 44940
rect 6549 44931 6607 44937
rect 6549 44928 6561 44931
rect 6236 44900 6561 44928
rect 6236 44888 6242 44900
rect 6549 44897 6561 44900
rect 6595 44928 6607 44931
rect 7515 44931 7573 44937
rect 7515 44928 7527 44931
rect 6595 44900 7527 44928
rect 6595 44897 6607 44900
rect 6549 44891 6607 44897
rect 7515 44897 7527 44900
rect 7561 44897 7573 44931
rect 7515 44891 7573 44897
rect 7653 44931 7711 44937
rect 7653 44897 7665 44931
rect 7699 44928 7711 44931
rect 8294 44928 8300 44940
rect 7699 44900 8300 44928
rect 7699 44897 7711 44900
rect 7653 44891 7711 44897
rect 4120 44832 4752 44860
rect 5169 44863 5227 44869
rect 4120 44820 4126 44832
rect 5169 44829 5181 44863
rect 5215 44860 5227 44863
rect 5258 44860 5264 44872
rect 5215 44832 5264 44860
rect 5215 44829 5227 44832
rect 5169 44823 5227 44829
rect 5258 44820 5264 44832
rect 5316 44820 5322 44872
rect 6914 44820 6920 44872
rect 6972 44860 6978 44872
rect 7282 44860 7288 44872
rect 6972 44832 7288 44860
rect 6972 44820 6978 44832
rect 7282 44820 7288 44832
rect 7340 44860 7346 44872
rect 7377 44863 7435 44869
rect 7377 44860 7389 44863
rect 7340 44832 7389 44860
rect 7340 44820 7346 44832
rect 7377 44829 7389 44832
rect 7423 44829 7435 44863
rect 7377 44823 7435 44829
rect 5629 44795 5687 44801
rect 5629 44761 5641 44795
rect 5675 44792 5687 44795
rect 6086 44792 6092 44804
rect 5675 44764 6092 44792
rect 5675 44761 5687 44764
rect 5629 44755 5687 44761
rect 6086 44752 6092 44764
rect 6144 44752 6150 44804
rect 7098 44752 7104 44804
rect 7156 44792 7162 44804
rect 7668 44792 7696 44891
rect 8294 44888 8300 44900
rect 8352 44888 8358 44940
rect 9232 44937 9260 44968
rect 11517 44965 11529 44999
rect 11563 44996 11575 44999
rect 12894 44996 12900 45008
rect 11563 44968 12900 44996
rect 11563 44965 11575 44968
rect 11517 44959 11575 44965
rect 12894 44956 12900 44968
rect 12952 44956 12958 45008
rect 14826 44956 14832 45008
rect 14884 44996 14890 45008
rect 15930 44996 15936 45008
rect 14884 44968 15936 44996
rect 14884 44956 14890 44968
rect 15930 44956 15936 44968
rect 15988 44996 15994 45008
rect 16224 44996 16252 45024
rect 15988 44968 16068 44996
rect 16224 44968 16988 44996
rect 15988 44956 15994 44968
rect 9033 44931 9091 44937
rect 9033 44897 9045 44931
rect 9079 44897 9091 44931
rect 9033 44891 9091 44897
rect 9217 44931 9275 44937
rect 9217 44897 9229 44931
rect 9263 44897 9275 44931
rect 9217 44891 9275 44897
rect 9048 44860 9076 44891
rect 9766 44888 9772 44940
rect 9824 44928 9830 44940
rect 10597 44931 10655 44937
rect 10597 44928 10609 44931
rect 9824 44900 10609 44928
rect 9824 44888 9830 44900
rect 10597 44897 10609 44900
rect 10643 44897 10655 44931
rect 10870 44928 10876 44940
rect 10831 44900 10876 44928
rect 10597 44891 10655 44897
rect 9493 44863 9551 44869
rect 9048 44832 9260 44860
rect 9232 44804 9260 44832
rect 9493 44829 9505 44863
rect 9539 44860 9551 44863
rect 9582 44860 9588 44872
rect 9539 44832 9588 44860
rect 9539 44829 9551 44832
rect 9493 44823 9551 44829
rect 9582 44820 9588 44832
rect 9640 44820 9646 44872
rect 10612 44860 10640 44891
rect 10870 44888 10876 44900
rect 10928 44888 10934 44940
rect 11333 44931 11391 44937
rect 11333 44897 11345 44931
rect 11379 44928 11391 44931
rect 11606 44928 11612 44940
rect 11379 44900 11612 44928
rect 11379 44897 11391 44900
rect 11333 44891 11391 44897
rect 11606 44888 11612 44900
rect 11664 44928 11670 44940
rect 12158 44928 12164 44940
rect 11664 44900 12164 44928
rect 11664 44888 11670 44900
rect 12158 44888 12164 44900
rect 12216 44888 12222 44940
rect 13449 44931 13507 44937
rect 13449 44897 13461 44931
rect 13495 44928 13507 44931
rect 13538 44928 13544 44940
rect 13495 44900 13544 44928
rect 13495 44897 13507 44900
rect 13449 44891 13507 44897
rect 13538 44888 13544 44900
rect 13596 44888 13602 44940
rect 15197 44931 15255 44937
rect 15197 44897 15209 44931
rect 15243 44928 15255 44931
rect 15746 44928 15752 44940
rect 15243 44900 15752 44928
rect 15243 44897 15255 44900
rect 15197 44891 15255 44897
rect 15746 44888 15752 44900
rect 15804 44888 15810 44940
rect 16040 44937 16068 44968
rect 16025 44931 16083 44937
rect 16025 44897 16037 44931
rect 16071 44897 16083 44931
rect 16666 44928 16672 44940
rect 16627 44900 16672 44928
rect 16025 44891 16083 44897
rect 16666 44888 16672 44900
rect 16724 44888 16730 44940
rect 16960 44937 16988 44968
rect 16945 44931 17003 44937
rect 16945 44897 16957 44931
rect 16991 44897 17003 44931
rect 16945 44891 17003 44897
rect 12434 44860 12440 44872
rect 10612 44832 12440 44860
rect 12434 44820 12440 44832
rect 12492 44820 12498 44872
rect 12526 44820 12532 44872
rect 12584 44860 12590 44872
rect 12894 44860 12900 44872
rect 12584 44832 12900 44860
rect 12584 44820 12590 44832
rect 12894 44820 12900 44832
rect 12952 44860 12958 44872
rect 13173 44863 13231 44869
rect 13173 44860 13185 44863
rect 12952 44832 13185 44860
rect 12952 44820 12958 44832
rect 13173 44829 13185 44832
rect 13219 44829 13231 44863
rect 13173 44823 13231 44829
rect 7156 44764 7696 44792
rect 7156 44752 7162 44764
rect 9214 44752 9220 44804
rect 9272 44752 9278 44804
rect 10962 44752 10968 44804
rect 11020 44792 11026 44804
rect 11514 44792 11520 44804
rect 11020 44764 11520 44792
rect 11020 44752 11026 44764
rect 11514 44752 11520 44764
rect 11572 44752 11578 44804
rect 1578 44724 1584 44736
rect 1539 44696 1584 44724
rect 1578 44684 1584 44696
rect 1636 44684 1642 44736
rect 5997 44727 6055 44733
rect 5997 44693 6009 44727
rect 6043 44724 6055 44727
rect 6270 44724 6276 44736
rect 6043 44696 6276 44724
rect 6043 44693 6055 44696
rect 5997 44687 6055 44693
rect 6270 44684 6276 44696
rect 6328 44684 6334 44736
rect 11790 44724 11796 44736
rect 11751 44696 11796 44724
rect 11790 44684 11796 44696
rect 11848 44684 11854 44736
rect 14550 44724 14556 44736
rect 14511 44696 14556 44724
rect 14550 44684 14556 44696
rect 14608 44684 14614 44736
rect 15749 44727 15807 44733
rect 15749 44693 15761 44727
rect 15795 44724 15807 44727
rect 15838 44724 15844 44736
rect 15795 44696 15844 44724
rect 15795 44693 15807 44696
rect 15749 44687 15807 44693
rect 15838 44684 15844 44696
rect 15896 44684 15902 44736
rect 1104 44634 18860 44656
rect 1104 44582 4315 44634
rect 4367 44582 4379 44634
rect 4431 44582 4443 44634
rect 4495 44582 4507 44634
rect 4559 44582 10982 44634
rect 11034 44582 11046 44634
rect 11098 44582 11110 44634
rect 11162 44582 11174 44634
rect 11226 44582 17648 44634
rect 17700 44582 17712 44634
rect 17764 44582 17776 44634
rect 17828 44582 17840 44634
rect 17892 44582 18860 44634
rect 1104 44560 18860 44582
rect 1670 44520 1676 44532
rect 1583 44492 1676 44520
rect 1670 44480 1676 44492
rect 1728 44520 1734 44532
rect 2314 44520 2320 44532
rect 1728 44492 2320 44520
rect 1728 44480 1734 44492
rect 2314 44480 2320 44492
rect 2372 44480 2378 44532
rect 3513 44523 3571 44529
rect 3513 44489 3525 44523
rect 3559 44520 3571 44523
rect 3970 44520 3976 44532
rect 3559 44492 3976 44520
rect 3559 44489 3571 44492
rect 3513 44483 3571 44489
rect 3970 44480 3976 44492
rect 4028 44480 4034 44532
rect 7190 44520 7196 44532
rect 7103 44492 7196 44520
rect 7190 44480 7196 44492
rect 7248 44520 7254 44532
rect 8110 44520 8116 44532
rect 7248 44492 8116 44520
rect 7248 44480 7254 44492
rect 8110 44480 8116 44492
rect 8168 44480 8174 44532
rect 9030 44480 9036 44532
rect 9088 44520 9094 44532
rect 9401 44523 9459 44529
rect 9401 44520 9413 44523
rect 9088 44492 9413 44520
rect 9088 44480 9094 44492
rect 9401 44489 9413 44492
rect 9447 44489 9459 44523
rect 9401 44483 9459 44489
rect 11057 44523 11115 44529
rect 11057 44489 11069 44523
rect 11103 44520 11115 44523
rect 11606 44520 11612 44532
rect 11103 44492 11612 44520
rect 11103 44489 11115 44492
rect 11057 44483 11115 44489
rect 3881 44455 3939 44461
rect 3881 44421 3893 44455
rect 3927 44452 3939 44455
rect 4062 44452 4068 44464
rect 3927 44424 4068 44452
rect 3927 44421 3939 44424
rect 3881 44415 3939 44421
rect 4062 44412 4068 44424
rect 4120 44452 4126 44464
rect 4246 44452 4252 44464
rect 4120 44424 4252 44452
rect 4120 44412 4126 44424
rect 4246 44412 4252 44424
rect 4304 44412 4310 44464
rect 5994 44412 6000 44464
rect 6052 44452 6058 44464
rect 6181 44455 6239 44461
rect 6181 44452 6193 44455
rect 6052 44424 6193 44452
rect 6052 44412 6058 44424
rect 6181 44421 6193 44424
rect 6227 44421 6239 44455
rect 7374 44452 7380 44464
rect 7335 44424 7380 44452
rect 6181 44415 6239 44421
rect 7374 44412 7380 44424
rect 7432 44412 7438 44464
rect 8849 44455 8907 44461
rect 8849 44421 8861 44455
rect 8895 44452 8907 44455
rect 9214 44452 9220 44464
rect 8895 44424 9220 44452
rect 8895 44421 8907 44424
rect 8849 44415 8907 44421
rect 9214 44412 9220 44424
rect 9272 44412 9278 44464
rect 4893 44387 4951 44393
rect 4893 44353 4905 44387
rect 4939 44384 4951 44387
rect 5537 44387 5595 44393
rect 5537 44384 5549 44387
rect 4939 44356 5549 44384
rect 4939 44353 4951 44356
rect 4893 44347 4951 44353
rect 5537 44353 5549 44356
rect 5583 44384 5595 44387
rect 8018 44384 8024 44396
rect 5583 44356 8024 44384
rect 5583 44353 5595 44356
rect 5537 44347 5595 44353
rect 3970 44276 3976 44328
rect 4028 44316 4034 44328
rect 4249 44319 4307 44325
rect 4249 44316 4261 44319
rect 4028 44288 4261 44316
rect 4028 44276 4034 44288
rect 4249 44285 4261 44288
rect 4295 44316 4307 44319
rect 5258 44316 5264 44328
rect 4295 44288 5264 44316
rect 4295 44285 4307 44288
rect 4249 44279 4307 44285
rect 5258 44276 5264 44288
rect 5316 44276 5322 44328
rect 5626 44276 5632 44328
rect 5684 44316 5690 44328
rect 5721 44319 5779 44325
rect 5721 44316 5733 44319
rect 5684 44288 5733 44316
rect 5684 44276 5690 44288
rect 5721 44285 5733 44288
rect 5767 44285 5779 44319
rect 6270 44316 6276 44328
rect 6231 44288 6276 44316
rect 5721 44279 5779 44285
rect 6270 44276 6276 44288
rect 6328 44276 6334 44328
rect 7944 44325 7972 44356
rect 8018 44344 8024 44356
rect 8076 44384 8082 44396
rect 8294 44384 8300 44396
rect 8076 44356 8300 44384
rect 8076 44344 8082 44356
rect 8294 44344 8300 44356
rect 8352 44344 8358 44396
rect 7469 44319 7527 44325
rect 7469 44285 7481 44319
rect 7515 44285 7527 44319
rect 7469 44279 7527 44285
rect 7929 44319 7987 44325
rect 7929 44285 7941 44319
rect 7975 44285 7987 44319
rect 8110 44316 8116 44328
rect 8071 44288 8116 44316
rect 7929 44279 7987 44285
rect 5169 44251 5227 44257
rect 5169 44217 5181 44251
rect 5215 44248 5227 44251
rect 5644 44248 5672 44276
rect 5215 44220 5672 44248
rect 5215 44217 5227 44220
rect 5169 44211 5227 44217
rect 5994 44208 6000 44260
rect 6052 44248 6058 44260
rect 6546 44248 6552 44260
rect 6052 44220 6552 44248
rect 6052 44208 6058 44220
rect 6546 44208 6552 44220
rect 6604 44208 6610 44260
rect 6825 44251 6883 44257
rect 6825 44217 6837 44251
rect 6871 44248 6883 44251
rect 7006 44248 7012 44260
rect 6871 44220 7012 44248
rect 6871 44217 6883 44220
rect 6825 44211 6883 44217
rect 7006 44208 7012 44220
rect 7064 44248 7070 44260
rect 7484 44248 7512 44279
rect 8110 44276 8116 44288
rect 8168 44276 8174 44328
rect 9416 44316 9444 44483
rect 11606 44480 11612 44492
rect 11664 44480 11670 44532
rect 13265 44523 13323 44529
rect 13265 44489 13277 44523
rect 13311 44520 13323 44523
rect 13538 44520 13544 44532
rect 13311 44492 13544 44520
rect 13311 44489 13323 44492
rect 13265 44483 13323 44489
rect 13538 44480 13544 44492
rect 13596 44480 13602 44532
rect 14737 44523 14795 44529
rect 14737 44489 14749 44523
rect 14783 44520 14795 44523
rect 14918 44520 14924 44532
rect 14783 44492 14924 44520
rect 14783 44489 14795 44492
rect 14737 44483 14795 44489
rect 11514 44452 11520 44464
rect 11475 44424 11520 44452
rect 11514 44412 11520 44424
rect 11572 44412 11578 44464
rect 12434 44412 12440 44464
rect 12492 44452 12498 44464
rect 14090 44452 14096 44464
rect 12492 44424 14096 44452
rect 12492 44412 12498 44424
rect 14090 44412 14096 44424
rect 14148 44412 14154 44464
rect 9674 44344 9680 44396
rect 9732 44384 9738 44396
rect 9732 44356 10548 44384
rect 9732 44344 9738 44356
rect 10226 44316 10232 44328
rect 9416 44288 10232 44316
rect 10226 44276 10232 44288
rect 10284 44276 10290 44328
rect 10520 44325 10548 44356
rect 10505 44319 10563 44325
rect 10505 44285 10517 44319
rect 10551 44285 10563 44319
rect 10505 44279 10563 44285
rect 10689 44319 10747 44325
rect 10689 44285 10701 44319
rect 10735 44285 10747 44319
rect 10689 44279 10747 44285
rect 8018 44248 8024 44260
rect 7064 44220 8024 44248
rect 7064 44208 7070 44220
rect 8018 44208 8024 44220
rect 8076 44208 8082 44260
rect 9677 44251 9735 44257
rect 9677 44217 9689 44251
rect 9723 44248 9735 44251
rect 9766 44248 9772 44260
rect 9723 44220 9772 44248
rect 9723 44217 9735 44220
rect 9677 44211 9735 44217
rect 9766 44208 9772 44220
rect 9824 44208 9830 44260
rect 9858 44208 9864 44260
rect 9916 44248 9922 44260
rect 10704 44248 10732 44279
rect 10870 44276 10876 44328
rect 10928 44316 10934 44328
rect 11532 44316 11560 44412
rect 12710 44384 12716 44396
rect 12671 44356 12716 44384
rect 12710 44344 12716 44356
rect 12768 44344 12774 44396
rect 11609 44319 11667 44325
rect 11609 44316 11621 44319
rect 10928 44288 11621 44316
rect 10928 44276 10934 44288
rect 11609 44285 11621 44288
rect 11655 44285 11667 44319
rect 11609 44279 11667 44285
rect 12253 44319 12311 44325
rect 12253 44285 12265 44319
rect 12299 44316 12311 44319
rect 12342 44316 12348 44328
rect 12299 44288 12348 44316
rect 12299 44285 12311 44288
rect 12253 44279 12311 44285
rect 12342 44276 12348 44288
rect 12400 44276 12406 44328
rect 12526 44276 12532 44328
rect 12584 44316 12590 44328
rect 12621 44319 12679 44325
rect 12621 44316 12633 44319
rect 12584 44288 12633 44316
rect 12584 44276 12590 44288
rect 12621 44285 12633 44288
rect 12667 44316 12679 44319
rect 13722 44316 13728 44328
rect 12667 44288 13728 44316
rect 12667 44285 12679 44288
rect 12621 44279 12679 44285
rect 13722 44276 13728 44288
rect 13780 44276 13786 44328
rect 13909 44319 13967 44325
rect 13909 44285 13921 44319
rect 13955 44285 13967 44319
rect 13909 44279 13967 44285
rect 14001 44319 14059 44325
rect 14001 44285 14013 44319
rect 14047 44316 14059 44319
rect 14090 44316 14096 44328
rect 14047 44288 14096 44316
rect 14047 44285 14059 44288
rect 14001 44279 14059 44285
rect 9916 44220 10732 44248
rect 9916 44208 9922 44220
rect 12710 44208 12716 44260
rect 12768 44248 12774 44260
rect 13354 44248 13360 44260
rect 12768 44220 13360 44248
rect 12768 44208 12774 44220
rect 13354 44208 13360 44220
rect 13412 44208 13418 44260
rect 13814 44208 13820 44260
rect 13872 44248 13878 44260
rect 13924 44248 13952 44279
rect 14090 44276 14096 44288
rect 14148 44276 14154 44328
rect 14369 44319 14427 44325
rect 14369 44285 14381 44319
rect 14415 44316 14427 44319
rect 14752 44316 14780 44483
rect 14918 44480 14924 44492
rect 14976 44480 14982 44532
rect 16942 44520 16948 44532
rect 15028 44492 16948 44520
rect 14918 44344 14924 44396
rect 14976 44384 14982 44396
rect 15028 44384 15056 44492
rect 16942 44480 16948 44492
rect 17000 44480 17006 44532
rect 15657 44455 15715 44461
rect 15657 44421 15669 44455
rect 15703 44452 15715 44455
rect 16666 44452 16672 44464
rect 15703 44424 16672 44452
rect 15703 44421 15715 44424
rect 15657 44415 15715 44421
rect 16666 44412 16672 44424
rect 16724 44452 16730 44464
rect 16724 44424 16896 44452
rect 16724 44412 16730 44424
rect 14976 44356 15056 44384
rect 16577 44387 16635 44393
rect 14976 44344 14982 44356
rect 16577 44353 16589 44387
rect 16623 44353 16635 44387
rect 16577 44347 16635 44353
rect 14415 44288 14780 44316
rect 14415 44285 14427 44288
rect 14369 44279 14427 44285
rect 15746 44276 15752 44328
rect 15804 44316 15810 44328
rect 16117 44319 16175 44325
rect 16117 44316 16129 44319
rect 15804 44288 16129 44316
rect 15804 44276 15810 44288
rect 16117 44285 16129 44288
rect 16163 44285 16175 44319
rect 16117 44279 16175 44285
rect 16485 44319 16543 44325
rect 16485 44285 16497 44319
rect 16531 44285 16543 44319
rect 16485 44279 16543 44285
rect 15013 44251 15071 44257
rect 15013 44248 15025 44251
rect 13872 44220 15025 44248
rect 13872 44208 13878 44220
rect 15013 44217 15025 44220
rect 15059 44217 15071 44251
rect 15013 44211 15071 44217
rect 15378 44208 15384 44260
rect 15436 44248 15442 44260
rect 15933 44251 15991 44257
rect 15933 44248 15945 44251
rect 15436 44220 15945 44248
rect 15436 44208 15442 44220
rect 15933 44217 15945 44220
rect 15979 44248 15991 44251
rect 16390 44248 16396 44260
rect 15979 44220 16396 44248
rect 15979 44217 15991 44220
rect 15933 44211 15991 44217
rect 16390 44208 16396 44220
rect 16448 44248 16454 44260
rect 16500 44248 16528 44279
rect 16448 44220 16528 44248
rect 16448 44208 16454 44220
rect 16592 44192 16620 44347
rect 16868 44325 16896 44424
rect 16853 44319 16911 44325
rect 16853 44285 16865 44319
rect 16899 44316 16911 44319
rect 17310 44316 17316 44328
rect 16899 44288 17316 44316
rect 16899 44285 16911 44288
rect 16853 44279 16911 44285
rect 17310 44276 17316 44288
rect 17368 44276 17374 44328
rect 17586 44316 17592 44328
rect 17547 44288 17592 44316
rect 17586 44276 17592 44288
rect 17644 44276 17650 44328
rect 17328 44248 17356 44276
rect 17865 44251 17923 44257
rect 17865 44248 17877 44251
rect 17328 44220 17877 44248
rect 17865 44217 17877 44220
rect 17911 44217 17923 44251
rect 17865 44211 17923 44217
rect 14734 44140 14740 44192
rect 14792 44180 14798 44192
rect 15654 44180 15660 44192
rect 14792 44152 15660 44180
rect 14792 44140 14798 44152
rect 15654 44140 15660 44152
rect 15712 44140 15718 44192
rect 16574 44140 16580 44192
rect 16632 44140 16638 44192
rect 1104 44090 18860 44112
rect 1104 44038 7648 44090
rect 7700 44038 7712 44090
rect 7764 44038 7776 44090
rect 7828 44038 7840 44090
rect 7892 44038 14315 44090
rect 14367 44038 14379 44090
rect 14431 44038 14443 44090
rect 14495 44038 14507 44090
rect 14559 44038 18860 44090
rect 1104 44016 18860 44038
rect 6273 43979 6331 43985
rect 6273 43945 6285 43979
rect 6319 43976 6331 43979
rect 7098 43976 7104 43988
rect 6319 43948 7104 43976
rect 6319 43945 6331 43948
rect 6273 43939 6331 43945
rect 7098 43936 7104 43948
rect 7156 43936 7162 43988
rect 8294 43976 8300 43988
rect 8255 43948 8300 43976
rect 8294 43936 8300 43948
rect 8352 43936 8358 43988
rect 10318 43976 10324 43988
rect 8864 43948 10324 43976
rect 3145 43911 3203 43917
rect 3145 43877 3157 43911
rect 3191 43908 3203 43911
rect 3234 43908 3240 43920
rect 3191 43880 3240 43908
rect 3191 43877 3203 43880
rect 3145 43871 3203 43877
rect 3234 43868 3240 43880
rect 3292 43868 3298 43920
rect 4154 43908 4160 43920
rect 4115 43880 4160 43908
rect 4154 43868 4160 43880
rect 4212 43868 4218 43920
rect 4982 43868 4988 43920
rect 5040 43868 5046 43920
rect 3970 43800 3976 43852
rect 4028 43840 4034 43852
rect 4893 43843 4951 43849
rect 4893 43840 4905 43843
rect 4028 43812 4905 43840
rect 4028 43800 4034 43812
rect 4893 43809 4905 43812
rect 4939 43840 4951 43843
rect 5000 43840 5028 43868
rect 6914 43840 6920 43852
rect 4939 43812 5028 43840
rect 6875 43812 6920 43840
rect 4939 43809 4951 43812
rect 4893 43803 4951 43809
rect 6914 43800 6920 43812
rect 6972 43800 6978 43852
rect 7098 43800 7104 43852
rect 7156 43840 7162 43852
rect 7285 43843 7343 43849
rect 7285 43840 7297 43843
rect 7156 43812 7297 43840
rect 7156 43800 7162 43812
rect 7285 43809 7297 43812
rect 7331 43809 7343 43843
rect 7285 43803 7343 43809
rect 7466 43800 7472 43852
rect 7524 43840 7530 43852
rect 7745 43843 7803 43849
rect 7745 43840 7757 43843
rect 7524 43812 7757 43840
rect 7524 43800 7530 43812
rect 7745 43809 7757 43812
rect 7791 43809 7803 43843
rect 7745 43803 7803 43809
rect 8294 43800 8300 43852
rect 8352 43840 8358 43852
rect 8864 43840 8892 43948
rect 10318 43936 10324 43948
rect 10376 43936 10382 43988
rect 11882 43936 11888 43988
rect 11940 43976 11946 43988
rect 12069 43979 12127 43985
rect 12069 43976 12081 43979
rect 11940 43948 12081 43976
rect 11940 43936 11946 43948
rect 12069 43945 12081 43948
rect 12115 43976 12127 43979
rect 12434 43976 12440 43988
rect 12115 43948 12440 43976
rect 12115 43945 12127 43948
rect 12069 43939 12127 43945
rect 12434 43936 12440 43948
rect 12492 43936 12498 43988
rect 12710 43936 12716 43988
rect 12768 43976 12774 43988
rect 12989 43979 13047 43985
rect 12989 43976 13001 43979
rect 12768 43948 13001 43976
rect 12768 43936 12774 43948
rect 12989 43945 13001 43948
rect 13035 43976 13047 43979
rect 13262 43976 13268 43988
rect 13035 43948 13268 43976
rect 13035 43945 13047 43948
rect 12989 43939 13047 43945
rect 13262 43936 13268 43948
rect 13320 43936 13326 43988
rect 15562 43976 15568 43988
rect 15523 43948 15568 43976
rect 15562 43936 15568 43948
rect 15620 43936 15626 43988
rect 9401 43911 9459 43917
rect 9401 43877 9413 43911
rect 9447 43908 9459 43911
rect 9447 43880 10364 43908
rect 9447 43877 9459 43880
rect 9401 43871 9459 43877
rect 10336 43852 10364 43880
rect 14182 43868 14188 43920
rect 14240 43908 14246 43920
rect 14366 43908 14372 43920
rect 14240 43880 14372 43908
rect 14240 43868 14246 43880
rect 14366 43868 14372 43880
rect 14424 43868 14430 43920
rect 15197 43911 15255 43917
rect 15197 43877 15209 43911
rect 15243 43908 15255 43911
rect 15580 43908 15608 43936
rect 17586 43908 17592 43920
rect 15243 43880 17592 43908
rect 15243 43877 15255 43880
rect 15197 43871 15255 43877
rect 16960 43852 16988 43880
rect 17586 43868 17592 43880
rect 17644 43868 17650 43920
rect 8352 43812 8892 43840
rect 8352 43800 8358 43812
rect 9674 43800 9680 43852
rect 9732 43840 9738 43852
rect 9953 43843 10011 43849
rect 9953 43840 9965 43843
rect 9732 43812 9965 43840
rect 9732 43800 9738 43812
rect 9953 43809 9965 43812
rect 9999 43809 10011 43843
rect 10318 43840 10324 43852
rect 10279 43812 10324 43840
rect 9953 43803 10011 43809
rect 10318 43800 10324 43812
rect 10376 43800 10382 43852
rect 10965 43843 11023 43849
rect 10965 43809 10977 43843
rect 11011 43840 11023 43843
rect 11514 43840 11520 43852
rect 11011 43812 11520 43840
rect 11011 43809 11023 43812
rect 10965 43803 11023 43809
rect 11514 43800 11520 43812
rect 11572 43800 11578 43852
rect 12713 43843 12771 43849
rect 12713 43809 12725 43843
rect 12759 43840 12771 43843
rect 13078 43840 13084 43852
rect 12759 43812 13084 43840
rect 12759 43809 12771 43812
rect 12713 43803 12771 43809
rect 13078 43800 13084 43812
rect 13136 43800 13142 43852
rect 13449 43843 13507 43849
rect 13449 43809 13461 43843
rect 13495 43840 13507 43843
rect 13538 43840 13544 43852
rect 13495 43812 13544 43840
rect 13495 43809 13507 43812
rect 13449 43803 13507 43809
rect 13538 43800 13544 43812
rect 13596 43800 13602 43852
rect 14274 43800 14280 43852
rect 14332 43840 14338 43852
rect 15746 43840 15752 43852
rect 14332 43812 15752 43840
rect 14332 43800 14338 43812
rect 15746 43800 15752 43812
rect 15804 43800 15810 43852
rect 16022 43840 16028 43852
rect 15983 43812 16028 43840
rect 16022 43800 16028 43812
rect 16080 43800 16086 43852
rect 16390 43840 16396 43852
rect 16351 43812 16396 43840
rect 16390 43800 16396 43812
rect 16448 43800 16454 43852
rect 16942 43840 16948 43852
rect 16855 43812 16948 43840
rect 16942 43800 16948 43812
rect 17000 43800 17006 43852
rect 1489 43775 1547 43781
rect 1489 43741 1501 43775
rect 1535 43772 1547 43775
rect 1670 43772 1676 43784
rect 1535 43744 1676 43772
rect 1535 43741 1547 43744
rect 1489 43735 1547 43741
rect 1670 43732 1676 43744
rect 1728 43732 1734 43784
rect 1765 43775 1823 43781
rect 1765 43741 1777 43775
rect 1811 43772 1823 43775
rect 1946 43772 1952 43784
rect 1811 43744 1952 43772
rect 1811 43741 1823 43744
rect 1765 43735 1823 43741
rect 1946 43732 1952 43744
rect 2004 43732 2010 43784
rect 4062 43772 4068 43784
rect 4023 43744 4068 43772
rect 4062 43732 4068 43744
rect 4120 43732 4126 43784
rect 4982 43772 4988 43784
rect 4895 43744 4988 43772
rect 3881 43707 3939 43713
rect 3881 43673 3893 43707
rect 3927 43704 3939 43707
rect 4908 43704 4936 43744
rect 4982 43732 4988 43744
rect 5040 43732 5046 43784
rect 9769 43775 9827 43781
rect 9769 43741 9781 43775
rect 9815 43772 9827 43775
rect 9858 43772 9864 43784
rect 9815 43744 9864 43772
rect 9815 43741 9827 43744
rect 9769 43735 9827 43741
rect 9858 43732 9864 43744
rect 9916 43732 9922 43784
rect 10410 43772 10416 43784
rect 10371 43744 10416 43772
rect 10410 43732 10416 43744
rect 10468 43732 10474 43784
rect 11701 43775 11759 43781
rect 11701 43741 11713 43775
rect 11747 43772 11759 43775
rect 12526 43772 12532 43784
rect 11747 43744 12532 43772
rect 11747 43741 11759 43744
rect 11701 43735 11759 43741
rect 12526 43732 12532 43744
rect 12584 43732 12590 43784
rect 12894 43732 12900 43784
rect 12952 43772 12958 43784
rect 13173 43775 13231 43781
rect 13173 43772 13185 43775
rect 12952 43744 13185 43772
rect 12952 43732 12958 43744
rect 13173 43741 13185 43744
rect 13219 43741 13231 43775
rect 16114 43772 16120 43784
rect 16075 43744 16120 43772
rect 13173 43735 13231 43741
rect 16114 43732 16120 43744
rect 16172 43732 16178 43784
rect 3927 43676 4936 43704
rect 5721 43707 5779 43713
rect 3927 43673 3939 43676
rect 3881 43667 3939 43673
rect 5721 43673 5733 43707
rect 5767 43704 5779 43707
rect 6638 43704 6644 43716
rect 5767 43676 6644 43704
rect 5767 43673 5779 43676
rect 5721 43667 5779 43673
rect 6638 43664 6644 43676
rect 6696 43664 6702 43716
rect 6914 43664 6920 43716
rect 6972 43704 6978 43716
rect 7745 43707 7803 43713
rect 7745 43704 7757 43707
rect 6972 43676 7757 43704
rect 6972 43664 6978 43676
rect 7745 43673 7757 43676
rect 7791 43673 7803 43707
rect 7745 43667 7803 43673
rect 3510 43636 3516 43648
rect 3471 43608 3516 43636
rect 3510 43596 3516 43608
rect 3568 43596 3574 43648
rect 6454 43596 6460 43648
rect 6512 43636 6518 43648
rect 6549 43639 6607 43645
rect 6549 43636 6561 43639
rect 6512 43608 6561 43636
rect 6512 43596 6518 43608
rect 6549 43605 6561 43608
rect 6595 43636 6607 43639
rect 6822 43636 6828 43648
rect 6595 43608 6828 43636
rect 6595 43605 6607 43608
rect 6549 43599 6607 43605
rect 6822 43596 6828 43608
rect 6880 43596 6886 43648
rect 8662 43596 8668 43648
rect 8720 43636 8726 43648
rect 8757 43639 8815 43645
rect 8757 43636 8769 43639
rect 8720 43608 8769 43636
rect 8720 43596 8726 43608
rect 8757 43605 8769 43608
rect 8803 43605 8815 43639
rect 8757 43599 8815 43605
rect 12710 43596 12716 43648
rect 12768 43636 12774 43648
rect 14553 43639 14611 43645
rect 14553 43636 14565 43639
rect 12768 43608 14565 43636
rect 12768 43596 12774 43608
rect 14553 43605 14565 43608
rect 14599 43605 14611 43639
rect 14553 43599 14611 43605
rect 14826 43596 14832 43648
rect 14884 43636 14890 43648
rect 15010 43636 15016 43648
rect 14884 43608 15016 43636
rect 14884 43596 14890 43608
rect 15010 43596 15016 43608
rect 15068 43596 15074 43648
rect 15930 43596 15936 43648
rect 15988 43636 15994 43648
rect 17405 43639 17463 43645
rect 17405 43636 17417 43639
rect 15988 43608 17417 43636
rect 15988 43596 15994 43608
rect 17405 43605 17417 43608
rect 17451 43605 17463 43639
rect 17405 43599 17463 43605
rect 1104 43546 18860 43568
rect 1104 43494 4315 43546
rect 4367 43494 4379 43546
rect 4431 43494 4443 43546
rect 4495 43494 4507 43546
rect 4559 43494 10982 43546
rect 11034 43494 11046 43546
rect 11098 43494 11110 43546
rect 11162 43494 11174 43546
rect 11226 43494 17648 43546
rect 17700 43494 17712 43546
rect 17764 43494 17776 43546
rect 17828 43494 17840 43546
rect 17892 43494 18860 43546
rect 1104 43472 18860 43494
rect 3513 43435 3571 43441
rect 3513 43401 3525 43435
rect 3559 43432 3571 43435
rect 3694 43432 3700 43444
rect 3559 43404 3700 43432
rect 3559 43401 3571 43404
rect 3513 43395 3571 43401
rect 3694 43392 3700 43404
rect 3752 43392 3758 43444
rect 3881 43435 3939 43441
rect 3881 43401 3893 43435
rect 3927 43432 3939 43435
rect 3970 43432 3976 43444
rect 3927 43404 3976 43432
rect 3927 43401 3939 43404
rect 3881 43395 3939 43401
rect 3970 43392 3976 43404
rect 4028 43392 4034 43444
rect 4062 43392 4068 43444
rect 4120 43432 4126 43444
rect 4157 43435 4215 43441
rect 4157 43432 4169 43435
rect 4120 43404 4169 43432
rect 4120 43392 4126 43404
rect 4157 43401 4169 43404
rect 4203 43432 4215 43435
rect 5077 43435 5135 43441
rect 5077 43432 5089 43435
rect 4203 43404 5089 43432
rect 4203 43401 4215 43404
rect 4157 43395 4215 43401
rect 5077 43401 5089 43404
rect 5123 43401 5135 43435
rect 5077 43395 5135 43401
rect 7006 43392 7012 43444
rect 7064 43432 7070 43444
rect 7377 43435 7435 43441
rect 7377 43432 7389 43435
rect 7064 43404 7389 43432
rect 7064 43392 7070 43404
rect 7377 43401 7389 43404
rect 7423 43401 7435 43435
rect 7377 43395 7435 43401
rect 7466 43392 7472 43444
rect 7524 43432 7530 43444
rect 7745 43435 7803 43441
rect 7745 43432 7757 43435
rect 7524 43404 7757 43432
rect 7524 43392 7530 43404
rect 7745 43401 7757 43404
rect 7791 43401 7803 43435
rect 8294 43432 8300 43444
rect 8255 43404 8300 43432
rect 7745 43395 7803 43401
rect 8294 43392 8300 43404
rect 8352 43392 8358 43444
rect 8478 43392 8484 43444
rect 8536 43432 8542 43444
rect 9033 43435 9091 43441
rect 9033 43432 9045 43435
rect 8536 43404 9045 43432
rect 8536 43392 8542 43404
rect 9033 43401 9045 43404
rect 9079 43401 9091 43435
rect 9033 43395 9091 43401
rect 9493 43435 9551 43441
rect 9493 43401 9505 43435
rect 9539 43432 9551 43435
rect 10778 43432 10784 43444
rect 9539 43404 10784 43432
rect 9539 43401 9551 43404
rect 9493 43395 9551 43401
rect 4890 43324 4896 43376
rect 4948 43364 4954 43376
rect 5534 43364 5540 43376
rect 4948 43336 5540 43364
rect 4948 43324 4954 43336
rect 5534 43324 5540 43336
rect 5592 43324 5598 43376
rect 6178 43364 6184 43376
rect 5920 43336 6184 43364
rect 1489 43299 1547 43305
rect 1489 43265 1501 43299
rect 1535 43296 1547 43299
rect 1670 43296 1676 43308
rect 1535 43268 1676 43296
rect 1535 43265 1547 43268
rect 1489 43259 1547 43265
rect 1670 43256 1676 43268
rect 1728 43256 1734 43308
rect 3145 43299 3203 43305
rect 3145 43265 3157 43299
rect 3191 43296 3203 43299
rect 3602 43296 3608 43308
rect 3191 43268 3608 43296
rect 3191 43265 3203 43268
rect 3145 43259 3203 43265
rect 3602 43256 3608 43268
rect 3660 43256 3666 43308
rect 1578 43188 1584 43240
rect 1636 43228 1642 43240
rect 1765 43231 1823 43237
rect 1765 43228 1777 43231
rect 1636 43200 1777 43228
rect 1636 43188 1642 43200
rect 1765 43197 1777 43200
rect 1811 43197 1823 43231
rect 1765 43191 1823 43197
rect 3694 43188 3700 43240
rect 3752 43228 3758 43240
rect 4065 43231 4123 43237
rect 4065 43228 4077 43231
rect 3752 43200 4077 43228
rect 3752 43188 3758 43200
rect 4065 43197 4077 43200
rect 4111 43197 4123 43231
rect 4065 43191 4123 43197
rect 4801 43231 4859 43237
rect 4801 43197 4813 43231
rect 4847 43228 4859 43231
rect 4890 43228 4896 43240
rect 4847 43200 4896 43228
rect 4847 43197 4859 43200
rect 4801 43191 4859 43197
rect 4890 43188 4896 43200
rect 4948 43188 4954 43240
rect 5920 43237 5948 43336
rect 6178 43324 6184 43336
rect 6236 43324 6242 43376
rect 7282 43324 7288 43376
rect 7340 43364 7346 43376
rect 7484 43364 7512 43392
rect 7340 43336 7512 43364
rect 9048 43364 9076 43395
rect 9048 43336 9996 43364
rect 7340 43324 7346 43336
rect 6270 43296 6276 43308
rect 6231 43268 6276 43296
rect 6270 43256 6276 43268
rect 6328 43256 6334 43308
rect 9858 43296 9864 43308
rect 9819 43268 9864 43296
rect 9858 43256 9864 43268
rect 9916 43256 9922 43308
rect 5905 43231 5963 43237
rect 5905 43197 5917 43231
rect 5951 43197 5963 43231
rect 5905 43191 5963 43197
rect 5997 43231 6055 43237
rect 5997 43197 6009 43231
rect 6043 43197 6055 43231
rect 5997 43191 6055 43197
rect 5537 43095 5595 43101
rect 5537 43061 5549 43095
rect 5583 43092 5595 43095
rect 5810 43092 5816 43104
rect 5583 43064 5816 43092
rect 5583 43061 5595 43064
rect 5537 43055 5595 43061
rect 5810 43052 5816 43064
rect 5868 43092 5874 43104
rect 6012 43092 6040 43191
rect 6086 43188 6092 43240
rect 6144 43228 6150 43240
rect 6365 43231 6423 43237
rect 6365 43228 6377 43231
rect 6144 43200 6377 43228
rect 6144 43188 6150 43200
rect 6365 43197 6377 43200
rect 6411 43197 6423 43231
rect 6365 43191 6423 43197
rect 6638 43188 6644 43240
rect 6696 43228 6702 43240
rect 6917 43231 6975 43237
rect 6917 43228 6929 43231
rect 6696 43200 6929 43228
rect 6696 43188 6702 43200
rect 6917 43197 6929 43200
rect 6963 43197 6975 43231
rect 6917 43191 6975 43197
rect 7190 43188 7196 43240
rect 7248 43228 7254 43240
rect 8570 43228 8576 43240
rect 7248 43200 8576 43228
rect 7248 43188 7254 43200
rect 8570 43188 8576 43200
rect 8628 43188 8634 43240
rect 9769 43231 9827 43237
rect 9769 43197 9781 43231
rect 9815 43197 9827 43231
rect 9968 43228 9996 43336
rect 10045 43231 10103 43237
rect 10045 43228 10057 43231
rect 9968 43200 10057 43228
rect 9769 43191 9827 43197
rect 10045 43197 10057 43200
rect 10091 43197 10103 43231
rect 10045 43191 10103 43197
rect 9784 43160 9812 43191
rect 10318 43188 10324 43240
rect 10376 43228 10382 43240
rect 10428 43237 10456 43404
rect 10778 43392 10784 43404
rect 10836 43392 10842 43444
rect 11514 43432 11520 43444
rect 11475 43404 11520 43432
rect 11514 43392 11520 43404
rect 11572 43392 11578 43444
rect 12345 43435 12403 43441
rect 12345 43401 12357 43435
rect 12391 43432 12403 43435
rect 12618 43432 12624 43444
rect 12391 43404 12624 43432
rect 12391 43401 12403 43404
rect 12345 43395 12403 43401
rect 12544 43237 12572 43404
rect 12618 43392 12624 43404
rect 12676 43392 12682 43444
rect 13538 43432 13544 43444
rect 13499 43404 13544 43432
rect 13538 43392 13544 43404
rect 13596 43392 13602 43444
rect 13814 43392 13820 43444
rect 13872 43432 13878 43444
rect 14185 43435 14243 43441
rect 14185 43432 14197 43435
rect 13872 43404 14197 43432
rect 13872 43392 13878 43404
rect 14185 43401 14197 43404
rect 14231 43401 14243 43435
rect 14185 43395 14243 43401
rect 15105 43435 15163 43441
rect 15105 43401 15117 43435
rect 15151 43432 15163 43435
rect 16022 43432 16028 43444
rect 15151 43404 16028 43432
rect 15151 43401 15163 43404
rect 15105 43395 15163 43401
rect 16022 43392 16028 43404
rect 16080 43392 16086 43444
rect 13909 43367 13967 43373
rect 13909 43333 13921 43367
rect 13955 43364 13967 43367
rect 14274 43364 14280 43376
rect 13955 43336 14280 43364
rect 13955 43333 13967 43336
rect 13909 43327 13967 43333
rect 14274 43324 14280 43336
rect 14332 43324 14338 43376
rect 14384 43336 17448 43364
rect 13173 43299 13231 43305
rect 13173 43265 13185 43299
rect 13219 43296 13231 43299
rect 13722 43296 13728 43308
rect 13219 43268 13728 43296
rect 13219 43265 13231 43268
rect 13173 43259 13231 43265
rect 13722 43256 13728 43268
rect 13780 43256 13786 43308
rect 14182 43256 14188 43308
rect 14240 43296 14246 43308
rect 14384 43296 14412 43336
rect 14240 43268 14412 43296
rect 14240 43256 14246 43268
rect 16942 43256 16948 43308
rect 17000 43296 17006 43308
rect 17420 43305 17448 43336
rect 17405 43299 17463 43305
rect 17000 43268 17356 43296
rect 17000 43256 17006 43268
rect 10413 43231 10471 43237
rect 10413 43228 10425 43231
rect 10376 43200 10425 43228
rect 10376 43188 10382 43200
rect 10413 43197 10425 43200
rect 10459 43197 10471 43231
rect 10413 43191 10471 43197
rect 11977 43231 12035 43237
rect 11977 43197 11989 43231
rect 12023 43228 12035 43231
rect 12529 43231 12587 43237
rect 12023 43200 12480 43228
rect 12023 43197 12035 43200
rect 11977 43191 12035 43197
rect 10778 43160 10784 43172
rect 9784 43132 10784 43160
rect 10778 43120 10784 43132
rect 10836 43160 10842 43172
rect 12452 43160 12480 43200
rect 12529 43197 12541 43231
rect 12575 43197 12587 43231
rect 12897 43231 12955 43237
rect 12897 43228 12909 43231
rect 12529 43191 12587 43197
rect 12636 43200 12909 43228
rect 12636 43172 12664 43200
rect 12897 43197 12909 43200
rect 12943 43197 12955 43231
rect 12897 43191 12955 43197
rect 13814 43188 13820 43240
rect 13872 43228 13878 43240
rect 14001 43231 14059 43237
rect 14001 43228 14013 43231
rect 13872 43200 14013 43228
rect 13872 43188 13878 43200
rect 14001 43197 14013 43200
rect 14047 43228 14059 43231
rect 14461 43231 14519 43237
rect 14461 43228 14473 43231
rect 14047 43200 14473 43228
rect 14047 43197 14059 43200
rect 14001 43191 14059 43197
rect 14461 43197 14473 43200
rect 14507 43197 14519 43231
rect 14461 43191 14519 43197
rect 15930 43188 15936 43240
rect 15988 43228 15994 43240
rect 16025 43231 16083 43237
rect 16025 43228 16037 43231
rect 15988 43200 16037 43228
rect 15988 43188 15994 43200
rect 16025 43197 16037 43200
rect 16071 43197 16083 43231
rect 16666 43228 16672 43240
rect 16627 43200 16672 43228
rect 16025 43191 16083 43197
rect 16666 43188 16672 43200
rect 16724 43188 16730 43240
rect 17328 43237 17356 43268
rect 17405 43265 17417 43299
rect 17451 43296 17463 43299
rect 18414 43296 18420 43308
rect 17451 43268 18420 43296
rect 17451 43265 17463 43268
rect 17405 43259 17463 43265
rect 18414 43256 18420 43268
rect 18472 43256 18478 43308
rect 17037 43231 17095 43237
rect 17037 43197 17049 43231
rect 17083 43197 17095 43231
rect 17037 43191 17095 43197
rect 17313 43231 17371 43237
rect 17313 43197 17325 43231
rect 17359 43197 17371 43231
rect 17313 43191 17371 43197
rect 12618 43160 12624 43172
rect 10836 43132 12204 43160
rect 12452 43132 12624 43160
rect 10836 43120 10842 43132
rect 5868 43064 6040 43092
rect 11241 43095 11299 43101
rect 5868 43052 5874 43064
rect 11241 43061 11253 43095
rect 11287 43092 11299 43095
rect 12066 43092 12072 43104
rect 11287 43064 12072 43092
rect 11287 43061 11299 43064
rect 11241 43055 11299 43061
rect 12066 43052 12072 43064
rect 12124 43052 12130 43104
rect 12176 43092 12204 43132
rect 12618 43120 12624 43132
rect 12676 43120 12682 43172
rect 14366 43120 14372 43172
rect 14424 43160 14430 43172
rect 14826 43160 14832 43172
rect 14424 43132 14832 43160
rect 14424 43120 14430 43132
rect 14826 43120 14832 43132
rect 14884 43120 14890 43172
rect 17052 43160 17080 43191
rect 17052 43132 17908 43160
rect 17328 43104 17356 43132
rect 13078 43092 13084 43104
rect 12176 43064 13084 43092
rect 13078 43052 13084 43064
rect 13136 43052 13142 43104
rect 13538 43052 13544 43104
rect 13596 43092 13602 43104
rect 14918 43092 14924 43104
rect 13596 43064 14924 43092
rect 13596 43052 13602 43064
rect 14918 43052 14924 43064
rect 14976 43052 14982 43104
rect 15378 43052 15384 43104
rect 15436 43092 15442 43104
rect 15657 43095 15715 43101
rect 15657 43092 15669 43095
rect 15436 43064 15669 43092
rect 15436 43052 15442 43064
rect 15657 43061 15669 43064
rect 15703 43061 15715 43095
rect 15657 43055 15715 43061
rect 17310 43052 17316 43104
rect 17368 43052 17374 43104
rect 17880 43101 17908 43132
rect 17865 43095 17923 43101
rect 17865 43061 17877 43095
rect 17911 43092 17923 43095
rect 18046 43092 18052 43104
rect 17911 43064 18052 43092
rect 17911 43061 17923 43064
rect 17865 43055 17923 43061
rect 18046 43052 18052 43064
rect 18104 43052 18110 43104
rect 1104 43002 18860 43024
rect 1104 42950 7648 43002
rect 7700 42950 7712 43002
rect 7764 42950 7776 43002
rect 7828 42950 7840 43002
rect 7892 42950 14315 43002
rect 14367 42950 14379 43002
rect 14431 42950 14443 43002
rect 14495 42950 14507 43002
rect 14559 42950 18860 43002
rect 1104 42928 18860 42950
rect 1670 42848 1676 42900
rect 1728 42888 1734 42900
rect 2317 42891 2375 42897
rect 2317 42888 2329 42891
rect 1728 42860 2329 42888
rect 1728 42848 1734 42860
rect 2317 42857 2329 42860
rect 2363 42857 2375 42891
rect 2317 42851 2375 42857
rect 3786 42848 3792 42900
rect 3844 42888 3850 42900
rect 4062 42888 4068 42900
rect 3844 42860 4068 42888
rect 3844 42848 3850 42860
rect 4062 42848 4068 42860
rect 4120 42848 4126 42900
rect 4982 42888 4988 42900
rect 4943 42860 4988 42888
rect 4982 42848 4988 42860
rect 5040 42848 5046 42900
rect 6089 42891 6147 42897
rect 6089 42857 6101 42891
rect 6135 42888 6147 42891
rect 6178 42888 6184 42900
rect 6135 42860 6184 42888
rect 6135 42857 6147 42860
rect 6089 42851 6147 42857
rect 6178 42848 6184 42860
rect 6236 42848 6242 42900
rect 8386 42888 8392 42900
rect 7944 42860 8392 42888
rect 7944 42832 7972 42860
rect 8386 42848 8392 42860
rect 8444 42848 8450 42900
rect 8570 42848 8576 42900
rect 8628 42848 8634 42900
rect 10226 42848 10232 42900
rect 10284 42888 10290 42900
rect 10505 42891 10563 42897
rect 10505 42888 10517 42891
rect 10284 42860 10517 42888
rect 10284 42848 10290 42860
rect 10505 42857 10517 42860
rect 10551 42857 10563 42891
rect 10505 42851 10563 42857
rect 11885 42891 11943 42897
rect 11885 42857 11897 42891
rect 11931 42888 11943 42891
rect 12434 42888 12440 42900
rect 11931 42860 12440 42888
rect 11931 42857 11943 42860
rect 11885 42851 11943 42857
rect 12434 42848 12440 42860
rect 12492 42888 12498 42900
rect 12710 42888 12716 42900
rect 12492 42860 12716 42888
rect 12492 42848 12498 42860
rect 12710 42848 12716 42860
rect 12768 42848 12774 42900
rect 14277 42891 14335 42897
rect 14277 42857 14289 42891
rect 14323 42888 14335 42891
rect 15102 42888 15108 42900
rect 14323 42860 15108 42888
rect 14323 42857 14335 42860
rect 14277 42851 14335 42857
rect 15102 42848 15108 42860
rect 15160 42888 15166 42900
rect 16666 42888 16672 42900
rect 15160 42860 16068 42888
rect 16627 42860 16672 42888
rect 15160 42848 15166 42860
rect 6641 42823 6699 42829
rect 6641 42789 6653 42823
rect 6687 42820 6699 42823
rect 7190 42820 7196 42832
rect 6687 42792 7196 42820
rect 6687 42789 6699 42792
rect 6641 42783 6699 42789
rect 7190 42780 7196 42792
rect 7248 42780 7254 42832
rect 7926 42780 7932 42832
rect 7984 42780 7990 42832
rect 8110 42780 8116 42832
rect 8168 42820 8174 42832
rect 8588 42820 8616 42848
rect 10778 42820 10784 42832
rect 8168 42792 8524 42820
rect 8588 42792 9168 42820
rect 8168 42780 8174 42792
rect 8496 42764 8524 42792
rect 3510 42712 3516 42764
rect 3568 42752 3574 42764
rect 3697 42755 3755 42761
rect 3697 42752 3709 42755
rect 3568 42724 3709 42752
rect 3568 42712 3574 42724
rect 3697 42721 3709 42724
rect 3743 42752 3755 42755
rect 4890 42752 4896 42764
rect 3743 42724 4896 42752
rect 3743 42721 3755 42724
rect 3697 42715 3755 42721
rect 4890 42712 4896 42724
rect 4948 42712 4954 42764
rect 8205 42755 8263 42761
rect 8205 42721 8217 42755
rect 8251 42721 8263 42755
rect 8386 42752 8392 42764
rect 8347 42724 8392 42752
rect 8205 42715 8263 42721
rect 1946 42684 1952 42696
rect 1907 42656 1952 42684
rect 1946 42644 1952 42656
rect 2004 42644 2010 42696
rect 3418 42684 3424 42696
rect 3379 42656 3424 42684
rect 3418 42644 3424 42656
rect 3476 42644 3482 42696
rect 8220 42684 8248 42715
rect 8386 42712 8392 42724
rect 8444 42712 8450 42764
rect 8478 42712 8484 42764
rect 8536 42752 8542 42764
rect 9140 42761 9168 42792
rect 10060 42792 10784 42820
rect 8757 42755 8815 42761
rect 8757 42752 8769 42755
rect 8536 42724 8769 42752
rect 8536 42712 8542 42724
rect 8757 42721 8769 42724
rect 8803 42721 8815 42755
rect 8757 42715 8815 42721
rect 9125 42755 9183 42761
rect 9125 42721 9137 42755
rect 9171 42721 9183 42755
rect 9125 42715 9183 42721
rect 9582 42712 9588 42764
rect 9640 42752 9646 42764
rect 9677 42755 9735 42761
rect 9677 42752 9689 42755
rect 9640 42724 9689 42752
rect 9640 42712 9646 42724
rect 9677 42721 9689 42724
rect 9723 42721 9735 42755
rect 9677 42715 9735 42721
rect 8294 42684 8300 42696
rect 8207 42656 8300 42684
rect 8294 42644 8300 42656
rect 8352 42684 8358 42696
rect 9766 42684 9772 42696
rect 8352 42656 9772 42684
rect 8352 42644 8358 42656
rect 9766 42644 9772 42656
rect 9824 42644 9830 42696
rect 5721 42619 5779 42625
rect 5721 42585 5733 42619
rect 5767 42616 5779 42619
rect 6086 42616 6092 42628
rect 5767 42588 6092 42616
rect 5767 42585 5779 42588
rect 5721 42579 5779 42585
rect 6086 42576 6092 42588
rect 6144 42576 6150 42628
rect 8205 42619 8263 42625
rect 8205 42585 8217 42619
rect 8251 42616 8263 42619
rect 8662 42616 8668 42628
rect 8251 42588 8668 42616
rect 8251 42585 8263 42588
rect 8205 42579 8263 42585
rect 8662 42576 8668 42588
rect 8720 42576 8726 42628
rect 10060 42616 10088 42792
rect 10778 42780 10784 42792
rect 10836 42780 10842 42832
rect 11514 42820 11520 42832
rect 11475 42792 11520 42820
rect 11514 42780 11520 42792
rect 11572 42780 11578 42832
rect 13262 42780 13268 42832
rect 13320 42820 13326 42832
rect 15562 42820 15568 42832
rect 13320 42792 13860 42820
rect 13320 42780 13326 42792
rect 13832 42764 13860 42792
rect 15120 42792 15568 42820
rect 10226 42752 10232 42764
rect 10187 42724 10232 42752
rect 10226 42712 10232 42724
rect 10284 42712 10290 42764
rect 10686 42712 10692 42764
rect 10744 42752 10750 42764
rect 10965 42755 11023 42761
rect 10965 42752 10977 42755
rect 10744 42724 10977 42752
rect 10744 42712 10750 42724
rect 10965 42721 10977 42724
rect 11011 42721 11023 42755
rect 10965 42715 11023 42721
rect 11057 42755 11115 42761
rect 11057 42721 11069 42755
rect 11103 42721 11115 42755
rect 11057 42715 11115 42721
rect 12253 42755 12311 42761
rect 12253 42721 12265 42755
rect 12299 42752 12311 42755
rect 12897 42755 12955 42761
rect 12897 42752 12909 42755
rect 12299 42724 12909 42752
rect 12299 42721 12311 42724
rect 12253 42715 12311 42721
rect 12897 42721 12909 42724
rect 12943 42752 12955 42755
rect 13538 42752 13544 42764
rect 12943 42724 13544 42752
rect 12943 42721 12955 42724
rect 12897 42715 12955 42721
rect 10244 42684 10272 42712
rect 11072 42684 11100 42715
rect 13538 42712 13544 42724
rect 13596 42712 13602 42764
rect 13814 42752 13820 42764
rect 13727 42724 13820 42752
rect 13814 42712 13820 42724
rect 13872 42712 13878 42764
rect 14829 42755 14887 42761
rect 14829 42721 14841 42755
rect 14875 42752 14887 42755
rect 15120 42752 15148 42792
rect 15562 42780 15568 42792
rect 15620 42780 15626 42832
rect 14875 42724 15148 42752
rect 15197 42755 15255 42761
rect 14875 42721 14887 42724
rect 14829 42715 14887 42721
rect 15197 42721 15209 42755
rect 15243 42721 15255 42755
rect 15381 42755 15439 42761
rect 15381 42752 15393 42755
rect 15197 42715 15255 42721
rect 15304 42724 15393 42752
rect 10244 42656 11100 42684
rect 13078 42644 13084 42696
rect 13136 42684 13142 42696
rect 13173 42687 13231 42693
rect 13173 42684 13185 42687
rect 13136 42656 13185 42684
rect 13136 42644 13142 42656
rect 13173 42653 13185 42656
rect 13219 42684 13231 42687
rect 14182 42684 14188 42696
rect 13219 42656 14188 42684
rect 13219 42653 13231 42656
rect 13173 42647 13231 42653
rect 14182 42644 14188 42656
rect 14240 42644 14246 42696
rect 10502 42616 10508 42628
rect 8864 42588 10088 42616
rect 10463 42588 10508 42616
rect 1486 42508 1492 42560
rect 1544 42548 1550 42560
rect 1581 42551 1639 42557
rect 1581 42548 1593 42551
rect 1544 42520 1593 42548
rect 1544 42508 1550 42520
rect 1581 42517 1593 42520
rect 1627 42517 1639 42551
rect 7006 42548 7012 42560
rect 6967 42520 7012 42548
rect 1581 42511 1639 42517
rect 7006 42508 7012 42520
rect 7064 42508 7070 42560
rect 7742 42548 7748 42560
rect 7703 42520 7748 42548
rect 7742 42508 7748 42520
rect 7800 42508 7806 42560
rect 8110 42508 8116 42560
rect 8168 42548 8174 42560
rect 8864 42548 8892 42588
rect 10502 42576 10508 42588
rect 10560 42576 10566 42628
rect 10778 42616 10784 42628
rect 10739 42588 10784 42616
rect 10778 42576 10784 42588
rect 10836 42576 10842 42628
rect 13909 42619 13967 42625
rect 13909 42585 13921 42619
rect 13955 42616 13967 42619
rect 14918 42616 14924 42628
rect 13955 42588 14924 42616
rect 13955 42585 13967 42588
rect 13909 42579 13967 42585
rect 14918 42576 14924 42588
rect 14976 42576 14982 42628
rect 15212 42616 15240 42715
rect 15304 42696 15332 42724
rect 15381 42721 15393 42724
rect 15427 42721 15439 42755
rect 15930 42752 15936 42764
rect 15891 42724 15936 42752
rect 15381 42715 15439 42721
rect 15930 42712 15936 42724
rect 15988 42712 15994 42764
rect 16040 42752 16068 42860
rect 16666 42848 16672 42860
rect 16724 42848 16730 42900
rect 16209 42755 16267 42761
rect 16209 42752 16221 42755
rect 16040 42724 16221 42752
rect 16209 42721 16221 42724
rect 16255 42721 16267 42755
rect 16209 42715 16267 42721
rect 15286 42644 15292 42696
rect 15344 42644 15350 42696
rect 15562 42616 15568 42628
rect 15212 42588 15568 42616
rect 15562 42576 15568 42588
rect 15620 42616 15626 42628
rect 16666 42616 16672 42628
rect 15620 42588 16672 42616
rect 15620 42576 15626 42588
rect 16666 42576 16672 42588
rect 16724 42576 16730 42628
rect 8168 42520 8892 42548
rect 8168 42508 8174 42520
rect 9398 42508 9404 42560
rect 9456 42548 9462 42560
rect 9766 42548 9772 42560
rect 9456 42520 9772 42548
rect 9456 42508 9462 42520
rect 9766 42508 9772 42520
rect 9824 42508 9830 42560
rect 10686 42548 10692 42560
rect 10647 42520 10692 42548
rect 10686 42508 10692 42520
rect 10744 42508 10750 42560
rect 13170 42508 13176 42560
rect 13228 42548 13234 42560
rect 14277 42551 14335 42557
rect 14277 42548 14289 42551
rect 13228 42520 14289 42548
rect 13228 42508 13234 42520
rect 14277 42517 14289 42520
rect 14323 42517 14335 42551
rect 14277 42511 14335 42517
rect 14461 42551 14519 42557
rect 14461 42517 14473 42551
rect 14507 42548 14519 42551
rect 14826 42548 14832 42560
rect 14507 42520 14832 42548
rect 14507 42517 14519 42520
rect 14461 42511 14519 42517
rect 14826 42508 14832 42520
rect 14884 42548 14890 42560
rect 15930 42548 15936 42560
rect 14884 42520 15936 42548
rect 14884 42508 14890 42520
rect 15930 42508 15936 42520
rect 15988 42508 15994 42560
rect 16022 42508 16028 42560
rect 16080 42548 16086 42560
rect 16117 42551 16175 42557
rect 16117 42548 16129 42551
rect 16080 42520 16129 42548
rect 16080 42508 16086 42520
rect 16117 42517 16129 42520
rect 16163 42517 16175 42551
rect 16117 42511 16175 42517
rect 16390 42508 16396 42560
rect 16448 42548 16454 42560
rect 17037 42551 17095 42557
rect 17037 42548 17049 42551
rect 16448 42520 17049 42548
rect 16448 42508 16454 42520
rect 17037 42517 17049 42520
rect 17083 42548 17095 42551
rect 17405 42551 17463 42557
rect 17405 42548 17417 42551
rect 17083 42520 17417 42548
rect 17083 42517 17095 42520
rect 17037 42511 17095 42517
rect 17405 42517 17417 42520
rect 17451 42517 17463 42551
rect 17405 42511 17463 42517
rect 1104 42458 18860 42480
rect 1104 42406 4315 42458
rect 4367 42406 4379 42458
rect 4431 42406 4443 42458
rect 4495 42406 4507 42458
rect 4559 42406 10982 42458
rect 11034 42406 11046 42458
rect 11098 42406 11110 42458
rect 11162 42406 11174 42458
rect 11226 42406 17648 42458
rect 17700 42406 17712 42458
rect 17764 42406 17776 42458
rect 17828 42406 17840 42458
rect 17892 42406 18860 42458
rect 1104 42384 18860 42406
rect 2866 42344 2872 42356
rect 2827 42316 2872 42344
rect 2866 42304 2872 42316
rect 2924 42304 2930 42356
rect 3510 42344 3516 42356
rect 3471 42316 3516 42344
rect 3510 42304 3516 42316
rect 3568 42304 3574 42356
rect 4154 42304 4160 42356
rect 4212 42344 4218 42356
rect 4341 42347 4399 42353
rect 4341 42344 4353 42347
rect 4212 42316 4353 42344
rect 4212 42304 4218 42316
rect 4341 42313 4353 42316
rect 4387 42313 4399 42347
rect 4341 42307 4399 42313
rect 4801 42347 4859 42353
rect 4801 42313 4813 42347
rect 4847 42344 4859 42347
rect 5994 42344 6000 42356
rect 4847 42316 6000 42344
rect 4847 42313 4859 42316
rect 4801 42307 4859 42313
rect 1489 42211 1547 42217
rect 1489 42177 1501 42211
rect 1535 42208 1547 42211
rect 1670 42208 1676 42220
rect 1535 42180 1676 42208
rect 1535 42177 1547 42180
rect 1489 42171 1547 42177
rect 1670 42168 1676 42180
rect 1728 42168 1734 42220
rect 4356 42208 4384 42307
rect 5994 42304 6000 42316
rect 6052 42304 6058 42356
rect 7193 42347 7251 42353
rect 7193 42313 7205 42347
rect 7239 42344 7251 42347
rect 8386 42344 8392 42356
rect 7239 42316 8392 42344
rect 7239 42313 7251 42316
rect 7193 42307 7251 42313
rect 8386 42304 8392 42316
rect 8444 42304 8450 42356
rect 8938 42304 8944 42356
rect 8996 42344 9002 42356
rect 9398 42344 9404 42356
rect 8996 42316 9404 42344
rect 8996 42304 9002 42316
rect 9398 42304 9404 42316
rect 9456 42304 9462 42356
rect 9493 42347 9551 42353
rect 9493 42313 9505 42347
rect 9539 42344 9551 42347
rect 9582 42344 9588 42356
rect 9539 42316 9588 42344
rect 9539 42313 9551 42316
rect 9493 42307 9551 42313
rect 4890 42236 4896 42288
rect 4948 42276 4954 42288
rect 4985 42279 5043 42285
rect 4985 42276 4997 42279
rect 4948 42248 4997 42276
rect 4948 42236 4954 42248
rect 4985 42245 4997 42248
rect 5031 42245 5043 42279
rect 7558 42276 7564 42288
rect 7519 42248 7564 42276
rect 4985 42239 5043 42245
rect 7558 42236 7564 42248
rect 7616 42236 7622 42288
rect 7742 42208 7748 42220
rect 4356 42180 5764 42208
rect 7703 42180 7748 42208
rect 1578 42100 1584 42152
rect 1636 42140 1642 42152
rect 1765 42143 1823 42149
rect 1765 42140 1777 42143
rect 1636 42112 1777 42140
rect 1636 42100 1642 42112
rect 1765 42109 1777 42112
rect 1811 42109 1823 42143
rect 5166 42140 5172 42152
rect 5127 42112 5172 42140
rect 1765 42103 1823 42109
rect 5166 42100 5172 42112
rect 5224 42100 5230 42152
rect 5736 42149 5764 42180
rect 7742 42168 7748 42180
rect 7800 42168 7806 42220
rect 7837 42211 7895 42217
rect 7837 42177 7849 42211
rect 7883 42208 7895 42211
rect 9508 42208 9536 42307
rect 9582 42304 9588 42316
rect 9640 42304 9646 42356
rect 9861 42347 9919 42353
rect 9861 42313 9873 42347
rect 9907 42313 9919 42347
rect 10226 42344 10232 42356
rect 10187 42316 10232 42344
rect 9861 42307 9919 42313
rect 9876 42276 9904 42307
rect 10226 42304 10232 42316
rect 10284 42304 10290 42356
rect 10686 42304 10692 42356
rect 10744 42344 10750 42356
rect 10781 42347 10839 42353
rect 10781 42344 10793 42347
rect 10744 42316 10793 42344
rect 10744 42304 10750 42316
rect 10781 42313 10793 42316
rect 10827 42313 10839 42347
rect 10781 42307 10839 42313
rect 11422 42304 11428 42356
rect 11480 42344 11486 42356
rect 12161 42347 12219 42353
rect 12161 42344 12173 42347
rect 11480 42316 12173 42344
rect 11480 42304 11486 42316
rect 12161 42313 12173 42316
rect 12207 42313 12219 42347
rect 12161 42307 12219 42313
rect 13078 42304 13084 42356
rect 13136 42344 13142 42356
rect 13136 42316 13181 42344
rect 13136 42304 13142 42316
rect 13998 42304 14004 42356
rect 14056 42344 14062 42356
rect 14182 42344 14188 42356
rect 14056 42316 14188 42344
rect 14056 42304 14062 42316
rect 14182 42304 14188 42316
rect 14240 42304 14246 42356
rect 14826 42304 14832 42356
rect 14884 42344 14890 42356
rect 15013 42347 15071 42353
rect 15013 42344 15025 42347
rect 14884 42316 15025 42344
rect 14884 42304 14890 42316
rect 15013 42313 15025 42316
rect 15059 42344 15071 42347
rect 15286 42344 15292 42356
rect 15059 42316 15292 42344
rect 15059 42313 15071 42316
rect 15013 42307 15071 42313
rect 15286 42304 15292 42316
rect 15344 42304 15350 42356
rect 15562 42344 15568 42356
rect 15523 42316 15568 42344
rect 15562 42304 15568 42316
rect 15620 42304 15626 42356
rect 11440 42276 11468 42304
rect 9876 42248 11468 42276
rect 9858 42208 9864 42220
rect 7883 42180 9536 42208
rect 9600 42180 9864 42208
rect 7883 42177 7895 42180
rect 7837 42171 7895 42177
rect 5629 42143 5687 42149
rect 5629 42109 5641 42143
rect 5675 42109 5687 42143
rect 5629 42103 5687 42109
rect 5721 42143 5779 42149
rect 5721 42109 5733 42143
rect 5767 42109 5779 42143
rect 5721 42103 5779 42109
rect 3881 42075 3939 42081
rect 3881 42041 3893 42075
rect 3927 42072 3939 42075
rect 5644 42072 5672 42103
rect 5994 42100 6000 42152
rect 6052 42140 6058 42152
rect 6089 42143 6147 42149
rect 6089 42140 6101 42143
rect 6052 42112 6101 42140
rect 6052 42100 6058 42112
rect 6089 42109 6101 42112
rect 6135 42140 6147 42143
rect 6270 42140 6276 42152
rect 6135 42112 6276 42140
rect 6135 42109 6147 42112
rect 6089 42103 6147 42109
rect 6270 42100 6276 42112
rect 6328 42100 6334 42152
rect 6733 42143 6791 42149
rect 6733 42109 6745 42143
rect 6779 42140 6791 42143
rect 8573 42143 8631 42149
rect 8573 42140 8585 42143
rect 6779 42112 8585 42140
rect 6779 42109 6791 42112
rect 6733 42103 6791 42109
rect 8573 42109 8585 42112
rect 8619 42109 8631 42143
rect 8573 42103 8631 42109
rect 8665 42143 8723 42149
rect 8665 42109 8677 42143
rect 8711 42140 8723 42143
rect 8938 42140 8944 42152
rect 8711 42112 8944 42140
rect 8711 42109 8723 42112
rect 8665 42103 8723 42109
rect 7466 42072 7472 42084
rect 3927 42044 7472 42072
rect 3927 42041 3939 42044
rect 3881 42035 3939 42041
rect 7466 42032 7472 42044
rect 7524 42032 7530 42084
rect 7926 42032 7932 42084
rect 7984 42072 7990 42084
rect 8588 42072 8616 42103
rect 8938 42100 8944 42112
rect 8996 42140 9002 42152
rect 9125 42143 9183 42149
rect 9125 42140 9137 42143
rect 8996 42112 9137 42140
rect 8996 42100 9002 42112
rect 9125 42109 9137 42112
rect 9171 42140 9183 42143
rect 9600 42140 9628 42180
rect 9858 42168 9864 42180
rect 9916 42168 9922 42220
rect 9171 42112 9628 42140
rect 9677 42143 9735 42149
rect 9171 42109 9183 42112
rect 9125 42103 9183 42109
rect 9677 42109 9689 42143
rect 9723 42140 9735 42143
rect 10226 42140 10232 42152
rect 9723 42112 10232 42140
rect 9723 42109 9735 42112
rect 9677 42103 9735 42109
rect 10226 42100 10232 42112
rect 10284 42100 10290 42152
rect 10520 42140 10548 42248
rect 13538 42236 13544 42288
rect 13596 42236 13602 42288
rect 15304 42276 15332 42304
rect 15930 42276 15936 42288
rect 15304 42248 15936 42276
rect 15930 42236 15936 42248
rect 15988 42236 15994 42288
rect 17221 42279 17279 42285
rect 17221 42245 17233 42279
rect 17267 42276 17279 42279
rect 17770 42276 17776 42288
rect 17267 42248 17776 42276
rect 17267 42245 17279 42248
rect 17221 42239 17279 42245
rect 17770 42236 17776 42248
rect 17828 42276 17834 42288
rect 18322 42276 18328 42288
rect 17828 42248 18328 42276
rect 17828 42236 17834 42248
rect 18322 42236 18328 42248
rect 18380 42236 18386 42288
rect 10597 42211 10655 42217
rect 10597 42177 10609 42211
rect 10643 42208 10655 42211
rect 10643 42180 11652 42208
rect 10643 42177 10655 42180
rect 10597 42171 10655 42177
rect 11624 42152 11652 42180
rect 12158 42168 12164 42220
rect 12216 42208 12222 42220
rect 12986 42208 12992 42220
rect 12216 42180 12992 42208
rect 12216 42168 12222 42180
rect 12986 42168 12992 42180
rect 13044 42168 13050 42220
rect 13262 42168 13268 42220
rect 13320 42208 13326 42220
rect 13556 42208 13584 42236
rect 17310 42208 17316 42220
rect 13320 42180 13676 42208
rect 13320 42168 13326 42180
rect 10686 42140 10692 42152
rect 10520 42112 10692 42140
rect 10686 42100 10692 42112
rect 10744 42100 10750 42152
rect 11333 42143 11391 42149
rect 11333 42109 11345 42143
rect 11379 42109 11391 42143
rect 11333 42103 11391 42109
rect 9030 42072 9036 42084
rect 7984 42044 8524 42072
rect 8588 42044 9036 42072
rect 7984 42032 7990 42044
rect 4246 41964 4252 42016
rect 4304 42004 4310 42016
rect 5258 42004 5264 42016
rect 4304 41976 5264 42004
rect 4304 41964 4310 41976
rect 5258 41964 5264 41976
rect 5316 41964 5322 42016
rect 8496 42004 8524 42044
rect 9030 42032 9036 42044
rect 9088 42032 9094 42084
rect 11348 42072 11376 42103
rect 11606 42100 11612 42152
rect 11664 42140 11670 42152
rect 11701 42143 11759 42149
rect 11701 42140 11713 42143
rect 11664 42112 11713 42140
rect 11664 42100 11670 42112
rect 11701 42109 11713 42112
rect 11747 42140 11759 42143
rect 11974 42140 11980 42152
rect 11747 42112 11980 42140
rect 11747 42109 11759 42112
rect 11701 42103 11759 42109
rect 11974 42100 11980 42112
rect 12032 42100 12038 42152
rect 12176 42072 12204 42168
rect 13449 42143 13507 42149
rect 13449 42109 13461 42143
rect 13495 42140 13507 42143
rect 13538 42140 13544 42152
rect 13495 42112 13544 42140
rect 13495 42109 13507 42112
rect 13449 42103 13507 42109
rect 13538 42100 13544 42112
rect 13596 42100 13602 42152
rect 13648 42149 13676 42180
rect 16868 42180 17316 42208
rect 13633 42143 13691 42149
rect 13633 42109 13645 42143
rect 13679 42109 13691 42143
rect 13633 42103 13691 42109
rect 13814 42100 13820 42152
rect 13872 42140 13878 42152
rect 14093 42143 14151 42149
rect 14093 42140 14105 42143
rect 13872 42112 14105 42140
rect 13872 42100 13878 42112
rect 14093 42109 14105 42112
rect 14139 42109 14151 42143
rect 15838 42140 15844 42152
rect 15799 42112 15844 42140
rect 14093 42103 14151 42109
rect 15838 42100 15844 42112
rect 15896 42140 15902 42152
rect 16390 42140 16396 42152
rect 15896 42112 16396 42140
rect 15896 42100 15902 42112
rect 16390 42100 16396 42112
rect 16448 42100 16454 42152
rect 16868 42149 16896 42180
rect 17310 42168 17316 42180
rect 17368 42208 17374 42220
rect 17589 42211 17647 42217
rect 17589 42208 17601 42211
rect 17368 42180 17601 42208
rect 17368 42168 17374 42180
rect 17589 42177 17601 42180
rect 17635 42177 17647 42211
rect 17589 42171 17647 42177
rect 17954 42168 17960 42220
rect 18012 42168 18018 42220
rect 16485 42143 16543 42149
rect 16485 42109 16497 42143
rect 16531 42109 16543 42143
rect 16485 42103 16543 42109
rect 16853 42143 16911 42149
rect 16853 42109 16865 42143
rect 16899 42109 16911 42143
rect 16853 42103 16911 42109
rect 11348 42044 12204 42072
rect 14369 42075 14427 42081
rect 14369 42041 14381 42075
rect 14415 42072 14427 42075
rect 15102 42072 15108 42084
rect 14415 42044 15108 42072
rect 14415 42041 14427 42044
rect 14369 42035 14427 42041
rect 15102 42032 15108 42044
rect 15160 42032 15166 42084
rect 15746 42032 15752 42084
rect 15804 42072 15810 42084
rect 16500 42072 16528 42103
rect 16942 42100 16948 42152
rect 17000 42140 17006 42152
rect 17129 42143 17187 42149
rect 17129 42140 17141 42143
rect 17000 42112 17141 42140
rect 17000 42100 17006 42112
rect 17129 42109 17141 42112
rect 17175 42109 17187 42143
rect 17129 42103 17187 42109
rect 17972 42081 18000 42168
rect 17957 42075 18015 42081
rect 17957 42072 17969 42075
rect 15804 42044 17969 42072
rect 15804 42032 15810 42044
rect 17957 42041 17969 42044
rect 18003 42041 18015 42075
rect 17957 42035 18015 42041
rect 9490 42004 9496 42016
rect 8496 41976 9496 42004
rect 9490 41964 9496 41976
rect 9548 41964 9554 42016
rect 12526 42004 12532 42016
rect 12487 41976 12532 42004
rect 12526 41964 12532 41976
rect 12584 41964 12590 42016
rect 1104 41914 18860 41936
rect 1104 41862 7648 41914
rect 7700 41862 7712 41914
rect 7764 41862 7776 41914
rect 7828 41862 7840 41914
rect 7892 41862 14315 41914
rect 14367 41862 14379 41914
rect 14431 41862 14443 41914
rect 14495 41862 14507 41914
rect 14559 41862 18860 41914
rect 1104 41840 18860 41862
rect 1670 41760 1676 41812
rect 1728 41800 1734 41812
rect 1949 41803 2007 41809
rect 1949 41800 1961 41803
rect 1728 41772 1961 41800
rect 1728 41760 1734 41772
rect 1949 41769 1961 41772
rect 1995 41769 2007 41803
rect 3418 41800 3424 41812
rect 3379 41772 3424 41800
rect 1949 41763 2007 41769
rect 3418 41760 3424 41772
rect 3476 41760 3482 41812
rect 4341 41803 4399 41809
rect 4341 41769 4353 41803
rect 4387 41800 4399 41803
rect 5166 41800 5172 41812
rect 4387 41772 5172 41800
rect 4387 41769 4399 41772
rect 4341 41763 4399 41769
rect 5166 41760 5172 41772
rect 5224 41760 5230 41812
rect 6178 41800 6184 41812
rect 5276 41772 6184 41800
rect 4154 41692 4160 41744
rect 4212 41732 4218 41744
rect 4982 41732 4988 41744
rect 4212 41704 4988 41732
rect 4212 41692 4218 41704
rect 4982 41692 4988 41704
rect 5040 41692 5046 41744
rect 5276 41732 5304 41772
rect 5736 41744 5764 41772
rect 6178 41760 6184 41772
rect 6236 41760 6242 41812
rect 7190 41760 7196 41812
rect 7248 41800 7254 41812
rect 7561 41803 7619 41809
rect 7561 41800 7573 41803
rect 7248 41772 7573 41800
rect 7248 41760 7254 41772
rect 7561 41769 7573 41772
rect 7607 41769 7619 41803
rect 8294 41800 8300 41812
rect 8255 41772 8300 41800
rect 7561 41763 7619 41769
rect 8294 41760 8300 41772
rect 8352 41760 8358 41812
rect 8478 41760 8484 41812
rect 8536 41760 8542 41812
rect 10318 41800 10324 41812
rect 10279 41772 10324 41800
rect 10318 41760 10324 41772
rect 10376 41760 10382 41812
rect 10689 41803 10747 41809
rect 10689 41769 10701 41803
rect 10735 41800 10747 41803
rect 10778 41800 10784 41812
rect 10735 41772 10784 41800
rect 10735 41769 10747 41772
rect 10689 41763 10747 41769
rect 10778 41760 10784 41772
rect 10836 41760 10842 41812
rect 13814 41760 13820 41812
rect 13872 41800 13878 41812
rect 14277 41803 14335 41809
rect 14277 41800 14289 41803
rect 13872 41772 14289 41800
rect 13872 41760 13878 41772
rect 14277 41769 14289 41772
rect 14323 41769 14335 41803
rect 14277 41763 14335 41769
rect 15105 41803 15163 41809
rect 15105 41769 15117 41803
rect 15151 41800 15163 41803
rect 15562 41800 15568 41812
rect 15151 41772 15568 41800
rect 15151 41769 15163 41772
rect 15105 41763 15163 41769
rect 5092 41704 5304 41732
rect 4709 41599 4767 41605
rect 4709 41565 4721 41599
rect 4755 41596 4767 41599
rect 4985 41599 5043 41605
rect 4985 41596 4997 41599
rect 4755 41568 4997 41596
rect 4755 41565 4767 41568
rect 4709 41559 4767 41565
rect 4985 41565 4997 41568
rect 5031 41596 5043 41599
rect 5092 41596 5120 41704
rect 5718 41692 5724 41744
rect 5776 41692 5782 41744
rect 5905 41735 5963 41741
rect 5905 41701 5917 41735
rect 5951 41732 5963 41735
rect 7006 41732 7012 41744
rect 5951 41704 7012 41732
rect 5951 41701 5963 41704
rect 5905 41695 5963 41701
rect 7006 41692 7012 41704
rect 7064 41692 7070 41744
rect 8021 41735 8079 41741
rect 8021 41701 8033 41735
rect 8067 41732 8079 41735
rect 8496 41732 8524 41760
rect 14734 41732 14740 41744
rect 8067 41704 8524 41732
rect 11440 41704 14740 41732
rect 8067 41701 8079 41704
rect 8021 41695 8079 41701
rect 5169 41667 5227 41673
rect 5169 41633 5181 41667
rect 5215 41633 5227 41667
rect 5169 41627 5227 41633
rect 5031 41568 5120 41596
rect 5184 41596 5212 41627
rect 5258 41624 5264 41676
rect 5316 41664 5322 41676
rect 5629 41667 5687 41673
rect 5629 41664 5641 41667
rect 5316 41636 5641 41664
rect 5316 41624 5322 41636
rect 5629 41633 5641 41636
rect 5675 41664 5687 41667
rect 5994 41664 6000 41676
rect 5675 41636 6000 41664
rect 5675 41633 5687 41636
rect 5629 41627 5687 41633
rect 5994 41624 6000 41636
rect 6052 41624 6058 41676
rect 7098 41624 7104 41676
rect 7156 41664 7162 41676
rect 7285 41667 7343 41673
rect 7285 41664 7297 41667
rect 7156 41636 7297 41664
rect 7156 41624 7162 41636
rect 7285 41633 7297 41636
rect 7331 41664 7343 41667
rect 8110 41664 8116 41676
rect 7331 41636 8116 41664
rect 7331 41633 7343 41636
rect 7285 41627 7343 41633
rect 8110 41624 8116 41636
rect 8168 41664 8174 41676
rect 8481 41667 8539 41673
rect 8481 41664 8493 41667
rect 8168 41636 8493 41664
rect 8168 41624 8174 41636
rect 8481 41633 8493 41636
rect 8527 41633 8539 41667
rect 9125 41667 9183 41673
rect 9125 41664 9137 41667
rect 8481 41627 8539 41633
rect 8956 41636 9137 41664
rect 8956 41608 8984 41636
rect 9125 41633 9137 41636
rect 9171 41664 9183 41667
rect 9214 41664 9220 41676
rect 9171 41636 9220 41664
rect 9171 41633 9183 41636
rect 9125 41627 9183 41633
rect 9214 41624 9220 41636
rect 9272 41624 9278 41676
rect 9490 41664 9496 41676
rect 9451 41636 9496 41664
rect 9490 41624 9496 41636
rect 9548 41624 9554 41676
rect 9674 41624 9680 41676
rect 9732 41664 9738 41676
rect 11440 41673 11468 41704
rect 14734 41692 14740 41704
rect 14792 41692 14798 41744
rect 9769 41667 9827 41673
rect 9769 41664 9781 41667
rect 9732 41636 9781 41664
rect 9732 41624 9738 41636
rect 9769 41633 9781 41636
rect 9815 41633 9827 41667
rect 9769 41627 9827 41633
rect 11425 41667 11483 41673
rect 11425 41633 11437 41667
rect 11471 41633 11483 41667
rect 11425 41627 11483 41633
rect 11514 41624 11520 41676
rect 11572 41664 11578 41676
rect 11572 41636 11617 41664
rect 11572 41624 11578 41636
rect 11974 41624 11980 41676
rect 12032 41664 12038 41676
rect 12437 41667 12495 41673
rect 12437 41664 12449 41667
rect 12032 41636 12449 41664
rect 12032 41624 12038 41636
rect 12437 41633 12449 41636
rect 12483 41633 12495 41667
rect 12986 41664 12992 41676
rect 12947 41636 12992 41664
rect 12437 41627 12495 41633
rect 12986 41624 12992 41636
rect 13044 41624 13050 41676
rect 13449 41667 13507 41673
rect 13449 41633 13461 41667
rect 13495 41664 13507 41667
rect 13722 41664 13728 41676
rect 13495 41636 13728 41664
rect 13495 41633 13507 41636
rect 13449 41627 13507 41633
rect 13722 41624 13728 41636
rect 13780 41624 13786 41676
rect 15304 41673 15332 41772
rect 15562 41760 15568 41772
rect 15620 41800 15626 41812
rect 15838 41800 15844 41812
rect 15620 41772 15844 41800
rect 15620 41760 15626 41772
rect 15838 41760 15844 41772
rect 15896 41760 15902 41812
rect 16942 41800 16948 41812
rect 16903 41772 16948 41800
rect 16942 41760 16948 41772
rect 17000 41760 17006 41812
rect 15746 41692 15752 41744
rect 15804 41732 15810 41744
rect 17313 41735 17371 41741
rect 17313 41732 17325 41735
rect 15804 41704 17325 41732
rect 15804 41692 15810 41704
rect 17313 41701 17325 41704
rect 17359 41701 17371 41735
rect 17313 41695 17371 41701
rect 15289 41667 15347 41673
rect 15289 41633 15301 41667
rect 15335 41633 15347 41667
rect 15289 41627 15347 41633
rect 15378 41624 15384 41676
rect 15436 41664 15442 41676
rect 15565 41667 15623 41673
rect 15565 41664 15577 41667
rect 15436 41636 15577 41664
rect 15436 41624 15442 41636
rect 15565 41633 15577 41636
rect 15611 41633 15623 41667
rect 15930 41664 15936 41676
rect 15891 41636 15936 41664
rect 15565 41627 15623 41633
rect 15930 41624 15936 41636
rect 15988 41624 15994 41676
rect 16390 41624 16396 41676
rect 16448 41624 16454 41676
rect 16669 41667 16727 41673
rect 16669 41633 16681 41667
rect 16715 41664 16727 41667
rect 16758 41664 16764 41676
rect 16715 41636 16764 41664
rect 16715 41633 16727 41636
rect 16669 41627 16727 41633
rect 16758 41624 16764 41636
rect 16816 41624 16822 41676
rect 6178 41596 6184 41608
rect 5184 41568 6184 41596
rect 5031 41565 5043 41568
rect 4985 41559 5043 41565
rect 6178 41556 6184 41568
rect 6236 41556 6242 41608
rect 8938 41556 8944 41608
rect 8996 41556 9002 41608
rect 9030 41556 9036 41608
rect 9088 41596 9094 41608
rect 9508 41596 9536 41624
rect 9088 41568 9536 41596
rect 9088 41556 9094 41568
rect 12158 41556 12164 41608
rect 12216 41596 12222 41608
rect 12526 41596 12532 41608
rect 12216 41568 12532 41596
rect 12216 41556 12222 41568
rect 12526 41556 12532 41568
rect 12584 41556 12590 41608
rect 13170 41556 13176 41608
rect 13228 41596 13234 41608
rect 14645 41599 14703 41605
rect 14645 41596 14657 41599
rect 13228 41568 14657 41596
rect 13228 41556 13234 41568
rect 14645 41565 14657 41568
rect 14691 41565 14703 41599
rect 15746 41596 15752 41608
rect 15707 41568 15752 41596
rect 14645 41559 14703 41565
rect 15746 41556 15752 41568
rect 15804 41556 15810 41608
rect 5626 41488 5632 41540
rect 5684 41528 5690 41540
rect 5994 41528 6000 41540
rect 5684 41500 6000 41528
rect 5684 41488 5690 41500
rect 5994 41488 6000 41500
rect 6052 41488 6058 41540
rect 15930 41488 15936 41540
rect 15988 41528 15994 41540
rect 16408 41528 16436 41624
rect 15988 41500 16436 41528
rect 15988 41488 15994 41500
rect 17494 41488 17500 41540
rect 17552 41528 17558 41540
rect 18322 41528 18328 41540
rect 17552 41500 18328 41528
rect 17552 41488 17558 41500
rect 18322 41488 18328 41500
rect 18380 41488 18386 41540
rect 1578 41460 1584 41472
rect 1539 41432 1584 41460
rect 1578 41420 1584 41432
rect 1636 41420 1642 41472
rect 6641 41463 6699 41469
rect 6641 41429 6653 41463
rect 6687 41460 6699 41463
rect 6822 41460 6828 41472
rect 6687 41432 6828 41460
rect 6687 41429 6699 41432
rect 6641 41423 6699 41429
rect 6822 41420 6828 41432
rect 6880 41420 6886 41472
rect 8478 41420 8484 41472
rect 8536 41460 8542 41472
rect 8573 41463 8631 41469
rect 8573 41460 8585 41463
rect 8536 41432 8585 41460
rect 8536 41420 8542 41432
rect 8573 41429 8585 41432
rect 8619 41429 8631 41463
rect 8573 41423 8631 41429
rect 12069 41463 12127 41469
rect 12069 41429 12081 41463
rect 12115 41460 12127 41463
rect 12710 41460 12716 41472
rect 12115 41432 12716 41460
rect 12115 41429 12127 41432
rect 12069 41423 12127 41429
rect 12710 41420 12716 41432
rect 12768 41420 12774 41472
rect 13538 41420 13544 41472
rect 13596 41460 13602 41472
rect 13998 41460 14004 41472
rect 13596 41432 14004 41460
rect 13596 41420 13602 41432
rect 13998 41420 14004 41432
rect 14056 41420 14062 41472
rect 1104 41370 18860 41392
rect 1104 41318 4315 41370
rect 4367 41318 4379 41370
rect 4431 41318 4443 41370
rect 4495 41318 4507 41370
rect 4559 41318 10982 41370
rect 11034 41318 11046 41370
rect 11098 41318 11110 41370
rect 11162 41318 11174 41370
rect 11226 41318 17648 41370
rect 17700 41318 17712 41370
rect 17764 41318 17776 41370
rect 17828 41318 17840 41370
rect 17892 41318 18860 41370
rect 1104 41296 18860 41318
rect 1762 41216 1768 41268
rect 1820 41256 1826 41268
rect 2498 41256 2504 41268
rect 1820 41228 2504 41256
rect 1820 41216 1826 41228
rect 2498 41216 2504 41228
rect 2556 41216 2562 41268
rect 3053 41259 3111 41265
rect 3053 41225 3065 41259
rect 3099 41256 3111 41259
rect 3234 41256 3240 41268
rect 3099 41228 3240 41256
rect 3099 41225 3111 41228
rect 3053 41219 3111 41225
rect 3234 41216 3240 41228
rect 3292 41216 3298 41268
rect 4617 41259 4675 41265
rect 4617 41225 4629 41259
rect 4663 41256 4675 41259
rect 6178 41256 6184 41268
rect 4663 41228 6184 41256
rect 4663 41225 4675 41228
rect 4617 41219 4675 41225
rect 1489 41123 1547 41129
rect 1489 41089 1501 41123
rect 1535 41120 1547 41123
rect 1670 41120 1676 41132
rect 1535 41092 1676 41120
rect 1535 41089 1547 41092
rect 1489 41083 1547 41089
rect 1670 41080 1676 41092
rect 1728 41080 1734 41132
rect 4908 41129 4936 41228
rect 6178 41216 6184 41228
rect 6236 41256 6242 41268
rect 7006 41256 7012 41268
rect 6236 41228 7012 41256
rect 6236 41216 6242 41228
rect 7006 41216 7012 41228
rect 7064 41216 7070 41268
rect 8757 41259 8815 41265
rect 8757 41225 8769 41259
rect 8803 41256 8815 41259
rect 9214 41256 9220 41268
rect 8803 41228 9220 41256
rect 8803 41225 8815 41228
rect 8757 41219 8815 41225
rect 9214 41216 9220 41228
rect 9272 41216 9278 41268
rect 11882 41256 11888 41268
rect 11532 41228 11888 41256
rect 5534 41188 5540 41200
rect 5495 41160 5540 41188
rect 5534 41148 5540 41160
rect 5592 41148 5598 41200
rect 6822 41188 6828 41200
rect 6656 41160 6828 41188
rect 4893 41123 4951 41129
rect 4893 41089 4905 41123
rect 4939 41089 4951 41123
rect 4893 41083 4951 41089
rect 1578 41012 1584 41064
rect 1636 41052 1642 41064
rect 1765 41055 1823 41061
rect 1765 41052 1777 41055
rect 1636 41024 1777 41052
rect 1636 41012 1642 41024
rect 1765 41021 1777 41024
rect 1811 41021 1823 41055
rect 1765 41015 1823 41021
rect 3881 41055 3939 41061
rect 3881 41021 3893 41055
rect 3927 41052 3939 41055
rect 4614 41052 4620 41064
rect 3927 41024 4620 41052
rect 3927 41021 3939 41024
rect 3881 41015 3939 41021
rect 4614 41012 4620 41024
rect 4672 41052 4678 41064
rect 5074 41052 5080 41064
rect 4672 41024 5080 41052
rect 4672 41012 4678 41024
rect 5074 41012 5080 41024
rect 5132 41012 5138 41064
rect 5626 41052 5632 41064
rect 5587 41024 5632 41052
rect 5626 41012 5632 41024
rect 5684 41012 5690 41064
rect 6178 41012 6184 41064
rect 6236 41052 6242 41064
rect 6656 41061 6684 41160
rect 6822 41148 6828 41160
rect 6880 41148 6886 41200
rect 7466 41188 7472 41200
rect 7427 41160 7472 41188
rect 7466 41148 7472 41160
rect 7524 41148 7530 41200
rect 8570 41148 8576 41200
rect 8628 41148 8634 41200
rect 8938 41148 8944 41200
rect 8996 41188 9002 41200
rect 9033 41191 9091 41197
rect 9033 41188 9045 41191
rect 8996 41160 9045 41188
rect 8996 41148 9002 41160
rect 9033 41157 9045 41160
rect 9079 41188 9091 41191
rect 9401 41191 9459 41197
rect 9401 41188 9413 41191
rect 9079 41160 9413 41188
rect 9079 41157 9091 41160
rect 9033 41151 9091 41157
rect 9401 41157 9413 41160
rect 9447 41157 9459 41191
rect 9401 41151 9459 41157
rect 8588 41120 8616 41148
rect 9214 41120 9220 41132
rect 8588 41092 9220 41120
rect 9214 41080 9220 41092
rect 9272 41080 9278 41132
rect 6641 41055 6699 41061
rect 6641 41052 6653 41055
rect 6236 41024 6653 41052
rect 6236 41012 6242 41024
rect 6641 41021 6653 41024
rect 6687 41021 6699 41055
rect 6641 41015 6699 41021
rect 6914 41012 6920 41064
rect 6972 41052 6978 41064
rect 7009 41055 7067 41061
rect 7009 41052 7021 41055
rect 6972 41024 7021 41052
rect 6972 41012 6978 41024
rect 7009 41021 7021 41024
rect 7055 41021 7067 41055
rect 7009 41015 7067 41021
rect 7469 41055 7527 41061
rect 7469 41021 7481 41055
rect 7515 41021 7527 41055
rect 7469 41015 7527 41021
rect 7484 40984 7512 41015
rect 8294 41012 8300 41064
rect 8352 41052 8358 41064
rect 8573 41055 8631 41061
rect 8573 41052 8585 41055
rect 8352 41024 8585 41052
rect 8352 41012 8358 41024
rect 8573 41021 8585 41024
rect 8619 41021 8631 41055
rect 8573 41015 8631 41021
rect 8754 41012 8760 41064
rect 8812 41052 8818 41064
rect 8938 41052 8944 41064
rect 8812 41024 8944 41052
rect 8812 41012 8818 41024
rect 8938 41012 8944 41024
rect 8996 41012 9002 41064
rect 9416 41052 9444 41151
rect 9674 41148 9680 41200
rect 9732 41188 9738 41200
rect 9769 41191 9827 41197
rect 9769 41188 9781 41191
rect 9732 41160 9781 41188
rect 9732 41148 9738 41160
rect 9769 41157 9781 41160
rect 9815 41157 9827 41191
rect 9769 41151 9827 41157
rect 10226 41080 10232 41132
rect 10284 41120 10290 41132
rect 10284 41092 11376 41120
rect 10284 41080 10290 41092
rect 9677 41055 9735 41061
rect 9677 41052 9689 41055
rect 9416 41024 9689 41052
rect 9677 41021 9689 41024
rect 9723 41021 9735 41055
rect 10045 41055 10103 41061
rect 10045 41052 10057 41055
rect 9677 41015 9735 41021
rect 9784 41024 10057 41052
rect 7024 40956 7512 40984
rect 7024 40928 7052 40956
rect 6549 40919 6607 40925
rect 6549 40885 6561 40919
rect 6595 40916 6607 40919
rect 7006 40916 7012 40928
rect 6595 40888 7012 40916
rect 6595 40885 6607 40888
rect 6549 40879 6607 40885
rect 7006 40876 7012 40888
rect 7064 40876 7070 40928
rect 8110 40916 8116 40928
rect 8071 40888 8116 40916
rect 8110 40876 8116 40888
rect 8168 40876 8174 40928
rect 8481 40919 8539 40925
rect 8481 40885 8493 40919
rect 8527 40916 8539 40919
rect 8570 40916 8576 40928
rect 8527 40888 8576 40916
rect 8527 40885 8539 40888
rect 8481 40879 8539 40885
rect 8570 40876 8576 40888
rect 8628 40876 8634 40928
rect 9784 40916 9812 41024
rect 10045 41021 10057 41024
rect 10091 41021 10103 41055
rect 10045 41015 10103 41021
rect 10318 41012 10324 41064
rect 10376 41052 10382 41064
rect 10413 41055 10471 41061
rect 10413 41052 10425 41055
rect 10376 41024 10425 41052
rect 10376 41012 10382 41024
rect 10413 41021 10425 41024
rect 10459 41021 10471 41055
rect 10413 41015 10471 41021
rect 10965 41055 11023 41061
rect 10965 41021 10977 41055
rect 11011 41021 11023 41055
rect 11348 41052 11376 41092
rect 11422 41080 11428 41132
rect 11480 41120 11486 41132
rect 11532 41120 11560 41228
rect 11882 41216 11888 41228
rect 11940 41216 11946 41268
rect 12250 41216 12256 41268
rect 12308 41216 12314 41268
rect 14737 41259 14795 41265
rect 14737 41225 14749 41259
rect 14783 41256 14795 41259
rect 15378 41256 15384 41268
rect 14783 41228 15384 41256
rect 14783 41225 14795 41228
rect 14737 41219 14795 41225
rect 15378 41216 15384 41228
rect 15436 41216 15442 41268
rect 16390 41216 16396 41268
rect 16448 41256 16454 41268
rect 16942 41256 16948 41268
rect 16448 41228 16948 41256
rect 16448 41216 16454 41228
rect 16942 41216 16948 41228
rect 17000 41216 17006 41268
rect 17954 41256 17960 41268
rect 17915 41228 17960 41256
rect 17954 41216 17960 41228
rect 18012 41216 18018 41268
rect 12268 41188 12296 41216
rect 11716 41160 12296 41188
rect 11480 41092 11560 41120
rect 11480 41080 11486 41092
rect 11606 41080 11612 41132
rect 11664 41120 11670 41132
rect 11716 41120 11744 41160
rect 13998 41148 14004 41200
rect 14056 41188 14062 41200
rect 15654 41188 15660 41200
rect 14056 41160 15660 41188
rect 14056 41148 14062 41160
rect 15654 41148 15660 41160
rect 15712 41148 15718 41200
rect 16850 41188 16856 41200
rect 16408 41160 16856 41188
rect 16408 41132 16436 41160
rect 16850 41148 16856 41160
rect 16908 41148 16914 41200
rect 17402 41148 17408 41200
rect 17460 41188 17466 41200
rect 18322 41188 18328 41200
rect 17460 41160 18328 41188
rect 17460 41148 17466 41160
rect 18322 41148 18328 41160
rect 18380 41148 18386 41200
rect 11974 41120 11980 41132
rect 11664 41092 11744 41120
rect 11808 41092 11980 41120
rect 11664 41080 11670 41092
rect 11808 41061 11836 41092
rect 11974 41080 11980 41092
rect 12032 41080 12038 41132
rect 12618 41120 12624 41132
rect 12579 41092 12624 41120
rect 12618 41080 12624 41092
rect 12676 41080 12682 41132
rect 13814 41120 13820 41132
rect 13775 41092 13820 41120
rect 13814 41080 13820 41092
rect 13872 41080 13878 41132
rect 14550 41080 14556 41132
rect 14608 41120 14614 41132
rect 15470 41120 15476 41132
rect 14608 41092 15476 41120
rect 14608 41080 14614 41092
rect 15470 41080 15476 41092
rect 15528 41120 15534 41132
rect 15528 41092 16252 41120
rect 15528 41080 15534 41092
rect 11793 41055 11851 41061
rect 11793 41052 11805 41055
rect 11348 41024 11805 41052
rect 10965 41015 11023 41021
rect 11793 41021 11805 41024
rect 11839 41021 11851 41055
rect 12158 41052 12164 41064
rect 12119 41024 12164 41052
rect 11793 41015 11851 41021
rect 9858 40944 9864 40996
rect 9916 40984 9922 40996
rect 10870 40984 10876 40996
rect 9916 40956 10876 40984
rect 9916 40944 9922 40956
rect 10870 40944 10876 40956
rect 10928 40984 10934 40996
rect 10980 40984 11008 41015
rect 12158 41012 12164 41024
rect 12216 41012 12222 41064
rect 12345 41055 12403 41061
rect 12345 41021 12357 41055
rect 12391 41021 12403 41055
rect 12345 41015 12403 41021
rect 10928 40956 11008 40984
rect 11517 40987 11575 40993
rect 10928 40944 10934 40956
rect 11517 40953 11529 40987
rect 11563 40984 11575 40987
rect 11974 40984 11980 40996
rect 11563 40956 11980 40984
rect 11563 40953 11575 40956
rect 11517 40947 11575 40953
rect 11974 40944 11980 40956
rect 12032 40984 12038 40996
rect 12360 40984 12388 41015
rect 12710 41012 12716 41064
rect 12768 41052 12774 41064
rect 12986 41052 12992 41064
rect 12768 41024 12992 41052
rect 12768 41012 12774 41024
rect 12986 41012 12992 41024
rect 13044 41012 13050 41064
rect 13265 41055 13323 41061
rect 13265 41021 13277 41055
rect 13311 41021 13323 41055
rect 13265 41015 13323 41021
rect 14185 41055 14243 41061
rect 14185 41021 14197 41055
rect 14231 41052 14243 41055
rect 14734 41052 14740 41064
rect 14231 41024 14740 41052
rect 14231 41021 14243 41024
rect 14185 41015 14243 41021
rect 12032 40956 12388 40984
rect 12032 40944 12038 40956
rect 12618 40944 12624 40996
rect 12676 40984 12682 40996
rect 13280 40984 13308 41015
rect 14734 41012 14740 41024
rect 14792 41012 14798 41064
rect 15930 41012 15936 41064
rect 15988 41052 15994 41064
rect 16224 41061 16252 41092
rect 16390 41080 16396 41132
rect 16448 41080 16454 41132
rect 16761 41123 16819 41129
rect 16761 41120 16773 41123
rect 16684 41092 16773 41120
rect 16684 41064 16712 41092
rect 16761 41089 16773 41092
rect 16807 41089 16819 41123
rect 16761 41083 16819 41089
rect 16117 41055 16175 41061
rect 16117 41052 16129 41055
rect 15988 41024 16129 41052
rect 15988 41012 15994 41024
rect 16117 41021 16129 41024
rect 16163 41021 16175 41055
rect 16117 41015 16175 41021
rect 16209 41055 16267 41061
rect 16209 41021 16221 41055
rect 16255 41021 16267 41055
rect 16209 41015 16267 41021
rect 16577 41055 16635 41061
rect 16577 41021 16589 41055
rect 16623 41021 16635 41055
rect 16577 41015 16635 41021
rect 12676 40956 13308 40984
rect 16132 40984 16160 41015
rect 16298 40984 16304 40996
rect 16132 40956 16304 40984
rect 12676 40944 12682 40956
rect 16298 40944 16304 40956
rect 16356 40944 16362 40996
rect 10318 40916 10324 40928
rect 9784 40888 10324 40916
rect 10318 40876 10324 40888
rect 10376 40876 10382 40928
rect 14826 40876 14832 40928
rect 14884 40916 14890 40928
rect 15010 40916 15016 40928
rect 14884 40888 15016 40916
rect 14884 40876 14890 40888
rect 15010 40876 15016 40888
rect 15068 40876 15074 40928
rect 15470 40916 15476 40928
rect 15431 40888 15476 40916
rect 15470 40876 15476 40888
rect 15528 40876 15534 40928
rect 15654 40876 15660 40928
rect 15712 40916 15718 40928
rect 16592 40916 16620 41015
rect 16666 41012 16672 41064
rect 16724 41012 16730 41064
rect 17313 41055 17371 41061
rect 17313 41021 17325 41055
rect 17359 41052 17371 41055
rect 17586 41052 17592 41064
rect 17359 41024 17592 41052
rect 17359 41021 17371 41024
rect 17313 41015 17371 41021
rect 17586 41012 17592 41024
rect 17644 41012 17650 41064
rect 17310 40916 17316 40928
rect 15712 40888 17316 40916
rect 15712 40876 15718 40888
rect 17310 40876 17316 40888
rect 17368 40916 17374 40928
rect 17589 40919 17647 40925
rect 17589 40916 17601 40919
rect 17368 40888 17601 40916
rect 17368 40876 17374 40888
rect 17589 40885 17601 40888
rect 17635 40885 17647 40919
rect 17589 40879 17647 40885
rect 1104 40826 18860 40848
rect 1104 40774 7648 40826
rect 7700 40774 7712 40826
rect 7764 40774 7776 40826
rect 7828 40774 7840 40826
rect 7892 40774 14315 40826
rect 14367 40774 14379 40826
rect 14431 40774 14443 40826
rect 14495 40774 14507 40826
rect 14559 40774 18860 40826
rect 1104 40752 18860 40774
rect 4982 40672 4988 40724
rect 5040 40712 5046 40724
rect 5077 40715 5135 40721
rect 5077 40712 5089 40715
rect 5040 40684 5089 40712
rect 5040 40672 5046 40684
rect 5077 40681 5089 40684
rect 5123 40681 5135 40715
rect 5077 40675 5135 40681
rect 5905 40715 5963 40721
rect 5905 40681 5917 40715
rect 5951 40712 5963 40715
rect 6178 40712 6184 40724
rect 5951 40684 6184 40712
rect 5951 40681 5963 40684
rect 5905 40675 5963 40681
rect 6178 40672 6184 40684
rect 6236 40672 6242 40724
rect 6914 40672 6920 40724
rect 6972 40712 6978 40724
rect 7009 40715 7067 40721
rect 7009 40712 7021 40715
rect 6972 40684 7021 40712
rect 6972 40672 6978 40684
rect 7009 40681 7021 40684
rect 7055 40681 7067 40715
rect 7009 40675 7067 40681
rect 7466 40672 7472 40724
rect 7524 40712 7530 40724
rect 7561 40715 7619 40721
rect 7561 40712 7573 40715
rect 7524 40684 7573 40712
rect 7524 40672 7530 40684
rect 7561 40681 7573 40684
rect 7607 40681 7619 40715
rect 7561 40675 7619 40681
rect 9122 40672 9128 40724
rect 9180 40672 9186 40724
rect 11698 40712 11704 40724
rect 11532 40684 11704 40712
rect 4709 40647 4767 40653
rect 4709 40613 4721 40647
rect 4755 40644 4767 40647
rect 5258 40644 5264 40656
rect 4755 40616 5264 40644
rect 4755 40613 4767 40616
rect 4709 40607 4767 40613
rect 5258 40604 5264 40616
rect 5316 40604 5322 40656
rect 8110 40604 8116 40656
rect 8168 40644 8174 40656
rect 8297 40647 8355 40653
rect 8297 40644 8309 40647
rect 8168 40616 8309 40644
rect 8168 40604 8174 40616
rect 8297 40613 8309 40616
rect 8343 40644 8355 40647
rect 8343 40616 9076 40644
rect 8343 40613 8355 40616
rect 8297 40607 8355 40613
rect 9048 40588 9076 40616
rect 4246 40536 4252 40588
rect 4304 40576 4310 40588
rect 4893 40579 4951 40585
rect 4893 40576 4905 40579
rect 4304 40548 4905 40576
rect 4304 40536 4310 40548
rect 4893 40545 4905 40548
rect 4939 40545 4951 40579
rect 4893 40539 4951 40545
rect 6641 40579 6699 40585
rect 6641 40545 6653 40579
rect 6687 40576 6699 40579
rect 7377 40579 7435 40585
rect 7377 40576 7389 40579
rect 6687 40548 7389 40576
rect 6687 40545 6699 40548
rect 6641 40539 6699 40545
rect 7377 40545 7389 40548
rect 7423 40576 7435 40579
rect 7466 40576 7472 40588
rect 7423 40548 7472 40576
rect 7423 40545 7435 40548
rect 7377 40539 7435 40545
rect 4908 40508 4936 40539
rect 7466 40536 7472 40548
rect 7524 40536 7530 40588
rect 8665 40579 8723 40585
rect 8665 40545 8677 40579
rect 8711 40545 8723 40579
rect 9030 40576 9036 40588
rect 8991 40548 9036 40576
rect 8665 40539 8723 40545
rect 5258 40508 5264 40520
rect 4908 40480 5264 40508
rect 5258 40468 5264 40480
rect 5316 40468 5322 40520
rect 4341 40443 4399 40449
rect 4341 40409 4353 40443
rect 4387 40440 4399 40443
rect 5626 40440 5632 40452
rect 4387 40412 5632 40440
rect 4387 40409 4399 40412
rect 4341 40403 4399 40409
rect 5626 40400 5632 40412
rect 5684 40400 5690 40452
rect 6273 40443 6331 40449
rect 6273 40409 6285 40443
rect 6319 40440 6331 40443
rect 6914 40440 6920 40452
rect 6319 40412 6920 40440
rect 6319 40409 6331 40412
rect 6273 40403 6331 40409
rect 6914 40400 6920 40412
rect 6972 40400 6978 40452
rect 8680 40440 8708 40539
rect 9030 40536 9036 40548
rect 9088 40536 9094 40588
rect 9140 40576 9168 40672
rect 11532 40653 11560 40684
rect 11698 40672 11704 40684
rect 11756 40672 11762 40724
rect 16393 40715 16451 40721
rect 16393 40681 16405 40715
rect 16439 40712 16451 40715
rect 16758 40712 16764 40724
rect 16439 40684 16764 40712
rect 16439 40681 16451 40684
rect 16393 40675 16451 40681
rect 16758 40672 16764 40684
rect 16816 40712 16822 40724
rect 17586 40712 17592 40724
rect 16816 40684 17592 40712
rect 16816 40672 16822 40684
rect 17586 40672 17592 40684
rect 17644 40672 17650 40724
rect 11517 40647 11575 40653
rect 11517 40613 11529 40647
rect 11563 40613 11575 40647
rect 13541 40647 13599 40653
rect 13541 40644 13553 40647
rect 11517 40607 11575 40613
rect 12820 40616 13553 40644
rect 9217 40579 9275 40585
rect 9217 40576 9229 40579
rect 9140 40548 9229 40576
rect 9217 40545 9229 40548
rect 9263 40545 9275 40579
rect 9217 40539 9275 40545
rect 8846 40508 8852 40520
rect 8807 40480 8852 40508
rect 8846 40468 8852 40480
rect 8904 40468 8910 40520
rect 9232 40452 9260 40539
rect 9582 40536 9588 40588
rect 9640 40576 9646 40588
rect 9677 40579 9735 40585
rect 9677 40576 9689 40579
rect 9640 40548 9689 40576
rect 9640 40536 9646 40548
rect 9677 40545 9689 40548
rect 9723 40545 9735 40579
rect 9677 40539 9735 40545
rect 10318 40536 10324 40588
rect 10376 40576 10382 40588
rect 10505 40579 10563 40585
rect 10505 40576 10517 40579
rect 10376 40548 10517 40576
rect 10376 40536 10382 40548
rect 10505 40545 10517 40548
rect 10551 40545 10563 40579
rect 10778 40576 10784 40588
rect 10739 40548 10784 40576
rect 10505 40539 10563 40545
rect 10778 40536 10784 40548
rect 10836 40536 10842 40588
rect 10870 40536 10876 40588
rect 10928 40576 10934 40588
rect 11057 40579 11115 40585
rect 10928 40548 10973 40576
rect 10928 40536 10934 40548
rect 11057 40545 11069 40579
rect 11103 40576 11115 40579
rect 12158 40576 12164 40588
rect 11103 40548 12164 40576
rect 11103 40545 11115 40548
rect 11057 40539 11115 40545
rect 12158 40536 12164 40548
rect 12216 40536 12222 40588
rect 12434 40536 12440 40588
rect 12492 40576 12498 40588
rect 12820 40585 12848 40616
rect 13541 40613 13553 40616
rect 13587 40613 13599 40647
rect 15194 40644 15200 40656
rect 13541 40607 13599 40613
rect 13924 40616 15200 40644
rect 12805 40579 12863 40585
rect 12805 40576 12817 40579
rect 12492 40548 12817 40576
rect 12492 40536 12498 40548
rect 12805 40545 12817 40548
rect 12851 40545 12863 40579
rect 13078 40576 13084 40588
rect 13039 40548 13084 40576
rect 12805 40539 12863 40545
rect 13078 40536 13084 40548
rect 13136 40536 13142 40588
rect 13814 40536 13820 40588
rect 13872 40576 13878 40588
rect 13924 40585 13952 40616
rect 15194 40604 15200 40616
rect 15252 40644 15258 40656
rect 15252 40616 15424 40644
rect 15252 40604 15258 40616
rect 13909 40579 13967 40585
rect 13909 40576 13921 40579
rect 13872 40548 13921 40576
rect 13872 40536 13878 40548
rect 13909 40545 13921 40548
rect 13955 40545 13967 40579
rect 13909 40539 13967 40545
rect 14553 40579 14611 40585
rect 14553 40545 14565 40579
rect 14599 40545 14611 40579
rect 14553 40539 14611 40545
rect 13265 40511 13323 40517
rect 13265 40477 13277 40511
rect 13311 40508 13323 40511
rect 13630 40508 13636 40520
rect 13311 40480 13636 40508
rect 13311 40477 13323 40480
rect 13265 40471 13323 40477
rect 13630 40468 13636 40480
rect 13688 40508 13694 40520
rect 14093 40511 14151 40517
rect 14093 40508 14105 40511
rect 13688 40480 14105 40508
rect 13688 40468 13694 40480
rect 14093 40477 14105 40480
rect 14139 40477 14151 40511
rect 14093 40471 14151 40477
rect 9030 40440 9036 40452
rect 8680 40412 9036 40440
rect 9030 40400 9036 40412
rect 9088 40400 9094 40452
rect 9214 40400 9220 40452
rect 9272 40400 9278 40452
rect 13814 40400 13820 40452
rect 13872 40440 13878 40452
rect 14185 40443 14243 40449
rect 14185 40440 14197 40443
rect 13872 40412 14197 40440
rect 13872 40400 13878 40412
rect 14185 40409 14197 40412
rect 14231 40409 14243 40443
rect 14568 40440 14596 40539
rect 14642 40536 14648 40588
rect 14700 40576 14706 40588
rect 14918 40576 14924 40588
rect 14700 40548 14924 40576
rect 14700 40536 14706 40548
rect 14918 40536 14924 40548
rect 14976 40576 14982 40588
rect 15396 40585 15424 40616
rect 15013 40579 15071 40585
rect 15013 40576 15025 40579
rect 14976 40548 15025 40576
rect 14976 40536 14982 40548
rect 15013 40545 15025 40548
rect 15059 40545 15071 40579
rect 15013 40539 15071 40545
rect 15381 40579 15439 40585
rect 15381 40545 15393 40579
rect 15427 40545 15439 40579
rect 15838 40576 15844 40588
rect 15799 40548 15844 40576
rect 15381 40539 15439 40545
rect 15838 40536 15844 40548
rect 15896 40536 15902 40588
rect 16853 40579 16911 40585
rect 16853 40545 16865 40579
rect 16899 40576 16911 40579
rect 18138 40576 18144 40588
rect 16899 40548 18144 40576
rect 16899 40545 16911 40548
rect 16853 40539 16911 40545
rect 18138 40536 18144 40548
rect 18196 40536 18202 40588
rect 14642 40440 14648 40452
rect 14555 40412 14648 40440
rect 14185 40403 14243 40409
rect 14642 40400 14648 40412
rect 14700 40440 14706 40452
rect 15470 40440 15476 40452
rect 14700 40412 15476 40440
rect 14700 40400 14706 40412
rect 15470 40400 15476 40412
rect 15528 40440 15534 40452
rect 16850 40440 16856 40452
rect 15528 40412 16856 40440
rect 15528 40400 15534 40412
rect 16850 40400 16856 40412
rect 16908 40440 16914 40452
rect 17037 40443 17095 40449
rect 17037 40440 17049 40443
rect 16908 40412 17049 40440
rect 16908 40400 16914 40412
rect 17037 40409 17049 40412
rect 17083 40409 17095 40443
rect 17037 40403 17095 40409
rect 1578 40372 1584 40384
rect 1539 40344 1584 40372
rect 1578 40332 1584 40344
rect 1636 40332 1642 40384
rect 1670 40332 1676 40384
rect 1728 40372 1734 40384
rect 1949 40375 2007 40381
rect 1949 40372 1961 40375
rect 1728 40344 1961 40372
rect 1728 40332 1734 40344
rect 1949 40341 1961 40344
rect 1995 40341 2007 40375
rect 1949 40335 2007 40341
rect 7929 40375 7987 40381
rect 7929 40341 7941 40375
rect 7975 40372 7987 40375
rect 8294 40372 8300 40384
rect 7975 40344 8300 40372
rect 7975 40341 7987 40344
rect 7929 40335 7987 40341
rect 8294 40332 8300 40344
rect 8352 40332 8358 40384
rect 9858 40332 9864 40384
rect 9916 40372 9922 40384
rect 10137 40375 10195 40381
rect 10137 40372 10149 40375
rect 9916 40344 10149 40372
rect 9916 40332 9922 40344
rect 10137 40341 10149 40344
rect 10183 40341 10195 40375
rect 10137 40335 10195 40341
rect 12069 40375 12127 40381
rect 12069 40341 12081 40375
rect 12115 40372 12127 40375
rect 12618 40372 12624 40384
rect 12115 40344 12624 40372
rect 12115 40341 12127 40344
rect 12069 40335 12127 40341
rect 12618 40332 12624 40344
rect 12676 40332 12682 40384
rect 16298 40332 16304 40384
rect 16356 40372 16362 40384
rect 17310 40372 17316 40384
rect 16356 40344 17316 40372
rect 16356 40332 16362 40344
rect 17310 40332 17316 40344
rect 17368 40332 17374 40384
rect 1104 40282 18860 40304
rect 1104 40230 4315 40282
rect 4367 40230 4379 40282
rect 4431 40230 4443 40282
rect 4495 40230 4507 40282
rect 4559 40230 10982 40282
rect 11034 40230 11046 40282
rect 11098 40230 11110 40282
rect 11162 40230 11174 40282
rect 11226 40230 17648 40282
rect 17700 40230 17712 40282
rect 17764 40230 17776 40282
rect 17828 40230 17840 40282
rect 17892 40230 18860 40282
rect 1104 40208 18860 40230
rect 3694 40128 3700 40180
rect 3752 40168 3758 40180
rect 3789 40171 3847 40177
rect 3789 40168 3801 40171
rect 3752 40140 3801 40168
rect 3752 40128 3758 40140
rect 3789 40137 3801 40140
rect 3835 40137 3847 40171
rect 11974 40168 11980 40180
rect 11935 40140 11980 40168
rect 3789 40131 3847 40137
rect 3804 40032 3832 40131
rect 11974 40128 11980 40140
rect 12032 40128 12038 40180
rect 12158 40128 12164 40180
rect 12216 40168 12222 40180
rect 12342 40168 12348 40180
rect 12216 40140 12348 40168
rect 12216 40128 12222 40140
rect 12342 40128 12348 40140
rect 12400 40168 12406 40180
rect 13725 40171 13783 40177
rect 13725 40168 13737 40171
rect 12400 40140 13737 40168
rect 12400 40128 12406 40140
rect 13725 40137 13737 40140
rect 13771 40168 13783 40171
rect 14829 40171 14887 40177
rect 13771 40140 14228 40168
rect 13771 40137 13783 40140
rect 13725 40131 13783 40137
rect 4890 40060 4896 40112
rect 4948 40100 4954 40112
rect 4948 40072 5396 40100
rect 4948 40060 4954 40072
rect 5077 40035 5135 40041
rect 5077 40032 5089 40035
rect 3804 40004 5089 40032
rect 5077 40001 5089 40004
rect 5123 40001 5135 40035
rect 5368 40032 5396 40072
rect 7466 40060 7472 40112
rect 7524 40100 7530 40112
rect 9030 40100 9036 40112
rect 7524 40072 9036 40100
rect 7524 40060 7530 40072
rect 9030 40060 9036 40072
rect 9088 40060 9094 40112
rect 9769 40103 9827 40109
rect 9769 40100 9781 40103
rect 9324 40072 9781 40100
rect 6549 40035 6607 40041
rect 6549 40032 6561 40035
rect 5368 40004 6561 40032
rect 5077 39995 5135 40001
rect 6549 40001 6561 40004
rect 6595 40001 6607 40035
rect 6549 39995 6607 40001
rect 6914 39992 6920 40044
rect 6972 40032 6978 40044
rect 9324 40032 9352 40072
rect 9769 40069 9781 40072
rect 9815 40069 9827 40103
rect 9769 40063 9827 40069
rect 10042 40060 10048 40112
rect 10100 40100 10106 40112
rect 10226 40100 10232 40112
rect 10100 40072 10232 40100
rect 10100 40060 10106 40072
rect 10226 40060 10232 40072
rect 10284 40060 10290 40112
rect 10962 40060 10968 40112
rect 11020 40100 11026 40112
rect 14093 40103 14151 40109
rect 14093 40100 14105 40103
rect 11020 40072 14105 40100
rect 11020 40060 11026 40072
rect 14093 40069 14105 40072
rect 14139 40069 14151 40103
rect 14200 40100 14228 40140
rect 14829 40137 14841 40171
rect 14875 40168 14887 40171
rect 14918 40168 14924 40180
rect 14875 40140 14924 40168
rect 14875 40137 14887 40140
rect 14829 40131 14887 40137
rect 14918 40128 14924 40140
rect 14976 40128 14982 40180
rect 15194 40128 15200 40180
rect 15252 40168 15258 40180
rect 15473 40171 15531 40177
rect 15473 40168 15485 40171
rect 15252 40140 15485 40168
rect 15252 40128 15258 40140
rect 15473 40137 15485 40140
rect 15519 40168 15531 40171
rect 15930 40168 15936 40180
rect 15519 40140 15936 40168
rect 15519 40137 15531 40140
rect 15473 40131 15531 40137
rect 15930 40128 15936 40140
rect 15988 40128 15994 40180
rect 17218 40168 17224 40180
rect 17179 40140 17224 40168
rect 17218 40128 17224 40140
rect 17276 40128 17282 40180
rect 18138 40168 18144 40180
rect 17788 40140 18144 40168
rect 17788 40109 17816 40140
rect 18138 40128 18144 40140
rect 18196 40128 18202 40180
rect 17773 40103 17831 40109
rect 17773 40100 17785 40103
rect 14200 40072 17785 40100
rect 14093 40063 14151 40069
rect 17773 40069 17785 40072
rect 17819 40069 17831 40103
rect 17773 40063 17831 40069
rect 11422 40032 11428 40044
rect 6972 40004 9352 40032
rect 9968 40004 11428 40032
rect 6972 39992 6978 40004
rect 3513 39967 3571 39973
rect 3513 39933 3525 39967
rect 3559 39964 3571 39967
rect 4249 39967 4307 39973
rect 4249 39964 4261 39967
rect 3559 39936 4261 39964
rect 3559 39933 3571 39936
rect 3513 39927 3571 39933
rect 4249 39933 4261 39936
rect 4295 39964 4307 39967
rect 4614 39964 4620 39976
rect 4295 39936 4620 39964
rect 4295 39933 4307 39936
rect 4249 39927 4307 39933
rect 4614 39924 4620 39936
rect 4672 39924 4678 39976
rect 4801 39967 4859 39973
rect 4801 39933 4813 39967
rect 4847 39933 4859 39967
rect 5994 39964 6000 39976
rect 5907 39936 6000 39964
rect 4801 39927 4859 39933
rect 4430 39856 4436 39908
rect 4488 39896 4494 39908
rect 4816 39896 4844 39927
rect 5994 39924 6000 39936
rect 6052 39964 6058 39976
rect 6273 39967 6331 39973
rect 6273 39964 6285 39967
rect 6052 39936 6285 39964
rect 6052 39924 6058 39936
rect 6273 39933 6285 39936
rect 6319 39933 6331 39967
rect 6273 39927 6331 39933
rect 6641 39967 6699 39973
rect 6641 39933 6653 39967
rect 6687 39933 6699 39967
rect 7190 39964 7196 39976
rect 7151 39936 7196 39964
rect 6641 39927 6699 39933
rect 4890 39896 4896 39908
rect 4488 39868 4896 39896
rect 4488 39856 4494 39868
rect 4890 39856 4896 39868
rect 4948 39856 4954 39908
rect 4338 39828 4344 39840
rect 4299 39800 4344 39828
rect 4338 39788 4344 39800
rect 4396 39788 4402 39840
rect 5718 39828 5724 39840
rect 5679 39800 5724 39828
rect 5718 39788 5724 39800
rect 5776 39788 5782 39840
rect 6012 39828 6040 39924
rect 6089 39899 6147 39905
rect 6089 39865 6101 39899
rect 6135 39896 6147 39899
rect 6178 39896 6184 39908
rect 6135 39868 6184 39896
rect 6135 39865 6147 39868
rect 6089 39859 6147 39865
rect 6178 39856 6184 39868
rect 6236 39896 6242 39908
rect 6656 39896 6684 39927
rect 7190 39924 7196 39936
rect 7248 39924 7254 39976
rect 7484 39973 7512 40004
rect 9968 39973 9996 40004
rect 11422 39992 11428 40004
rect 11480 39992 11486 40044
rect 7469 39967 7527 39973
rect 7469 39933 7481 39967
rect 7515 39933 7527 39967
rect 7469 39927 7527 39933
rect 7837 39967 7895 39973
rect 7837 39933 7849 39967
rect 7883 39933 7895 39967
rect 7837 39927 7895 39933
rect 9953 39967 10011 39973
rect 9953 39933 9965 39967
rect 9999 39933 10011 39967
rect 9953 39927 10011 39933
rect 10229 39967 10287 39973
rect 10229 39933 10241 39967
rect 10275 39933 10287 39967
rect 10229 39927 10287 39933
rect 6236 39868 6684 39896
rect 6236 39856 6242 39868
rect 6914 39856 6920 39908
rect 6972 39896 6978 39908
rect 7852 39896 7880 39927
rect 9401 39899 9459 39905
rect 9401 39896 9413 39899
rect 6972 39868 7880 39896
rect 8588 39868 9413 39896
rect 6972 39856 6978 39868
rect 8588 39840 8616 39868
rect 9401 39865 9413 39868
rect 9447 39896 9459 39899
rect 9582 39896 9588 39908
rect 9447 39868 9588 39896
rect 9447 39865 9459 39868
rect 9401 39859 9459 39865
rect 9582 39856 9588 39868
rect 9640 39896 9646 39908
rect 10244 39896 10272 39927
rect 9640 39868 10272 39896
rect 9640 39856 9646 39868
rect 6638 39828 6644 39840
rect 6012 39800 6644 39828
rect 6638 39788 6644 39800
rect 6696 39788 6702 39840
rect 8481 39831 8539 39837
rect 8481 39797 8493 39831
rect 8527 39828 8539 39831
rect 8570 39828 8576 39840
rect 8527 39800 8576 39828
rect 8527 39797 8539 39800
rect 8481 39791 8539 39797
rect 8570 39788 8576 39800
rect 8628 39788 8634 39840
rect 8849 39831 8907 39837
rect 8849 39797 8861 39831
rect 8895 39828 8907 39831
rect 9214 39828 9220 39840
rect 8895 39800 9220 39828
rect 8895 39797 8907 39800
rect 8849 39791 8907 39797
rect 9214 39788 9220 39800
rect 9272 39828 9278 39840
rect 10042 39828 10048 39840
rect 9272 39800 10048 39828
rect 9272 39788 9278 39800
rect 10042 39788 10048 39800
rect 10100 39788 10106 39840
rect 10870 39828 10876 39840
rect 10831 39800 10876 39828
rect 10870 39788 10876 39800
rect 10928 39788 10934 39840
rect 11238 39828 11244 39840
rect 11199 39800 11244 39828
rect 11238 39788 11244 39800
rect 11296 39788 11302 39840
rect 11440 39828 11468 39992
rect 11698 39964 11704 39976
rect 11659 39936 11704 39964
rect 11698 39924 11704 39936
rect 11756 39924 11762 39976
rect 11882 39964 11888 39976
rect 11843 39936 11888 39964
rect 11882 39924 11888 39936
rect 11940 39924 11946 39976
rect 12526 39964 12532 39976
rect 12487 39936 12532 39964
rect 12526 39924 12532 39936
rect 12584 39924 12590 39976
rect 12621 39967 12679 39973
rect 12621 39933 12633 39967
rect 12667 39933 12679 39967
rect 12621 39927 12679 39933
rect 11716 39896 11744 39924
rect 12636 39896 12664 39927
rect 13538 39924 13544 39976
rect 13596 39964 13602 39976
rect 13909 39967 13967 39973
rect 13909 39964 13921 39967
rect 13596 39936 13921 39964
rect 13596 39924 13602 39936
rect 13909 39933 13921 39936
rect 13955 39964 13967 39967
rect 14369 39967 14427 39973
rect 14369 39964 14381 39967
rect 13955 39936 14381 39964
rect 13955 39933 13967 39936
rect 13909 39927 13967 39933
rect 14369 39933 14381 39936
rect 14415 39933 14427 39967
rect 16298 39964 16304 39976
rect 16259 39936 16304 39964
rect 14369 39927 14427 39933
rect 16298 39924 16304 39936
rect 16356 39924 16362 39976
rect 16393 39967 16451 39973
rect 16393 39933 16405 39967
rect 16439 39933 16451 39967
rect 16758 39964 16764 39976
rect 16719 39936 16764 39964
rect 16393 39927 16451 39933
rect 11716 39868 12664 39896
rect 15194 39856 15200 39908
rect 15252 39896 15258 39908
rect 15838 39896 15844 39908
rect 15252 39868 15844 39896
rect 15252 39856 15258 39868
rect 15838 39856 15844 39868
rect 15896 39896 15902 39908
rect 16408 39896 16436 39927
rect 16758 39924 16764 39936
rect 16816 39924 16822 39976
rect 16850 39924 16856 39976
rect 16908 39964 16914 39976
rect 17313 39967 17371 39973
rect 17313 39964 17325 39967
rect 16908 39936 17325 39964
rect 16908 39924 16914 39936
rect 17313 39933 17325 39936
rect 17359 39933 17371 39967
rect 17313 39927 17371 39933
rect 15896 39868 16436 39896
rect 15896 39856 15902 39868
rect 12158 39828 12164 39840
rect 11440 39800 12164 39828
rect 12158 39788 12164 39800
rect 12216 39788 12222 39840
rect 13078 39788 13084 39840
rect 13136 39828 13142 39840
rect 13262 39828 13268 39840
rect 13136 39800 13268 39828
rect 13136 39788 13142 39800
rect 13262 39788 13268 39800
rect 13320 39828 13326 39840
rect 13357 39831 13415 39837
rect 13357 39828 13369 39831
rect 13320 39800 13369 39828
rect 13320 39788 13326 39800
rect 13357 39797 13369 39800
rect 13403 39797 13415 39831
rect 13357 39791 13415 39797
rect 17126 39788 17132 39840
rect 17184 39828 17190 39840
rect 18414 39828 18420 39840
rect 17184 39800 18420 39828
rect 17184 39788 17190 39800
rect 18414 39788 18420 39800
rect 18472 39788 18478 39840
rect 1104 39738 18860 39760
rect 1104 39686 7648 39738
rect 7700 39686 7712 39738
rect 7764 39686 7776 39738
rect 7828 39686 7840 39738
rect 7892 39686 14315 39738
rect 14367 39686 14379 39738
rect 14431 39686 14443 39738
rect 14495 39686 14507 39738
rect 14559 39686 18860 39738
rect 1104 39664 18860 39686
rect 2130 39584 2136 39636
rect 2188 39624 2194 39636
rect 2314 39624 2320 39636
rect 2188 39596 2320 39624
rect 2188 39584 2194 39596
rect 2314 39584 2320 39596
rect 2372 39584 2378 39636
rect 4341 39627 4399 39633
rect 4341 39593 4353 39627
rect 4387 39624 4399 39627
rect 4430 39624 4436 39636
rect 4387 39596 4436 39624
rect 4387 39593 4399 39596
rect 4341 39587 4399 39593
rect 4430 39584 4436 39596
rect 4488 39584 4494 39636
rect 4614 39624 4620 39636
rect 4575 39596 4620 39624
rect 4614 39584 4620 39596
rect 4672 39584 4678 39636
rect 5258 39584 5264 39636
rect 5316 39624 5322 39636
rect 5537 39627 5595 39633
rect 5537 39624 5549 39627
rect 5316 39596 5549 39624
rect 5316 39584 5322 39596
rect 5537 39593 5549 39596
rect 5583 39593 5595 39627
rect 5537 39587 5595 39593
rect 6273 39627 6331 39633
rect 6273 39593 6285 39627
rect 6319 39624 6331 39627
rect 7190 39624 7196 39636
rect 6319 39596 7196 39624
rect 6319 39593 6331 39596
rect 6273 39587 6331 39593
rect 7190 39584 7196 39596
rect 7248 39584 7254 39636
rect 8297 39627 8355 39633
rect 8297 39593 8309 39627
rect 8343 39624 8355 39627
rect 9582 39624 9588 39636
rect 8343 39596 9588 39624
rect 8343 39593 8355 39596
rect 8297 39587 8355 39593
rect 9582 39584 9588 39596
rect 9640 39584 9646 39636
rect 10045 39627 10103 39633
rect 10045 39593 10057 39627
rect 10091 39593 10103 39627
rect 11882 39624 11888 39636
rect 11843 39596 11888 39624
rect 10045 39587 10103 39593
rect 2958 39516 2964 39568
rect 3016 39556 3022 39568
rect 3326 39556 3332 39568
rect 3016 39528 3332 39556
rect 3016 39516 3022 39528
rect 3326 39516 3332 39528
rect 3384 39516 3390 39568
rect 3602 39556 3608 39568
rect 3436 39528 3608 39556
rect 3234 39488 3240 39500
rect 3147 39460 3240 39488
rect 3234 39448 3240 39460
rect 3292 39488 3298 39500
rect 3436 39488 3464 39528
rect 3602 39516 3608 39528
rect 3660 39516 3666 39568
rect 7837 39559 7895 39565
rect 7837 39525 7849 39559
rect 7883 39556 7895 39559
rect 8110 39556 8116 39568
rect 7883 39528 8116 39556
rect 7883 39525 7895 39528
rect 7837 39519 7895 39525
rect 8110 39516 8116 39528
rect 8168 39516 8174 39568
rect 9398 39516 9404 39568
rect 9456 39556 9462 39568
rect 10060 39556 10088 39587
rect 11882 39584 11888 39596
rect 11940 39584 11946 39636
rect 12342 39584 12348 39636
rect 12400 39624 12406 39636
rect 14553 39627 14611 39633
rect 12400 39596 14412 39624
rect 12400 39584 12406 39596
rect 14384 39568 14412 39596
rect 14553 39593 14565 39627
rect 14599 39624 14611 39627
rect 14642 39624 14648 39636
rect 14599 39596 14648 39624
rect 14599 39593 14611 39596
rect 14553 39587 14611 39593
rect 14642 39584 14648 39596
rect 14700 39584 14706 39636
rect 17310 39624 17316 39636
rect 17271 39596 17316 39624
rect 17310 39584 17316 39596
rect 17368 39584 17374 39636
rect 12434 39556 12440 39568
rect 9456 39528 10088 39556
rect 11624 39528 12440 39556
rect 9456 39516 9462 39528
rect 3694 39488 3700 39500
rect 3292 39460 3464 39488
rect 3655 39460 3700 39488
rect 3292 39448 3298 39460
rect 3694 39448 3700 39460
rect 3752 39448 3758 39500
rect 4614 39488 4620 39500
rect 4575 39460 4620 39488
rect 4614 39448 4620 39460
rect 4672 39448 4678 39500
rect 5077 39491 5135 39497
rect 5077 39457 5089 39491
rect 5123 39488 5135 39491
rect 5350 39488 5356 39500
rect 5123 39460 5356 39488
rect 5123 39457 5135 39460
rect 5077 39451 5135 39457
rect 5350 39448 5356 39460
rect 5408 39448 5414 39500
rect 7377 39491 7435 39497
rect 7377 39457 7389 39491
rect 7423 39457 7435 39491
rect 7650 39488 7656 39500
rect 7611 39460 7656 39488
rect 7377 39451 7435 39457
rect 3326 39420 3332 39432
rect 3287 39392 3332 39420
rect 3326 39380 3332 39392
rect 3384 39380 3390 39432
rect 7392 39420 7420 39451
rect 7650 39448 7656 39460
rect 7708 39448 7714 39500
rect 8757 39491 8815 39497
rect 8757 39457 8769 39491
rect 8803 39457 8815 39491
rect 10870 39488 10876 39500
rect 10831 39460 10876 39488
rect 8757 39451 8815 39457
rect 7558 39420 7564 39432
rect 7392 39392 7564 39420
rect 7558 39380 7564 39392
rect 7616 39380 7622 39432
rect 6638 39284 6644 39296
rect 6599 39256 6644 39284
rect 6638 39244 6644 39256
rect 6696 39244 6702 39296
rect 8665 39287 8723 39293
rect 8665 39253 8677 39287
rect 8711 39284 8723 39287
rect 8772 39284 8800 39451
rect 10870 39448 10876 39460
rect 10928 39448 10934 39500
rect 11238 39448 11244 39500
rect 11296 39488 11302 39500
rect 11333 39491 11391 39497
rect 11333 39488 11345 39491
rect 11296 39460 11345 39488
rect 11296 39448 11302 39460
rect 11333 39457 11345 39460
rect 11379 39457 11391 39491
rect 11333 39451 11391 39457
rect 11624 39432 11652 39528
rect 12434 39516 12440 39528
rect 12492 39516 12498 39568
rect 14182 39556 14188 39568
rect 14143 39528 14188 39556
rect 14182 39516 14188 39528
rect 14240 39516 14246 39568
rect 14366 39516 14372 39568
rect 14424 39516 14430 39568
rect 15286 39516 15292 39568
rect 15344 39556 15350 39568
rect 15344 39528 16344 39556
rect 15344 39516 15350 39528
rect 16316 39500 16344 39528
rect 11974 39448 11980 39500
rect 12032 39488 12038 39500
rect 12805 39491 12863 39497
rect 12805 39488 12817 39491
rect 12032 39460 12817 39488
rect 12032 39448 12038 39460
rect 12805 39457 12817 39460
rect 12851 39457 12863 39491
rect 12805 39451 12863 39457
rect 13170 39448 13176 39500
rect 13228 39488 13234 39500
rect 13446 39488 13452 39500
rect 13228 39460 13452 39488
rect 13228 39448 13234 39460
rect 13446 39448 13452 39460
rect 13504 39448 13510 39500
rect 15565 39491 15623 39497
rect 15565 39488 15577 39491
rect 15304 39460 15577 39488
rect 15304 39432 15332 39460
rect 15565 39457 15577 39460
rect 15611 39488 15623 39491
rect 15654 39488 15660 39500
rect 15611 39460 15660 39488
rect 15611 39457 15623 39460
rect 15565 39451 15623 39457
rect 15654 39448 15660 39460
rect 15712 39448 15718 39500
rect 15930 39488 15936 39500
rect 15891 39460 15936 39488
rect 15930 39448 15936 39460
rect 15988 39448 15994 39500
rect 16298 39488 16304 39500
rect 16211 39460 16304 39488
rect 16298 39448 16304 39460
rect 16356 39448 16362 39500
rect 16850 39488 16856 39500
rect 16811 39460 16856 39488
rect 16850 39448 16856 39460
rect 16908 39448 16914 39500
rect 11149 39423 11207 39429
rect 11149 39389 11161 39423
rect 11195 39420 11207 39423
rect 11606 39420 11612 39432
rect 11195 39392 11612 39420
rect 11195 39389 11207 39392
rect 11149 39383 11207 39389
rect 11606 39380 11612 39392
rect 11664 39380 11670 39432
rect 12529 39423 12587 39429
rect 12529 39389 12541 39423
rect 12575 39420 12587 39423
rect 12710 39420 12716 39432
rect 12575 39392 12716 39420
rect 12575 39389 12587 39392
rect 12529 39383 12587 39389
rect 12710 39380 12716 39392
rect 12768 39420 12774 39432
rect 12894 39420 12900 39432
rect 12768 39392 12900 39420
rect 12768 39380 12774 39392
rect 12894 39380 12900 39392
rect 12952 39380 12958 39432
rect 15286 39380 15292 39432
rect 15344 39380 15350 39432
rect 15473 39423 15531 39429
rect 15473 39389 15485 39423
rect 15519 39420 15531 39423
rect 16758 39420 16764 39432
rect 15519 39392 16764 39420
rect 15519 39389 15531 39392
rect 15473 39383 15531 39389
rect 16758 39380 16764 39392
rect 16816 39380 16822 39432
rect 11238 39312 11244 39364
rect 11296 39312 11302 39364
rect 9490 39284 9496 39296
rect 8711 39256 9496 39284
rect 8711 39253 8723 39256
rect 8665 39247 8723 39253
rect 9490 39244 9496 39256
rect 9548 39244 9554 39296
rect 11256 39284 11284 39312
rect 13446 39284 13452 39296
rect 11256 39256 13452 39284
rect 13446 39244 13452 39256
rect 13504 39244 13510 39296
rect 14921 39287 14979 39293
rect 14921 39253 14933 39287
rect 14967 39284 14979 39287
rect 15194 39284 15200 39296
rect 14967 39256 15200 39284
rect 14967 39253 14979 39256
rect 14921 39247 14979 39253
rect 15194 39244 15200 39256
rect 15252 39244 15258 39296
rect 15470 39244 15476 39296
rect 15528 39284 15534 39296
rect 15657 39287 15715 39293
rect 15657 39284 15669 39287
rect 15528 39256 15669 39284
rect 15528 39244 15534 39256
rect 15657 39253 15669 39256
rect 15703 39253 15715 39287
rect 15657 39247 15715 39253
rect 1104 39194 18860 39216
rect 1104 39142 4315 39194
rect 4367 39142 4379 39194
rect 4431 39142 4443 39194
rect 4495 39142 4507 39194
rect 4559 39142 10982 39194
rect 11034 39142 11046 39194
rect 11098 39142 11110 39194
rect 11162 39142 11174 39194
rect 11226 39142 17648 39194
rect 17700 39142 17712 39194
rect 17764 39142 17776 39194
rect 17828 39142 17840 39194
rect 17892 39142 18860 39194
rect 1104 39120 18860 39142
rect 2682 39080 2688 39092
rect 2643 39052 2688 39080
rect 2682 39040 2688 39052
rect 2740 39040 2746 39092
rect 3053 39083 3111 39089
rect 3053 39049 3065 39083
rect 3099 39080 3111 39083
rect 3234 39080 3240 39092
rect 3099 39052 3240 39080
rect 3099 39049 3111 39052
rect 3053 39043 3111 39049
rect 3234 39040 3240 39052
rect 3292 39040 3298 39092
rect 3326 39040 3332 39092
rect 3384 39080 3390 39092
rect 3421 39083 3479 39089
rect 3421 39080 3433 39083
rect 3384 39052 3433 39080
rect 3384 39040 3390 39052
rect 3421 39049 3433 39052
rect 3467 39049 3479 39083
rect 3786 39080 3792 39092
rect 3747 39052 3792 39080
rect 3421 39043 3479 39049
rect 3436 38944 3464 39043
rect 3786 39040 3792 39052
rect 3844 39040 3850 39092
rect 5350 39040 5356 39092
rect 5408 39080 5414 39092
rect 5445 39083 5503 39089
rect 5445 39080 5457 39083
rect 5408 39052 5457 39080
rect 5408 39040 5414 39052
rect 5445 39049 5457 39052
rect 5491 39049 5503 39083
rect 5445 39043 5503 39049
rect 5718 39040 5724 39092
rect 5776 39080 5782 39092
rect 6914 39080 6920 39092
rect 5776 39052 6920 39080
rect 5776 39040 5782 39052
rect 6914 39040 6920 39052
rect 6972 39040 6978 39092
rect 8386 39080 8392 39092
rect 7208 39052 7604 39080
rect 8347 39052 8392 39080
rect 5626 38972 5632 39024
rect 5684 39012 5690 39024
rect 6273 39015 6331 39021
rect 6273 39012 6285 39015
rect 5684 38984 6285 39012
rect 5684 38972 5690 38984
rect 6273 38981 6285 38984
rect 6319 39012 6331 39015
rect 7208 39012 7236 39052
rect 6319 38984 7236 39012
rect 6319 38981 6331 38984
rect 6273 38975 6331 38981
rect 4157 38947 4215 38953
rect 4157 38944 4169 38947
rect 3436 38916 4169 38944
rect 4157 38913 4169 38916
rect 4203 38913 4215 38947
rect 4157 38907 4215 38913
rect 4249 38947 4307 38953
rect 4249 38913 4261 38947
rect 4295 38944 4307 38947
rect 4706 38944 4712 38956
rect 4295 38916 4712 38944
rect 4295 38913 4307 38916
rect 4249 38907 4307 38913
rect 4706 38904 4712 38916
rect 4764 38904 4770 38956
rect 3326 38836 3332 38888
rect 3384 38876 3390 38888
rect 3786 38876 3792 38888
rect 3384 38848 3792 38876
rect 3384 38836 3390 38848
rect 3786 38836 3792 38848
rect 3844 38876 3850 38888
rect 4985 38879 5043 38885
rect 4985 38876 4997 38879
rect 3844 38848 4997 38876
rect 3844 38836 3850 38848
rect 4985 38845 4997 38848
rect 5031 38845 5043 38879
rect 4985 38839 5043 38845
rect 5074 38836 5080 38888
rect 5132 38876 5138 38888
rect 5132 38848 5177 38876
rect 5132 38836 5138 38848
rect 6178 38836 6184 38888
rect 6236 38876 6242 38888
rect 6825 38879 6883 38885
rect 6825 38876 6837 38879
rect 6236 38848 6837 38876
rect 6236 38836 6242 38848
rect 6825 38845 6837 38848
rect 6871 38845 6883 38879
rect 7466 38876 7472 38888
rect 7427 38848 7472 38876
rect 6825 38839 6883 38845
rect 7466 38836 7472 38848
rect 7524 38836 7530 38888
rect 7576 38885 7604 39052
rect 8386 39040 8392 39052
rect 8444 39040 8450 39092
rect 10318 39040 10324 39092
rect 10376 39080 10382 39092
rect 10376 39052 10824 39080
rect 10376 39040 10382 39052
rect 10226 38972 10232 39024
rect 10284 39012 10290 39024
rect 10284 38984 10732 39012
rect 10284 38972 10290 38984
rect 10594 38944 10600 38956
rect 10555 38916 10600 38944
rect 10594 38904 10600 38916
rect 10652 38904 10658 38956
rect 7561 38879 7619 38885
rect 7561 38845 7573 38879
rect 7607 38845 7619 38879
rect 8478 38876 8484 38888
rect 8439 38848 8484 38876
rect 7561 38839 7619 38845
rect 8478 38836 8484 38848
rect 8536 38836 8542 38888
rect 8846 38876 8852 38888
rect 8807 38848 8852 38876
rect 8846 38836 8852 38848
rect 8904 38836 8910 38888
rect 9309 38879 9367 38885
rect 9309 38845 9321 38879
rect 9355 38876 9367 38879
rect 9582 38876 9588 38888
rect 9355 38848 9588 38876
rect 9355 38845 9367 38848
rect 9309 38839 9367 38845
rect 9582 38836 9588 38848
rect 9640 38836 9646 38888
rect 9950 38836 9956 38888
rect 10008 38876 10014 38888
rect 10045 38879 10103 38885
rect 10045 38876 10057 38879
rect 10008 38848 10057 38876
rect 10008 38836 10014 38848
rect 10045 38845 10057 38848
rect 10091 38876 10103 38879
rect 10226 38876 10232 38888
rect 10091 38848 10232 38876
rect 10091 38845 10103 38848
rect 10045 38839 10103 38845
rect 10226 38836 10232 38848
rect 10284 38836 10290 38888
rect 10410 38876 10416 38888
rect 10371 38848 10416 38876
rect 10410 38836 10416 38848
rect 10468 38836 10474 38888
rect 2317 38811 2375 38817
rect 2317 38777 2329 38811
rect 2363 38808 2375 38811
rect 3694 38808 3700 38820
rect 2363 38780 3700 38808
rect 2363 38777 2375 38780
rect 2317 38771 2375 38777
rect 3694 38768 3700 38780
rect 3752 38768 3758 38820
rect 5997 38811 6055 38817
rect 5997 38777 6009 38811
rect 6043 38808 6055 38811
rect 6730 38808 6736 38820
rect 6043 38780 6736 38808
rect 6043 38777 6055 38780
rect 5997 38771 6055 38777
rect 6730 38768 6736 38780
rect 6788 38808 6794 38820
rect 7484 38808 7512 38836
rect 6788 38780 7512 38808
rect 6788 38768 6794 38780
rect 7650 38768 7656 38820
rect 7708 38768 7714 38820
rect 8110 38768 8116 38820
rect 8168 38808 8174 38820
rect 8864 38808 8892 38836
rect 8168 38780 8892 38808
rect 8168 38768 8174 38780
rect 10594 38768 10600 38820
rect 10652 38808 10658 38820
rect 10704 38808 10732 38984
rect 10796 38944 10824 39052
rect 12526 39040 12532 39092
rect 12584 39080 12590 39092
rect 12710 39080 12716 39092
rect 12584 39052 12716 39080
rect 12584 39040 12590 39052
rect 12710 39040 12716 39052
rect 12768 39040 12774 39092
rect 13630 39080 13636 39092
rect 13591 39052 13636 39080
rect 13630 39040 13636 39052
rect 13688 39040 13694 39092
rect 14366 39080 14372 39092
rect 14327 39052 14372 39080
rect 14366 39040 14372 39052
rect 14424 39040 14430 39092
rect 15378 39040 15384 39092
rect 15436 39080 15442 39092
rect 15933 39083 15991 39089
rect 15933 39080 15945 39083
rect 15436 39052 15945 39080
rect 15436 39040 15442 39052
rect 15933 39049 15945 39052
rect 15979 39080 15991 39083
rect 16482 39080 16488 39092
rect 15979 39052 16488 39080
rect 15979 39049 15991 39052
rect 15933 39043 15991 39049
rect 16482 39040 16488 39052
rect 16540 39040 16546 39092
rect 18230 39080 18236 39092
rect 18191 39052 18236 39080
rect 18230 39040 18236 39052
rect 18288 39040 18294 39092
rect 12342 38972 12348 39024
rect 12400 39012 12406 39024
rect 12400 38984 13216 39012
rect 12400 38972 12406 38984
rect 10962 38944 10968 38956
rect 10796 38916 10968 38944
rect 10796 38885 10824 38916
rect 10962 38904 10968 38916
rect 11020 38904 11026 38956
rect 12986 38944 12992 38956
rect 12947 38916 12992 38944
rect 12986 38904 12992 38916
rect 13044 38904 13050 38956
rect 10781 38879 10839 38885
rect 10781 38845 10793 38879
rect 10827 38845 10839 38879
rect 11054 38876 11060 38888
rect 11015 38848 11060 38876
rect 10781 38839 10839 38845
rect 11054 38836 11060 38848
rect 11112 38836 11118 38888
rect 11974 38876 11980 38888
rect 11935 38848 11980 38876
rect 11974 38836 11980 38848
rect 12032 38836 12038 38888
rect 12158 38876 12164 38888
rect 12119 38848 12164 38876
rect 12158 38836 12164 38848
rect 12216 38836 12222 38888
rect 13188 38885 13216 38984
rect 13630 38904 13636 38956
rect 13688 38944 13694 38956
rect 14384 38944 14412 39040
rect 16206 39012 16212 39024
rect 16167 38984 16212 39012
rect 16206 38972 16212 38984
rect 16264 38972 16270 39024
rect 13688 38916 14412 38944
rect 15657 38947 15715 38953
rect 13688 38904 13694 38916
rect 15657 38913 15669 38947
rect 15703 38944 15715 38947
rect 15703 38916 16988 38944
rect 15703 38913 15715 38916
rect 15657 38907 15715 38913
rect 16960 38888 16988 38916
rect 12805 38879 12863 38885
rect 12805 38845 12817 38879
rect 12851 38845 12863 38879
rect 12805 38839 12863 38845
rect 13173 38879 13231 38885
rect 13173 38845 13185 38879
rect 13219 38876 13231 38879
rect 13538 38876 13544 38888
rect 13219 38848 13544 38876
rect 13219 38845 13231 38848
rect 13173 38839 13231 38845
rect 10652 38780 10732 38808
rect 11701 38811 11759 38817
rect 10652 38768 10658 38780
rect 11701 38777 11713 38811
rect 11747 38808 11759 38811
rect 12820 38808 12848 38839
rect 13538 38836 13544 38848
rect 13596 38836 13602 38888
rect 14185 38879 14243 38885
rect 14185 38876 14197 38879
rect 13832 38848 14197 38876
rect 13722 38808 13728 38820
rect 11747 38780 13728 38808
rect 11747 38777 11759 38780
rect 11701 38771 11759 38777
rect 13722 38768 13728 38780
rect 13780 38768 13786 38820
rect 6641 38743 6699 38749
rect 6641 38709 6653 38743
rect 6687 38740 6699 38743
rect 7668 38740 7696 38768
rect 6687 38712 7696 38740
rect 6687 38709 6699 38712
rect 6641 38703 6699 38709
rect 8846 38700 8852 38752
rect 8904 38740 8910 38752
rect 12434 38740 12440 38752
rect 8904 38712 12440 38740
rect 8904 38700 8910 38712
rect 12434 38700 12440 38712
rect 12492 38700 12498 38752
rect 13446 38700 13452 38752
rect 13504 38740 13510 38752
rect 13832 38740 13860 38848
rect 14185 38845 14197 38848
rect 14231 38876 14243 38879
rect 14645 38879 14703 38885
rect 14645 38876 14657 38879
rect 14231 38848 14657 38876
rect 14231 38845 14243 38848
rect 14185 38839 14243 38845
rect 14645 38845 14657 38848
rect 14691 38845 14703 38879
rect 14645 38839 14703 38845
rect 15105 38879 15163 38885
rect 15105 38845 15117 38879
rect 15151 38876 15163 38879
rect 15286 38876 15292 38888
rect 15151 38848 15292 38876
rect 15151 38845 15163 38848
rect 15105 38839 15163 38845
rect 15286 38836 15292 38848
rect 15344 38876 15350 38888
rect 16298 38876 16304 38888
rect 15344 38848 16304 38876
rect 15344 38836 15350 38848
rect 16298 38836 16304 38848
rect 16356 38836 16362 38888
rect 16482 38876 16488 38888
rect 16443 38848 16488 38876
rect 16482 38836 16488 38848
rect 16540 38836 16546 38888
rect 16853 38879 16911 38885
rect 16853 38845 16865 38879
rect 16899 38845 16911 38879
rect 16853 38839 16911 38845
rect 14093 38811 14151 38817
rect 14093 38777 14105 38811
rect 14139 38808 14151 38811
rect 15930 38808 15936 38820
rect 14139 38780 15936 38808
rect 14139 38777 14151 38780
rect 14093 38771 14151 38777
rect 15930 38768 15936 38780
rect 15988 38768 15994 38820
rect 16758 38768 16764 38820
rect 16816 38808 16822 38820
rect 16868 38808 16896 38839
rect 16942 38836 16948 38888
rect 17000 38876 17006 38888
rect 17405 38879 17463 38885
rect 17405 38876 17417 38879
rect 17000 38848 17417 38876
rect 17000 38836 17006 38848
rect 17405 38845 17417 38848
rect 17451 38845 17463 38879
rect 17405 38839 17463 38845
rect 17865 38811 17923 38817
rect 17865 38808 17877 38811
rect 16816 38780 17877 38808
rect 16816 38768 16822 38780
rect 17865 38777 17877 38780
rect 17911 38808 17923 38811
rect 18046 38808 18052 38820
rect 17911 38780 18052 38808
rect 17911 38777 17923 38780
rect 17865 38771 17923 38777
rect 18046 38768 18052 38780
rect 18104 38768 18110 38820
rect 13504 38712 13860 38740
rect 13504 38700 13510 38712
rect 1104 38650 18860 38672
rect 1104 38598 7648 38650
rect 7700 38598 7712 38650
rect 7764 38598 7776 38650
rect 7828 38598 7840 38650
rect 7892 38598 14315 38650
rect 14367 38598 14379 38650
rect 14431 38598 14443 38650
rect 14495 38598 14507 38650
rect 14559 38598 18860 38650
rect 1104 38576 18860 38598
rect 3881 38539 3939 38545
rect 3881 38505 3893 38539
rect 3927 38536 3939 38539
rect 4614 38536 4620 38548
rect 3927 38508 4620 38536
rect 3927 38505 3939 38508
rect 3881 38499 3939 38505
rect 4614 38496 4620 38508
rect 4672 38536 4678 38548
rect 5353 38539 5411 38545
rect 5353 38536 5365 38539
rect 4672 38508 5365 38536
rect 4672 38496 4678 38508
rect 5353 38505 5365 38508
rect 5399 38505 5411 38539
rect 5353 38499 5411 38505
rect 5534 38496 5540 38548
rect 5592 38536 5598 38548
rect 6549 38539 6607 38545
rect 6549 38536 6561 38539
rect 5592 38508 6561 38536
rect 5592 38496 5598 38508
rect 6549 38505 6561 38508
rect 6595 38505 6607 38539
rect 6549 38499 6607 38505
rect 3145 38471 3203 38477
rect 3145 38437 3157 38471
rect 3191 38468 3203 38471
rect 3970 38468 3976 38480
rect 3191 38440 3976 38468
rect 3191 38437 3203 38440
rect 3145 38431 3203 38437
rect 3970 38428 3976 38440
rect 4028 38428 4034 38480
rect 1578 38360 1584 38412
rect 1636 38400 1642 38412
rect 1765 38403 1823 38409
rect 1765 38400 1777 38403
rect 1636 38372 1777 38400
rect 1636 38360 1642 38372
rect 1765 38369 1777 38372
rect 1811 38369 1823 38403
rect 1765 38363 1823 38369
rect 3510 38360 3516 38412
rect 3568 38400 3574 38412
rect 4249 38403 4307 38409
rect 4249 38400 4261 38403
rect 3568 38372 4261 38400
rect 3568 38360 3574 38372
rect 4249 38369 4261 38372
rect 4295 38400 4307 38403
rect 5350 38400 5356 38412
rect 4295 38372 5356 38400
rect 4295 38369 4307 38372
rect 4249 38363 4307 38369
rect 5350 38360 5356 38372
rect 5408 38400 5414 38412
rect 5552 38400 5580 38496
rect 5408 38372 5580 38400
rect 5408 38360 5414 38372
rect 1489 38335 1547 38341
rect 1489 38301 1501 38335
rect 1535 38332 1547 38335
rect 1670 38332 1676 38344
rect 1535 38304 1676 38332
rect 1535 38301 1547 38304
rect 1489 38295 1547 38301
rect 1670 38292 1676 38304
rect 1728 38292 1734 38344
rect 3970 38332 3976 38344
rect 3931 38304 3976 38332
rect 3970 38292 3976 38304
rect 4028 38292 4034 38344
rect 6564 38332 6592 38499
rect 6822 38496 6828 38548
rect 6880 38536 6886 38548
rect 7009 38539 7067 38545
rect 7009 38536 7021 38539
rect 6880 38508 7021 38536
rect 6880 38496 6886 38508
rect 7009 38505 7021 38508
rect 7055 38505 7067 38539
rect 7009 38499 7067 38505
rect 7929 38539 7987 38545
rect 7929 38505 7941 38539
rect 7975 38536 7987 38539
rect 8110 38536 8116 38548
rect 7975 38508 8116 38536
rect 7975 38505 7987 38508
rect 7929 38499 7987 38505
rect 8110 38496 8116 38508
rect 8168 38496 8174 38548
rect 9306 38496 9312 38548
rect 9364 38496 9370 38548
rect 10502 38496 10508 38548
rect 10560 38536 10566 38548
rect 10778 38536 10784 38548
rect 10560 38508 10784 38536
rect 10560 38496 10566 38508
rect 10778 38496 10784 38508
rect 10836 38496 10842 38548
rect 10870 38496 10876 38548
rect 10928 38536 10934 38548
rect 11793 38539 11851 38545
rect 11793 38536 11805 38539
rect 10928 38508 11805 38536
rect 10928 38496 10934 38508
rect 11793 38505 11805 38508
rect 11839 38536 11851 38539
rect 12434 38536 12440 38548
rect 11839 38508 12440 38536
rect 11839 38505 11851 38508
rect 11793 38499 11851 38505
rect 12434 38496 12440 38508
rect 12492 38496 12498 38548
rect 12802 38496 12808 38548
rect 12860 38536 12866 38548
rect 13449 38539 13507 38545
rect 13449 38536 13461 38539
rect 12860 38508 13461 38536
rect 12860 38496 12866 38508
rect 13449 38505 13461 38508
rect 13495 38505 13507 38539
rect 13449 38499 13507 38505
rect 13722 38496 13728 38548
rect 13780 38536 13786 38548
rect 14001 38539 14059 38545
rect 14001 38536 14013 38539
rect 13780 38508 14013 38536
rect 13780 38496 13786 38508
rect 14001 38505 14013 38508
rect 14047 38505 14059 38539
rect 14001 38499 14059 38505
rect 14461 38539 14519 38545
rect 14461 38505 14473 38539
rect 14507 38536 14519 38539
rect 15286 38536 15292 38548
rect 14507 38508 15292 38536
rect 14507 38505 14519 38508
rect 14461 38499 14519 38505
rect 7561 38471 7619 38477
rect 7561 38437 7573 38471
rect 7607 38468 7619 38471
rect 8478 38468 8484 38480
rect 7607 38440 8484 38468
rect 7607 38437 7619 38440
rect 7561 38431 7619 38437
rect 8478 38428 8484 38440
rect 8536 38428 8542 38480
rect 9324 38468 9352 38496
rect 8680 38440 9352 38468
rect 10045 38471 10103 38477
rect 6822 38400 6828 38412
rect 6783 38372 6828 38400
rect 6822 38360 6828 38372
rect 6880 38360 6886 38412
rect 8680 38409 8708 38440
rect 10045 38437 10057 38471
rect 10091 38468 10103 38471
rect 10597 38471 10655 38477
rect 10597 38468 10609 38471
rect 10091 38440 10609 38468
rect 10091 38437 10103 38440
rect 10045 38431 10103 38437
rect 10597 38437 10609 38440
rect 10643 38468 10655 38471
rect 10962 38468 10968 38480
rect 10643 38440 10968 38468
rect 10643 38437 10655 38440
rect 10597 38431 10655 38437
rect 10962 38428 10968 38440
rect 11020 38428 11026 38480
rect 11517 38471 11575 38477
rect 11517 38437 11529 38471
rect 11563 38468 11575 38471
rect 12161 38471 12219 38477
rect 12161 38468 12173 38471
rect 11563 38440 12173 38468
rect 11563 38437 11575 38440
rect 11517 38431 11575 38437
rect 12161 38437 12173 38440
rect 12207 38468 12219 38471
rect 12342 38468 12348 38480
rect 12207 38440 12348 38468
rect 12207 38437 12219 38440
rect 12161 38431 12219 38437
rect 12342 38428 12348 38440
rect 12400 38428 12406 38480
rect 8021 38403 8079 38409
rect 8021 38369 8033 38403
rect 8067 38369 8079 38403
rect 8021 38363 8079 38369
rect 8665 38403 8723 38409
rect 8665 38369 8677 38403
rect 8711 38369 8723 38403
rect 8665 38363 8723 38369
rect 8757 38403 8815 38409
rect 8757 38369 8769 38403
rect 8803 38400 8815 38403
rect 8938 38400 8944 38412
rect 8803 38372 8944 38400
rect 8803 38369 8815 38372
rect 8757 38363 8815 38369
rect 8036 38332 8064 38363
rect 6564 38304 8064 38332
rect 8386 38292 8392 38344
rect 8444 38332 8450 38344
rect 8772 38332 8800 38363
rect 8938 38360 8944 38372
rect 8996 38360 9002 38412
rect 9309 38403 9367 38409
rect 9309 38400 9321 38403
rect 9140 38372 9321 38400
rect 8444 38304 8800 38332
rect 8444 38292 8450 38304
rect 8570 38224 8576 38276
rect 8628 38264 8634 38276
rect 9140 38264 9168 38372
rect 9309 38369 9321 38372
rect 9355 38369 9367 38403
rect 9309 38363 9367 38369
rect 9766 38360 9772 38412
rect 9824 38400 9830 38412
rect 10778 38400 10784 38412
rect 9824 38372 10784 38400
rect 9824 38360 9830 38372
rect 10778 38360 10784 38372
rect 10836 38360 10842 38412
rect 10870 38360 10876 38412
rect 10928 38400 10934 38412
rect 11241 38403 11299 38409
rect 11241 38400 11253 38403
rect 10928 38372 11253 38400
rect 10928 38360 10934 38372
rect 11241 38369 11253 38372
rect 11287 38369 11299 38403
rect 11241 38363 11299 38369
rect 12989 38403 13047 38409
rect 12989 38369 13001 38403
rect 13035 38369 13047 38403
rect 12989 38363 13047 38369
rect 13265 38403 13323 38409
rect 13265 38369 13277 38403
rect 13311 38400 13323 38403
rect 13630 38400 13636 38412
rect 13311 38372 13636 38400
rect 13311 38369 13323 38372
rect 13265 38363 13323 38369
rect 10229 38335 10287 38341
rect 10229 38301 10241 38335
rect 10275 38332 10287 38335
rect 10410 38332 10416 38344
rect 10275 38304 10416 38332
rect 10275 38301 10287 38304
rect 10229 38295 10287 38301
rect 10410 38292 10416 38304
rect 10468 38332 10474 38344
rect 10888 38332 10916 38360
rect 10468 38304 10916 38332
rect 13004 38332 13032 38363
rect 13630 38360 13636 38372
rect 13688 38360 13694 38412
rect 13722 38332 13728 38344
rect 13004 38304 13728 38332
rect 10468 38292 10474 38304
rect 13722 38292 13728 38304
rect 13780 38292 13786 38344
rect 14016 38332 14044 38499
rect 14734 38400 14740 38412
rect 14695 38372 14740 38400
rect 14734 38360 14740 38372
rect 14792 38360 14798 38412
rect 14936 38409 14964 38508
rect 15286 38496 15292 38508
rect 15344 38536 15350 38548
rect 15838 38536 15844 38548
rect 15344 38508 15844 38536
rect 15344 38496 15350 38508
rect 15838 38496 15844 38508
rect 15896 38496 15902 38548
rect 16393 38539 16451 38545
rect 16393 38505 16405 38539
rect 16439 38536 16451 38539
rect 16761 38539 16819 38545
rect 16761 38536 16773 38539
rect 16439 38508 16773 38536
rect 16439 38505 16451 38508
rect 16393 38499 16451 38505
rect 16761 38505 16773 38508
rect 16807 38536 16819 38539
rect 16850 38536 16856 38548
rect 16807 38508 16856 38536
rect 16807 38505 16819 38508
rect 16761 38499 16819 38505
rect 16850 38496 16856 38508
rect 16908 38536 16914 38548
rect 17037 38539 17095 38545
rect 17037 38536 17049 38539
rect 16908 38508 17049 38536
rect 16908 38496 16914 38508
rect 17037 38505 17049 38508
rect 17083 38536 17095 38539
rect 17310 38536 17316 38548
rect 17083 38508 17316 38536
rect 17083 38505 17095 38508
rect 17037 38499 17095 38505
rect 17310 38496 17316 38508
rect 17368 38496 17374 38548
rect 14921 38403 14979 38409
rect 14921 38369 14933 38403
rect 14967 38369 14979 38403
rect 15562 38400 15568 38412
rect 15523 38372 15568 38400
rect 14921 38363 14979 38369
rect 15562 38360 15568 38372
rect 15620 38360 15626 38412
rect 15841 38403 15899 38409
rect 15841 38369 15853 38403
rect 15887 38400 15899 38403
rect 16850 38400 16856 38412
rect 15887 38372 16856 38400
rect 15887 38369 15899 38372
rect 15841 38363 15899 38369
rect 15856 38332 15884 38363
rect 16850 38360 16856 38372
rect 16908 38360 16914 38412
rect 14016 38304 15884 38332
rect 16298 38292 16304 38344
rect 16356 38332 16362 38344
rect 17313 38335 17371 38341
rect 17313 38332 17325 38335
rect 16356 38304 17325 38332
rect 16356 38292 16362 38304
rect 17313 38301 17325 38304
rect 17359 38301 17371 38335
rect 17313 38295 17371 38301
rect 8628 38236 9168 38264
rect 8628 38224 8634 38236
rect 9766 38224 9772 38276
rect 9824 38264 9830 38276
rect 10045 38267 10103 38273
rect 10045 38264 10057 38267
rect 9824 38236 10057 38264
rect 9824 38224 9830 38236
rect 10045 38233 10057 38236
rect 10091 38233 10103 38267
rect 10045 38227 10103 38233
rect 11238 38224 11244 38276
rect 11296 38224 11302 38276
rect 12802 38224 12808 38276
rect 12860 38264 12866 38276
rect 12897 38267 12955 38273
rect 12897 38264 12909 38267
rect 12860 38236 12909 38264
rect 12860 38224 12866 38236
rect 12897 38233 12909 38236
rect 12943 38264 12955 38267
rect 13081 38267 13139 38273
rect 13081 38264 13093 38267
rect 12943 38236 13093 38264
rect 12943 38233 12955 38236
rect 12897 38227 12955 38233
rect 13081 38233 13093 38236
rect 13127 38233 13139 38267
rect 13081 38227 13139 38233
rect 13538 38224 13544 38276
rect 13596 38264 13602 38276
rect 15654 38264 15660 38276
rect 13596 38236 15660 38264
rect 13596 38224 13602 38236
rect 15654 38224 15660 38236
rect 15712 38224 15718 38276
rect 3513 38199 3571 38205
rect 3513 38165 3525 38199
rect 3559 38196 3571 38199
rect 5074 38196 5080 38208
rect 3559 38168 5080 38196
rect 3559 38165 3571 38168
rect 3513 38159 3571 38165
rect 5074 38156 5080 38168
rect 5132 38156 5138 38208
rect 6178 38196 6184 38208
rect 6139 38168 6184 38196
rect 6178 38156 6184 38168
rect 6236 38156 6242 38208
rect 9214 38196 9220 38208
rect 9175 38168 9220 38196
rect 9214 38156 9220 38168
rect 9272 38156 9278 38208
rect 9861 38199 9919 38205
rect 9861 38165 9873 38199
rect 9907 38196 9919 38199
rect 9950 38196 9956 38208
rect 9907 38168 9956 38196
rect 9907 38165 9919 38168
rect 9861 38159 9919 38165
rect 9950 38156 9956 38168
rect 10008 38156 10014 38208
rect 10410 38156 10416 38208
rect 10468 38196 10474 38208
rect 11256 38196 11284 38224
rect 14642 38196 14648 38208
rect 10468 38168 11284 38196
rect 14603 38168 14648 38196
rect 10468 38156 10474 38168
rect 14642 38156 14648 38168
rect 14700 38156 14706 38208
rect 1104 38106 18860 38128
rect 1104 38054 4315 38106
rect 4367 38054 4379 38106
rect 4431 38054 4443 38106
rect 4495 38054 4507 38106
rect 4559 38054 10982 38106
rect 11034 38054 11046 38106
rect 11098 38054 11110 38106
rect 11162 38054 11174 38106
rect 11226 38054 17648 38106
rect 17700 38054 17712 38106
rect 17764 38054 17776 38106
rect 17828 38054 17840 38106
rect 17892 38054 18860 38106
rect 1104 38032 18860 38054
rect 1670 37992 1676 38004
rect 1504 37964 1676 37992
rect 1504 37797 1532 37964
rect 1670 37952 1676 37964
rect 1728 37952 1734 38004
rect 3053 37995 3111 38001
rect 3053 37961 3065 37995
rect 3099 37992 3111 37995
rect 3234 37992 3240 38004
rect 3099 37964 3240 37992
rect 3099 37961 3111 37964
rect 3053 37955 3111 37961
rect 3234 37952 3240 37964
rect 3292 37952 3298 38004
rect 3510 37992 3516 38004
rect 3471 37964 3516 37992
rect 3510 37952 3516 37964
rect 3568 37952 3574 38004
rect 9125 37995 9183 38001
rect 9125 37961 9137 37995
rect 9171 37992 9183 37995
rect 9306 37992 9312 38004
rect 9171 37964 9312 37992
rect 9171 37961 9183 37964
rect 9125 37955 9183 37961
rect 9306 37952 9312 37964
rect 9364 37952 9370 38004
rect 13630 37952 13636 38004
rect 13688 37992 13694 38004
rect 13817 37995 13875 38001
rect 13817 37992 13829 37995
rect 13688 37964 13829 37992
rect 13688 37952 13694 37964
rect 13817 37961 13829 37964
rect 13863 37961 13875 37995
rect 13817 37955 13875 37961
rect 14369 37995 14427 38001
rect 14369 37961 14381 37995
rect 14415 37992 14427 37995
rect 15010 37992 15016 38004
rect 14415 37964 15016 37992
rect 14415 37961 14427 37964
rect 14369 37955 14427 37961
rect 15010 37952 15016 37964
rect 15068 37952 15074 38004
rect 15105 37995 15163 38001
rect 15105 37961 15117 37995
rect 15151 37992 15163 37995
rect 15562 37992 15568 38004
rect 15151 37964 15568 37992
rect 15151 37961 15163 37964
rect 15105 37955 15163 37961
rect 7374 37924 7380 37936
rect 7335 37896 7380 37924
rect 7374 37884 7380 37896
rect 7432 37884 7438 37936
rect 7466 37884 7472 37936
rect 7524 37924 7530 37936
rect 8110 37924 8116 37936
rect 7524 37896 8116 37924
rect 7524 37884 7530 37896
rect 8110 37884 8116 37896
rect 8168 37884 8174 37936
rect 10410 37884 10416 37936
rect 10468 37924 10474 37936
rect 10468 37896 10548 37924
rect 10468 37884 10474 37896
rect 5534 37816 5540 37868
rect 5592 37856 5598 37868
rect 5994 37856 6000 37868
rect 5592 37828 6000 37856
rect 5592 37816 5598 37828
rect 5994 37816 6000 37828
rect 6052 37816 6058 37868
rect 9677 37859 9735 37865
rect 6932 37828 8524 37856
rect 6932 37800 6960 37828
rect 1489 37791 1547 37797
rect 1489 37757 1501 37791
rect 1535 37757 1547 37791
rect 1489 37751 1547 37757
rect 1765 37791 1823 37797
rect 1765 37757 1777 37791
rect 1811 37788 1823 37791
rect 1854 37788 1860 37800
rect 1811 37760 1860 37788
rect 1811 37757 1823 37760
rect 1765 37751 1823 37757
rect 1504 37652 1532 37751
rect 1854 37748 1860 37760
rect 1912 37748 1918 37800
rect 3602 37748 3608 37800
rect 3660 37788 3666 37800
rect 3970 37788 3976 37800
rect 3660 37760 3976 37788
rect 3660 37748 3666 37760
rect 3970 37748 3976 37760
rect 4028 37788 4034 37800
rect 4065 37791 4123 37797
rect 4065 37788 4077 37791
rect 4028 37760 4077 37788
rect 4028 37748 4034 37760
rect 4065 37757 4077 37760
rect 4111 37757 4123 37791
rect 4341 37791 4399 37797
rect 4341 37788 4353 37791
rect 4065 37751 4123 37757
rect 4172 37760 4353 37788
rect 1762 37652 1768 37664
rect 1504 37624 1768 37652
rect 1762 37612 1768 37624
rect 1820 37612 1826 37664
rect 3786 37652 3792 37664
rect 3747 37624 3792 37652
rect 3786 37612 3792 37624
rect 3844 37652 3850 37664
rect 4172 37652 4200 37760
rect 4341 37757 4353 37760
rect 4387 37757 4399 37791
rect 6730 37788 6736 37800
rect 6691 37760 6736 37788
rect 4341 37751 4399 37757
rect 6730 37748 6736 37760
rect 6788 37748 6794 37800
rect 6914 37788 6920 37800
rect 6875 37760 6920 37788
rect 6914 37748 6920 37760
rect 6972 37748 6978 37800
rect 7466 37788 7472 37800
rect 7427 37760 7472 37788
rect 7466 37748 7472 37760
rect 7524 37748 7530 37800
rect 8496 37797 8524 37828
rect 9677 37825 9689 37859
rect 9723 37856 9735 37859
rect 10134 37856 10140 37868
rect 9723 37828 10140 37856
rect 9723 37825 9735 37828
rect 9677 37819 9735 37825
rect 10134 37816 10140 37828
rect 10192 37816 10198 37868
rect 8481 37791 8539 37797
rect 8481 37757 8493 37791
rect 8527 37757 8539 37791
rect 8481 37751 8539 37757
rect 9122 37748 9128 37800
rect 9180 37788 9186 37800
rect 10413 37791 10471 37797
rect 10413 37788 10425 37791
rect 9180 37760 10425 37788
rect 9180 37748 9186 37760
rect 10413 37757 10425 37760
rect 10459 37757 10471 37791
rect 10413 37751 10471 37757
rect 5721 37723 5779 37729
rect 5721 37689 5733 37723
rect 5767 37720 5779 37723
rect 5994 37720 6000 37732
rect 5767 37692 6000 37720
rect 5767 37689 5779 37692
rect 5721 37683 5779 37689
rect 5994 37680 6000 37692
rect 6052 37680 6058 37732
rect 6089 37723 6147 37729
rect 6089 37689 6101 37723
rect 6135 37720 6147 37723
rect 6822 37720 6828 37732
rect 6135 37692 6828 37720
rect 6135 37689 6147 37692
rect 6089 37683 6147 37689
rect 6822 37680 6828 37692
rect 6880 37680 6886 37732
rect 9493 37723 9551 37729
rect 9493 37689 9505 37723
rect 9539 37720 9551 37723
rect 9858 37720 9864 37732
rect 9539 37692 9864 37720
rect 9539 37689 9551 37692
rect 9493 37683 9551 37689
rect 9858 37680 9864 37692
rect 9916 37680 9922 37732
rect 10045 37723 10103 37729
rect 10045 37689 10057 37723
rect 10091 37720 10103 37723
rect 10520 37720 10548 37896
rect 11422 37816 11428 37868
rect 11480 37856 11486 37868
rect 11882 37856 11888 37868
rect 11480 37828 11888 37856
rect 11480 37816 11486 37828
rect 11882 37816 11888 37828
rect 11940 37856 11946 37868
rect 12618 37856 12624 37868
rect 11940 37828 12480 37856
rect 12579 37828 12624 37856
rect 11940 37816 11946 37828
rect 11974 37788 11980 37800
rect 11935 37760 11980 37788
rect 11974 37748 11980 37760
rect 12032 37748 12038 37800
rect 12066 37748 12072 37800
rect 12124 37788 12130 37800
rect 12345 37791 12403 37797
rect 12345 37788 12357 37791
rect 12124 37760 12357 37788
rect 12124 37748 12130 37760
rect 12345 37757 12357 37760
rect 12391 37757 12403 37791
rect 12452 37788 12480 37828
rect 12618 37816 12624 37828
rect 12676 37816 12682 37868
rect 12713 37791 12771 37797
rect 12713 37788 12725 37791
rect 12452 37760 12725 37788
rect 12345 37751 12403 37757
rect 12713 37757 12725 37760
rect 12759 37757 12771 37791
rect 12713 37751 12771 37757
rect 14185 37791 14243 37797
rect 14185 37757 14197 37791
rect 14231 37757 14243 37791
rect 14185 37751 14243 37757
rect 10962 37720 10968 37732
rect 10091 37692 10968 37720
rect 10091 37689 10103 37692
rect 10045 37683 10103 37689
rect 10962 37680 10968 37692
rect 11020 37680 11026 37732
rect 12434 37680 12440 37732
rect 12492 37720 12498 37732
rect 14200 37720 14228 37751
rect 14918 37748 14924 37800
rect 14976 37788 14982 37800
rect 15120 37788 15148 37955
rect 15562 37952 15568 37964
rect 15620 37952 15626 38004
rect 15933 37995 15991 38001
rect 15933 37961 15945 37995
rect 15979 37992 15991 37995
rect 16482 37992 16488 38004
rect 15979 37964 16488 37992
rect 15979 37961 15991 37964
rect 15933 37955 15991 37961
rect 16482 37952 16488 37964
rect 16540 37952 16546 38004
rect 16850 37952 16856 38004
rect 16908 37992 16914 38004
rect 17773 37995 17831 38001
rect 17773 37992 17785 37995
rect 16908 37964 17785 37992
rect 16908 37952 16914 37964
rect 17773 37961 17785 37964
rect 17819 37992 17831 37995
rect 17954 37992 17960 38004
rect 17819 37964 17960 37992
rect 17819 37961 17831 37964
rect 17773 37955 17831 37961
rect 17954 37952 17960 37964
rect 18012 37952 18018 38004
rect 16850 37856 16856 37868
rect 16811 37828 16856 37856
rect 16850 37816 16856 37828
rect 16908 37816 16914 37868
rect 14976 37760 15148 37788
rect 14976 37748 14982 37760
rect 15562 37748 15568 37800
rect 15620 37788 15626 37800
rect 15930 37788 15936 37800
rect 15620 37760 15936 37788
rect 15620 37748 15626 37760
rect 15930 37748 15936 37760
rect 15988 37788 15994 37800
rect 16025 37791 16083 37797
rect 16025 37788 16037 37791
rect 15988 37760 16037 37788
rect 15988 37748 15994 37760
rect 16025 37757 16037 37760
rect 16071 37757 16083 37791
rect 16025 37751 16083 37757
rect 16393 37791 16451 37797
rect 16393 37757 16405 37791
rect 16439 37757 16451 37791
rect 16393 37751 16451 37757
rect 14645 37723 14703 37729
rect 14645 37720 14657 37723
rect 12492 37692 14657 37720
rect 12492 37680 12498 37692
rect 14645 37689 14657 37692
rect 14691 37689 14703 37723
rect 14645 37683 14703 37689
rect 14734 37680 14740 37732
rect 14792 37720 14798 37732
rect 15473 37723 15531 37729
rect 15473 37720 15485 37723
rect 14792 37692 15485 37720
rect 14792 37680 14798 37692
rect 15473 37689 15485 37692
rect 15519 37689 15531 37723
rect 15473 37683 15531 37689
rect 15654 37680 15660 37732
rect 15712 37720 15718 37732
rect 16298 37720 16304 37732
rect 15712 37692 16304 37720
rect 15712 37680 15718 37692
rect 16298 37680 16304 37692
rect 16356 37720 16362 37732
rect 16408 37720 16436 37751
rect 16482 37748 16488 37800
rect 16540 37788 16546 37800
rect 16761 37791 16819 37797
rect 16761 37788 16773 37791
rect 16540 37760 16773 37788
rect 16540 37748 16546 37760
rect 16761 37757 16773 37760
rect 16807 37757 16819 37791
rect 17310 37788 17316 37800
rect 17271 37760 17316 37788
rect 16761 37751 16819 37757
rect 17310 37748 17316 37760
rect 17368 37748 17374 37800
rect 16356 37692 16436 37720
rect 16356 37680 16362 37692
rect 3844 37624 4200 37652
rect 6457 37655 6515 37661
rect 3844 37612 3850 37624
rect 6457 37621 6469 37655
rect 6503 37652 6515 37655
rect 7006 37652 7012 37664
rect 6503 37624 7012 37652
rect 6503 37621 6515 37624
rect 6457 37615 6515 37621
rect 7006 37612 7012 37624
rect 7064 37652 7070 37664
rect 7466 37652 7472 37664
rect 7064 37624 7472 37652
rect 7064 37612 7070 37624
rect 7466 37612 7472 37624
rect 7524 37612 7530 37664
rect 8113 37655 8171 37661
rect 8113 37621 8125 37655
rect 8159 37652 8171 37655
rect 8386 37652 8392 37664
rect 8159 37624 8392 37652
rect 8159 37621 8171 37624
rect 8113 37615 8171 37621
rect 8386 37612 8392 37624
rect 8444 37612 8450 37664
rect 8478 37612 8484 37664
rect 8536 37652 8542 37664
rect 8665 37655 8723 37661
rect 8665 37652 8677 37655
rect 8536 37624 8677 37652
rect 8536 37612 8542 37624
rect 8665 37621 8677 37624
rect 8711 37621 8723 37655
rect 8665 37615 8723 37621
rect 9306 37612 9312 37664
rect 9364 37652 9370 37664
rect 9953 37655 10011 37661
rect 9953 37652 9965 37655
rect 9364 37624 9965 37652
rect 9364 37612 9370 37624
rect 9953 37621 9965 37624
rect 9999 37621 10011 37655
rect 9953 37615 10011 37621
rect 10410 37612 10416 37664
rect 10468 37652 10474 37664
rect 10778 37652 10784 37664
rect 10468 37624 10784 37652
rect 10468 37612 10474 37624
rect 10778 37612 10784 37624
rect 10836 37612 10842 37664
rect 10870 37612 10876 37664
rect 10928 37652 10934 37664
rect 11149 37655 11207 37661
rect 11149 37652 11161 37655
rect 10928 37624 11161 37652
rect 10928 37612 10934 37624
rect 11149 37621 11161 37624
rect 11195 37621 11207 37655
rect 11882 37652 11888 37664
rect 11843 37624 11888 37652
rect 11149 37615 11207 37621
rect 11882 37612 11888 37624
rect 11940 37612 11946 37664
rect 13541 37655 13599 37661
rect 13541 37621 13553 37655
rect 13587 37652 13599 37655
rect 13722 37652 13728 37664
rect 13587 37624 13728 37652
rect 13587 37621 13599 37624
rect 13541 37615 13599 37621
rect 13722 37612 13728 37624
rect 13780 37612 13786 37664
rect 14090 37612 14096 37664
rect 14148 37652 14154 37664
rect 15930 37652 15936 37664
rect 14148 37624 15936 37652
rect 14148 37612 14154 37624
rect 15930 37612 15936 37624
rect 15988 37612 15994 37664
rect 1104 37562 18860 37584
rect 1104 37510 7648 37562
rect 7700 37510 7712 37562
rect 7764 37510 7776 37562
rect 7828 37510 7840 37562
rect 7892 37510 14315 37562
rect 14367 37510 14379 37562
rect 14431 37510 14443 37562
rect 14495 37510 14507 37562
rect 14559 37510 18860 37562
rect 1104 37488 18860 37510
rect 4985 37451 5043 37457
rect 4985 37417 4997 37451
rect 5031 37448 5043 37451
rect 5074 37448 5080 37460
rect 5031 37420 5080 37448
rect 5031 37417 5043 37420
rect 4985 37411 5043 37417
rect 5074 37408 5080 37420
rect 5132 37408 5138 37460
rect 6641 37451 6699 37457
rect 6641 37417 6653 37451
rect 6687 37448 6699 37451
rect 6914 37448 6920 37460
rect 6687 37420 6920 37448
rect 6687 37417 6699 37420
rect 6641 37411 6699 37417
rect 6914 37408 6920 37420
rect 6972 37448 6978 37460
rect 7285 37451 7343 37457
rect 7285 37448 7297 37451
rect 6972 37420 7297 37448
rect 6972 37408 6978 37420
rect 7285 37417 7297 37420
rect 7331 37417 7343 37451
rect 7285 37411 7343 37417
rect 7745 37451 7803 37457
rect 7745 37417 7757 37451
rect 7791 37448 7803 37451
rect 9306 37448 9312 37460
rect 7791 37420 9312 37448
rect 7791 37417 7803 37420
rect 7745 37411 7803 37417
rect 9306 37408 9312 37420
rect 9364 37408 9370 37460
rect 11238 37408 11244 37460
rect 11296 37448 11302 37460
rect 11425 37451 11483 37457
rect 11425 37448 11437 37451
rect 11296 37420 11437 37448
rect 11296 37408 11302 37420
rect 11425 37417 11437 37420
rect 11471 37417 11483 37451
rect 11425 37411 11483 37417
rect 12342 37408 12348 37460
rect 12400 37448 12406 37460
rect 13725 37451 13783 37457
rect 12400 37420 12664 37448
rect 12400 37408 12406 37420
rect 6273 37383 6331 37389
rect 6273 37349 6285 37383
rect 6319 37380 6331 37383
rect 6730 37380 6736 37392
rect 6319 37352 6736 37380
rect 6319 37349 6331 37352
rect 6273 37343 6331 37349
rect 6730 37340 6736 37352
rect 6788 37340 6794 37392
rect 8481 37383 8539 37389
rect 8481 37349 8493 37383
rect 8527 37380 8539 37383
rect 9030 37380 9036 37392
rect 8527 37352 9036 37380
rect 8527 37349 8539 37352
rect 8481 37343 8539 37349
rect 9030 37340 9036 37352
rect 9088 37340 9094 37392
rect 11974 37380 11980 37392
rect 9692 37352 11980 37380
rect 1486 37272 1492 37324
rect 1544 37312 1550 37324
rect 1581 37315 1639 37321
rect 1581 37312 1593 37315
rect 1544 37284 1593 37312
rect 1544 37272 1550 37284
rect 1581 37281 1593 37284
rect 1627 37281 1639 37315
rect 1581 37275 1639 37281
rect 1854 37272 1860 37324
rect 1912 37312 1918 37324
rect 1949 37315 2007 37321
rect 1949 37312 1961 37315
rect 1912 37284 1961 37312
rect 1912 37272 1918 37284
rect 1949 37281 1961 37284
rect 1995 37281 2007 37315
rect 1949 37275 2007 37281
rect 3694 37272 3700 37324
rect 3752 37272 3758 37324
rect 6178 37272 6184 37324
rect 6236 37312 6242 37324
rect 6822 37312 6828 37324
rect 6236 37284 6684 37312
rect 6783 37284 6828 37312
rect 6236 37272 6242 37284
rect 3602 37244 3608 37256
rect 3436 37216 3608 37244
rect 1762 37068 1768 37120
rect 1820 37108 1826 37120
rect 2317 37111 2375 37117
rect 2317 37108 2329 37111
rect 1820 37080 2329 37108
rect 1820 37068 1826 37080
rect 2317 37077 2329 37080
rect 2363 37077 2375 37111
rect 2317 37071 2375 37077
rect 3145 37111 3203 37117
rect 3145 37077 3157 37111
rect 3191 37108 3203 37111
rect 3234 37108 3240 37120
rect 3191 37080 3240 37108
rect 3191 37077 3203 37080
rect 3145 37071 3203 37077
rect 3234 37068 3240 37080
rect 3292 37108 3298 37120
rect 3436 37117 3464 37216
rect 3602 37204 3608 37216
rect 3660 37204 3666 37256
rect 3712 37244 3740 37272
rect 3881 37247 3939 37253
rect 3881 37244 3893 37247
rect 3712 37216 3893 37244
rect 3881 37213 3893 37216
rect 3927 37244 3939 37247
rect 3970 37244 3976 37256
rect 3927 37216 3976 37244
rect 3927 37213 3939 37216
rect 3881 37207 3939 37213
rect 3970 37204 3976 37216
rect 4028 37204 4034 37256
rect 6656 37244 6684 37284
rect 6822 37272 6828 37284
rect 6880 37272 6886 37324
rect 6914 37272 6920 37324
rect 6972 37312 6978 37324
rect 7190 37312 7196 37324
rect 6972 37284 7196 37312
rect 6972 37272 6978 37284
rect 7190 37272 7196 37284
rect 7248 37272 7254 37324
rect 8113 37315 8171 37321
rect 8113 37281 8125 37315
rect 8159 37312 8171 37315
rect 8570 37312 8576 37324
rect 8159 37284 8576 37312
rect 8159 37281 8171 37284
rect 8113 37275 8171 37281
rect 8570 37272 8576 37284
rect 8628 37272 8634 37324
rect 8754 37312 8760 37324
rect 8715 37284 8760 37312
rect 8754 37272 8760 37284
rect 8812 37272 8818 37324
rect 9122 37312 9128 37324
rect 9083 37284 9128 37312
rect 9122 37272 9128 37284
rect 9180 37272 9186 37324
rect 9306 37312 9312 37324
rect 9267 37284 9312 37312
rect 9306 37272 9312 37284
rect 9364 37272 9370 37324
rect 9582 37272 9588 37324
rect 9640 37312 9646 37324
rect 9692 37321 9720 37352
rect 11974 37340 11980 37352
rect 12032 37340 12038 37392
rect 12434 37340 12440 37392
rect 12492 37380 12498 37392
rect 12529 37383 12587 37389
rect 12529 37380 12541 37383
rect 12492 37352 12541 37380
rect 12492 37340 12498 37352
rect 12529 37349 12541 37352
rect 12575 37349 12587 37383
rect 12636 37380 12664 37420
rect 13725 37417 13737 37451
rect 13771 37448 13783 37451
rect 14918 37448 14924 37460
rect 13771 37420 14924 37448
rect 13771 37417 13783 37420
rect 13725 37411 13783 37417
rect 14918 37408 14924 37420
rect 14976 37408 14982 37460
rect 15378 37448 15384 37460
rect 15028 37420 15384 37448
rect 12636 37352 12756 37380
rect 12529 37343 12587 37349
rect 9677 37315 9735 37321
rect 9677 37312 9689 37315
rect 9640 37284 9689 37312
rect 9640 37272 9646 37284
rect 9677 37281 9689 37284
rect 9723 37281 9735 37315
rect 10045 37315 10103 37321
rect 10045 37312 10057 37315
rect 9677 37275 9735 37281
rect 9784 37284 10057 37312
rect 7374 37244 7380 37256
rect 6656 37216 7380 37244
rect 7374 37204 7380 37216
rect 7432 37204 7438 37256
rect 8294 37204 8300 37256
rect 8352 37244 8358 37256
rect 9784 37244 9812 37284
rect 10045 37281 10057 37284
rect 10091 37281 10103 37315
rect 10045 37275 10103 37281
rect 10781 37315 10839 37321
rect 10781 37281 10793 37315
rect 10827 37312 10839 37315
rect 11241 37315 11299 37321
rect 10827 37284 11008 37312
rect 10827 37281 10839 37284
rect 10781 37275 10839 37281
rect 8352 37216 9812 37244
rect 10980 37244 11008 37284
rect 11241 37281 11253 37315
rect 11287 37312 11299 37315
rect 11330 37312 11336 37324
rect 11287 37284 11336 37312
rect 11287 37281 11299 37284
rect 11241 37275 11299 37281
rect 11330 37272 11336 37284
rect 11388 37272 11394 37324
rect 12066 37312 12072 37324
rect 12027 37284 12072 37312
rect 12066 37272 12072 37284
rect 12124 37272 12130 37324
rect 12728 37321 12756 37352
rect 12713 37315 12771 37321
rect 12713 37281 12725 37315
rect 12759 37281 12771 37315
rect 12713 37275 12771 37281
rect 13078 37272 13084 37324
rect 13136 37312 13142 37324
rect 14090 37312 14096 37324
rect 13136 37284 14096 37312
rect 13136 37272 13142 37284
rect 14090 37272 14096 37284
rect 14148 37312 14154 37324
rect 14461 37315 14519 37321
rect 14461 37312 14473 37315
rect 14148 37284 14473 37312
rect 14148 37272 14154 37284
rect 14461 37281 14473 37284
rect 14507 37312 14519 37315
rect 14550 37312 14556 37324
rect 14507 37284 14556 37312
rect 14507 37281 14519 37284
rect 14461 37275 14519 37281
rect 14550 37272 14556 37284
rect 14608 37272 14614 37324
rect 15028 37321 15056 37420
rect 15378 37408 15384 37420
rect 15436 37408 15442 37460
rect 17402 37448 17408 37460
rect 17363 37420 17408 37448
rect 17402 37408 17408 37420
rect 17460 37408 17466 37460
rect 15013 37315 15071 37321
rect 15013 37281 15025 37315
rect 15059 37281 15071 37315
rect 15013 37275 15071 37281
rect 12158 37244 12164 37256
rect 10980 37216 12164 37244
rect 8352 37204 8358 37216
rect 12158 37204 12164 37216
rect 12216 37204 12222 37256
rect 14277 37247 14335 37253
rect 14277 37213 14289 37247
rect 14323 37244 14335 37247
rect 14642 37244 14648 37256
rect 14323 37216 14648 37244
rect 14323 37213 14335 37216
rect 14277 37207 14335 37213
rect 14642 37204 14648 37216
rect 14700 37204 14706 37256
rect 15102 37244 15108 37256
rect 15063 37216 15108 37244
rect 15102 37204 15108 37216
rect 15160 37204 15166 37256
rect 15396 37244 15424 37408
rect 15930 37340 15936 37392
rect 15988 37380 15994 37392
rect 15988 37352 16436 37380
rect 15988 37340 15994 37352
rect 15562 37312 15568 37324
rect 15523 37284 15568 37312
rect 15562 37272 15568 37284
rect 15620 37272 15626 37324
rect 15654 37272 15660 37324
rect 15712 37312 15718 37324
rect 16408 37321 16436 37352
rect 15841 37315 15899 37321
rect 15841 37312 15853 37315
rect 15712 37284 15853 37312
rect 15712 37272 15718 37284
rect 15841 37281 15853 37284
rect 15887 37281 15899 37315
rect 16393 37315 16451 37321
rect 16393 37312 16405 37315
rect 16303 37284 16405 37312
rect 15841 37275 15899 37281
rect 16393 37281 16405 37284
rect 16439 37281 16451 37315
rect 16393 37275 16451 37281
rect 16945 37315 17003 37321
rect 16945 37281 16957 37315
rect 16991 37312 17003 37315
rect 17420 37312 17448 37408
rect 16991 37284 17448 37312
rect 16991 37281 17003 37284
rect 16945 37275 17003 37281
rect 15930 37244 15936 37256
rect 15396 37216 15936 37244
rect 15930 37204 15936 37216
rect 15988 37204 15994 37256
rect 16114 37244 16120 37256
rect 16075 37216 16120 37244
rect 16114 37204 16120 37216
rect 16172 37204 16178 37256
rect 6270 37136 6276 37188
rect 6328 37176 6334 37188
rect 7009 37179 7067 37185
rect 7009 37176 7021 37179
rect 6328 37148 7021 37176
rect 6328 37136 6334 37148
rect 7009 37145 7021 37148
rect 7055 37145 7067 37179
rect 7009 37139 7067 37145
rect 10962 37136 10968 37188
rect 11020 37136 11026 37188
rect 3421 37111 3479 37117
rect 3421 37108 3433 37111
rect 3292 37080 3433 37108
rect 3292 37068 3298 37080
rect 3421 37077 3433 37080
rect 3467 37077 3479 37111
rect 5626 37108 5632 37120
rect 5587 37080 5632 37108
rect 3421 37071 3479 37077
rect 5626 37068 5632 37080
rect 5684 37068 5690 37120
rect 8110 37068 8116 37120
rect 8168 37108 8174 37120
rect 8478 37108 8484 37120
rect 8168 37080 8484 37108
rect 8168 37068 8174 37080
rect 8478 37068 8484 37080
rect 8536 37068 8542 37120
rect 10778 37068 10784 37120
rect 10836 37108 10842 37120
rect 10980 37108 11008 37136
rect 11057 37111 11115 37117
rect 11057 37108 11069 37111
rect 10836 37080 11069 37108
rect 10836 37068 10842 37080
rect 11057 37077 11069 37080
rect 11103 37077 11115 37111
rect 11057 37071 11115 37077
rect 14182 37068 14188 37120
rect 14240 37108 14246 37120
rect 15102 37108 15108 37120
rect 14240 37080 15108 37108
rect 14240 37068 14246 37080
rect 15102 37068 15108 37080
rect 15160 37068 15166 37120
rect 16408 37108 16436 37275
rect 17126 37244 17132 37256
rect 17087 37216 17132 37244
rect 17126 37204 17132 37216
rect 17184 37204 17190 37256
rect 17420 37188 17448 37284
rect 17402 37136 17408 37188
rect 17460 37136 17466 37188
rect 18046 37108 18052 37120
rect 16408 37080 18052 37108
rect 18046 37068 18052 37080
rect 18104 37068 18110 37120
rect 1104 37018 18860 37040
rect 1104 36966 4315 37018
rect 4367 36966 4379 37018
rect 4431 36966 4443 37018
rect 4495 36966 4507 37018
rect 4559 36966 10982 37018
rect 11034 36966 11046 37018
rect 11098 36966 11110 37018
rect 11162 36966 11174 37018
rect 11226 36966 17648 37018
rect 17700 36966 17712 37018
rect 17764 36966 17776 37018
rect 17828 36966 17840 37018
rect 17892 36966 18860 37018
rect 1104 36944 18860 36966
rect 4433 36907 4491 36913
rect 4433 36873 4445 36907
rect 4479 36904 4491 36907
rect 4890 36904 4896 36916
rect 4479 36876 4896 36904
rect 4479 36873 4491 36876
rect 4433 36867 4491 36873
rect 4890 36864 4896 36876
rect 4948 36864 4954 36916
rect 6270 36904 6276 36916
rect 5092 36876 6276 36904
rect 3697 36839 3755 36845
rect 3697 36805 3709 36839
rect 3743 36836 3755 36839
rect 3970 36836 3976 36848
rect 3743 36808 3976 36836
rect 3743 36805 3755 36808
rect 3697 36799 3755 36805
rect 3970 36796 3976 36808
rect 4028 36836 4034 36848
rect 4985 36839 5043 36845
rect 4985 36836 4997 36839
rect 4028 36808 4997 36836
rect 4028 36796 4034 36808
rect 4985 36805 4997 36808
rect 5031 36805 5043 36839
rect 4985 36799 5043 36805
rect 4801 36771 4859 36777
rect 4801 36737 4813 36771
rect 4847 36768 4859 36771
rect 5092 36768 5120 36876
rect 6270 36864 6276 36876
rect 6328 36864 6334 36916
rect 8294 36864 8300 36916
rect 8352 36904 8358 36916
rect 8481 36907 8539 36913
rect 8481 36904 8493 36907
rect 8352 36876 8493 36904
rect 8352 36864 8358 36876
rect 8481 36873 8493 36876
rect 8527 36873 8539 36907
rect 8481 36867 8539 36873
rect 8941 36907 8999 36913
rect 8941 36873 8953 36907
rect 8987 36904 8999 36907
rect 9306 36904 9312 36916
rect 8987 36876 9312 36904
rect 8987 36873 8999 36876
rect 8941 36867 8999 36873
rect 9306 36864 9312 36876
rect 9364 36864 9370 36916
rect 10226 36904 10232 36916
rect 10187 36876 10232 36904
rect 10226 36864 10232 36876
rect 10284 36864 10290 36916
rect 10502 36864 10508 36916
rect 10560 36864 10566 36916
rect 10870 36904 10876 36916
rect 10831 36876 10876 36904
rect 10870 36864 10876 36876
rect 10928 36864 10934 36916
rect 12161 36907 12219 36913
rect 12161 36873 12173 36907
rect 12207 36904 12219 36907
rect 12342 36904 12348 36916
rect 12207 36876 12348 36904
rect 12207 36873 12219 36876
rect 12161 36867 12219 36873
rect 12342 36864 12348 36876
rect 12400 36864 12406 36916
rect 12802 36904 12808 36916
rect 12763 36876 12808 36904
rect 12802 36864 12808 36876
rect 12860 36864 12866 36916
rect 13541 36907 13599 36913
rect 13541 36873 13553 36907
rect 13587 36904 13599 36907
rect 13630 36904 13636 36916
rect 13587 36876 13636 36904
rect 13587 36873 13599 36876
rect 13541 36867 13599 36873
rect 13630 36864 13636 36876
rect 13688 36864 13694 36916
rect 14550 36864 14556 36916
rect 14608 36904 14614 36916
rect 15013 36907 15071 36913
rect 15013 36904 15025 36907
rect 14608 36876 15025 36904
rect 14608 36864 14614 36876
rect 15013 36873 15025 36876
rect 15059 36873 15071 36907
rect 15013 36867 15071 36873
rect 15194 36864 15200 36916
rect 15252 36904 15258 36916
rect 15473 36907 15531 36913
rect 15473 36904 15485 36907
rect 15252 36876 15485 36904
rect 15252 36864 15258 36876
rect 15473 36873 15485 36876
rect 15519 36873 15531 36907
rect 18046 36904 18052 36916
rect 18007 36876 18052 36904
rect 15473 36867 15531 36873
rect 18046 36864 18052 36876
rect 18104 36864 18110 36916
rect 5626 36836 5632 36848
rect 5539 36808 5632 36836
rect 4847 36740 5120 36768
rect 4847 36737 4859 36740
rect 4801 36731 4859 36737
rect 5169 36703 5227 36709
rect 5169 36669 5181 36703
rect 5215 36700 5227 36703
rect 5258 36700 5264 36712
rect 5215 36672 5264 36700
rect 5215 36669 5227 36672
rect 5169 36663 5227 36669
rect 5258 36660 5264 36672
rect 5316 36660 5322 36712
rect 5552 36709 5580 36808
rect 5626 36796 5632 36808
rect 5684 36836 5690 36848
rect 5684 36808 5764 36836
rect 5684 36796 5690 36808
rect 5736 36768 5764 36808
rect 5902 36796 5908 36848
rect 5960 36836 5966 36848
rect 6178 36836 6184 36848
rect 5960 36808 6184 36836
rect 5960 36796 5966 36808
rect 6178 36796 6184 36808
rect 6236 36796 6242 36848
rect 9122 36796 9128 36848
rect 9180 36836 9186 36848
rect 9217 36839 9275 36845
rect 9217 36836 9229 36839
rect 9180 36808 9229 36836
rect 9180 36796 9186 36808
rect 9217 36805 9229 36808
rect 9263 36805 9275 36839
rect 9217 36799 9275 36805
rect 9953 36839 10011 36845
rect 9953 36805 9965 36839
rect 9999 36836 10011 36839
rect 10134 36836 10140 36848
rect 9999 36808 10140 36836
rect 9999 36805 10011 36808
rect 9953 36799 10011 36805
rect 10134 36796 10140 36808
rect 10192 36796 10198 36848
rect 10520 36836 10548 36864
rect 10244 36808 10548 36836
rect 12529 36839 12587 36845
rect 10244 36780 10272 36808
rect 12529 36805 12541 36839
rect 12575 36836 12587 36839
rect 12894 36836 12900 36848
rect 12575 36808 12900 36836
rect 12575 36805 12587 36808
rect 12529 36799 12587 36805
rect 12894 36796 12900 36808
rect 12952 36796 12958 36848
rect 7193 36771 7251 36777
rect 7193 36768 7205 36771
rect 5736 36740 7205 36768
rect 7193 36737 7205 36740
rect 7239 36737 7251 36771
rect 7193 36731 7251 36737
rect 10226 36728 10232 36780
rect 10284 36728 10290 36780
rect 13648 36777 13676 36864
rect 14461 36839 14519 36845
rect 14461 36805 14473 36839
rect 14507 36836 14519 36839
rect 14737 36839 14795 36845
rect 14737 36836 14749 36839
rect 14507 36808 14749 36836
rect 14507 36805 14519 36808
rect 14461 36799 14519 36805
rect 14737 36805 14749 36808
rect 14783 36836 14795 36839
rect 15286 36836 15292 36848
rect 14783 36808 15292 36836
rect 14783 36805 14795 36808
rect 14737 36799 14795 36805
rect 15286 36796 15292 36808
rect 15344 36796 15350 36848
rect 16482 36796 16488 36848
rect 16540 36836 16546 36848
rect 16758 36836 16764 36848
rect 16540 36808 16764 36836
rect 16540 36796 16546 36808
rect 16758 36796 16764 36808
rect 16816 36796 16822 36848
rect 17402 36796 17408 36848
rect 17460 36796 17466 36848
rect 13633 36771 13691 36777
rect 13633 36737 13645 36771
rect 13679 36737 13691 36771
rect 13633 36731 13691 36737
rect 13998 36728 14004 36780
rect 14056 36768 14062 36780
rect 14369 36771 14427 36777
rect 14369 36768 14381 36771
rect 14056 36740 14381 36768
rect 14056 36728 14062 36740
rect 14369 36737 14381 36740
rect 14415 36737 14427 36771
rect 14369 36731 14427 36737
rect 16390 36728 16396 36780
rect 16448 36768 16454 36780
rect 17420 36768 17448 36796
rect 16448 36740 17540 36768
rect 16448 36728 16454 36740
rect 5537 36703 5595 36709
rect 5537 36669 5549 36703
rect 5583 36669 5595 36703
rect 5537 36663 5595 36669
rect 5721 36703 5779 36709
rect 5721 36669 5733 36703
rect 5767 36669 5779 36703
rect 6270 36700 6276 36712
rect 6231 36672 6276 36700
rect 5721 36663 5779 36669
rect 5736 36632 5764 36663
rect 6270 36660 6276 36672
rect 6328 36660 6334 36712
rect 7466 36700 7472 36712
rect 7024 36672 7472 36700
rect 4908 36604 5764 36632
rect 4908 36576 4936 36604
rect 7024 36576 7052 36672
rect 7466 36660 7472 36672
rect 7524 36700 7530 36712
rect 7653 36703 7711 36709
rect 7653 36700 7665 36703
rect 7524 36672 7665 36700
rect 7524 36660 7530 36672
rect 7653 36669 7665 36672
rect 7699 36669 7711 36703
rect 7653 36663 7711 36669
rect 7926 36660 7932 36712
rect 7984 36709 7990 36712
rect 7984 36703 8033 36709
rect 7984 36669 7987 36703
rect 8021 36669 8033 36703
rect 8110 36700 8116 36712
rect 8071 36672 8116 36700
rect 7984 36663 8033 36669
rect 7984 36660 7990 36663
rect 8110 36660 8116 36672
rect 8168 36660 8174 36712
rect 9950 36660 9956 36712
rect 10008 36700 10014 36712
rect 10134 36700 10140 36712
rect 10008 36672 10140 36700
rect 10008 36660 10014 36672
rect 10134 36660 10140 36672
rect 10192 36660 10198 36712
rect 10502 36660 10508 36712
rect 10560 36700 10566 36712
rect 10689 36703 10747 36709
rect 10689 36700 10701 36703
rect 10560 36672 10701 36700
rect 10560 36660 10566 36672
rect 10689 36669 10701 36672
rect 10735 36669 10747 36703
rect 10689 36663 10747 36669
rect 12434 36660 12440 36712
rect 12492 36700 12498 36712
rect 12621 36703 12679 36709
rect 12621 36700 12633 36703
rect 12492 36672 12633 36700
rect 12492 36660 12498 36672
rect 12621 36669 12633 36672
rect 12667 36700 12679 36703
rect 13081 36703 13139 36709
rect 13081 36700 13093 36703
rect 12667 36672 13093 36700
rect 12667 36669 12679 36672
rect 12621 36663 12679 36669
rect 13081 36669 13093 36672
rect 13127 36669 13139 36703
rect 14090 36700 14096 36712
rect 13081 36663 13139 36669
rect 13924 36672 14096 36700
rect 11514 36592 11520 36644
rect 11572 36632 11578 36644
rect 11974 36632 11980 36644
rect 11572 36604 11980 36632
rect 11572 36592 11578 36604
rect 11974 36592 11980 36604
rect 12032 36592 12038 36644
rect 12250 36592 12256 36644
rect 12308 36632 12314 36644
rect 13924 36641 13952 36672
rect 14090 36660 14096 36672
rect 14148 36700 14154 36712
rect 15289 36703 15347 36709
rect 15289 36700 15301 36703
rect 14148 36672 15301 36700
rect 14148 36660 14154 36672
rect 15289 36669 15301 36672
rect 15335 36700 15347 36703
rect 15749 36703 15807 36709
rect 15749 36700 15761 36703
rect 15335 36672 15761 36700
rect 15335 36669 15347 36672
rect 15289 36663 15347 36669
rect 15749 36669 15761 36672
rect 15795 36700 15807 36703
rect 15838 36700 15844 36712
rect 15795 36672 15844 36700
rect 15795 36669 15807 36672
rect 15749 36663 15807 36669
rect 15838 36660 15844 36672
rect 15896 36660 15902 36712
rect 16853 36703 16911 36709
rect 16853 36669 16865 36703
rect 16899 36669 16911 36703
rect 16853 36663 16911 36669
rect 17221 36703 17279 36709
rect 17221 36669 17233 36703
rect 17267 36700 17279 36703
rect 17402 36700 17408 36712
rect 17267 36672 17408 36700
rect 17267 36669 17279 36672
rect 17221 36663 17279 36669
rect 13909 36635 13967 36641
rect 13909 36632 13921 36635
rect 12308 36604 13921 36632
rect 12308 36592 12314 36604
rect 13909 36601 13921 36604
rect 13955 36601 13967 36635
rect 13909 36595 13967 36601
rect 14001 36635 14059 36641
rect 14001 36601 14013 36635
rect 14047 36632 14059 36635
rect 14461 36635 14519 36641
rect 14461 36632 14473 36635
rect 14047 36604 14473 36632
rect 14047 36601 14059 36604
rect 14001 36595 14059 36601
rect 14461 36601 14473 36604
rect 14507 36601 14519 36635
rect 16574 36632 16580 36644
rect 16487 36604 16580 36632
rect 14461 36595 14519 36601
rect 16574 36592 16580 36604
rect 16632 36632 16638 36644
rect 16868 36632 16896 36663
rect 17402 36660 17408 36672
rect 17460 36660 17466 36712
rect 17512 36709 17540 36740
rect 17497 36703 17555 36709
rect 17497 36669 17509 36703
rect 17543 36669 17555 36703
rect 17497 36663 17555 36669
rect 17678 36632 17684 36644
rect 16632 36604 17684 36632
rect 16632 36592 16638 36604
rect 17678 36592 17684 36604
rect 17736 36592 17742 36644
rect 17773 36635 17831 36641
rect 17773 36601 17785 36635
rect 17819 36632 17831 36635
rect 17862 36632 17868 36644
rect 17819 36604 17868 36632
rect 17819 36601 17831 36604
rect 17773 36595 17831 36601
rect 17862 36592 17868 36604
rect 17920 36592 17926 36644
rect 1673 36567 1731 36573
rect 1673 36533 1685 36567
rect 1719 36564 1731 36567
rect 1762 36564 1768 36576
rect 1719 36536 1768 36564
rect 1719 36533 1731 36536
rect 1673 36527 1731 36533
rect 1762 36524 1768 36536
rect 1820 36524 1826 36576
rect 3234 36564 3240 36576
rect 3195 36536 3240 36564
rect 3234 36524 3240 36536
rect 3292 36524 3298 36576
rect 4890 36524 4896 36576
rect 4948 36524 4954 36576
rect 5534 36524 5540 36576
rect 5592 36564 5598 36576
rect 5810 36564 5816 36576
rect 5592 36536 5816 36564
rect 5592 36524 5598 36536
rect 5810 36524 5816 36536
rect 5868 36524 5874 36576
rect 6270 36524 6276 36576
rect 6328 36564 6334 36576
rect 6641 36567 6699 36573
rect 6641 36564 6653 36567
rect 6328 36536 6653 36564
rect 6328 36524 6334 36536
rect 6641 36533 6653 36536
rect 6687 36564 6699 36567
rect 6822 36564 6828 36576
rect 6687 36536 6828 36564
rect 6687 36533 6699 36536
rect 6641 36527 6699 36533
rect 6822 36524 6828 36536
rect 6880 36524 6886 36576
rect 7006 36564 7012 36576
rect 6967 36536 7012 36564
rect 7006 36524 7012 36536
rect 7064 36524 7070 36576
rect 11330 36524 11336 36576
rect 11388 36564 11394 36576
rect 11609 36567 11667 36573
rect 11609 36564 11621 36567
rect 11388 36536 11621 36564
rect 11388 36524 11394 36536
rect 11609 36533 11621 36536
rect 11655 36533 11667 36567
rect 11609 36527 11667 36533
rect 13817 36567 13875 36573
rect 13817 36533 13829 36567
rect 13863 36564 13875 36567
rect 14918 36564 14924 36576
rect 13863 36536 14924 36564
rect 13863 36533 13875 36536
rect 13817 36527 13875 36533
rect 14918 36524 14924 36536
rect 14976 36524 14982 36576
rect 16114 36564 16120 36576
rect 16075 36536 16120 36564
rect 16114 36524 16120 36536
rect 16172 36524 16178 36576
rect 1104 36474 18860 36496
rect 1104 36422 7648 36474
rect 7700 36422 7712 36474
rect 7764 36422 7776 36474
rect 7828 36422 7840 36474
rect 7892 36422 14315 36474
rect 14367 36422 14379 36474
rect 14431 36422 14443 36474
rect 14495 36422 14507 36474
rect 14559 36422 18860 36474
rect 1104 36400 18860 36422
rect 4801 36363 4859 36369
rect 4801 36329 4813 36363
rect 4847 36360 4859 36363
rect 5258 36360 5264 36372
rect 4847 36332 5264 36360
rect 4847 36329 4859 36332
rect 4801 36323 4859 36329
rect 5258 36320 5264 36332
rect 5316 36320 5322 36372
rect 6641 36363 6699 36369
rect 6641 36329 6653 36363
rect 6687 36360 6699 36363
rect 6730 36360 6736 36372
rect 6687 36332 6736 36360
rect 6687 36329 6699 36332
rect 6641 36323 6699 36329
rect 6730 36320 6736 36332
rect 6788 36320 6794 36372
rect 8573 36363 8631 36369
rect 8573 36329 8585 36363
rect 8619 36360 8631 36363
rect 8754 36360 8760 36372
rect 8619 36332 8760 36360
rect 8619 36329 8631 36332
rect 8573 36323 8631 36329
rect 8754 36320 8760 36332
rect 8812 36320 8818 36372
rect 9306 36360 9312 36372
rect 9267 36332 9312 36360
rect 9306 36320 9312 36332
rect 9364 36320 9370 36372
rect 10502 36320 10508 36372
rect 10560 36360 10566 36372
rect 10597 36363 10655 36369
rect 10597 36360 10609 36363
rect 10560 36332 10609 36360
rect 10560 36320 10566 36332
rect 10597 36329 10609 36332
rect 10643 36360 10655 36363
rect 10870 36360 10876 36372
rect 10643 36332 10876 36360
rect 10643 36329 10655 36332
rect 10597 36323 10655 36329
rect 10870 36320 10876 36332
rect 10928 36320 10934 36372
rect 12158 36360 12164 36372
rect 12119 36332 12164 36360
rect 12158 36320 12164 36332
rect 12216 36320 12222 36372
rect 12710 36360 12716 36372
rect 12671 36332 12716 36360
rect 12710 36320 12716 36332
rect 12768 36320 12774 36372
rect 13446 36360 13452 36372
rect 13407 36332 13452 36360
rect 13446 36320 13452 36332
rect 13504 36320 13510 36372
rect 14090 36360 14096 36372
rect 14051 36332 14096 36360
rect 14090 36320 14096 36332
rect 14148 36320 14154 36372
rect 14461 36363 14519 36369
rect 14461 36329 14473 36363
rect 14507 36360 14519 36363
rect 14642 36360 14648 36372
rect 14507 36332 14648 36360
rect 14507 36329 14519 36332
rect 14461 36323 14519 36329
rect 14642 36320 14648 36332
rect 14700 36360 14706 36372
rect 15194 36360 15200 36372
rect 14700 36332 15200 36360
rect 14700 36320 14706 36332
rect 15194 36320 15200 36332
rect 15252 36320 15258 36372
rect 16390 36360 16396 36372
rect 16351 36332 16396 36360
rect 16390 36320 16396 36332
rect 16448 36320 16454 36372
rect 16574 36320 16580 36372
rect 16632 36360 16638 36372
rect 17037 36363 17095 36369
rect 17037 36360 17049 36363
rect 16632 36332 17049 36360
rect 16632 36320 16638 36332
rect 17037 36329 17049 36332
rect 17083 36329 17095 36363
rect 17402 36360 17408 36372
rect 17363 36332 17408 36360
rect 17037 36323 17095 36329
rect 17402 36320 17408 36332
rect 17460 36320 17466 36372
rect 4890 36292 4896 36304
rect 4851 36264 4896 36292
rect 4890 36252 4896 36264
rect 4948 36252 4954 36304
rect 6273 36295 6331 36301
rect 6273 36261 6285 36295
rect 6319 36292 6331 36295
rect 8021 36295 8079 36301
rect 8021 36292 8033 36295
rect 6319 36264 8033 36292
rect 6319 36261 6331 36264
rect 6273 36255 6331 36261
rect 8021 36261 8033 36264
rect 8067 36292 8079 36295
rect 8110 36292 8116 36304
rect 8067 36264 8116 36292
rect 8067 36261 8079 36264
rect 8021 36255 8079 36261
rect 8110 36252 8116 36264
rect 8168 36252 8174 36304
rect 11517 36295 11575 36301
rect 11517 36261 11529 36295
rect 11563 36292 11575 36295
rect 11790 36292 11796 36304
rect 11563 36264 11796 36292
rect 11563 36261 11575 36264
rect 11517 36255 11575 36261
rect 11790 36252 11796 36264
rect 11848 36252 11854 36304
rect 12802 36252 12808 36304
rect 12860 36292 12866 36304
rect 14550 36292 14556 36304
rect 12860 36264 14556 36292
rect 12860 36252 12866 36264
rect 14550 36252 14556 36264
rect 14608 36292 14614 36304
rect 16482 36292 16488 36304
rect 14608 36264 16488 36292
rect 14608 36252 14614 36264
rect 5350 36224 5356 36236
rect 5311 36196 5356 36224
rect 5350 36184 5356 36196
rect 5408 36184 5414 36236
rect 7009 36227 7067 36233
rect 7009 36193 7021 36227
rect 7055 36193 7067 36227
rect 7190 36224 7196 36236
rect 7151 36196 7196 36224
rect 7009 36187 7067 36193
rect 7024 36156 7052 36187
rect 7190 36184 7196 36196
rect 7248 36184 7254 36236
rect 7282 36184 7288 36236
rect 7340 36224 7346 36236
rect 7561 36227 7619 36233
rect 7561 36224 7573 36227
rect 7340 36196 7573 36224
rect 7340 36184 7346 36196
rect 7561 36193 7573 36196
rect 7607 36193 7619 36227
rect 9214 36224 9220 36236
rect 9175 36196 9220 36224
rect 7561 36187 7619 36193
rect 9214 36184 9220 36196
rect 9272 36184 9278 36236
rect 11330 36224 11336 36236
rect 11291 36196 11336 36224
rect 11330 36184 11336 36196
rect 11388 36184 11394 36236
rect 13078 36224 13084 36236
rect 13039 36196 13084 36224
rect 13078 36184 13084 36196
rect 13136 36184 13142 36236
rect 14734 36224 14740 36236
rect 14695 36196 14740 36224
rect 14734 36184 14740 36196
rect 14792 36184 14798 36236
rect 14918 36224 14924 36236
rect 14879 36196 14924 36224
rect 14918 36184 14924 36196
rect 14976 36184 14982 36236
rect 15304 36233 15332 36264
rect 16482 36252 16488 36264
rect 16540 36292 16546 36304
rect 16540 36264 16896 36292
rect 16540 36252 16546 36264
rect 16868 36233 16896 36264
rect 15289 36227 15347 36233
rect 15289 36193 15301 36227
rect 15335 36193 15347 36227
rect 15289 36187 15347 36193
rect 16025 36227 16083 36233
rect 16025 36193 16037 36227
rect 16071 36193 16083 36227
rect 16025 36187 16083 36193
rect 16853 36227 16911 36233
rect 16853 36193 16865 36227
rect 16899 36193 16911 36227
rect 16853 36187 16911 36193
rect 8294 36156 8300 36168
rect 7024 36128 8300 36156
rect 8294 36116 8300 36128
rect 8352 36116 8358 36168
rect 14274 36116 14280 36168
rect 14332 36156 14338 36168
rect 16040 36156 16068 36187
rect 17954 36184 17960 36236
rect 18012 36184 18018 36236
rect 16390 36156 16396 36168
rect 14332 36128 16396 36156
rect 14332 36116 14338 36128
rect 16390 36116 16396 36128
rect 16448 36156 16454 36168
rect 17972 36156 18000 36184
rect 16448 36128 18000 36156
rect 16448 36116 16454 36128
rect 1673 36023 1731 36029
rect 1673 35989 1685 36023
rect 1719 36020 1731 36023
rect 1854 36020 1860 36032
rect 1719 35992 1860 36020
rect 1719 35989 1731 35992
rect 1673 35983 1731 35989
rect 1854 35980 1860 35992
rect 1912 35980 1918 36032
rect 2038 35980 2044 36032
rect 2096 36020 2102 36032
rect 2314 36020 2320 36032
rect 2096 35992 2320 36020
rect 2096 35980 2102 35992
rect 2314 35980 2320 35992
rect 2372 35980 2378 36032
rect 5902 35980 5908 36032
rect 5960 36020 5966 36032
rect 6454 36020 6460 36032
rect 5960 35992 6460 36020
rect 5960 35980 5966 35992
rect 6454 35980 6460 35992
rect 6512 35980 6518 36032
rect 15933 36023 15991 36029
rect 15933 35989 15945 36023
rect 15979 36020 15991 36023
rect 16574 36020 16580 36032
rect 15979 35992 16580 36020
rect 15979 35989 15991 35992
rect 15933 35983 15991 35989
rect 16574 35980 16580 35992
rect 16632 36020 16638 36032
rect 16669 36023 16727 36029
rect 16669 36020 16681 36023
rect 16632 35992 16681 36020
rect 16632 35980 16638 35992
rect 16669 35989 16681 35992
rect 16715 35989 16727 36023
rect 16669 35983 16727 35989
rect 1104 35930 18860 35952
rect 1104 35878 4315 35930
rect 4367 35878 4379 35930
rect 4431 35878 4443 35930
rect 4495 35878 4507 35930
rect 4559 35878 10982 35930
rect 11034 35878 11046 35930
rect 11098 35878 11110 35930
rect 11162 35878 11174 35930
rect 11226 35878 17648 35930
rect 17700 35878 17712 35930
rect 17764 35878 17776 35930
rect 17828 35878 17840 35930
rect 17892 35878 18860 35930
rect 1104 35856 18860 35878
rect 3053 35819 3111 35825
rect 3053 35785 3065 35819
rect 3099 35816 3111 35819
rect 3878 35816 3884 35828
rect 3099 35788 3884 35816
rect 3099 35785 3111 35788
rect 3053 35779 3111 35785
rect 3878 35776 3884 35788
rect 3936 35776 3942 35828
rect 4985 35819 5043 35825
rect 4985 35785 4997 35819
rect 5031 35816 5043 35819
rect 5350 35816 5356 35828
rect 5031 35788 5356 35816
rect 5031 35785 5043 35788
rect 4985 35779 5043 35785
rect 5350 35776 5356 35788
rect 5408 35776 5414 35828
rect 6362 35816 6368 35828
rect 6323 35788 6368 35816
rect 6362 35776 6368 35788
rect 6420 35776 6426 35828
rect 7282 35776 7288 35828
rect 7340 35816 7346 35828
rect 7469 35819 7527 35825
rect 7469 35816 7481 35819
rect 7340 35788 7481 35816
rect 7340 35776 7346 35788
rect 7469 35785 7481 35788
rect 7515 35785 7527 35819
rect 7469 35779 7527 35785
rect 7837 35819 7895 35825
rect 7837 35785 7849 35819
rect 7883 35816 7895 35819
rect 8478 35816 8484 35828
rect 7883 35788 8484 35816
rect 7883 35785 7895 35788
rect 7837 35779 7895 35785
rect 8478 35776 8484 35788
rect 8536 35776 8542 35828
rect 8941 35819 8999 35825
rect 8941 35785 8953 35819
rect 8987 35816 8999 35819
rect 9214 35816 9220 35828
rect 8987 35788 9220 35816
rect 8987 35785 8999 35788
rect 8941 35779 8999 35785
rect 9214 35776 9220 35788
rect 9272 35776 9278 35828
rect 9309 35819 9367 35825
rect 9309 35785 9321 35819
rect 9355 35816 9367 35819
rect 9582 35816 9588 35828
rect 9355 35788 9588 35816
rect 9355 35785 9367 35788
rect 9309 35779 9367 35785
rect 9582 35776 9588 35788
rect 9640 35776 9646 35828
rect 10505 35819 10563 35825
rect 10505 35785 10517 35819
rect 10551 35816 10563 35819
rect 11057 35819 11115 35825
rect 11057 35816 11069 35819
rect 10551 35788 11069 35816
rect 10551 35785 10563 35788
rect 10505 35779 10563 35785
rect 11057 35785 11069 35788
rect 11103 35816 11115 35819
rect 11330 35816 11336 35828
rect 11103 35788 11336 35816
rect 11103 35785 11115 35788
rect 11057 35779 11115 35785
rect 11330 35776 11336 35788
rect 11388 35776 11394 35828
rect 12526 35816 12532 35828
rect 12487 35788 12532 35816
rect 12526 35776 12532 35788
rect 12584 35776 12590 35828
rect 13078 35816 13084 35828
rect 13039 35788 13084 35816
rect 13078 35776 13084 35788
rect 13136 35776 13142 35828
rect 14093 35819 14151 35825
rect 14093 35785 14105 35819
rect 14139 35816 14151 35819
rect 14274 35816 14280 35828
rect 14139 35788 14280 35816
rect 14139 35785 14151 35788
rect 14093 35779 14151 35785
rect 14274 35776 14280 35788
rect 14332 35776 14338 35828
rect 14737 35819 14795 35825
rect 14737 35785 14749 35819
rect 14783 35816 14795 35819
rect 14918 35816 14924 35828
rect 14783 35788 14924 35816
rect 14783 35785 14795 35788
rect 14737 35779 14795 35785
rect 14918 35776 14924 35788
rect 14976 35776 14982 35828
rect 15565 35819 15623 35825
rect 15565 35785 15577 35819
rect 15611 35816 15623 35819
rect 15654 35816 15660 35828
rect 15611 35788 15660 35816
rect 15611 35785 15623 35788
rect 15565 35779 15623 35785
rect 15654 35776 15660 35788
rect 15712 35776 15718 35828
rect 15838 35816 15844 35828
rect 15799 35788 15844 35816
rect 15838 35776 15844 35788
rect 15896 35776 15902 35828
rect 16482 35776 16488 35828
rect 16540 35816 16546 35828
rect 16577 35819 16635 35825
rect 16577 35816 16589 35819
rect 16540 35788 16589 35816
rect 16540 35776 16546 35788
rect 16577 35785 16589 35788
rect 16623 35785 16635 35819
rect 18138 35816 18144 35828
rect 18099 35788 18144 35816
rect 16577 35779 16635 35785
rect 18138 35776 18144 35788
rect 18196 35776 18202 35828
rect 8294 35708 8300 35760
rect 8352 35748 8358 35760
rect 8573 35751 8631 35757
rect 8573 35748 8585 35751
rect 8352 35720 8585 35748
rect 8352 35708 8358 35720
rect 8573 35717 8585 35720
rect 8619 35748 8631 35751
rect 9398 35748 9404 35760
rect 8619 35720 9404 35748
rect 8619 35717 8631 35720
rect 8573 35711 8631 35717
rect 9398 35708 9404 35720
rect 9456 35708 9462 35760
rect 10137 35751 10195 35757
rect 10137 35717 10149 35751
rect 10183 35717 10195 35751
rect 10137 35711 10195 35717
rect 1489 35683 1547 35689
rect 1489 35649 1501 35683
rect 1535 35680 1547 35683
rect 1854 35680 1860 35692
rect 1535 35652 1860 35680
rect 1535 35649 1547 35652
rect 1489 35643 1547 35649
rect 1854 35640 1860 35652
rect 1912 35680 1918 35692
rect 2498 35680 2504 35692
rect 1912 35652 2504 35680
rect 1912 35640 1918 35652
rect 2498 35640 2504 35652
rect 2556 35640 2562 35692
rect 1578 35572 1584 35624
rect 1636 35612 1642 35624
rect 1765 35615 1823 35621
rect 1765 35612 1777 35615
rect 1636 35584 1777 35612
rect 1636 35572 1642 35584
rect 1765 35581 1777 35584
rect 1811 35581 1823 35615
rect 1765 35575 1823 35581
rect 5997 35615 6055 35621
rect 5997 35581 6009 35615
rect 6043 35612 6055 35615
rect 6733 35615 6791 35621
rect 6733 35612 6745 35615
rect 6043 35584 6745 35612
rect 6043 35581 6055 35584
rect 5997 35575 6055 35581
rect 6733 35581 6745 35584
rect 6779 35612 6791 35615
rect 6822 35612 6828 35624
rect 6779 35584 6828 35612
rect 6779 35581 6791 35584
rect 6733 35575 6791 35581
rect 6822 35572 6828 35584
rect 6880 35572 6886 35624
rect 7653 35615 7711 35621
rect 7653 35612 7665 35615
rect 7208 35584 7665 35612
rect 7208 35488 7236 35584
rect 7653 35581 7665 35584
rect 7699 35612 7711 35615
rect 8113 35615 8171 35621
rect 8113 35612 8125 35615
rect 7699 35584 8125 35612
rect 7699 35581 7711 35584
rect 7653 35575 7711 35581
rect 8113 35581 8125 35584
rect 8159 35581 8171 35615
rect 9950 35612 9956 35624
rect 9911 35584 9956 35612
rect 8113 35575 8171 35581
rect 9950 35572 9956 35584
rect 10008 35572 10014 35624
rect 10152 35612 10180 35711
rect 12158 35708 12164 35760
rect 12216 35748 12222 35760
rect 13538 35748 13544 35760
rect 12216 35720 13544 35748
rect 12216 35708 12222 35720
rect 13538 35708 13544 35720
rect 13596 35708 13602 35760
rect 14369 35751 14427 35757
rect 14369 35717 14381 35751
rect 14415 35748 14427 35751
rect 15286 35748 15292 35760
rect 14415 35720 15292 35748
rect 14415 35717 14427 35720
rect 14369 35711 14427 35717
rect 15286 35708 15292 35720
rect 15344 35708 15350 35760
rect 17494 35748 17500 35760
rect 17455 35720 17500 35748
rect 17494 35708 17500 35720
rect 17552 35708 17558 35760
rect 12342 35640 12348 35692
rect 12400 35680 12406 35692
rect 18156 35680 18184 35776
rect 12400 35652 14228 35680
rect 12400 35640 12406 35652
rect 14200 35624 14228 35652
rect 17236 35652 18184 35680
rect 10873 35615 10931 35621
rect 10873 35612 10885 35615
rect 10152 35584 10885 35612
rect 10873 35581 10885 35584
rect 10919 35612 10931 35615
rect 11241 35615 11299 35621
rect 11241 35612 11253 35615
rect 10919 35584 11253 35612
rect 10919 35581 10931 35584
rect 10873 35575 10931 35581
rect 11241 35581 11253 35584
rect 11287 35612 11299 35615
rect 11422 35612 11428 35624
rect 11287 35584 11428 35612
rect 11287 35581 11299 35584
rect 11241 35575 11299 35581
rect 11422 35572 11428 35584
rect 11480 35572 11486 35624
rect 11701 35615 11759 35621
rect 11701 35581 11713 35615
rect 11747 35612 11759 35615
rect 11790 35612 11796 35624
rect 11747 35584 11796 35612
rect 11747 35581 11759 35584
rect 11701 35575 11759 35581
rect 11790 35572 11796 35584
rect 11848 35612 11854 35624
rect 11974 35612 11980 35624
rect 11848 35584 11980 35612
rect 11848 35572 11854 35584
rect 11974 35572 11980 35584
rect 12032 35572 12038 35624
rect 13173 35615 13231 35621
rect 13173 35581 13185 35615
rect 13219 35612 13231 35615
rect 14182 35612 14188 35624
rect 13219 35584 13768 35612
rect 14095 35584 14188 35612
rect 13219 35581 13231 35584
rect 13173 35575 13231 35581
rect 13740 35488 13768 35584
rect 14182 35572 14188 35584
rect 14240 35572 14246 35624
rect 15381 35615 15439 35621
rect 15381 35581 15393 35615
rect 15427 35612 15439 35615
rect 15838 35612 15844 35624
rect 15427 35584 15844 35612
rect 15427 35581 15439 35584
rect 15381 35575 15439 35581
rect 15838 35572 15844 35584
rect 15896 35572 15902 35624
rect 16574 35572 16580 35624
rect 16632 35612 16638 35624
rect 17236 35621 17264 35652
rect 16669 35615 16727 35621
rect 16669 35612 16681 35615
rect 16632 35584 16681 35612
rect 16632 35572 16638 35584
rect 16669 35581 16681 35584
rect 16715 35581 16727 35615
rect 16669 35575 16727 35581
rect 17221 35615 17279 35621
rect 17221 35581 17233 35615
rect 17267 35581 17279 35615
rect 17221 35575 17279 35581
rect 17589 35615 17647 35621
rect 17589 35581 17601 35615
rect 17635 35612 17647 35615
rect 18417 35615 18475 35621
rect 18417 35612 18429 35615
rect 17635 35584 18429 35612
rect 17635 35581 17647 35584
rect 17589 35575 17647 35581
rect 18417 35581 18429 35584
rect 18463 35581 18475 35615
rect 18417 35575 18475 35581
rect 14550 35504 14556 35556
rect 14608 35544 14614 35556
rect 14918 35544 14924 35556
rect 14608 35516 14924 35544
rect 14608 35504 14614 35516
rect 14918 35504 14924 35516
rect 14976 35504 14982 35556
rect 15930 35504 15936 35556
rect 15988 35544 15994 35556
rect 17604 35544 17632 35575
rect 15988 35516 17632 35544
rect 15988 35504 15994 35516
rect 5718 35436 5724 35488
rect 5776 35476 5782 35488
rect 5994 35476 6000 35488
rect 5776 35448 6000 35476
rect 5776 35436 5782 35448
rect 5994 35436 6000 35448
rect 6052 35436 6058 35488
rect 7190 35476 7196 35488
rect 7151 35448 7196 35476
rect 7190 35436 7196 35448
rect 7248 35436 7254 35488
rect 13262 35436 13268 35488
rect 13320 35476 13326 35488
rect 13357 35479 13415 35485
rect 13357 35476 13369 35479
rect 13320 35448 13369 35476
rect 13320 35436 13326 35448
rect 13357 35445 13369 35448
rect 13403 35476 13415 35479
rect 13538 35476 13544 35488
rect 13403 35448 13544 35476
rect 13403 35445 13415 35448
rect 13357 35439 13415 35445
rect 13538 35436 13544 35448
rect 13596 35436 13602 35488
rect 13722 35476 13728 35488
rect 13683 35448 13728 35476
rect 13722 35436 13728 35448
rect 13780 35436 13786 35488
rect 14734 35436 14740 35488
rect 14792 35476 14798 35488
rect 15013 35479 15071 35485
rect 15013 35476 15025 35479
rect 14792 35448 15025 35476
rect 14792 35436 14798 35448
rect 15013 35445 15025 35448
rect 15059 35445 15071 35479
rect 15013 35439 15071 35445
rect 1104 35386 18860 35408
rect 1104 35334 7648 35386
rect 7700 35334 7712 35386
rect 7764 35334 7776 35386
rect 7828 35334 7840 35386
rect 7892 35334 14315 35386
rect 14367 35334 14379 35386
rect 14431 35334 14443 35386
rect 14495 35334 14507 35386
rect 14559 35334 18860 35386
rect 1104 35312 18860 35334
rect 5997 35275 6055 35281
rect 5997 35241 6009 35275
rect 6043 35272 6055 35275
rect 6178 35272 6184 35284
rect 6043 35244 6184 35272
rect 6043 35241 6055 35244
rect 5997 35235 6055 35241
rect 6178 35232 6184 35244
rect 6236 35232 6242 35284
rect 14182 35272 14188 35284
rect 14143 35244 14188 35272
rect 14182 35232 14188 35244
rect 14240 35232 14246 35284
rect 14645 35275 14703 35281
rect 14645 35241 14657 35275
rect 14691 35272 14703 35275
rect 14918 35272 14924 35284
rect 14691 35244 14924 35272
rect 14691 35241 14703 35244
rect 14645 35235 14703 35241
rect 14918 35232 14924 35244
rect 14976 35232 14982 35284
rect 17402 35272 17408 35284
rect 17363 35244 17408 35272
rect 17402 35232 17408 35244
rect 17460 35232 17466 35284
rect 2314 35164 2320 35216
rect 2372 35164 2378 35216
rect 6012 35176 7558 35204
rect 2332 35136 2360 35164
rect 6012 35148 6040 35176
rect 2593 35139 2651 35145
rect 2593 35136 2605 35139
rect 2332 35108 2605 35136
rect 2593 35105 2605 35108
rect 2639 35105 2651 35139
rect 2593 35099 2651 35105
rect 5994 35096 6000 35148
rect 6052 35096 6058 35148
rect 6914 35096 6920 35148
rect 6972 35136 6978 35148
rect 7530 35145 7558 35176
rect 9674 35164 9680 35216
rect 9732 35204 9738 35216
rect 10597 35207 10655 35213
rect 10597 35204 10609 35207
rect 9732 35176 10609 35204
rect 9732 35164 9738 35176
rect 10597 35173 10609 35176
rect 10643 35173 10655 35207
rect 10597 35167 10655 35173
rect 13078 35164 13084 35216
rect 13136 35204 13142 35216
rect 17420 35204 17448 35232
rect 13136 35176 14780 35204
rect 13136 35164 13142 35176
rect 14752 35148 14780 35176
rect 16592 35176 17448 35204
rect 7377 35139 7435 35145
rect 7377 35136 7389 35139
rect 6972 35108 7389 35136
rect 6972 35096 6978 35108
rect 7377 35105 7389 35108
rect 7423 35105 7435 35139
rect 7377 35099 7435 35105
rect 7515 35139 7573 35145
rect 7515 35105 7527 35139
rect 7561 35105 7573 35139
rect 7515 35099 7573 35105
rect 7653 35139 7711 35145
rect 7653 35105 7665 35139
rect 7699 35136 7711 35139
rect 8478 35136 8484 35148
rect 7699 35108 8484 35136
rect 7699 35105 7711 35108
rect 7653 35099 7711 35105
rect 2317 35071 2375 35077
rect 2317 35037 2329 35071
rect 2363 35068 2375 35071
rect 2498 35068 2504 35080
rect 2363 35040 2504 35068
rect 2363 35037 2375 35040
rect 2317 35031 2375 35037
rect 2498 35028 2504 35040
rect 2556 35028 2562 35080
rect 3970 35068 3976 35080
rect 3931 35040 3976 35068
rect 3970 35028 3976 35040
rect 4028 35028 4034 35080
rect 6825 35071 6883 35077
rect 6825 35037 6837 35071
rect 6871 35068 6883 35071
rect 7282 35068 7288 35080
rect 6871 35040 7288 35068
rect 6871 35037 6883 35040
rect 6825 35031 6883 35037
rect 7282 35028 7288 35040
rect 7340 35028 7346 35080
rect 4433 35003 4491 35009
rect 4433 34969 4445 35003
rect 4479 35000 4491 35003
rect 4614 35000 4620 35012
rect 4479 34972 4620 35000
rect 4479 34969 4491 34972
rect 4433 34963 4491 34969
rect 4614 34960 4620 34972
rect 4672 35000 4678 35012
rect 7668 35000 7696 35099
rect 8478 35096 8484 35108
rect 8536 35096 8542 35148
rect 9950 35136 9956 35148
rect 9863 35108 9956 35136
rect 9950 35096 9956 35108
rect 10008 35136 10014 35148
rect 10689 35139 10747 35145
rect 10689 35136 10701 35139
rect 10008 35108 10701 35136
rect 10008 35096 10014 35108
rect 10689 35105 10701 35108
rect 10735 35105 10747 35139
rect 10689 35099 10747 35105
rect 13630 35096 13636 35148
rect 13688 35136 13694 35148
rect 13725 35139 13783 35145
rect 13725 35136 13737 35139
rect 13688 35108 13737 35136
rect 13688 35096 13694 35108
rect 13725 35105 13737 35108
rect 13771 35105 13783 35139
rect 14734 35136 14740 35148
rect 14647 35108 14740 35136
rect 13725 35099 13783 35105
rect 14734 35096 14740 35108
rect 14792 35096 14798 35148
rect 16206 35136 16212 35148
rect 16167 35108 16212 35136
rect 16206 35096 16212 35108
rect 16264 35096 16270 35148
rect 16482 35096 16488 35148
rect 16540 35136 16546 35148
rect 16592 35145 16620 35176
rect 16577 35139 16635 35145
rect 16577 35136 16589 35139
rect 16540 35108 16589 35136
rect 16540 35096 16546 35108
rect 16577 35105 16589 35108
rect 16623 35105 16635 35139
rect 16577 35099 16635 35105
rect 16853 35139 16911 35145
rect 16853 35105 16865 35139
rect 16899 35105 16911 35139
rect 16853 35099 16911 35105
rect 4672 34972 7696 35000
rect 4672 34960 4678 34972
rect 1578 34932 1584 34944
rect 1539 34904 1584 34932
rect 1578 34892 1584 34904
rect 1636 34892 1642 34944
rect 4801 34935 4859 34941
rect 4801 34901 4813 34935
rect 4847 34932 4859 34935
rect 5074 34932 5080 34944
rect 4847 34904 5080 34932
rect 4847 34901 4859 34904
rect 4801 34895 4859 34901
rect 5074 34892 5080 34904
rect 5132 34892 5138 34944
rect 6365 34935 6423 34941
rect 6365 34901 6377 34935
rect 6411 34932 6423 34935
rect 6730 34932 6736 34944
rect 6411 34904 6736 34932
rect 6411 34901 6423 34904
rect 6365 34895 6423 34901
rect 6730 34892 6736 34904
rect 6788 34892 6794 34944
rect 9766 34892 9772 34944
rect 9824 34932 9830 34944
rect 9968 34941 9996 35096
rect 15933 35071 15991 35077
rect 15933 35037 15945 35071
rect 15979 35068 15991 35071
rect 16298 35068 16304 35080
rect 15979 35040 16304 35068
rect 15979 35037 15991 35040
rect 15933 35031 15991 35037
rect 16298 35028 16304 35040
rect 16356 35068 16362 35080
rect 16868 35068 16896 35099
rect 17126 35068 17132 35080
rect 16356 35040 16896 35068
rect 17087 35040 17132 35068
rect 16356 35028 16362 35040
rect 17126 35028 17132 35040
rect 17184 35028 17190 35080
rect 13909 35003 13967 35009
rect 13909 34969 13921 35003
rect 13955 35000 13967 35003
rect 14642 35000 14648 35012
rect 13955 34972 14648 35000
rect 13955 34969 13967 34972
rect 13909 34963 13967 34969
rect 14642 34960 14648 34972
rect 14700 34960 14706 35012
rect 14921 35003 14979 35009
rect 14921 34969 14933 35003
rect 14967 35000 14979 35003
rect 16390 35000 16396 35012
rect 14967 34972 16396 35000
rect 14967 34969 14979 34972
rect 14921 34963 14979 34969
rect 15948 34944 15976 34972
rect 16390 34960 16396 34972
rect 16448 34960 16454 35012
rect 9953 34935 10011 34941
rect 9953 34932 9965 34935
rect 9824 34904 9965 34932
rect 9824 34892 9830 34904
rect 9953 34901 9965 34904
rect 9999 34901 10011 34935
rect 9953 34895 10011 34901
rect 15930 34892 15936 34944
rect 15988 34892 15994 34944
rect 1104 34842 18860 34864
rect 1104 34790 4315 34842
rect 4367 34790 4379 34842
rect 4431 34790 4443 34842
rect 4495 34790 4507 34842
rect 4559 34790 10982 34842
rect 11034 34790 11046 34842
rect 11098 34790 11110 34842
rect 11162 34790 11174 34842
rect 11226 34790 17648 34842
rect 17700 34790 17712 34842
rect 17764 34790 17776 34842
rect 17828 34790 17840 34842
rect 17892 34790 18860 34842
rect 1104 34768 18860 34790
rect 5813 34731 5871 34737
rect 5813 34697 5825 34731
rect 5859 34728 5871 34731
rect 5994 34728 6000 34740
rect 5859 34700 6000 34728
rect 5859 34697 5871 34700
rect 5813 34691 5871 34697
rect 5994 34688 6000 34700
rect 6052 34688 6058 34740
rect 6181 34731 6239 34737
rect 6181 34697 6193 34731
rect 6227 34728 6239 34731
rect 7926 34728 7932 34740
rect 6227 34700 7932 34728
rect 6227 34697 6239 34700
rect 6181 34691 6239 34697
rect 7926 34688 7932 34700
rect 7984 34688 7990 34740
rect 14734 34728 14740 34740
rect 14695 34700 14740 34728
rect 14734 34688 14740 34700
rect 14792 34688 14798 34740
rect 15562 34728 15568 34740
rect 15523 34700 15568 34728
rect 15562 34688 15568 34700
rect 15620 34688 15626 34740
rect 16206 34728 16212 34740
rect 16167 34700 16212 34728
rect 16206 34688 16212 34700
rect 16264 34688 16270 34740
rect 16298 34688 16304 34740
rect 16356 34688 16362 34740
rect 2314 34660 2320 34672
rect 2275 34632 2320 34660
rect 2314 34620 2320 34632
rect 2372 34620 2378 34672
rect 15286 34620 15292 34672
rect 15344 34660 15350 34672
rect 15841 34663 15899 34669
rect 15841 34660 15853 34663
rect 15344 34632 15853 34660
rect 15344 34620 15350 34632
rect 4525 34595 4583 34601
rect 4525 34561 4537 34595
rect 4571 34592 4583 34595
rect 4614 34592 4620 34604
rect 4571 34564 4620 34592
rect 4571 34561 4583 34564
rect 4525 34555 4583 34561
rect 4614 34552 4620 34564
rect 4672 34552 4678 34604
rect 4982 34592 4988 34604
rect 4895 34564 4988 34592
rect 1486 34484 1492 34536
rect 1544 34524 1550 34536
rect 2498 34524 2504 34536
rect 1544 34496 2504 34524
rect 1544 34484 1550 34496
rect 2498 34484 2504 34496
rect 2556 34524 2562 34536
rect 4908 34533 4936 34564
rect 4982 34552 4988 34564
rect 5040 34592 5046 34604
rect 5442 34592 5448 34604
rect 5040 34564 5304 34592
rect 5403 34564 5448 34592
rect 5040 34552 5046 34564
rect 2685 34527 2743 34533
rect 2685 34524 2697 34527
rect 2556 34496 2697 34524
rect 2556 34484 2562 34496
rect 2685 34493 2697 34496
rect 2731 34493 2743 34527
rect 2685 34487 2743 34493
rect 3881 34527 3939 34533
rect 3881 34493 3893 34527
rect 3927 34524 3939 34527
rect 4893 34527 4951 34533
rect 4893 34524 4905 34527
rect 3927 34496 4905 34524
rect 3927 34493 3939 34496
rect 3881 34487 3939 34493
rect 4893 34493 4905 34496
rect 4939 34493 4951 34527
rect 4893 34487 4951 34493
rect 5074 34484 5080 34536
rect 5132 34524 5138 34536
rect 5169 34527 5227 34533
rect 5169 34524 5181 34527
rect 5132 34496 5181 34524
rect 5132 34484 5138 34496
rect 5169 34493 5181 34496
rect 5215 34493 5227 34527
rect 5276 34524 5304 34564
rect 5442 34552 5448 34564
rect 5500 34552 5506 34604
rect 6178 34552 6184 34604
rect 6236 34592 6242 34604
rect 6236 34564 7512 34592
rect 6236 34552 6242 34564
rect 5276 34496 5580 34524
rect 5169 34487 5227 34493
rect 5552 34456 5580 34496
rect 5810 34484 5816 34536
rect 5868 34524 5874 34536
rect 6273 34527 6331 34533
rect 6273 34524 6285 34527
rect 5868 34496 6285 34524
rect 5868 34484 5874 34496
rect 6273 34493 6285 34496
rect 6319 34524 6331 34527
rect 6362 34524 6368 34536
rect 6319 34496 6368 34524
rect 6319 34493 6331 34496
rect 6273 34487 6331 34493
rect 6362 34484 6368 34496
rect 6420 34484 6426 34536
rect 6730 34524 6736 34536
rect 6691 34496 6736 34524
rect 6730 34484 6736 34496
rect 6788 34484 6794 34536
rect 7484 34533 7512 34564
rect 14642 34552 14648 34604
rect 14700 34592 14706 34604
rect 14918 34592 14924 34604
rect 14700 34564 14924 34592
rect 14700 34552 14706 34564
rect 14918 34552 14924 34564
rect 14976 34552 14982 34604
rect 7469 34527 7527 34533
rect 7469 34493 7481 34527
rect 7515 34493 7527 34527
rect 7926 34524 7932 34536
rect 7887 34496 7932 34524
rect 7469 34487 7527 34493
rect 7926 34484 7932 34496
rect 7984 34484 7990 34536
rect 8478 34524 8484 34536
rect 8391 34496 8484 34524
rect 8478 34484 8484 34496
rect 8536 34524 8542 34536
rect 8938 34524 8944 34536
rect 8536 34496 8944 34524
rect 8536 34484 8542 34496
rect 8938 34484 8944 34496
rect 8996 34484 9002 34536
rect 9766 34484 9772 34536
rect 9824 34524 9830 34536
rect 10597 34527 10655 34533
rect 10597 34524 10609 34527
rect 9824 34496 10609 34524
rect 9824 34484 9830 34496
rect 10597 34493 10609 34496
rect 10643 34493 10655 34527
rect 10597 34487 10655 34493
rect 13630 34484 13636 34536
rect 13688 34524 13694 34536
rect 13817 34527 13875 34533
rect 13817 34524 13829 34527
rect 13688 34496 13829 34524
rect 13688 34484 13694 34496
rect 13817 34493 13829 34496
rect 13863 34524 13875 34527
rect 14734 34524 14740 34536
rect 13863 34496 14740 34524
rect 13863 34493 13875 34496
rect 13817 34487 13875 34493
rect 14734 34484 14740 34496
rect 14792 34484 14798 34536
rect 15396 34533 15424 34632
rect 15841 34629 15853 34632
rect 15887 34629 15899 34663
rect 16316 34660 16344 34688
rect 17494 34660 17500 34672
rect 16316 34632 17356 34660
rect 17455 34632 17500 34660
rect 15841 34623 15899 34629
rect 16850 34592 16856 34604
rect 16811 34564 16856 34592
rect 16850 34552 16856 34564
rect 16908 34552 16914 34604
rect 17328 34592 17356 34632
rect 17494 34620 17500 34632
rect 17552 34620 17558 34672
rect 18049 34595 18107 34601
rect 18049 34592 18061 34595
rect 17328 34564 18061 34592
rect 15381 34527 15439 34533
rect 15381 34493 15393 34527
rect 15427 34493 15439 34527
rect 15381 34487 15439 34493
rect 17221 34527 17279 34533
rect 17221 34493 17233 34527
rect 17267 34524 17279 34527
rect 17402 34524 17408 34536
rect 17267 34496 17408 34524
rect 17267 34493 17279 34496
rect 17221 34487 17279 34493
rect 17402 34484 17408 34496
rect 17460 34484 17466 34536
rect 17512 34533 17540 34564
rect 18049 34561 18061 34564
rect 18095 34561 18107 34595
rect 18049 34555 18107 34561
rect 17497 34527 17555 34533
rect 17497 34493 17509 34527
rect 17543 34493 17555 34527
rect 17497 34487 17555 34493
rect 6822 34456 6828 34468
rect 5552 34428 6828 34456
rect 6822 34416 6828 34428
rect 6880 34416 6886 34468
rect 8294 34416 8300 34468
rect 8352 34456 8358 34468
rect 8570 34456 8576 34468
rect 8352 34428 8576 34456
rect 8352 34416 8358 34428
rect 8570 34416 8576 34428
rect 8628 34416 8634 34468
rect 7193 34391 7251 34397
rect 7193 34357 7205 34391
rect 7239 34388 7251 34391
rect 7466 34388 7472 34400
rect 7239 34360 7472 34388
rect 7239 34357 7251 34360
rect 7193 34351 7251 34357
rect 7466 34348 7472 34360
rect 7524 34348 7530 34400
rect 1104 34298 18860 34320
rect 1104 34246 7648 34298
rect 7700 34246 7712 34298
rect 7764 34246 7776 34298
rect 7828 34246 7840 34298
rect 7892 34246 14315 34298
rect 14367 34246 14379 34298
rect 14431 34246 14443 34298
rect 14495 34246 14507 34298
rect 14559 34246 18860 34298
rect 1104 34224 18860 34246
rect 5997 34187 6055 34193
rect 5997 34153 6009 34187
rect 6043 34184 6055 34187
rect 6914 34184 6920 34196
rect 6043 34156 6920 34184
rect 6043 34153 6055 34156
rect 5997 34147 6055 34153
rect 6914 34144 6920 34156
rect 6972 34144 6978 34196
rect 14185 34187 14243 34193
rect 14185 34153 14197 34187
rect 14231 34184 14243 34187
rect 14826 34184 14832 34196
rect 14231 34156 14832 34184
rect 14231 34153 14243 34156
rect 14185 34147 14243 34153
rect 14826 34144 14832 34156
rect 14884 34144 14890 34196
rect 15565 34187 15623 34193
rect 15565 34153 15577 34187
rect 15611 34184 15623 34187
rect 15654 34184 15660 34196
rect 15611 34156 15660 34184
rect 15611 34153 15623 34156
rect 15565 34147 15623 34153
rect 15654 34144 15660 34156
rect 15712 34144 15718 34196
rect 16850 34144 16856 34196
rect 16908 34184 16914 34196
rect 17405 34187 17463 34193
rect 17405 34184 17417 34187
rect 16908 34156 17417 34184
rect 16908 34144 16914 34156
rect 17405 34153 17417 34156
rect 17451 34153 17463 34187
rect 17405 34147 17463 34153
rect 6362 34116 6368 34128
rect 6323 34088 6368 34116
rect 6362 34076 6368 34088
rect 6420 34076 6426 34128
rect 15672 34116 15700 34144
rect 16298 34116 16304 34128
rect 15672 34088 16304 34116
rect 16298 34076 16304 34088
rect 16356 34116 16362 34128
rect 16356 34088 16896 34116
rect 16356 34076 16362 34088
rect 3510 34048 3516 34060
rect 3471 34020 3516 34048
rect 3510 34008 3516 34020
rect 3568 34008 3574 34060
rect 6822 34048 6828 34060
rect 6783 34020 6828 34048
rect 6822 34008 6828 34020
rect 6880 34008 6886 34060
rect 7282 34008 7288 34060
rect 7340 34048 7346 34060
rect 7377 34051 7435 34057
rect 7377 34048 7389 34051
rect 7340 34020 7389 34048
rect 7340 34008 7346 34020
rect 7377 34017 7389 34020
rect 7423 34017 7435 34051
rect 7377 34011 7435 34017
rect 7466 34008 7472 34060
rect 7524 34048 7530 34060
rect 7653 34051 7711 34057
rect 7653 34048 7665 34051
rect 7524 34020 7665 34048
rect 7524 34008 7530 34020
rect 7653 34017 7665 34020
rect 7699 34017 7711 34051
rect 9582 34048 9588 34060
rect 9543 34020 9588 34048
rect 7653 34011 7711 34017
rect 9582 34008 9588 34020
rect 9640 34008 9646 34060
rect 9674 34008 9680 34060
rect 9732 34048 9738 34060
rect 10042 34048 10048 34060
rect 9732 34020 9777 34048
rect 10003 34020 10048 34048
rect 9732 34008 9738 34020
rect 10042 34008 10048 34020
rect 10100 34048 10106 34060
rect 10226 34048 10232 34060
rect 10100 34020 10232 34048
rect 10100 34008 10106 34020
rect 10226 34008 10232 34020
rect 10284 34008 10290 34060
rect 14182 34048 14188 34060
rect 14143 34020 14188 34048
rect 14182 34008 14188 34020
rect 14240 34008 14246 34060
rect 14826 34048 14832 34060
rect 14787 34020 14832 34048
rect 14826 34008 14832 34020
rect 14884 34008 14890 34060
rect 15838 34008 15844 34060
rect 15896 34048 15902 34060
rect 15933 34051 15991 34057
rect 15933 34048 15945 34051
rect 15896 34020 15945 34048
rect 15896 34008 15902 34020
rect 15933 34017 15945 34020
rect 15979 34048 15991 34051
rect 16482 34048 16488 34060
rect 15979 34020 16488 34048
rect 15979 34017 15991 34020
rect 15933 34011 15991 34017
rect 16482 34008 16488 34020
rect 16540 34008 16546 34060
rect 16868 34057 16896 34088
rect 16853 34051 16911 34057
rect 16853 34017 16865 34051
rect 16899 34017 16911 34051
rect 16853 34011 16911 34017
rect 3234 33980 3240 33992
rect 3195 33952 3240 33980
rect 3234 33940 3240 33952
rect 3292 33940 3298 33992
rect 4890 33980 4896 33992
rect 4851 33952 4896 33980
rect 4890 33940 4896 33952
rect 4948 33940 4954 33992
rect 9122 33940 9128 33992
rect 9180 33980 9186 33992
rect 9692 33980 9720 34008
rect 9180 33952 9720 33980
rect 9769 33983 9827 33989
rect 9180 33940 9186 33952
rect 9769 33949 9781 33983
rect 9815 33949 9827 33983
rect 14918 33980 14924 33992
rect 14879 33952 14924 33980
rect 9769 33943 9827 33949
rect 6730 33872 6736 33924
rect 6788 33912 6794 33924
rect 6917 33915 6975 33921
rect 6917 33912 6929 33915
rect 6788 33884 6929 33912
rect 6788 33872 6794 33884
rect 6917 33881 6929 33884
rect 6963 33881 6975 33915
rect 6917 33875 6975 33881
rect 9674 33872 9680 33924
rect 9732 33912 9738 33924
rect 9784 33912 9812 33943
rect 14918 33940 14924 33952
rect 14976 33940 14982 33992
rect 16206 33980 16212 33992
rect 16167 33952 16212 33980
rect 16206 33940 16212 33952
rect 16264 33940 16270 33992
rect 17126 33980 17132 33992
rect 17087 33952 17132 33980
rect 17126 33940 17132 33952
rect 17184 33940 17190 33992
rect 9732 33884 9812 33912
rect 9732 33872 9738 33884
rect 1104 33754 18860 33776
rect 1104 33702 4315 33754
rect 4367 33702 4379 33754
rect 4431 33702 4443 33754
rect 4495 33702 4507 33754
rect 4559 33702 10982 33754
rect 11034 33702 11046 33754
rect 11098 33702 11110 33754
rect 11162 33702 11174 33754
rect 11226 33702 17648 33754
rect 17700 33702 17712 33754
rect 17764 33702 17776 33754
rect 17828 33702 17840 33754
rect 17892 33702 18860 33754
rect 1104 33680 18860 33702
rect 2590 33640 2596 33652
rect 1688 33612 2596 33640
rect 1688 33584 1716 33612
rect 2590 33600 2596 33612
rect 2648 33600 2654 33652
rect 3329 33643 3387 33649
rect 3329 33609 3341 33643
rect 3375 33640 3387 33643
rect 3510 33640 3516 33652
rect 3375 33612 3516 33640
rect 3375 33609 3387 33612
rect 3329 33603 3387 33609
rect 3510 33600 3516 33612
rect 3568 33600 3574 33652
rect 5626 33600 5632 33652
rect 5684 33640 5690 33652
rect 5994 33640 6000 33652
rect 5684 33612 6000 33640
rect 5684 33600 5690 33612
rect 5994 33600 6000 33612
rect 6052 33600 6058 33652
rect 6641 33643 6699 33649
rect 6641 33609 6653 33643
rect 6687 33640 6699 33643
rect 6822 33640 6828 33652
rect 6687 33612 6828 33640
rect 6687 33609 6699 33612
rect 6641 33603 6699 33609
rect 6822 33600 6828 33612
rect 6880 33600 6886 33652
rect 8294 33640 8300 33652
rect 8255 33612 8300 33640
rect 8294 33600 8300 33612
rect 8352 33600 8358 33652
rect 8754 33600 8760 33652
rect 8812 33640 8818 33652
rect 9033 33643 9091 33649
rect 9033 33640 9045 33643
rect 8812 33612 9045 33640
rect 8812 33600 8818 33612
rect 9033 33609 9045 33612
rect 9079 33640 9091 33643
rect 9122 33640 9128 33652
rect 9079 33612 9128 33640
rect 9079 33609 9091 33612
rect 9033 33603 9091 33609
rect 9122 33600 9128 33612
rect 9180 33600 9186 33652
rect 9401 33643 9459 33649
rect 9401 33609 9413 33643
rect 9447 33640 9459 33643
rect 10042 33640 10048 33652
rect 9447 33612 10048 33640
rect 9447 33609 9459 33612
rect 9401 33603 9459 33609
rect 10042 33600 10048 33612
rect 10100 33600 10106 33652
rect 10413 33643 10471 33649
rect 10413 33609 10425 33643
rect 10459 33640 10471 33643
rect 10502 33640 10508 33652
rect 10459 33612 10508 33640
rect 10459 33609 10471 33612
rect 10413 33603 10471 33609
rect 1670 33532 1676 33584
rect 1728 33532 1734 33584
rect 5626 33464 5632 33516
rect 5684 33504 5690 33516
rect 6089 33507 6147 33513
rect 6089 33504 6101 33507
rect 5684 33476 6101 33504
rect 5684 33464 5690 33476
rect 6089 33473 6101 33476
rect 6135 33504 6147 33507
rect 6135 33476 6960 33504
rect 6135 33473 6147 33476
rect 6089 33467 6147 33473
rect 2774 33396 2780 33448
rect 2832 33436 2838 33448
rect 3970 33436 3976 33448
rect 2832 33408 3976 33436
rect 2832 33396 2838 33408
rect 3970 33396 3976 33408
rect 4028 33396 4034 33448
rect 4065 33439 4123 33445
rect 4065 33405 4077 33439
rect 4111 33405 4123 33439
rect 4341 33439 4399 33445
rect 4341 33436 4353 33439
rect 4065 33399 4123 33405
rect 4172 33408 4353 33436
rect 2041 33371 2099 33377
rect 2041 33337 2053 33371
rect 2087 33368 2099 33371
rect 2682 33368 2688 33380
rect 2087 33340 2688 33368
rect 2087 33337 2099 33340
rect 2041 33331 2099 33337
rect 2682 33328 2688 33340
rect 2740 33368 2746 33380
rect 2869 33371 2927 33377
rect 2869 33368 2881 33371
rect 2740 33340 2881 33368
rect 2740 33328 2746 33340
rect 2869 33337 2881 33340
rect 2915 33368 2927 33371
rect 3234 33368 3240 33380
rect 2915 33340 3240 33368
rect 2915 33337 2927 33340
rect 2869 33331 2927 33337
rect 3234 33328 3240 33340
rect 3292 33368 3298 33380
rect 4080 33368 4108 33399
rect 3292 33340 4108 33368
rect 3292 33328 3298 33340
rect 1673 33303 1731 33309
rect 1673 33269 1685 33303
rect 1719 33300 1731 33303
rect 1762 33300 1768 33312
rect 1719 33272 1768 33300
rect 1719 33269 1731 33272
rect 1673 33263 1731 33269
rect 1762 33260 1768 33272
rect 1820 33260 1826 33312
rect 3786 33300 3792 33312
rect 3747 33272 3792 33300
rect 3786 33260 3792 33272
rect 3844 33300 3850 33312
rect 4172 33300 4200 33408
rect 4341 33405 4353 33408
rect 4387 33405 4399 33439
rect 6546 33436 6552 33448
rect 6507 33408 6552 33436
rect 4341 33399 4399 33405
rect 6546 33396 6552 33408
rect 6604 33396 6610 33448
rect 6932 33445 6960 33476
rect 6917 33439 6975 33445
rect 6917 33405 6929 33439
rect 6963 33405 6975 33439
rect 6917 33399 6975 33405
rect 7285 33439 7343 33445
rect 7285 33405 7297 33439
rect 7331 33405 7343 33439
rect 7285 33399 7343 33405
rect 7837 33439 7895 33445
rect 7837 33405 7849 33439
rect 7883 33405 7895 33439
rect 7837 33399 7895 33405
rect 9861 33439 9919 33445
rect 9861 33405 9873 33439
rect 9907 33436 9919 33439
rect 10428 33436 10456 33603
rect 10502 33600 10508 33612
rect 10560 33600 10566 33652
rect 14826 33640 14832 33652
rect 14787 33612 14832 33640
rect 14826 33600 14832 33612
rect 14884 33600 14890 33652
rect 15562 33640 15568 33652
rect 15523 33612 15568 33640
rect 15562 33600 15568 33612
rect 15620 33600 15626 33652
rect 15838 33640 15844 33652
rect 15799 33612 15844 33640
rect 15838 33600 15844 33612
rect 15896 33600 15902 33652
rect 17494 33572 17500 33584
rect 17455 33544 17500 33572
rect 17494 33532 17500 33544
rect 17552 33532 17558 33584
rect 18417 33507 18475 33513
rect 18417 33504 18429 33507
rect 17052 33476 18429 33504
rect 17052 33448 17080 33476
rect 18417 33473 18429 33476
rect 18463 33473 18475 33507
rect 18417 33467 18475 33473
rect 9907 33408 10456 33436
rect 9907 33405 9919 33408
rect 9861 33399 9919 33405
rect 5718 33368 5724 33380
rect 5679 33340 5724 33368
rect 5718 33328 5724 33340
rect 5776 33328 5782 33380
rect 5810 33328 5816 33380
rect 5868 33368 5874 33380
rect 6457 33371 6515 33377
rect 6457 33368 6469 33371
rect 5868 33340 6469 33368
rect 5868 33328 5874 33340
rect 6457 33337 6469 33340
rect 6503 33368 6515 33371
rect 7300 33368 7328 33399
rect 6503 33340 7328 33368
rect 6503 33337 6515 33340
rect 6457 33331 6515 33337
rect 3844 33272 4200 33300
rect 3844 33260 3850 33272
rect 6914 33260 6920 33312
rect 6972 33300 6978 33312
rect 7852 33300 7880 33399
rect 15562 33396 15568 33448
rect 15620 33436 15626 33448
rect 15657 33439 15715 33445
rect 15657 33436 15669 33439
rect 15620 33408 15669 33436
rect 15620 33396 15626 33408
rect 15657 33405 15669 33408
rect 15703 33405 15715 33439
rect 15657 33399 15715 33405
rect 16669 33439 16727 33445
rect 16669 33405 16681 33439
rect 16715 33405 16727 33439
rect 17034 33436 17040 33448
rect 16995 33408 17040 33436
rect 16669 33399 16727 33405
rect 9582 33328 9588 33380
rect 9640 33368 9646 33380
rect 10689 33371 10747 33377
rect 10689 33368 10701 33371
rect 9640 33340 10701 33368
rect 9640 33328 9646 33340
rect 10689 33337 10701 33340
rect 10735 33337 10747 33371
rect 10689 33331 10747 33337
rect 6972 33272 7880 33300
rect 6972 33260 6978 33272
rect 9950 33260 9956 33312
rect 10008 33300 10014 33312
rect 10045 33303 10103 33309
rect 10045 33300 10057 33303
rect 10008 33272 10057 33300
rect 10008 33260 10014 33272
rect 10045 33269 10057 33272
rect 10091 33269 10103 33303
rect 14090 33300 14096 33312
rect 14051 33272 14096 33300
rect 10045 33263 10103 33269
rect 14090 33260 14096 33272
rect 14148 33260 14154 33312
rect 14182 33260 14188 33312
rect 14240 33300 14246 33312
rect 14461 33303 14519 33309
rect 14461 33300 14473 33303
rect 14240 33272 14473 33300
rect 14240 33260 14246 33272
rect 14461 33269 14473 33272
rect 14507 33269 14519 33303
rect 14461 33263 14519 33269
rect 14826 33260 14832 33312
rect 14884 33300 14890 33312
rect 15930 33300 15936 33312
rect 14884 33272 15936 33300
rect 14884 33260 14890 33272
rect 15930 33260 15936 33272
rect 15988 33260 15994 33312
rect 16206 33300 16212 33312
rect 16167 33272 16212 33300
rect 16206 33260 16212 33272
rect 16264 33260 16270 33312
rect 16574 33300 16580 33312
rect 16535 33272 16580 33300
rect 16574 33260 16580 33272
rect 16632 33300 16638 33312
rect 16684 33300 16712 33399
rect 17034 33396 17040 33408
rect 17092 33396 17098 33448
rect 17589 33439 17647 33445
rect 17589 33405 17601 33439
rect 17635 33436 17647 33439
rect 17635 33408 18092 33436
rect 17635 33405 17647 33408
rect 17589 33399 17647 33405
rect 18064 33312 18092 33408
rect 18046 33300 18052 33312
rect 16632 33272 16712 33300
rect 18007 33272 18052 33300
rect 16632 33260 16638 33272
rect 18046 33260 18052 33272
rect 18104 33260 18110 33312
rect 1104 33210 18860 33232
rect 1104 33158 7648 33210
rect 7700 33158 7712 33210
rect 7764 33158 7776 33210
rect 7828 33158 7840 33210
rect 7892 33158 14315 33210
rect 14367 33158 14379 33210
rect 14431 33158 14443 33210
rect 14495 33158 14507 33210
rect 14559 33158 18860 33210
rect 1104 33136 18860 33158
rect 2958 33096 2964 33108
rect 2919 33068 2964 33096
rect 2958 33056 2964 33068
rect 3016 33056 3022 33108
rect 6273 33099 6331 33105
rect 6273 33065 6285 33099
rect 6319 33096 6331 33099
rect 6546 33096 6552 33108
rect 6319 33068 6552 33096
rect 6319 33065 6331 33068
rect 6273 33059 6331 33065
rect 6546 33056 6552 33068
rect 6604 33056 6610 33108
rect 6641 33099 6699 33105
rect 6641 33065 6653 33099
rect 6687 33096 6699 33099
rect 6822 33096 6828 33108
rect 6687 33068 6828 33096
rect 6687 33065 6699 33068
rect 6641 33059 6699 33065
rect 5810 33028 5816 33040
rect 5460 33000 5816 33028
rect 4341 32963 4399 32969
rect 4341 32929 4353 32963
rect 4387 32960 4399 32963
rect 4706 32960 4712 32972
rect 4387 32932 4712 32960
rect 4387 32929 4399 32932
rect 4341 32923 4399 32929
rect 4706 32920 4712 32932
rect 4764 32920 4770 32972
rect 5460 32969 5488 33000
rect 5810 32988 5816 33000
rect 5868 32988 5874 33040
rect 5077 32963 5135 32969
rect 5077 32929 5089 32963
rect 5123 32929 5135 32963
rect 5077 32923 5135 32929
rect 5445 32963 5503 32969
rect 5445 32929 5457 32963
rect 5491 32929 5503 32963
rect 5445 32923 5503 32929
rect 5905 32963 5963 32969
rect 5905 32929 5917 32963
rect 5951 32960 5963 32963
rect 6362 32960 6368 32972
rect 5951 32932 6368 32960
rect 5951 32929 5963 32932
rect 5905 32923 5963 32929
rect 1394 32892 1400 32904
rect 1355 32864 1400 32892
rect 1394 32852 1400 32864
rect 1452 32852 1458 32904
rect 1673 32895 1731 32901
rect 1673 32861 1685 32895
rect 1719 32892 1731 32895
rect 1854 32892 1860 32904
rect 1719 32864 1860 32892
rect 1719 32861 1731 32864
rect 1673 32855 1731 32861
rect 1854 32852 1860 32864
rect 1912 32852 1918 32904
rect 4154 32852 4160 32904
rect 4212 32892 4218 32904
rect 4525 32895 4583 32901
rect 4525 32892 4537 32895
rect 4212 32864 4537 32892
rect 4212 32852 4218 32864
rect 4525 32861 4537 32864
rect 4571 32861 4583 32895
rect 5092 32892 5120 32923
rect 6362 32920 6368 32932
rect 6420 32960 6426 32972
rect 6656 32960 6684 33059
rect 6822 33056 6828 33068
rect 6880 33056 6886 33108
rect 7101 33099 7159 33105
rect 7101 33065 7113 33099
rect 7147 33096 7159 33099
rect 7282 33096 7288 33108
rect 7147 33068 7288 33096
rect 7147 33065 7159 33068
rect 7101 33059 7159 33065
rect 7282 33056 7288 33068
rect 7340 33056 7346 33108
rect 7466 33096 7472 33108
rect 7427 33068 7472 33096
rect 7466 33056 7472 33068
rect 7524 33056 7530 33108
rect 15194 33056 15200 33108
rect 15252 33096 15258 33108
rect 15381 33099 15439 33105
rect 15381 33096 15393 33099
rect 15252 33068 15393 33096
rect 15252 33056 15258 33068
rect 15381 33065 15393 33068
rect 15427 33065 15439 33099
rect 15838 33096 15844 33108
rect 15799 33068 15844 33096
rect 15381 33059 15439 33065
rect 15838 33056 15844 33068
rect 15896 33056 15902 33108
rect 17773 33099 17831 33105
rect 17773 33096 17785 33099
rect 16408 33068 17785 33096
rect 9122 32988 9128 33040
rect 9180 33028 9186 33040
rect 9858 33028 9864 33040
rect 9180 33000 9864 33028
rect 9180 32988 9186 33000
rect 9858 32988 9864 33000
rect 9916 32988 9922 33040
rect 10318 33028 10324 33040
rect 10060 33000 10324 33028
rect 9582 32960 9588 32972
rect 6420 32932 6684 32960
rect 9543 32932 9588 32960
rect 6420 32920 6426 32932
rect 9582 32920 9588 32932
rect 9640 32920 9646 32972
rect 9953 32963 10011 32969
rect 9953 32929 9965 32963
rect 9999 32960 10011 32963
rect 10060 32960 10088 33000
rect 10318 32988 10324 33000
rect 10376 32988 10382 33040
rect 14090 32988 14096 33040
rect 14148 33028 14154 33040
rect 14918 33028 14924 33040
rect 14148 33000 14924 33028
rect 14148 32988 14154 33000
rect 9999 32932 10088 32960
rect 10137 32963 10195 32969
rect 9999 32929 10011 32932
rect 9953 32923 10011 32929
rect 10137 32929 10149 32963
rect 10183 32929 10195 32963
rect 10137 32923 10195 32929
rect 5350 32892 5356 32904
rect 5092 32864 5356 32892
rect 4525 32855 4583 32861
rect 5350 32852 5356 32864
rect 5408 32892 5414 32904
rect 5626 32892 5632 32904
rect 5408 32864 5632 32892
rect 5408 32852 5414 32864
rect 5626 32852 5632 32864
rect 5684 32852 5690 32904
rect 9858 32892 9864 32904
rect 9819 32864 9864 32892
rect 9858 32852 9864 32864
rect 9916 32852 9922 32904
rect 9306 32784 9312 32836
rect 9364 32824 9370 32836
rect 10152 32824 10180 32923
rect 10226 32920 10232 32972
rect 10284 32960 10290 32972
rect 10597 32963 10655 32969
rect 10597 32960 10609 32963
rect 10284 32932 10609 32960
rect 10284 32920 10290 32932
rect 10597 32929 10609 32932
rect 10643 32929 10655 32963
rect 10597 32923 10655 32929
rect 13630 32920 13636 32972
rect 13688 32960 13694 32972
rect 14001 32963 14059 32969
rect 14001 32960 14013 32963
rect 13688 32932 14013 32960
rect 13688 32920 13694 32932
rect 14001 32929 14013 32932
rect 14047 32960 14059 32963
rect 14182 32960 14188 32972
rect 14047 32932 14188 32960
rect 14047 32929 14059 32932
rect 14001 32923 14059 32929
rect 14182 32920 14188 32932
rect 14240 32920 14246 32972
rect 14642 32960 14648 32972
rect 14603 32932 14648 32960
rect 14642 32920 14648 32932
rect 14700 32920 14706 32972
rect 14844 32969 14872 33000
rect 14918 32988 14924 33000
rect 14976 32988 14982 33040
rect 15856 33028 15884 33056
rect 16408 33028 16436 33068
rect 17773 33065 17785 33068
rect 17819 33065 17831 33099
rect 17773 33059 17831 33065
rect 17126 33028 17132 33040
rect 15856 33000 16436 33028
rect 17087 33000 17132 33028
rect 14829 32963 14887 32969
rect 14829 32929 14841 32963
rect 14875 32929 14887 32963
rect 14829 32923 14887 32929
rect 15746 32920 15752 32972
rect 15804 32960 15810 32972
rect 16408 32969 16436 33000
rect 17126 32988 17132 33000
rect 17184 32988 17190 33040
rect 17402 33028 17408 33040
rect 17363 33000 17408 33028
rect 17402 32988 17408 33000
rect 17460 32988 17466 33040
rect 16025 32963 16083 32969
rect 16025 32960 16037 32963
rect 15804 32932 16037 32960
rect 15804 32920 15810 32932
rect 16025 32929 16037 32932
rect 16071 32929 16083 32963
rect 16025 32923 16083 32929
rect 16393 32963 16451 32969
rect 16393 32929 16405 32963
rect 16439 32929 16451 32963
rect 16393 32923 16451 32929
rect 16853 32963 16911 32969
rect 16853 32929 16865 32963
rect 16899 32929 16911 32963
rect 16853 32923 16911 32929
rect 16298 32852 16304 32904
rect 16356 32892 16362 32904
rect 16868 32892 16896 32923
rect 18414 32892 18420 32904
rect 16356 32864 18420 32892
rect 16356 32852 16362 32864
rect 18414 32852 18420 32864
rect 18472 32852 18478 32904
rect 9364 32796 10180 32824
rect 9364 32784 9370 32796
rect 13906 32784 13912 32836
rect 13964 32824 13970 32836
rect 14182 32824 14188 32836
rect 13964 32796 14188 32824
rect 13964 32784 13970 32796
rect 14182 32784 14188 32796
rect 14240 32784 14246 32836
rect 14277 32827 14335 32833
rect 14277 32793 14289 32827
rect 14323 32824 14335 32827
rect 15930 32824 15936 32836
rect 14323 32796 15936 32824
rect 14323 32793 14335 32796
rect 14277 32787 14335 32793
rect 15930 32784 15936 32796
rect 15988 32784 15994 32836
rect 3510 32716 3516 32768
rect 3568 32756 3574 32768
rect 3881 32759 3939 32765
rect 3881 32756 3893 32759
rect 3568 32728 3893 32756
rect 3568 32716 3574 32728
rect 3881 32725 3893 32728
rect 3927 32725 3939 32759
rect 9122 32756 9128 32768
rect 9083 32728 9128 32756
rect 3881 32719 3939 32725
rect 9122 32716 9128 32728
rect 9180 32716 9186 32768
rect 9766 32716 9772 32768
rect 9824 32756 9830 32768
rect 9950 32756 9956 32768
rect 9824 32728 9956 32756
rect 9824 32716 9830 32728
rect 9950 32716 9956 32728
rect 10008 32716 10014 32768
rect 10226 32716 10232 32768
rect 10284 32756 10290 32768
rect 11057 32759 11115 32765
rect 11057 32756 11069 32759
rect 10284 32728 11069 32756
rect 10284 32716 10290 32728
rect 11057 32725 11069 32728
rect 11103 32725 11115 32759
rect 11057 32719 11115 32725
rect 11330 32716 11336 32768
rect 11388 32756 11394 32768
rect 11425 32759 11483 32765
rect 11425 32756 11437 32759
rect 11388 32728 11437 32756
rect 11388 32716 11394 32728
rect 11425 32725 11437 32728
rect 11471 32725 11483 32759
rect 11425 32719 11483 32725
rect 1104 32666 18860 32688
rect 1104 32614 4315 32666
rect 4367 32614 4379 32666
rect 4431 32614 4443 32666
rect 4495 32614 4507 32666
rect 4559 32614 10982 32666
rect 11034 32614 11046 32666
rect 11098 32614 11110 32666
rect 11162 32614 11174 32666
rect 11226 32614 17648 32666
rect 17700 32614 17712 32666
rect 17764 32614 17776 32666
rect 17828 32614 17840 32666
rect 17892 32614 18860 32666
rect 1104 32592 18860 32614
rect 2866 32552 2872 32564
rect 2827 32524 2872 32552
rect 2866 32512 2872 32524
rect 2924 32512 2930 32564
rect 3510 32552 3516 32564
rect 3471 32524 3516 32552
rect 3510 32512 3516 32524
rect 3568 32512 3574 32564
rect 5074 32552 5080 32564
rect 5035 32524 5080 32552
rect 5074 32512 5080 32524
rect 5132 32512 5138 32564
rect 8018 32552 8024 32564
rect 7979 32524 8024 32552
rect 8018 32512 8024 32524
rect 8076 32512 8082 32564
rect 8294 32512 8300 32564
rect 8352 32552 8358 32564
rect 8389 32555 8447 32561
rect 8389 32552 8401 32555
rect 8352 32524 8401 32552
rect 8352 32512 8358 32524
rect 8389 32521 8401 32524
rect 8435 32552 8447 32555
rect 8570 32552 8576 32564
rect 8435 32524 8576 32552
rect 8435 32521 8447 32524
rect 8389 32515 8447 32521
rect 8570 32512 8576 32524
rect 8628 32512 8634 32564
rect 9033 32555 9091 32561
rect 9033 32521 9045 32555
rect 9079 32552 9091 32555
rect 10318 32552 10324 32564
rect 9079 32524 10324 32552
rect 9079 32521 9091 32524
rect 9033 32515 9091 32521
rect 10318 32512 10324 32524
rect 10376 32512 10382 32564
rect 14461 32555 14519 32561
rect 14461 32521 14473 32555
rect 14507 32552 14519 32555
rect 14642 32552 14648 32564
rect 14507 32524 14648 32552
rect 14507 32521 14519 32524
rect 14461 32515 14519 32521
rect 14642 32512 14648 32524
rect 14700 32512 14706 32564
rect 15746 32512 15752 32564
rect 15804 32552 15810 32564
rect 16117 32555 16175 32561
rect 16117 32552 16129 32555
rect 15804 32524 16129 32552
rect 15804 32512 15810 32524
rect 16117 32521 16129 32524
rect 16163 32521 16175 32555
rect 18414 32552 18420 32564
rect 18375 32524 18420 32552
rect 16117 32515 16175 32521
rect 18414 32512 18420 32524
rect 18472 32512 18478 32564
rect 8478 32444 8484 32496
rect 8536 32484 8542 32496
rect 8846 32484 8852 32496
rect 8536 32456 8852 32484
rect 8536 32444 8542 32456
rect 8846 32444 8852 32456
rect 8904 32444 8910 32496
rect 9306 32484 9312 32496
rect 9267 32456 9312 32484
rect 9306 32444 9312 32456
rect 9364 32444 9370 32496
rect 1762 32416 1768 32428
rect 1723 32388 1768 32416
rect 1762 32376 1768 32388
rect 1820 32376 1826 32428
rect 4525 32419 4583 32425
rect 4525 32385 4537 32419
rect 4571 32416 4583 32419
rect 4893 32419 4951 32425
rect 4893 32416 4905 32419
rect 4571 32388 4905 32416
rect 4571 32385 4583 32388
rect 4525 32379 4583 32385
rect 4893 32385 4905 32388
rect 4939 32416 4951 32419
rect 5626 32416 5632 32428
rect 4939 32388 5632 32416
rect 4939 32385 4951 32388
rect 4893 32379 4951 32385
rect 5626 32376 5632 32388
rect 5684 32416 5690 32428
rect 10137 32419 10195 32425
rect 5684 32388 5856 32416
rect 5684 32376 5690 32388
rect 5828 32360 5856 32388
rect 10137 32385 10149 32419
rect 10183 32416 10195 32419
rect 11054 32416 11060 32428
rect 10183 32388 10916 32416
rect 11015 32388 11060 32416
rect 10183 32385 10195 32388
rect 10137 32379 10195 32385
rect 1394 32308 1400 32360
rect 1452 32348 1458 32360
rect 1489 32351 1547 32357
rect 1489 32348 1501 32351
rect 1452 32320 1501 32348
rect 1452 32308 1458 32320
rect 1489 32317 1501 32320
rect 1535 32348 1547 32351
rect 2682 32348 2688 32360
rect 1535 32320 2688 32348
rect 1535 32317 1547 32320
rect 1489 32311 1547 32317
rect 2682 32308 2688 32320
rect 2740 32308 2746 32360
rect 4982 32348 4988 32360
rect 4943 32320 4988 32348
rect 4982 32308 4988 32320
rect 5040 32308 5046 32360
rect 5350 32348 5356 32360
rect 5311 32320 5356 32348
rect 5350 32308 5356 32320
rect 5408 32308 5414 32360
rect 5810 32348 5816 32360
rect 5771 32320 5816 32348
rect 5810 32308 5816 32320
rect 5868 32308 5874 32360
rect 6362 32348 6368 32360
rect 6323 32320 6368 32348
rect 6362 32308 6368 32320
rect 6420 32308 6426 32360
rect 8018 32308 8024 32360
rect 8076 32348 8082 32360
rect 8205 32351 8263 32357
rect 8205 32348 8217 32351
rect 8076 32320 8217 32348
rect 8076 32308 8082 32320
rect 8205 32317 8217 32320
rect 8251 32317 8263 32351
rect 8205 32311 8263 32317
rect 9122 32308 9128 32360
rect 9180 32348 9186 32360
rect 9306 32348 9312 32360
rect 9180 32320 9312 32348
rect 9180 32308 9186 32320
rect 9306 32308 9312 32320
rect 9364 32308 9370 32360
rect 10226 32308 10232 32360
rect 10284 32348 10290 32360
rect 10597 32351 10655 32357
rect 10597 32348 10609 32351
rect 10284 32320 10609 32348
rect 10284 32308 10290 32320
rect 10597 32317 10609 32320
rect 10643 32317 10655 32351
rect 10888 32348 10916 32388
rect 11054 32376 11060 32388
rect 11112 32376 11118 32428
rect 11882 32416 11888 32428
rect 11164 32388 11888 32416
rect 11164 32357 11192 32388
rect 11882 32376 11888 32388
rect 11940 32376 11946 32428
rect 11149 32351 11207 32357
rect 11149 32348 11161 32351
rect 10888 32320 11161 32348
rect 10597 32311 10655 32317
rect 11149 32317 11161 32320
rect 11195 32317 11207 32351
rect 11149 32311 11207 32317
rect 11609 32351 11667 32357
rect 11609 32317 11621 32351
rect 11655 32348 11667 32351
rect 11698 32348 11704 32360
rect 11655 32320 11704 32348
rect 11655 32317 11667 32320
rect 11609 32311 11667 32317
rect 3881 32283 3939 32289
rect 3881 32249 3893 32283
rect 3927 32280 3939 32283
rect 5368 32280 5396 32308
rect 3927 32252 5396 32280
rect 3927 32249 3939 32252
rect 3881 32243 3939 32249
rect 10318 32240 10324 32292
rect 10376 32280 10382 32292
rect 10505 32283 10563 32289
rect 10505 32280 10517 32283
rect 10376 32252 10517 32280
rect 10376 32240 10382 32252
rect 10505 32249 10517 32252
rect 10551 32280 10563 32283
rect 11624 32280 11652 32311
rect 11698 32308 11704 32320
rect 11756 32308 11762 32360
rect 11793 32351 11851 32357
rect 11793 32317 11805 32351
rect 11839 32317 11851 32351
rect 11793 32311 11851 32317
rect 11808 32280 11836 32311
rect 15194 32308 15200 32360
rect 15252 32348 15258 32360
rect 15378 32348 15384 32360
rect 15252 32320 15384 32348
rect 15252 32308 15258 32320
rect 15378 32308 15384 32320
rect 15436 32348 15442 32360
rect 15473 32351 15531 32357
rect 15473 32348 15485 32351
rect 15436 32320 15485 32348
rect 15436 32308 15442 32320
rect 15473 32317 15485 32320
rect 15519 32317 15531 32351
rect 15473 32311 15531 32317
rect 16669 32351 16727 32357
rect 16669 32317 16681 32351
rect 16715 32317 16727 32351
rect 16669 32311 16727 32317
rect 17221 32351 17279 32357
rect 17221 32317 17233 32351
rect 17267 32348 17279 32351
rect 17402 32348 17408 32360
rect 17267 32320 17408 32348
rect 17267 32317 17279 32320
rect 17221 32311 17279 32317
rect 10551 32252 11652 32280
rect 11716 32252 11836 32280
rect 10551 32249 10563 32252
rect 10505 32243 10563 32249
rect 2682 32172 2688 32224
rect 2740 32212 2746 32224
rect 3510 32212 3516 32224
rect 2740 32184 3516 32212
rect 2740 32172 2746 32184
rect 3510 32172 3516 32184
rect 3568 32172 3574 32224
rect 11330 32172 11336 32224
rect 11388 32212 11394 32224
rect 11716 32212 11744 32252
rect 13262 32240 13268 32292
rect 13320 32280 13326 32292
rect 14001 32283 14059 32289
rect 14001 32280 14013 32283
rect 13320 32252 14013 32280
rect 13320 32240 13326 32252
rect 14001 32249 14013 32252
rect 14047 32280 14059 32283
rect 14090 32280 14096 32292
rect 14047 32252 14096 32280
rect 14047 32249 14059 32252
rect 14001 32243 14059 32249
rect 14090 32240 14096 32252
rect 14148 32240 14154 32292
rect 15105 32283 15163 32289
rect 15105 32249 15117 32283
rect 15151 32280 15163 32283
rect 15286 32280 15292 32292
rect 15151 32252 15292 32280
rect 15151 32249 15163 32252
rect 15105 32243 15163 32249
rect 15286 32240 15292 32252
rect 15344 32240 15350 32292
rect 11388 32184 11744 32212
rect 11388 32172 11394 32184
rect 12894 32172 12900 32224
rect 12952 32212 12958 32224
rect 13630 32212 13636 32224
rect 12952 32184 13636 32212
rect 12952 32172 12958 32184
rect 13630 32172 13636 32184
rect 13688 32172 13694 32224
rect 15562 32212 15568 32224
rect 15523 32184 15568 32212
rect 15562 32172 15568 32184
rect 15620 32172 15626 32224
rect 16574 32212 16580 32224
rect 16535 32184 16580 32212
rect 16574 32172 16580 32184
rect 16632 32212 16638 32224
rect 16684 32212 16712 32311
rect 17402 32308 17408 32320
rect 17460 32308 17466 32360
rect 17497 32351 17555 32357
rect 17497 32317 17509 32351
rect 17543 32348 17555 32351
rect 18046 32348 18052 32360
rect 17543 32320 18052 32348
rect 17543 32317 17555 32320
rect 17497 32311 17555 32317
rect 16850 32240 16856 32292
rect 16908 32280 16914 32292
rect 17512 32280 17540 32311
rect 18046 32308 18052 32320
rect 18104 32308 18110 32360
rect 17770 32280 17776 32292
rect 16908 32252 17540 32280
rect 17731 32252 17776 32280
rect 16908 32240 16914 32252
rect 17770 32240 17776 32252
rect 17828 32240 17834 32292
rect 16632 32184 16712 32212
rect 16632 32172 16638 32184
rect 17402 32172 17408 32224
rect 17460 32212 17466 32224
rect 17954 32212 17960 32224
rect 17460 32184 17960 32212
rect 17460 32172 17466 32184
rect 17954 32172 17960 32184
rect 18012 32172 18018 32224
rect 1104 32122 18860 32144
rect 1104 32070 7648 32122
rect 7700 32070 7712 32122
rect 7764 32070 7776 32122
rect 7828 32070 7840 32122
rect 7892 32070 14315 32122
rect 14367 32070 14379 32122
rect 14431 32070 14443 32122
rect 14495 32070 14507 32122
rect 14559 32070 18860 32122
rect 1104 32048 18860 32070
rect 3326 31968 3332 32020
rect 3384 32008 3390 32020
rect 3510 32008 3516 32020
rect 3384 31980 3516 32008
rect 3384 31968 3390 31980
rect 3510 31968 3516 31980
rect 3568 31968 3574 32020
rect 5350 32008 5356 32020
rect 5311 31980 5356 32008
rect 5350 31968 5356 31980
rect 5408 31968 5414 32020
rect 5905 32011 5963 32017
rect 5905 31977 5917 32011
rect 5951 32008 5963 32011
rect 6638 32008 6644 32020
rect 5951 31980 6644 32008
rect 5951 31977 5963 31980
rect 5905 31971 5963 31977
rect 6638 31968 6644 31980
rect 6696 31968 6702 32020
rect 7282 31968 7288 32020
rect 7340 32008 7346 32020
rect 7653 32011 7711 32017
rect 7653 32008 7665 32011
rect 7340 31980 7665 32008
rect 7340 31968 7346 31980
rect 7653 31977 7665 31980
rect 7699 31977 7711 32011
rect 7653 31971 7711 31977
rect 9401 32011 9459 32017
rect 9401 31977 9413 32011
rect 9447 32008 9459 32011
rect 9582 32008 9588 32020
rect 9447 31980 9588 32008
rect 9447 31977 9459 31980
rect 9401 31971 9459 31977
rect 9582 31968 9588 31980
rect 9640 31968 9646 32020
rect 9858 32008 9864 32020
rect 9819 31980 9864 32008
rect 9858 31968 9864 31980
rect 9916 31968 9922 32020
rect 12618 32008 12624 32020
rect 12579 31980 12624 32008
rect 12618 31968 12624 31980
rect 12676 31968 12682 32020
rect 15470 31968 15476 32020
rect 15528 32008 15534 32020
rect 15565 32011 15623 32017
rect 15565 32008 15577 32011
rect 15528 31980 15577 32008
rect 15528 31968 15534 31980
rect 15565 31977 15577 31980
rect 15611 32008 15623 32011
rect 15746 32008 15752 32020
rect 15611 31980 15752 32008
rect 15611 31977 15623 31980
rect 15565 31971 15623 31977
rect 15746 31968 15752 31980
rect 15804 32008 15810 32020
rect 15804 31980 16528 32008
rect 15804 31968 15810 31980
rect 3142 31940 3148 31952
rect 3103 31912 3148 31940
rect 3142 31900 3148 31912
rect 3200 31900 3206 31952
rect 4525 31943 4583 31949
rect 4525 31909 4537 31943
rect 4571 31940 4583 31943
rect 5077 31943 5135 31949
rect 5077 31940 5089 31943
rect 4571 31912 5089 31940
rect 4571 31909 4583 31912
rect 4525 31903 4583 31909
rect 5077 31909 5089 31912
rect 5123 31940 5135 31943
rect 6362 31940 6368 31952
rect 5123 31912 6368 31940
rect 5123 31909 5135 31912
rect 5077 31903 5135 31909
rect 6362 31900 6368 31912
rect 6420 31900 6426 31952
rect 15838 31900 15844 31952
rect 15896 31940 15902 31952
rect 16500 31949 16528 31980
rect 16025 31943 16083 31949
rect 16025 31940 16037 31943
rect 15896 31912 16037 31940
rect 15896 31900 15902 31912
rect 16025 31909 16037 31912
rect 16071 31940 16083 31943
rect 16393 31943 16451 31949
rect 16393 31940 16405 31943
rect 16071 31912 16405 31940
rect 16071 31909 16083 31912
rect 16025 31903 16083 31909
rect 16393 31909 16405 31912
rect 16439 31909 16451 31943
rect 16393 31903 16451 31909
rect 16485 31943 16543 31949
rect 16485 31909 16497 31943
rect 16531 31909 16543 31943
rect 16485 31903 16543 31909
rect 16853 31943 16911 31949
rect 16853 31909 16865 31943
rect 16899 31940 16911 31943
rect 17221 31943 17279 31949
rect 17221 31940 17233 31943
rect 16899 31912 17233 31940
rect 16899 31909 16911 31912
rect 16853 31903 16911 31909
rect 17221 31909 17233 31912
rect 17267 31940 17279 31943
rect 17494 31940 17500 31952
rect 17267 31912 17500 31940
rect 17267 31909 17279 31912
rect 17221 31903 17279 31909
rect 17494 31900 17500 31912
rect 17552 31900 17558 31952
rect 1578 31832 1584 31884
rect 1636 31872 1642 31884
rect 1765 31875 1823 31881
rect 1765 31872 1777 31875
rect 1636 31844 1777 31872
rect 1636 31832 1642 31844
rect 1765 31841 1777 31844
rect 1811 31841 1823 31875
rect 1765 31835 1823 31841
rect 4982 31832 4988 31884
rect 5040 31872 5046 31884
rect 5810 31872 5816 31884
rect 5040 31844 5816 31872
rect 5040 31832 5046 31844
rect 5810 31832 5816 31844
rect 5868 31832 5874 31884
rect 5994 31832 6000 31884
rect 6052 31872 6058 31884
rect 6089 31875 6147 31881
rect 6089 31872 6101 31875
rect 6052 31844 6101 31872
rect 6052 31832 6058 31844
rect 6089 31841 6101 31844
rect 6135 31841 6147 31875
rect 6089 31835 6147 31841
rect 7745 31875 7803 31881
rect 7745 31841 7757 31875
rect 7791 31872 7803 31875
rect 8018 31872 8024 31884
rect 7791 31844 8024 31872
rect 7791 31841 7803 31844
rect 7745 31835 7803 31841
rect 8018 31832 8024 31844
rect 8076 31832 8082 31884
rect 8205 31875 8263 31881
rect 8205 31841 8217 31875
rect 8251 31872 8263 31875
rect 8754 31872 8760 31884
rect 8251 31844 8760 31872
rect 8251 31841 8263 31844
rect 8205 31835 8263 31841
rect 1486 31804 1492 31816
rect 1447 31776 1492 31804
rect 1486 31764 1492 31776
rect 1544 31764 1550 31816
rect 7466 31764 7472 31816
rect 7524 31804 7530 31816
rect 8220 31804 8248 31835
rect 8754 31832 8760 31844
rect 8812 31832 8818 31884
rect 10229 31875 10287 31881
rect 10229 31841 10241 31875
rect 10275 31872 10287 31875
rect 10594 31872 10600 31884
rect 10275 31844 10600 31872
rect 10275 31841 10287 31844
rect 10229 31835 10287 31841
rect 10594 31832 10600 31844
rect 10652 31832 10658 31884
rect 11054 31872 11060 31884
rect 11015 31844 11060 31872
rect 11054 31832 11060 31844
rect 11112 31832 11118 31884
rect 11425 31875 11483 31881
rect 11425 31841 11437 31875
rect 11471 31872 11483 31875
rect 11514 31872 11520 31884
rect 11471 31844 11520 31872
rect 11471 31841 11483 31844
rect 11425 31835 11483 31841
rect 11514 31832 11520 31844
rect 11572 31832 11578 31884
rect 12434 31832 12440 31884
rect 12492 31872 12498 31884
rect 12492 31844 12537 31872
rect 12492 31832 12498 31844
rect 13722 31832 13728 31884
rect 13780 31872 13786 31884
rect 14550 31872 14556 31884
rect 13780 31844 14556 31872
rect 13780 31832 13786 31844
rect 14550 31832 14556 31844
rect 14608 31832 14614 31884
rect 14642 31832 14648 31884
rect 14700 31872 14706 31884
rect 14826 31872 14832 31884
rect 14700 31844 14745 31872
rect 14787 31844 14832 31872
rect 14700 31832 14706 31844
rect 14826 31832 14832 31844
rect 14884 31832 14890 31884
rect 15289 31875 15347 31881
rect 15289 31841 15301 31875
rect 15335 31872 15347 31875
rect 16298 31872 16304 31884
rect 15335 31844 16304 31872
rect 15335 31841 15347 31844
rect 15289 31835 15347 31841
rect 16298 31832 16304 31844
rect 16356 31832 16362 31884
rect 7524 31776 8248 31804
rect 8573 31807 8631 31813
rect 7524 31764 7530 31776
rect 8573 31773 8585 31807
rect 8619 31804 8631 31807
rect 8846 31804 8852 31816
rect 8619 31776 8852 31804
rect 8619 31773 8631 31776
rect 8573 31767 8631 31773
rect 8846 31764 8852 31776
rect 8904 31764 8910 31816
rect 11072 31804 11100 31832
rect 10980 31776 11100 31804
rect 3326 31696 3332 31748
rect 3384 31736 3390 31748
rect 4062 31736 4068 31748
rect 3384 31708 4068 31736
rect 3384 31696 3390 31708
rect 4062 31696 4068 31708
rect 4120 31696 4126 31748
rect 9858 31696 9864 31748
rect 9916 31736 9922 31748
rect 10505 31739 10563 31745
rect 10505 31736 10517 31739
rect 9916 31708 10517 31736
rect 9916 31696 9922 31708
rect 10505 31705 10517 31708
rect 10551 31705 10563 31739
rect 10505 31699 10563 31705
rect 10686 31696 10692 31748
rect 10744 31736 10750 31748
rect 10980 31736 11008 31776
rect 15930 31764 15936 31816
rect 15988 31804 15994 31816
rect 16117 31807 16175 31813
rect 16117 31804 16129 31807
rect 15988 31776 16129 31804
rect 15988 31764 15994 31776
rect 16117 31773 16129 31776
rect 16163 31773 16175 31807
rect 16117 31767 16175 31773
rect 17310 31764 17316 31816
rect 17368 31804 17374 31816
rect 17497 31807 17555 31813
rect 17497 31804 17509 31807
rect 17368 31776 17509 31804
rect 17368 31764 17374 31776
rect 17497 31773 17509 31776
rect 17543 31773 17555 31807
rect 17497 31767 17555 31773
rect 10744 31708 11008 31736
rect 10744 31696 10750 31708
rect 10870 31628 10876 31680
rect 10928 31668 10934 31680
rect 11330 31668 11336 31680
rect 10928 31640 11336 31668
rect 10928 31628 10934 31640
rect 11330 31628 11336 31640
rect 11388 31628 11394 31680
rect 1104 31578 18860 31600
rect 1104 31526 4315 31578
rect 4367 31526 4379 31578
rect 4431 31526 4443 31578
rect 4495 31526 4507 31578
rect 4559 31526 10982 31578
rect 11034 31526 11046 31578
rect 11098 31526 11110 31578
rect 11162 31526 11174 31578
rect 11226 31526 17648 31578
rect 17700 31526 17712 31578
rect 17764 31526 17776 31578
rect 17828 31526 17840 31578
rect 17892 31526 18860 31578
rect 1104 31504 18860 31526
rect 1854 31424 1860 31476
rect 1912 31464 1918 31476
rect 1949 31467 2007 31473
rect 1949 31464 1961 31467
rect 1912 31436 1961 31464
rect 1912 31424 1918 31436
rect 1949 31433 1961 31436
rect 1995 31433 2007 31467
rect 1949 31427 2007 31433
rect 5813 31467 5871 31473
rect 5813 31433 5825 31467
rect 5859 31464 5871 31467
rect 5994 31464 6000 31476
rect 5859 31436 6000 31464
rect 5859 31433 5871 31436
rect 5813 31427 5871 31433
rect 5994 31424 6000 31436
rect 6052 31424 6058 31476
rect 6457 31467 6515 31473
rect 6457 31433 6469 31467
rect 6503 31464 6515 31467
rect 6546 31464 6552 31476
rect 6503 31436 6552 31464
rect 6503 31433 6515 31436
rect 6457 31427 6515 31433
rect 6546 31424 6552 31436
rect 6604 31424 6610 31476
rect 7466 31464 7472 31476
rect 7427 31436 7472 31464
rect 7466 31424 7472 31436
rect 7524 31424 7530 31476
rect 8665 31467 8723 31473
rect 8665 31433 8677 31467
rect 8711 31464 8723 31467
rect 8754 31464 8760 31476
rect 8711 31436 8760 31464
rect 8711 31433 8723 31436
rect 8665 31427 8723 31433
rect 8754 31424 8760 31436
rect 8812 31424 8818 31476
rect 14642 31424 14648 31476
rect 14700 31464 14706 31476
rect 14921 31467 14979 31473
rect 14921 31464 14933 31467
rect 14700 31436 14933 31464
rect 14700 31424 14706 31436
rect 14921 31433 14933 31436
rect 14967 31433 14979 31467
rect 14921 31427 14979 31433
rect 15930 31424 15936 31476
rect 15988 31464 15994 31476
rect 16485 31467 16543 31473
rect 16485 31464 16497 31467
rect 15988 31436 16497 31464
rect 15988 31424 15994 31436
rect 16485 31433 16497 31436
rect 16531 31433 16543 31467
rect 16485 31427 16543 31433
rect 1486 31356 1492 31408
rect 1544 31396 1550 31408
rect 2317 31399 2375 31405
rect 2317 31396 2329 31399
rect 1544 31368 2329 31396
rect 1544 31356 1550 31368
rect 2317 31365 2329 31368
rect 2363 31365 2375 31399
rect 2317 31359 2375 31365
rect 8018 31356 8024 31408
rect 8076 31356 8082 31408
rect 14277 31399 14335 31405
rect 14277 31365 14289 31399
rect 14323 31396 14335 31399
rect 14826 31396 14832 31408
rect 14323 31368 14832 31396
rect 14323 31365 14335 31368
rect 14277 31359 14335 31365
rect 14826 31356 14832 31368
rect 14884 31356 14890 31408
rect 8036 31328 8064 31356
rect 8113 31331 8171 31337
rect 8113 31328 8125 31331
rect 8036 31300 8125 31328
rect 8113 31297 8125 31300
rect 8159 31297 8171 31331
rect 8113 31291 8171 31297
rect 9125 31331 9183 31337
rect 9125 31297 9137 31331
rect 9171 31328 9183 31331
rect 10778 31328 10784 31340
rect 9171 31300 10784 31328
rect 9171 31297 9183 31300
rect 9125 31291 9183 31297
rect 2130 31220 2136 31272
rect 2188 31260 2194 31272
rect 2314 31260 2320 31272
rect 2188 31232 2320 31260
rect 2188 31220 2194 31232
rect 2314 31220 2320 31232
rect 2372 31220 2378 31272
rect 6270 31260 6276 31272
rect 6104 31232 6276 31260
rect 1578 31192 1584 31204
rect 1539 31164 1584 31192
rect 1578 31152 1584 31164
rect 1636 31152 1642 31204
rect 5994 31084 6000 31136
rect 6052 31124 6058 31136
rect 6104 31133 6132 31232
rect 6270 31220 6276 31232
rect 6328 31220 6334 31272
rect 7101 31263 7159 31269
rect 7101 31229 7113 31263
rect 7147 31260 7159 31263
rect 7837 31263 7895 31269
rect 7837 31260 7849 31263
rect 7147 31232 7849 31260
rect 7147 31229 7159 31232
rect 7101 31223 7159 31229
rect 7837 31229 7849 31232
rect 7883 31260 7895 31263
rect 7926 31260 7932 31272
rect 7883 31232 7932 31260
rect 7883 31229 7895 31232
rect 7837 31223 7895 31229
rect 7926 31220 7932 31232
rect 7984 31220 7990 31272
rect 8021 31263 8079 31269
rect 8021 31229 8033 31263
rect 8067 31229 8079 31263
rect 9490 31260 9496 31272
rect 9451 31232 9496 31260
rect 8021 31223 8079 31229
rect 7466 31152 7472 31204
rect 7524 31192 7530 31204
rect 8036 31192 8064 31223
rect 9490 31220 9496 31232
rect 9548 31220 9554 31272
rect 9858 31260 9864 31272
rect 9819 31232 9864 31260
rect 9858 31220 9864 31232
rect 9916 31220 9922 31272
rect 9950 31220 9956 31272
rect 10008 31260 10014 31272
rect 10704 31269 10732 31300
rect 10778 31288 10784 31300
rect 10836 31288 10842 31340
rect 15286 31288 15292 31340
rect 15344 31288 15350 31340
rect 15838 31328 15844 31340
rect 15799 31300 15844 31328
rect 15838 31288 15844 31300
rect 15896 31288 15902 31340
rect 10321 31263 10379 31269
rect 10321 31260 10333 31263
rect 10008 31232 10333 31260
rect 10008 31220 10014 31232
rect 10321 31229 10333 31232
rect 10367 31229 10379 31263
rect 10321 31223 10379 31229
rect 10689 31263 10747 31269
rect 10689 31229 10701 31263
rect 10735 31229 10747 31263
rect 10689 31223 10747 31229
rect 11330 31220 11336 31272
rect 11388 31260 11394 31272
rect 11793 31263 11851 31269
rect 11793 31260 11805 31263
rect 11388 31232 11805 31260
rect 11388 31220 11394 31232
rect 11793 31229 11805 31232
rect 11839 31229 11851 31263
rect 11793 31223 11851 31229
rect 12253 31263 12311 31269
rect 12253 31229 12265 31263
rect 12299 31229 12311 31263
rect 12253 31223 12311 31229
rect 12268 31192 12296 31223
rect 12434 31192 12440 31204
rect 7524 31164 8064 31192
rect 11624 31164 12440 31192
rect 7524 31152 7530 31164
rect 6089 31127 6147 31133
rect 6089 31124 6101 31127
rect 6052 31096 6101 31124
rect 6052 31084 6058 31096
rect 6089 31093 6101 31096
rect 6135 31093 6147 31127
rect 9950 31124 9956 31136
rect 9911 31096 9956 31124
rect 6089 31087 6147 31093
rect 9950 31084 9956 31096
rect 10008 31084 10014 31136
rect 11054 31084 11060 31136
rect 11112 31124 11118 31136
rect 11624 31133 11652 31164
rect 12434 31152 12440 31164
rect 12492 31192 12498 31204
rect 15304 31201 15332 31288
rect 15378 31220 15384 31272
rect 15436 31260 15442 31272
rect 15473 31263 15531 31269
rect 15473 31260 15485 31263
rect 15436 31232 15485 31260
rect 15436 31220 15442 31232
rect 15473 31229 15485 31232
rect 15519 31229 15531 31263
rect 15473 31223 15531 31229
rect 16114 31220 16120 31272
rect 16172 31220 16178 31272
rect 16574 31220 16580 31272
rect 16632 31260 16638 31272
rect 16669 31263 16727 31269
rect 16669 31260 16681 31263
rect 16632 31232 16681 31260
rect 16632 31220 16638 31232
rect 16669 31229 16681 31232
rect 16715 31229 16727 31263
rect 16669 31223 16727 31229
rect 17221 31263 17279 31269
rect 17221 31229 17233 31263
rect 17267 31260 17279 31263
rect 17310 31260 17316 31272
rect 17267 31232 17316 31260
rect 17267 31229 17279 31232
rect 17221 31223 17279 31229
rect 17310 31220 17316 31232
rect 17368 31220 17374 31272
rect 17494 31260 17500 31272
rect 17455 31232 17500 31260
rect 17494 31220 17500 31232
rect 17552 31220 17558 31272
rect 12805 31195 12863 31201
rect 12805 31192 12817 31195
rect 12492 31164 12817 31192
rect 12492 31152 12498 31164
rect 12805 31161 12817 31164
rect 12851 31161 12863 31195
rect 12805 31155 12863 31161
rect 15289 31195 15347 31201
rect 15289 31161 15301 31195
rect 15335 31161 15347 31195
rect 15289 31155 15347 31161
rect 11609 31127 11667 31133
rect 11609 31124 11621 31127
rect 11112 31096 11621 31124
rect 11112 31084 11118 31096
rect 11609 31093 11621 31096
rect 11655 31093 11667 31127
rect 12066 31124 12072 31136
rect 12027 31096 12072 31124
rect 11609 31087 11667 31093
rect 12066 31084 12072 31096
rect 12124 31084 12130 31136
rect 14642 31124 14648 31136
rect 14603 31096 14648 31124
rect 14642 31084 14648 31096
rect 14700 31084 14706 31136
rect 15304 31124 15332 31155
rect 15838 31152 15844 31204
rect 15896 31192 15902 31204
rect 16132 31192 16160 31220
rect 17770 31192 17776 31204
rect 15896 31164 16160 31192
rect 17731 31164 17776 31192
rect 15896 31152 15902 31164
rect 17770 31152 17776 31164
rect 17828 31152 17834 31204
rect 16114 31124 16120 31136
rect 15304 31096 16120 31124
rect 16114 31084 16120 31096
rect 16172 31084 16178 31136
rect 1104 31034 18860 31056
rect 1104 30982 7648 31034
rect 7700 30982 7712 31034
rect 7764 30982 7776 31034
rect 7828 30982 7840 31034
rect 7892 30982 14315 31034
rect 14367 30982 14379 31034
rect 14431 30982 14443 31034
rect 14495 30982 14507 31034
rect 14559 30982 18860 31034
rect 1104 30960 18860 30982
rect 4709 30923 4767 30929
rect 4709 30889 4721 30923
rect 4755 30920 4767 30923
rect 6546 30920 6552 30932
rect 4755 30892 6552 30920
rect 4755 30889 4767 30892
rect 4709 30883 4767 30889
rect 3329 30855 3387 30861
rect 3329 30821 3341 30855
rect 3375 30852 3387 30855
rect 3418 30852 3424 30864
rect 3375 30824 3424 30852
rect 3375 30821 3387 30824
rect 3329 30815 3387 30821
rect 3418 30812 3424 30824
rect 3476 30812 3482 30864
rect 1762 30744 1768 30796
rect 1820 30784 1826 30796
rect 5368 30793 5396 30892
rect 6546 30880 6552 30892
rect 6604 30880 6610 30932
rect 8018 30920 8024 30932
rect 7979 30892 8024 30920
rect 8018 30880 8024 30892
rect 8076 30880 8082 30932
rect 9858 30920 9864 30932
rect 9819 30892 9864 30920
rect 9858 30880 9864 30892
rect 9916 30880 9922 30932
rect 10594 30920 10600 30932
rect 10555 30892 10600 30920
rect 10594 30880 10600 30892
rect 10652 30880 10658 30932
rect 15562 30880 15568 30932
rect 15620 30880 15626 30932
rect 16025 30923 16083 30929
rect 16025 30889 16037 30923
rect 16071 30920 16083 30923
rect 16298 30920 16304 30932
rect 16071 30892 16304 30920
rect 16071 30889 16083 30892
rect 16025 30883 16083 30889
rect 16298 30880 16304 30892
rect 16356 30880 16362 30932
rect 16942 30880 16948 30932
rect 17000 30920 17006 30932
rect 17497 30923 17555 30929
rect 17497 30920 17509 30923
rect 17000 30892 17509 30920
rect 17000 30880 17006 30892
rect 17497 30889 17509 30892
rect 17543 30889 17555 30923
rect 17497 30883 17555 30889
rect 5905 30855 5963 30861
rect 5905 30821 5917 30855
rect 5951 30852 5963 30855
rect 6178 30852 6184 30864
rect 5951 30824 6184 30852
rect 5951 30821 5963 30824
rect 5905 30815 5963 30821
rect 6178 30812 6184 30824
rect 6236 30812 6242 30864
rect 10321 30855 10379 30861
rect 10321 30821 10333 30855
rect 10367 30852 10379 30855
rect 10686 30852 10692 30864
rect 10367 30824 10692 30852
rect 10367 30821 10379 30824
rect 10321 30815 10379 30821
rect 10686 30812 10692 30824
rect 10744 30812 10750 30864
rect 11330 30812 11336 30864
rect 11388 30852 11394 30864
rect 11793 30855 11851 30861
rect 11793 30852 11805 30855
rect 11388 30824 11805 30852
rect 11388 30812 11394 30824
rect 11793 30821 11805 30824
rect 11839 30821 11851 30855
rect 11793 30815 11851 30821
rect 1949 30787 2007 30793
rect 1949 30784 1961 30787
rect 1820 30756 1961 30784
rect 1820 30744 1826 30756
rect 1949 30753 1961 30756
rect 1995 30753 2007 30787
rect 1949 30747 2007 30753
rect 5353 30787 5411 30793
rect 5353 30753 5365 30787
rect 5399 30753 5411 30787
rect 5626 30784 5632 30796
rect 5587 30756 5632 30784
rect 5353 30747 5411 30753
rect 5626 30744 5632 30756
rect 5684 30744 5690 30796
rect 15580 30784 15608 30880
rect 15746 30812 15752 30864
rect 15804 30852 15810 30864
rect 15841 30855 15899 30861
rect 15841 30852 15853 30855
rect 15804 30824 15853 30852
rect 15804 30812 15810 30824
rect 15841 30821 15853 30824
rect 15887 30852 15899 30855
rect 16485 30855 16543 30861
rect 16485 30852 16497 30855
rect 15887 30824 16497 30852
rect 15887 30821 15899 30824
rect 15841 30815 15899 30821
rect 16485 30821 16497 30824
rect 16531 30821 16543 30855
rect 16850 30852 16856 30864
rect 16811 30824 16856 30852
rect 16485 30815 16543 30821
rect 16850 30812 16856 30824
rect 16908 30812 16914 30864
rect 16393 30787 16451 30793
rect 16393 30784 16405 30787
rect 15488 30756 16405 30784
rect 15488 30728 15516 30756
rect 16393 30753 16405 30756
rect 16439 30753 16451 30787
rect 16393 30747 16451 30753
rect 1673 30719 1731 30725
rect 1673 30685 1685 30719
rect 1719 30716 1731 30719
rect 2130 30716 2136 30728
rect 1719 30688 2136 30716
rect 1719 30685 1731 30688
rect 1673 30679 1731 30685
rect 2130 30676 2136 30688
rect 2188 30716 2194 30728
rect 2682 30716 2688 30728
rect 2188 30688 2688 30716
rect 2188 30676 2194 30688
rect 2682 30676 2688 30688
rect 2740 30676 2746 30728
rect 4982 30716 4988 30728
rect 4943 30688 4988 30716
rect 4982 30676 4988 30688
rect 5040 30676 5046 30728
rect 15470 30676 15476 30728
rect 15528 30676 15534 30728
rect 15930 30676 15936 30728
rect 15988 30716 15994 30728
rect 16117 30719 16175 30725
rect 16117 30716 16129 30719
rect 15988 30688 16129 30716
rect 15988 30676 15994 30688
rect 16117 30685 16129 30688
rect 16163 30685 16175 30719
rect 16117 30679 16175 30685
rect 11330 30608 11336 30660
rect 11388 30648 11394 30660
rect 11606 30648 11612 30660
rect 11388 30620 11612 30648
rect 11388 30608 11394 30620
rect 11606 30608 11612 30620
rect 11664 30608 11670 30660
rect 15378 30648 15384 30660
rect 15291 30620 15384 30648
rect 15378 30608 15384 30620
rect 15436 30648 15442 30660
rect 16482 30648 16488 30660
rect 15436 30620 16488 30648
rect 15436 30608 15442 30620
rect 16482 30608 16488 30620
rect 16540 30648 16546 30660
rect 16850 30648 16856 30660
rect 16540 30620 16856 30648
rect 16540 30608 16546 30620
rect 16850 30608 16856 30620
rect 16908 30608 16914 30660
rect 7650 30580 7656 30592
rect 7611 30552 7656 30580
rect 7650 30540 7656 30552
rect 7708 30540 7714 30592
rect 12710 30580 12716 30592
rect 12671 30552 12716 30580
rect 12710 30540 12716 30552
rect 12768 30540 12774 30592
rect 15194 30540 15200 30592
rect 15252 30580 15258 30592
rect 15841 30583 15899 30589
rect 15841 30580 15853 30583
rect 15252 30552 15853 30580
rect 15252 30540 15258 30552
rect 15841 30549 15853 30552
rect 15887 30549 15899 30583
rect 15841 30543 15899 30549
rect 16574 30540 16580 30592
rect 16632 30580 16638 30592
rect 17129 30583 17187 30589
rect 17129 30580 17141 30583
rect 16632 30552 17141 30580
rect 16632 30540 16638 30552
rect 17129 30549 17141 30552
rect 17175 30549 17187 30583
rect 17129 30543 17187 30549
rect 1104 30490 18860 30512
rect 1104 30438 4315 30490
rect 4367 30438 4379 30490
rect 4431 30438 4443 30490
rect 4495 30438 4507 30490
rect 4559 30438 10982 30490
rect 11034 30438 11046 30490
rect 11098 30438 11110 30490
rect 11162 30438 11174 30490
rect 11226 30438 17648 30490
rect 17700 30438 17712 30490
rect 17764 30438 17776 30490
rect 17828 30438 17840 30490
rect 17892 30438 18860 30490
rect 1104 30416 18860 30438
rect 4617 30379 4675 30385
rect 4617 30345 4629 30379
rect 4663 30376 4675 30379
rect 4982 30376 4988 30388
rect 4663 30348 4988 30376
rect 4663 30345 4675 30348
rect 4617 30339 4675 30345
rect 4982 30336 4988 30348
rect 5040 30336 5046 30388
rect 15470 30376 15476 30388
rect 14936 30348 15476 30376
rect 6914 30268 6920 30320
rect 6972 30308 6978 30320
rect 7561 30311 7619 30317
rect 7561 30308 7573 30311
rect 6972 30280 7573 30308
rect 6972 30268 6978 30280
rect 7561 30277 7573 30280
rect 7607 30277 7619 30311
rect 12894 30308 12900 30320
rect 12855 30280 12900 30308
rect 7561 30271 7619 30277
rect 12894 30268 12900 30280
rect 12952 30268 12958 30320
rect 14737 30311 14795 30317
rect 14737 30277 14749 30311
rect 14783 30308 14795 30311
rect 14936 30308 14964 30348
rect 15470 30336 15476 30348
rect 15528 30336 15534 30388
rect 15565 30379 15623 30385
rect 15565 30345 15577 30379
rect 15611 30376 15623 30379
rect 16298 30376 16304 30388
rect 15611 30348 16304 30376
rect 15611 30345 15623 30348
rect 15565 30339 15623 30345
rect 16298 30336 16304 30348
rect 16356 30336 16362 30388
rect 15102 30308 15108 30320
rect 14783 30280 14964 30308
rect 15063 30280 15108 30308
rect 14783 30277 14795 30280
rect 14737 30271 14795 30277
rect 15102 30268 15108 30280
rect 15160 30268 15166 30320
rect 15838 30308 15844 30320
rect 15799 30280 15844 30308
rect 15838 30268 15844 30280
rect 15896 30268 15902 30320
rect 15930 30268 15936 30320
rect 15988 30308 15994 30320
rect 16485 30311 16543 30317
rect 16485 30308 16497 30311
rect 15988 30280 16497 30308
rect 15988 30268 15994 30280
rect 16485 30277 16497 30280
rect 16531 30277 16543 30311
rect 16485 30271 16543 30277
rect 4430 30200 4436 30252
rect 4488 30240 4494 30252
rect 5169 30243 5227 30249
rect 5169 30240 5181 30243
rect 4488 30212 5181 30240
rect 4488 30200 4494 30212
rect 5169 30209 5181 30212
rect 5215 30240 5227 30243
rect 5626 30240 5632 30252
rect 5215 30212 5632 30240
rect 5215 30209 5227 30212
rect 5169 30203 5227 30209
rect 5626 30200 5632 30212
rect 5684 30200 5690 30252
rect 8938 30200 8944 30252
rect 8996 30240 9002 30252
rect 9677 30243 9735 30249
rect 9677 30240 9689 30243
rect 8996 30212 9689 30240
rect 8996 30200 9002 30212
rect 9677 30209 9689 30212
rect 9723 30209 9735 30243
rect 9677 30203 9735 30209
rect 17773 30243 17831 30249
rect 17773 30209 17785 30243
rect 17819 30240 17831 30243
rect 17862 30240 17868 30252
rect 17819 30212 17868 30240
rect 17819 30209 17831 30212
rect 17773 30203 17831 30209
rect 17862 30200 17868 30212
rect 17920 30200 17926 30252
rect 4890 30132 4896 30184
rect 4948 30172 4954 30184
rect 5077 30175 5135 30181
rect 5077 30172 5089 30175
rect 4948 30144 5089 30172
rect 4948 30132 4954 30144
rect 5077 30141 5089 30144
rect 5123 30172 5135 30175
rect 5350 30172 5356 30184
rect 5123 30144 5356 30172
rect 5123 30141 5135 30144
rect 5077 30135 5135 30141
rect 5350 30132 5356 30144
rect 5408 30132 5414 30184
rect 5442 30132 5448 30184
rect 5500 30172 5506 30184
rect 5500 30144 5545 30172
rect 5500 30132 5506 30144
rect 5718 30132 5724 30184
rect 5776 30172 5782 30184
rect 5813 30175 5871 30181
rect 5813 30172 5825 30175
rect 5776 30144 5825 30172
rect 5776 30132 5782 30144
rect 5813 30141 5825 30144
rect 5859 30141 5871 30175
rect 5813 30135 5871 30141
rect 5902 30132 5908 30184
rect 5960 30172 5966 30184
rect 6549 30175 6607 30181
rect 6549 30172 6561 30175
rect 5960 30144 6561 30172
rect 5960 30132 5966 30144
rect 6549 30141 6561 30144
rect 6595 30172 6607 30175
rect 6914 30172 6920 30184
rect 6595 30144 6920 30172
rect 6595 30141 6607 30144
rect 6549 30135 6607 30141
rect 6914 30132 6920 30144
rect 6972 30132 6978 30184
rect 7190 30132 7196 30184
rect 7248 30172 7254 30184
rect 7377 30175 7435 30181
rect 7377 30172 7389 30175
rect 7248 30144 7389 30172
rect 7248 30132 7254 30144
rect 7377 30141 7389 30144
rect 7423 30172 7435 30175
rect 7837 30175 7895 30181
rect 7837 30172 7849 30175
rect 7423 30144 7849 30172
rect 7423 30141 7435 30144
rect 7377 30135 7435 30141
rect 7837 30141 7849 30144
rect 7883 30141 7895 30175
rect 8386 30172 8392 30184
rect 8347 30144 8392 30172
rect 7837 30135 7895 30141
rect 4985 30107 5043 30113
rect 4985 30073 4997 30107
rect 5031 30104 5043 30107
rect 5460 30104 5488 30132
rect 5031 30076 5488 30104
rect 5031 30073 5043 30076
rect 4985 30067 5043 30073
rect 1670 30036 1676 30048
rect 1631 30008 1676 30036
rect 1670 29996 1676 30008
rect 1728 29996 1734 30048
rect 2130 30036 2136 30048
rect 2091 30008 2136 30036
rect 2130 29996 2136 30008
rect 2188 29996 2194 30048
rect 6546 29996 6552 30048
rect 6604 30036 6610 30048
rect 6825 30039 6883 30045
rect 6825 30036 6837 30039
rect 6604 30008 6837 30036
rect 6604 29996 6610 30008
rect 6825 30005 6837 30008
rect 6871 30005 6883 30039
rect 7852 30036 7880 30135
rect 8386 30132 8392 30144
rect 8444 30172 8450 30184
rect 8754 30172 8760 30184
rect 8444 30144 8760 30172
rect 8444 30132 8450 30144
rect 8754 30132 8760 30144
rect 8812 30172 8818 30184
rect 8849 30175 8907 30181
rect 8849 30172 8861 30175
rect 8812 30144 8861 30172
rect 8812 30132 8818 30144
rect 8849 30141 8861 30144
rect 8895 30141 8907 30175
rect 8849 30135 8907 30141
rect 9122 30132 9128 30184
rect 9180 30172 9186 30184
rect 9493 30175 9551 30181
rect 9493 30172 9505 30175
rect 9180 30144 9505 30172
rect 9180 30132 9186 30144
rect 9493 30141 9505 30144
rect 9539 30172 9551 30175
rect 10321 30175 10379 30181
rect 10321 30172 10333 30175
rect 9539 30144 10333 30172
rect 9539 30141 9551 30144
rect 9493 30135 9551 30141
rect 10321 30141 10333 30144
rect 10367 30172 10379 30175
rect 10502 30172 10508 30184
rect 10367 30144 10508 30172
rect 10367 30141 10379 30144
rect 10321 30135 10379 30141
rect 10502 30132 10508 30144
rect 10560 30132 10566 30184
rect 12710 30132 12716 30184
rect 12768 30172 12774 30184
rect 13081 30175 13139 30181
rect 13081 30172 13093 30175
rect 12768 30144 13093 30172
rect 12768 30132 12774 30144
rect 13081 30141 13093 30144
rect 13127 30141 13139 30175
rect 13081 30135 13139 30141
rect 13170 30132 13176 30184
rect 13228 30172 13234 30184
rect 13265 30175 13323 30181
rect 13265 30172 13277 30175
rect 13228 30144 13277 30172
rect 13228 30132 13234 30144
rect 13265 30141 13277 30144
rect 13311 30141 13323 30175
rect 13265 30135 13323 30141
rect 13449 30175 13507 30181
rect 13449 30141 13461 30175
rect 13495 30141 13507 30175
rect 13449 30135 13507 30141
rect 8294 30036 8300 30048
rect 7852 30008 8300 30036
rect 6825 29999 6883 30005
rect 8294 29996 8300 30008
rect 8352 30036 8358 30048
rect 8573 30039 8631 30045
rect 8573 30036 8585 30039
rect 8352 30008 8585 30036
rect 8352 29996 8358 30008
rect 8573 30005 8585 30008
rect 8619 30005 8631 30039
rect 12066 30036 12072 30048
rect 12027 30008 12072 30036
rect 8573 29999 8631 30005
rect 12066 29996 12072 30008
rect 12124 29996 12130 30048
rect 12526 30036 12532 30048
rect 12487 30008 12532 30036
rect 12526 29996 12532 30008
rect 12584 30036 12590 30048
rect 13464 30036 13492 30135
rect 15194 30132 15200 30184
rect 15252 30172 15258 30184
rect 15657 30175 15715 30181
rect 15657 30172 15669 30175
rect 15252 30144 15669 30172
rect 15252 30132 15258 30144
rect 15657 30141 15669 30144
rect 15703 30172 15715 30175
rect 16114 30172 16120 30184
rect 15703 30144 16120 30172
rect 15703 30141 15715 30144
rect 15657 30135 15715 30141
rect 16114 30132 16120 30144
rect 16172 30132 16178 30184
rect 16574 30132 16580 30184
rect 16632 30172 16638 30184
rect 16669 30175 16727 30181
rect 16669 30172 16681 30175
rect 16632 30144 16681 30172
rect 16632 30132 16638 30144
rect 16669 30141 16681 30144
rect 16715 30141 16727 30175
rect 16669 30135 16727 30141
rect 16942 30132 16948 30184
rect 17000 30172 17006 30184
rect 17037 30175 17095 30181
rect 17037 30172 17049 30175
rect 17000 30144 17049 30172
rect 17000 30132 17006 30144
rect 17037 30141 17049 30144
rect 17083 30141 17095 30175
rect 17494 30172 17500 30184
rect 17455 30144 17500 30172
rect 17037 30135 17095 30141
rect 17494 30132 17500 30144
rect 17552 30172 17558 30184
rect 18049 30175 18107 30181
rect 18049 30172 18061 30175
rect 17552 30144 18061 30172
rect 17552 30132 17558 30144
rect 18049 30141 18061 30144
rect 18095 30141 18107 30175
rect 18049 30135 18107 30141
rect 12584 30008 13492 30036
rect 12584 29996 12590 30008
rect 1104 29946 18860 29968
rect 1104 29894 7648 29946
rect 7700 29894 7712 29946
rect 7764 29894 7776 29946
rect 7828 29894 7840 29946
rect 7892 29894 14315 29946
rect 14367 29894 14379 29946
rect 14431 29894 14443 29946
rect 14495 29894 14507 29946
rect 14559 29894 18860 29946
rect 1104 29872 18860 29894
rect 1673 29835 1731 29841
rect 1673 29801 1685 29835
rect 1719 29832 1731 29835
rect 2038 29832 2044 29844
rect 1719 29804 2044 29832
rect 1719 29801 1731 29804
rect 1673 29795 1731 29801
rect 2038 29792 2044 29804
rect 2096 29792 2102 29844
rect 4522 29832 4528 29844
rect 4483 29804 4528 29832
rect 4522 29792 4528 29804
rect 4580 29792 4586 29844
rect 5169 29835 5227 29841
rect 5169 29801 5181 29835
rect 5215 29832 5227 29835
rect 5537 29835 5595 29841
rect 5537 29832 5549 29835
rect 5215 29804 5549 29832
rect 5215 29801 5227 29804
rect 5169 29795 5227 29801
rect 5537 29801 5549 29804
rect 5583 29832 5595 29835
rect 5718 29832 5724 29844
rect 5583 29804 5724 29832
rect 5583 29801 5595 29804
rect 5537 29795 5595 29801
rect 5718 29792 5724 29804
rect 5776 29832 5782 29844
rect 7009 29835 7067 29841
rect 7009 29832 7021 29835
rect 5776 29804 7021 29832
rect 5776 29792 5782 29804
rect 7009 29801 7021 29804
rect 7055 29801 7067 29835
rect 7009 29795 7067 29801
rect 13262 29792 13268 29844
rect 13320 29832 13326 29844
rect 13357 29835 13415 29841
rect 13357 29832 13369 29835
rect 13320 29804 13369 29832
rect 13320 29792 13326 29804
rect 13357 29801 13369 29804
rect 13403 29801 13415 29835
rect 15286 29832 15292 29844
rect 15247 29804 15292 29832
rect 13357 29795 13415 29801
rect 15286 29792 15292 29804
rect 15344 29792 15350 29844
rect 16022 29792 16028 29844
rect 16080 29792 16086 29844
rect 17126 29832 17132 29844
rect 17087 29804 17132 29832
rect 17126 29792 17132 29804
rect 17184 29792 17190 29844
rect 3694 29764 3700 29776
rect 3655 29736 3700 29764
rect 3694 29724 3700 29736
rect 3752 29724 3758 29776
rect 4430 29764 4436 29776
rect 4391 29736 4436 29764
rect 4430 29724 4436 29736
rect 4488 29724 4494 29776
rect 5626 29724 5632 29776
rect 5684 29764 5690 29776
rect 5902 29764 5908 29776
rect 5684 29736 5908 29764
rect 5684 29724 5690 29736
rect 5902 29724 5908 29736
rect 5960 29724 5966 29776
rect 8205 29767 8263 29773
rect 8205 29733 8217 29767
rect 8251 29764 8263 29767
rect 15933 29767 15991 29773
rect 8251 29736 9168 29764
rect 8251 29733 8263 29736
rect 8205 29727 8263 29733
rect 9140 29708 9168 29736
rect 15933 29733 15945 29767
rect 15979 29764 15991 29767
rect 16040 29764 16068 29792
rect 15979 29736 16068 29764
rect 15979 29733 15991 29736
rect 15933 29727 15991 29733
rect 1486 29656 1492 29708
rect 1544 29696 1550 29708
rect 2041 29699 2099 29705
rect 2041 29696 2053 29699
rect 1544 29668 2053 29696
rect 1544 29656 1550 29668
rect 2041 29665 2053 29668
rect 2087 29665 2099 29699
rect 2041 29659 2099 29665
rect 2130 29656 2136 29708
rect 2188 29696 2194 29708
rect 2317 29699 2375 29705
rect 2317 29696 2329 29699
rect 2188 29668 2329 29696
rect 2188 29656 2194 29668
rect 2317 29665 2329 29668
rect 2363 29665 2375 29699
rect 4706 29696 4712 29708
rect 4667 29668 4712 29696
rect 2317 29659 2375 29665
rect 4706 29656 4712 29668
rect 4764 29656 4770 29708
rect 6822 29696 6828 29708
rect 6783 29668 6828 29696
rect 6822 29656 6828 29668
rect 6880 29656 6886 29708
rect 8294 29696 8300 29708
rect 8255 29668 8300 29696
rect 8294 29656 8300 29668
rect 8352 29656 8358 29708
rect 9122 29696 9128 29708
rect 9083 29668 9128 29696
rect 9122 29656 9128 29668
rect 9180 29656 9186 29708
rect 9309 29699 9367 29705
rect 9309 29665 9321 29699
rect 9355 29696 9367 29699
rect 9490 29696 9496 29708
rect 9355 29668 9496 29696
rect 9355 29665 9367 29668
rect 9309 29659 9367 29665
rect 9490 29656 9496 29668
rect 9548 29696 9554 29708
rect 10134 29696 10140 29708
rect 9548 29668 10140 29696
rect 9548 29656 9554 29668
rect 10134 29656 10140 29668
rect 10192 29656 10198 29708
rect 10226 29656 10232 29708
rect 10284 29696 10290 29708
rect 10873 29699 10931 29705
rect 10873 29696 10885 29699
rect 10284 29668 10885 29696
rect 10284 29656 10290 29668
rect 10873 29665 10885 29668
rect 10919 29696 10931 29699
rect 10962 29696 10968 29708
rect 10919 29668 10968 29696
rect 10919 29665 10931 29668
rect 10873 29659 10931 29665
rect 10962 29656 10968 29668
rect 11020 29656 11026 29708
rect 12437 29699 12495 29705
rect 12437 29665 12449 29699
rect 12483 29665 12495 29699
rect 13265 29699 13323 29705
rect 13265 29696 13277 29699
rect 12437 29659 12495 29665
rect 12820 29668 13277 29696
rect 7745 29631 7803 29637
rect 7745 29597 7757 29631
rect 7791 29628 7803 29631
rect 8386 29628 8392 29640
rect 7791 29600 8392 29628
rect 7791 29597 7803 29600
rect 7745 29591 7803 29597
rect 8386 29588 8392 29600
rect 8444 29628 8450 29640
rect 10244 29628 10272 29656
rect 8444 29600 10272 29628
rect 12452 29628 12480 29659
rect 12618 29628 12624 29640
rect 12452 29600 12624 29628
rect 8444 29588 8450 29600
rect 12618 29588 12624 29600
rect 12676 29588 12682 29640
rect 12434 29520 12440 29572
rect 12492 29560 12498 29572
rect 12820 29560 12848 29668
rect 13265 29665 13277 29668
rect 13311 29696 13323 29699
rect 14366 29696 14372 29708
rect 13311 29668 14372 29696
rect 13311 29665 13323 29668
rect 13265 29659 13323 29665
rect 14366 29656 14372 29668
rect 14424 29656 14430 29708
rect 16025 29699 16083 29705
rect 16025 29665 16037 29699
rect 16071 29696 16083 29699
rect 16298 29696 16304 29708
rect 16071 29668 16304 29696
rect 16071 29665 16083 29668
rect 16025 29659 16083 29665
rect 16298 29656 16304 29668
rect 16356 29656 16362 29708
rect 13170 29628 13176 29640
rect 13131 29600 13176 29628
rect 13170 29588 13176 29600
rect 13228 29588 13234 29640
rect 15749 29631 15807 29637
rect 15749 29597 15761 29631
rect 15795 29628 15807 29631
rect 15930 29628 15936 29640
rect 15795 29600 15936 29628
rect 15795 29597 15807 29600
rect 15749 29591 15807 29597
rect 15930 29588 15936 29600
rect 15988 29588 15994 29640
rect 12492 29532 12848 29560
rect 12492 29520 12498 29532
rect 9398 29452 9404 29504
rect 9456 29492 9462 29504
rect 10686 29492 10692 29504
rect 9456 29464 9501 29492
rect 10647 29464 10692 29492
rect 9456 29452 9462 29464
rect 10686 29452 10692 29464
rect 10744 29452 10750 29504
rect 12250 29492 12256 29504
rect 12211 29464 12256 29492
rect 12250 29452 12256 29464
rect 12308 29452 12314 29504
rect 13630 29452 13636 29504
rect 13688 29492 13694 29504
rect 14553 29495 14611 29501
rect 14553 29492 14565 29495
rect 13688 29464 14565 29492
rect 13688 29452 13694 29464
rect 14553 29461 14565 29464
rect 14599 29461 14611 29495
rect 16206 29492 16212 29504
rect 16167 29464 16212 29492
rect 14553 29455 14611 29461
rect 16206 29452 16212 29464
rect 16264 29452 16270 29504
rect 16574 29452 16580 29504
rect 16632 29492 16638 29504
rect 16761 29495 16819 29501
rect 16761 29492 16773 29495
rect 16632 29464 16773 29492
rect 16632 29452 16638 29464
rect 16761 29461 16773 29464
rect 16807 29461 16819 29495
rect 17494 29492 17500 29504
rect 17455 29464 17500 29492
rect 16761 29455 16819 29461
rect 17494 29452 17500 29464
rect 17552 29452 17558 29504
rect 1104 29402 18860 29424
rect 1104 29350 4315 29402
rect 4367 29350 4379 29402
rect 4431 29350 4443 29402
rect 4495 29350 4507 29402
rect 4559 29350 10982 29402
rect 11034 29350 11046 29402
rect 11098 29350 11110 29402
rect 11162 29350 11174 29402
rect 11226 29350 17648 29402
rect 17700 29350 17712 29402
rect 17764 29350 17776 29402
rect 17828 29350 17840 29402
rect 17892 29350 18860 29402
rect 1104 29328 18860 29350
rect 7190 29248 7196 29300
rect 7248 29288 7254 29300
rect 7469 29291 7527 29297
rect 7469 29288 7481 29291
rect 7248 29260 7481 29288
rect 7248 29248 7254 29260
rect 7469 29257 7481 29260
rect 7515 29257 7527 29291
rect 9490 29288 9496 29300
rect 9451 29260 9496 29288
rect 7469 29251 7527 29257
rect 1486 29152 1492 29164
rect 1447 29124 1492 29152
rect 1486 29112 1492 29124
rect 1544 29152 1550 29164
rect 2590 29152 2596 29164
rect 1544 29124 2596 29152
rect 1544 29112 1550 29124
rect 2590 29112 2596 29124
rect 2648 29112 2654 29164
rect 5445 29155 5503 29161
rect 5445 29121 5457 29155
rect 5491 29152 5503 29155
rect 5718 29152 5724 29164
rect 5491 29124 5724 29152
rect 5491 29121 5503 29124
rect 5445 29115 5503 29121
rect 5718 29112 5724 29124
rect 5776 29112 5782 29164
rect 6178 29112 6184 29164
rect 6236 29152 6242 29164
rect 6822 29152 6828 29164
rect 6236 29124 6828 29152
rect 6236 29112 6242 29124
rect 6822 29112 6828 29124
rect 6880 29112 6886 29164
rect 7484 29152 7512 29251
rect 9490 29248 9496 29260
rect 9548 29248 9554 29300
rect 10137 29291 10195 29297
rect 10137 29257 10149 29291
rect 10183 29288 10195 29291
rect 10226 29288 10232 29300
rect 10183 29260 10232 29288
rect 10183 29257 10195 29260
rect 10137 29251 10195 29257
rect 10226 29248 10232 29260
rect 10284 29248 10290 29300
rect 10689 29291 10747 29297
rect 10689 29257 10701 29291
rect 10735 29288 10747 29291
rect 10870 29288 10876 29300
rect 10735 29260 10876 29288
rect 10735 29257 10747 29260
rect 10689 29251 10747 29257
rect 10870 29248 10876 29260
rect 10928 29248 10934 29300
rect 14366 29288 14372 29300
rect 14327 29260 14372 29288
rect 14366 29248 14372 29260
rect 14424 29248 14430 29300
rect 15930 29248 15936 29300
rect 15988 29288 15994 29300
rect 16117 29291 16175 29297
rect 16117 29288 16129 29291
rect 15988 29260 16129 29288
rect 15988 29248 15994 29260
rect 16117 29257 16129 29260
rect 16163 29257 16175 29291
rect 16117 29251 16175 29257
rect 9033 29155 9091 29161
rect 9033 29152 9045 29155
rect 7484 29124 9045 29152
rect 1765 29087 1823 29093
rect 1765 29053 1777 29087
rect 1811 29084 1823 29087
rect 2038 29084 2044 29096
rect 1811 29056 2044 29084
rect 1811 29053 1823 29056
rect 1765 29047 1823 29053
rect 2038 29044 2044 29056
rect 2096 29044 2102 29096
rect 5353 29087 5411 29093
rect 5353 29053 5365 29087
rect 5399 29084 5411 29087
rect 6362 29084 6368 29096
rect 5399 29056 6368 29084
rect 5399 29053 5411 29056
rect 5353 29047 5411 29053
rect 3142 29016 3148 29028
rect 3103 28988 3148 29016
rect 3142 28976 3148 28988
rect 3200 28976 3206 29028
rect 4617 29019 4675 29025
rect 4617 28985 4629 29019
rect 4663 29016 4675 29019
rect 4890 29016 4896 29028
rect 4663 28988 4896 29016
rect 4663 28985 4675 28988
rect 4617 28979 4675 28985
rect 4890 28976 4896 28988
rect 4948 28976 4954 29028
rect 4985 29019 5043 29025
rect 4985 28985 4997 29019
rect 5031 29016 5043 29019
rect 5626 29016 5632 29028
rect 5031 28988 5632 29016
rect 5031 28985 5043 28988
rect 4985 28979 5043 28985
rect 5626 28976 5632 28988
rect 5684 28976 5690 29028
rect 5828 29025 5856 29056
rect 6362 29044 6368 29056
rect 6420 29044 6426 29096
rect 7484 29084 7512 29124
rect 9033 29121 9045 29124
rect 9079 29121 9091 29155
rect 9033 29115 9091 29121
rect 12250 29112 12256 29164
rect 12308 29152 12314 29164
rect 13817 29155 13875 29161
rect 12308 29124 13676 29152
rect 12308 29112 12314 29124
rect 13648 29096 13676 29124
rect 13817 29121 13829 29155
rect 13863 29152 13875 29155
rect 14642 29152 14648 29164
rect 13863 29124 14648 29152
rect 13863 29121 13875 29124
rect 13817 29115 13875 29121
rect 14642 29112 14648 29124
rect 14700 29112 14706 29164
rect 15105 29155 15163 29161
rect 15105 29121 15117 29155
rect 15151 29152 15163 29155
rect 15289 29155 15347 29161
rect 15289 29152 15301 29155
rect 15151 29124 15301 29152
rect 15151 29121 15163 29124
rect 15105 29115 15163 29121
rect 15289 29121 15301 29124
rect 15335 29152 15347 29155
rect 15948 29152 15976 29248
rect 15335 29124 15976 29152
rect 15335 29121 15347 29124
rect 15289 29115 15347 29121
rect 7653 29087 7711 29093
rect 7653 29084 7665 29087
rect 7484 29056 7665 29084
rect 7653 29053 7665 29056
rect 7699 29053 7711 29087
rect 7653 29047 7711 29053
rect 8297 29087 8355 29093
rect 8297 29053 8309 29087
rect 8343 29084 8355 29087
rect 8386 29084 8392 29096
rect 8343 29056 8392 29084
rect 8343 29053 8355 29056
rect 8297 29047 8355 29053
rect 8386 29044 8392 29056
rect 8444 29044 8450 29096
rect 8481 29087 8539 29093
rect 8481 29053 8493 29087
rect 8527 29084 8539 29087
rect 9490 29084 9496 29096
rect 8527 29056 9496 29084
rect 8527 29053 8539 29056
rect 8481 29047 8539 29053
rect 5721 29019 5779 29025
rect 5721 28985 5733 29019
rect 5767 28985 5779 29019
rect 5721 28979 5779 28985
rect 5813 29019 5871 29025
rect 5813 28985 5825 29019
rect 5859 28985 5871 29019
rect 5813 28979 5871 28985
rect 3418 28948 3424 28960
rect 3379 28920 3424 28948
rect 3418 28908 3424 28920
rect 3476 28908 3482 28960
rect 4908 28948 4936 28976
rect 5736 28948 5764 28979
rect 5902 28976 5908 29028
rect 5960 29016 5966 29028
rect 6181 29019 6239 29025
rect 6181 29016 6193 29019
rect 5960 28988 6193 29016
rect 5960 28976 5966 28988
rect 6181 28985 6193 28988
rect 6227 28985 6239 29019
rect 6546 29016 6552 29028
rect 6181 28979 6239 28985
rect 6288 28988 6552 29016
rect 6288 28948 6316 28988
rect 6546 28976 6552 28988
rect 6604 28976 6610 29028
rect 8496 29016 8524 29047
rect 9490 29044 9496 29056
rect 9548 29044 9554 29096
rect 10134 29044 10140 29096
rect 10192 29084 10198 29096
rect 10321 29087 10379 29093
rect 10321 29084 10333 29087
rect 10192 29056 10333 29084
rect 10192 29044 10198 29056
rect 10321 29053 10333 29056
rect 10367 29053 10379 29087
rect 12618 29084 12624 29096
rect 12579 29056 12624 29084
rect 10321 29047 10379 29053
rect 12618 29044 12624 29056
rect 12676 29044 12682 29096
rect 12989 29087 13047 29093
rect 12989 29053 13001 29087
rect 13035 29053 13047 29087
rect 13630 29084 13636 29096
rect 13591 29056 13636 29084
rect 12989 29047 13047 29053
rect 11790 29016 11796 29028
rect 8220 28988 8524 29016
rect 11703 28988 11796 29016
rect 4908 28920 6316 28948
rect 7929 28951 7987 28957
rect 7929 28917 7941 28951
rect 7975 28948 7987 28951
rect 8018 28948 8024 28960
rect 7975 28920 8024 28948
rect 7975 28917 7987 28920
rect 7929 28911 7987 28917
rect 8018 28908 8024 28920
rect 8076 28908 8082 28960
rect 8110 28908 8116 28960
rect 8168 28948 8174 28960
rect 8220 28948 8248 28988
rect 11790 28976 11796 28988
rect 11848 29016 11854 29028
rect 13004 29016 13032 29047
rect 13630 29044 13636 29056
rect 13688 29044 13694 29096
rect 15378 29044 15384 29096
rect 15436 29084 15442 29096
rect 16669 29087 16727 29093
rect 15436 29056 15481 29084
rect 15436 29044 15442 29056
rect 16669 29053 16681 29087
rect 16715 29053 16727 29087
rect 17126 29084 17132 29096
rect 17087 29056 17132 29084
rect 16669 29047 16727 29053
rect 15838 29016 15844 29028
rect 11848 28988 13032 29016
rect 15799 28988 15844 29016
rect 11848 28976 11854 28988
rect 15838 28976 15844 28988
rect 15896 28976 15902 29028
rect 8168 28920 8248 28948
rect 11425 28951 11483 28957
rect 8168 28908 8174 28920
rect 11425 28917 11437 28951
rect 11471 28948 11483 28951
rect 12066 28948 12072 28960
rect 11471 28920 12072 28948
rect 11471 28917 11483 28920
rect 11425 28911 11483 28917
rect 12066 28908 12072 28920
rect 12124 28908 12130 28960
rect 12161 28951 12219 28957
rect 12161 28917 12173 28951
rect 12207 28948 12219 28951
rect 12529 28951 12587 28957
rect 12529 28948 12541 28951
rect 12207 28920 12541 28948
rect 12207 28917 12219 28920
rect 12161 28911 12219 28917
rect 12529 28917 12541 28920
rect 12575 28948 12587 28951
rect 12618 28948 12624 28960
rect 12575 28920 12624 28948
rect 12575 28917 12587 28920
rect 12529 28911 12587 28917
rect 12618 28908 12624 28920
rect 12676 28908 12682 28960
rect 16574 28948 16580 28960
rect 16535 28920 16580 28948
rect 16574 28908 16580 28920
rect 16632 28948 16638 28960
rect 16684 28948 16712 29047
rect 17126 29044 17132 29056
rect 17184 29044 17190 29096
rect 17494 29084 17500 29096
rect 17455 29056 17500 29084
rect 17494 29044 17500 29056
rect 17552 29044 17558 29096
rect 17770 29084 17776 29096
rect 17731 29056 17776 29084
rect 17770 29044 17776 29056
rect 17828 29044 17834 29096
rect 16632 28920 16712 28948
rect 16632 28908 16638 28920
rect 1104 28858 18860 28880
rect 1104 28806 7648 28858
rect 7700 28806 7712 28858
rect 7764 28806 7776 28858
rect 7828 28806 7840 28858
rect 7892 28806 14315 28858
rect 14367 28806 14379 28858
rect 14431 28806 14443 28858
rect 14495 28806 14507 28858
rect 14559 28806 18860 28858
rect 1104 28784 18860 28806
rect 2130 28704 2136 28756
rect 2188 28744 2194 28756
rect 2225 28747 2283 28753
rect 2225 28744 2237 28747
rect 2188 28716 2237 28744
rect 2188 28704 2194 28716
rect 2225 28713 2237 28716
rect 2271 28713 2283 28747
rect 2590 28744 2596 28756
rect 2551 28716 2596 28744
rect 2225 28707 2283 28713
rect 2590 28704 2596 28716
rect 2648 28744 2654 28756
rect 3418 28744 3424 28756
rect 2648 28716 3424 28744
rect 2648 28704 2654 28716
rect 3418 28704 3424 28716
rect 3476 28704 3482 28756
rect 6273 28747 6331 28753
rect 6273 28713 6285 28747
rect 6319 28744 6331 28747
rect 6730 28744 6736 28756
rect 6319 28716 6736 28744
rect 6319 28713 6331 28716
rect 6273 28707 6331 28713
rect 6730 28704 6736 28716
rect 6788 28704 6794 28756
rect 7098 28744 7104 28756
rect 7059 28716 7104 28744
rect 7098 28704 7104 28716
rect 7156 28704 7162 28756
rect 7745 28747 7803 28753
rect 7745 28713 7757 28747
rect 7791 28744 7803 28747
rect 8110 28744 8116 28756
rect 7791 28716 8116 28744
rect 7791 28713 7803 28716
rect 7745 28707 7803 28713
rect 8110 28704 8116 28716
rect 8168 28704 8174 28756
rect 10321 28747 10379 28753
rect 10321 28713 10333 28747
rect 10367 28744 10379 28747
rect 10410 28744 10416 28756
rect 10367 28716 10416 28744
rect 10367 28713 10379 28716
rect 10321 28707 10379 28713
rect 10410 28704 10416 28716
rect 10468 28704 10474 28756
rect 12253 28747 12311 28753
rect 12253 28713 12265 28747
rect 12299 28744 12311 28747
rect 12342 28744 12348 28756
rect 12299 28716 12348 28744
rect 12299 28713 12311 28716
rect 12253 28707 12311 28713
rect 12342 28704 12348 28716
rect 12400 28704 12406 28756
rect 12710 28744 12716 28756
rect 12671 28716 12716 28744
rect 12710 28704 12716 28716
rect 12768 28744 12774 28756
rect 13078 28744 13084 28756
rect 12768 28716 13084 28744
rect 12768 28704 12774 28716
rect 13078 28704 13084 28716
rect 13136 28704 13142 28756
rect 13906 28744 13912 28756
rect 13819 28716 13912 28744
rect 13906 28704 13912 28716
rect 13964 28744 13970 28756
rect 14734 28744 14740 28756
rect 13964 28716 14740 28744
rect 13964 28704 13970 28716
rect 14734 28704 14740 28716
rect 14792 28704 14798 28756
rect 15841 28747 15899 28753
rect 15841 28713 15853 28747
rect 15887 28744 15899 28747
rect 16022 28744 16028 28756
rect 15887 28716 16028 28744
rect 15887 28713 15899 28716
rect 15841 28707 15899 28713
rect 16022 28704 16028 28716
rect 16080 28704 16086 28756
rect 16574 28744 16580 28756
rect 16408 28716 16580 28744
rect 1397 28679 1455 28685
rect 1397 28645 1409 28679
rect 1443 28676 1455 28679
rect 1670 28676 1676 28688
rect 1443 28648 1676 28676
rect 1443 28645 1455 28648
rect 1397 28639 1455 28645
rect 1670 28636 1676 28648
rect 1728 28636 1734 28688
rect 12618 28676 12624 28688
rect 11348 28648 12624 28676
rect 1578 28608 1584 28620
rect 1539 28580 1584 28608
rect 1578 28568 1584 28580
rect 1636 28568 1642 28620
rect 3602 28608 3608 28620
rect 3515 28580 3608 28608
rect 3602 28568 3608 28580
rect 3660 28608 3666 28620
rect 4706 28608 4712 28620
rect 3660 28580 4712 28608
rect 3660 28568 3666 28580
rect 1946 28540 1952 28552
rect 1907 28512 1952 28540
rect 1946 28500 1952 28512
rect 2004 28500 2010 28552
rect 4632 28481 4660 28580
rect 4706 28568 4712 28580
rect 4764 28568 4770 28620
rect 5258 28608 5264 28620
rect 5219 28580 5264 28608
rect 5258 28568 5264 28580
rect 5316 28608 5322 28620
rect 5810 28608 5816 28620
rect 5316 28580 5816 28608
rect 5316 28568 5322 28580
rect 5810 28568 5816 28580
rect 5868 28568 5874 28620
rect 5905 28611 5963 28617
rect 5905 28577 5917 28611
rect 5951 28608 5963 28611
rect 6917 28611 6975 28617
rect 6917 28608 6929 28611
rect 5951 28580 6929 28608
rect 5951 28577 5963 28580
rect 5905 28571 5963 28577
rect 6917 28577 6929 28580
rect 6963 28608 6975 28611
rect 7006 28608 7012 28620
rect 6963 28580 7012 28608
rect 6963 28577 6975 28580
rect 6917 28571 6975 28577
rect 7006 28568 7012 28580
rect 7064 28568 7070 28620
rect 8018 28608 8024 28620
rect 7979 28580 8024 28608
rect 8018 28568 8024 28580
rect 8076 28568 8082 28620
rect 8481 28611 8539 28617
rect 8481 28577 8493 28611
rect 8527 28608 8539 28611
rect 8662 28608 8668 28620
rect 8527 28580 8668 28608
rect 8527 28577 8539 28580
rect 8481 28571 8539 28577
rect 8662 28568 8668 28580
rect 8720 28568 8726 28620
rect 8846 28608 8852 28620
rect 8807 28580 8852 28608
rect 8846 28568 8852 28580
rect 8904 28568 8910 28620
rect 10134 28608 10140 28620
rect 10095 28580 10140 28608
rect 10134 28568 10140 28580
rect 10192 28608 10198 28620
rect 11348 28617 11376 28648
rect 12618 28636 12624 28648
rect 12676 28636 12682 28688
rect 13170 28636 13176 28688
rect 13228 28636 13234 28688
rect 15102 28676 15108 28688
rect 15063 28648 15108 28676
rect 15102 28636 15108 28648
rect 15160 28636 15166 28688
rect 15473 28679 15531 28685
rect 15473 28645 15485 28679
rect 15519 28676 15531 28679
rect 16298 28676 16304 28688
rect 15519 28648 16304 28676
rect 15519 28645 15531 28648
rect 15473 28639 15531 28645
rect 16298 28636 16304 28648
rect 16356 28636 16362 28688
rect 10597 28611 10655 28617
rect 10597 28608 10609 28611
rect 10192 28580 10609 28608
rect 10192 28568 10198 28580
rect 10597 28577 10609 28580
rect 10643 28577 10655 28611
rect 10597 28571 10655 28577
rect 11333 28611 11391 28617
rect 11333 28577 11345 28611
rect 11379 28577 11391 28611
rect 11333 28571 11391 28577
rect 12434 28568 12440 28620
rect 12492 28608 12498 28620
rect 12636 28608 12664 28636
rect 12897 28611 12955 28617
rect 12897 28608 12909 28611
rect 12492 28580 12537 28608
rect 12636 28580 12909 28608
rect 12492 28568 12498 28580
rect 12897 28577 12909 28580
rect 12943 28577 12955 28611
rect 13188 28608 13216 28636
rect 13265 28611 13323 28617
rect 13265 28608 13277 28611
rect 12897 28571 12955 28577
rect 13004 28580 13277 28608
rect 12066 28500 12072 28552
rect 12124 28540 12130 28552
rect 13004 28540 13032 28580
rect 13265 28577 13277 28580
rect 13311 28577 13323 28611
rect 14642 28608 14648 28620
rect 14603 28580 14648 28608
rect 13265 28571 13323 28577
rect 14642 28568 14648 28580
rect 14700 28568 14706 28620
rect 12124 28512 13032 28540
rect 16209 28543 16267 28549
rect 12124 28500 12130 28512
rect 16209 28509 16221 28543
rect 16255 28540 16267 28543
rect 16298 28540 16304 28552
rect 16255 28512 16304 28540
rect 16255 28509 16267 28512
rect 16209 28503 16267 28509
rect 16298 28500 16304 28512
rect 16356 28540 16362 28552
rect 16408 28540 16436 28716
rect 16574 28704 16580 28716
rect 16632 28704 16638 28756
rect 17773 28747 17831 28753
rect 17773 28744 17785 28747
rect 16684 28716 17785 28744
rect 16684 28688 16712 28716
rect 17773 28713 17785 28716
rect 17819 28713 17831 28747
rect 17773 28707 17831 28713
rect 16666 28676 16672 28688
rect 16500 28648 16672 28676
rect 16500 28617 16528 28648
rect 16666 28636 16672 28648
rect 16724 28636 16730 28688
rect 17129 28679 17187 28685
rect 17129 28645 17141 28679
rect 17175 28676 17187 28679
rect 17218 28676 17224 28688
rect 17175 28648 17224 28676
rect 17175 28645 17187 28648
rect 17129 28639 17187 28645
rect 17218 28636 17224 28648
rect 17276 28636 17282 28688
rect 16485 28611 16543 28617
rect 16485 28577 16497 28611
rect 16531 28577 16543 28611
rect 16485 28571 16543 28577
rect 16574 28568 16580 28620
rect 16632 28608 16638 28620
rect 16853 28611 16911 28617
rect 16853 28608 16865 28611
rect 16632 28580 16865 28608
rect 16632 28568 16638 28580
rect 16853 28577 16865 28580
rect 16899 28608 16911 28611
rect 17494 28608 17500 28620
rect 16899 28580 17500 28608
rect 16899 28577 16911 28580
rect 16853 28571 16911 28577
rect 17494 28568 17500 28580
rect 17552 28568 17558 28620
rect 16356 28512 16436 28540
rect 16356 28500 16362 28512
rect 4617 28475 4675 28481
rect 4617 28441 4629 28475
rect 4663 28472 4675 28475
rect 5718 28472 5724 28484
rect 4663 28444 5724 28472
rect 4663 28441 4675 28444
rect 4617 28435 4675 28441
rect 5718 28432 5724 28444
rect 5776 28432 5782 28484
rect 8294 28432 8300 28484
rect 8352 28472 8358 28484
rect 8757 28475 8815 28481
rect 8757 28472 8769 28475
rect 8352 28444 8769 28472
rect 8352 28432 8358 28444
rect 8757 28441 8769 28444
rect 8803 28441 8815 28475
rect 8757 28435 8815 28441
rect 11517 28475 11575 28481
rect 11517 28441 11529 28475
rect 11563 28472 11575 28475
rect 12526 28472 12532 28484
rect 11563 28444 12532 28472
rect 11563 28441 11575 28444
rect 11517 28435 11575 28441
rect 12526 28432 12532 28444
rect 12584 28432 12590 28484
rect 11885 28407 11943 28413
rect 11885 28373 11897 28407
rect 11931 28404 11943 28407
rect 12066 28404 12072 28416
rect 11931 28376 12072 28404
rect 11931 28373 11943 28376
rect 11885 28367 11943 28373
rect 12066 28364 12072 28376
rect 12124 28364 12130 28416
rect 17402 28404 17408 28416
rect 17363 28376 17408 28404
rect 17402 28364 17408 28376
rect 17460 28364 17466 28416
rect 1104 28314 18860 28336
rect 1104 28262 4315 28314
rect 4367 28262 4379 28314
rect 4431 28262 4443 28314
rect 4495 28262 4507 28314
rect 4559 28262 10982 28314
rect 11034 28262 11046 28314
rect 11098 28262 11110 28314
rect 11162 28262 11174 28314
rect 11226 28262 17648 28314
rect 17700 28262 17712 28314
rect 17764 28262 17776 28314
rect 17828 28262 17840 28314
rect 17892 28262 18860 28314
rect 1104 28240 18860 28262
rect 1578 28160 1584 28212
rect 1636 28200 1642 28212
rect 1949 28203 2007 28209
rect 1949 28200 1961 28203
rect 1636 28172 1961 28200
rect 1636 28160 1642 28172
rect 1949 28169 1961 28172
rect 1995 28169 2007 28203
rect 1949 28163 2007 28169
rect 2409 28203 2467 28209
rect 2409 28169 2421 28203
rect 2455 28200 2467 28203
rect 2590 28200 2596 28212
rect 2455 28172 2596 28200
rect 2455 28169 2467 28172
rect 2409 28163 2467 28169
rect 2590 28160 2596 28172
rect 2648 28160 2654 28212
rect 3513 28203 3571 28209
rect 3513 28169 3525 28203
rect 3559 28200 3571 28203
rect 3602 28200 3608 28212
rect 3559 28172 3608 28200
rect 3559 28169 3571 28172
rect 3513 28163 3571 28169
rect 3602 28160 3608 28172
rect 3660 28160 3666 28212
rect 7653 28203 7711 28209
rect 7653 28169 7665 28203
rect 7699 28200 7711 28203
rect 8018 28200 8024 28212
rect 7699 28172 8024 28200
rect 7699 28169 7711 28172
rect 7653 28163 7711 28169
rect 8018 28160 8024 28172
rect 8076 28160 8082 28212
rect 8662 28200 8668 28212
rect 8128 28172 8668 28200
rect 7285 28135 7343 28141
rect 7285 28101 7297 28135
rect 7331 28132 7343 28135
rect 8128 28132 8156 28172
rect 8662 28160 8668 28172
rect 8720 28160 8726 28212
rect 8846 28160 8852 28212
rect 8904 28200 8910 28212
rect 9033 28203 9091 28209
rect 9033 28200 9045 28203
rect 8904 28172 9045 28200
rect 8904 28160 8910 28172
rect 9033 28169 9045 28172
rect 9079 28169 9091 28203
rect 9398 28200 9404 28212
rect 9359 28172 9404 28200
rect 9033 28163 9091 28169
rect 9398 28160 9404 28172
rect 9456 28160 9462 28212
rect 15930 28160 15936 28212
rect 15988 28200 15994 28212
rect 16117 28203 16175 28209
rect 16117 28200 16129 28203
rect 15988 28172 16129 28200
rect 15988 28160 15994 28172
rect 16117 28169 16129 28172
rect 16163 28169 16175 28203
rect 16117 28163 16175 28169
rect 8386 28132 8392 28144
rect 7331 28104 8156 28132
rect 8299 28104 8392 28132
rect 7331 28101 7343 28104
rect 7285 28095 7343 28101
rect 1670 28064 1676 28076
rect 1631 28036 1676 28064
rect 1670 28024 1676 28036
rect 1728 28024 1734 28076
rect 6641 28067 6699 28073
rect 6641 28033 6653 28067
rect 6687 28064 6699 28067
rect 6730 28064 6736 28076
rect 6687 28036 6736 28064
rect 6687 28033 6699 28036
rect 6641 28027 6699 28033
rect 6730 28024 6736 28036
rect 6788 28024 6794 28076
rect 8312 28073 8340 28104
rect 8386 28092 8392 28104
rect 8444 28132 8450 28144
rect 8864 28132 8892 28160
rect 8444 28104 8892 28132
rect 8444 28092 8450 28104
rect 8297 28067 8355 28073
rect 8297 28033 8309 28067
rect 8343 28033 8355 28067
rect 8297 28027 8355 28033
rect 8757 28067 8815 28073
rect 8757 28033 8769 28067
rect 8803 28064 8815 28067
rect 9416 28064 9444 28160
rect 8803 28036 9444 28064
rect 12069 28067 12127 28073
rect 8803 28033 8815 28036
rect 8757 28027 8815 28033
rect 12069 28033 12081 28067
rect 12115 28064 12127 28067
rect 12342 28064 12348 28076
rect 12115 28036 12348 28064
rect 12115 28033 12127 28036
rect 12069 28027 12127 28033
rect 12342 28024 12348 28036
rect 12400 28024 12406 28076
rect 13354 28064 13360 28076
rect 13188 28036 13360 28064
rect 3881 27999 3939 28005
rect 3881 27965 3893 27999
rect 3927 27996 3939 27999
rect 4706 27996 4712 28008
rect 3927 27968 4712 27996
rect 3927 27965 3939 27968
rect 3881 27959 3939 27965
rect 4706 27956 4712 27968
rect 4764 27956 4770 28008
rect 5813 27999 5871 28005
rect 5813 27965 5825 27999
rect 5859 27996 5871 27999
rect 5902 27996 5908 28008
rect 5859 27968 5908 27996
rect 5859 27965 5871 27968
rect 5813 27959 5871 27965
rect 5902 27956 5908 27968
rect 5960 27956 5966 28008
rect 6086 27956 6092 28008
rect 6144 27996 6150 28008
rect 6181 27999 6239 28005
rect 6181 27996 6193 27999
rect 6144 27968 6193 27996
rect 6144 27956 6150 27968
rect 6181 27965 6193 27968
rect 6227 27965 6239 27999
rect 6181 27959 6239 27965
rect 8573 27999 8631 28005
rect 8573 27965 8585 27999
rect 8619 27996 8631 27999
rect 9030 27996 9036 28008
rect 8619 27968 9036 27996
rect 8619 27965 8631 27968
rect 8573 27959 8631 27965
rect 9030 27956 9036 27968
rect 9088 27956 9094 28008
rect 10873 27999 10931 28005
rect 10873 27965 10885 27999
rect 10919 27996 10931 27999
rect 11882 27996 11888 28008
rect 10919 27968 11888 27996
rect 10919 27965 10931 27968
rect 10873 27959 10931 27965
rect 11882 27956 11888 27968
rect 11940 27996 11946 28008
rect 12434 27996 12440 28008
rect 11940 27968 12440 27996
rect 11940 27956 11946 27968
rect 12434 27956 12440 27968
rect 12492 27956 12498 28008
rect 12894 27996 12900 28008
rect 12855 27968 12900 27996
rect 12894 27956 12900 27968
rect 12952 27956 12958 28008
rect 13188 28005 13216 28036
rect 13354 28024 13360 28036
rect 13412 28024 13418 28076
rect 14645 28067 14703 28073
rect 14645 28064 14657 28067
rect 13464 28036 14657 28064
rect 13173 27999 13231 28005
rect 13173 27965 13185 27999
rect 13219 27965 13231 27999
rect 13173 27959 13231 27965
rect 13262 27956 13268 28008
rect 13320 27996 13326 28008
rect 13464 28005 13492 28036
rect 14645 28033 14657 28036
rect 14691 28033 14703 28067
rect 14645 28027 14703 28033
rect 15289 28067 15347 28073
rect 15289 28033 15301 28067
rect 15335 28064 15347 28067
rect 15948 28064 15976 28160
rect 17770 28064 17776 28076
rect 15335 28036 15976 28064
rect 17731 28036 17776 28064
rect 15335 28033 15347 28036
rect 15289 28027 15347 28033
rect 17770 28024 17776 28036
rect 17828 28024 17834 28076
rect 13449 27999 13507 28005
rect 13449 27996 13461 27999
rect 13320 27968 13461 27996
rect 13320 27956 13326 27968
rect 13449 27965 13461 27968
rect 13495 27965 13507 27999
rect 13449 27959 13507 27965
rect 13633 27999 13691 28005
rect 13633 27965 13645 27999
rect 13679 27965 13691 27999
rect 13906 27996 13912 28008
rect 13867 27968 13912 27996
rect 13633 27959 13691 27965
rect 7466 27888 7472 27940
rect 7524 27928 7530 27940
rect 7745 27931 7803 27937
rect 7745 27928 7757 27931
rect 7524 27900 7757 27928
rect 7524 27888 7530 27900
rect 7745 27897 7757 27900
rect 7791 27897 7803 27931
rect 13648 27928 13676 27959
rect 13906 27956 13912 27968
rect 13964 27956 13970 28008
rect 14369 27999 14427 28005
rect 14369 27965 14381 27999
rect 14415 27996 14427 27999
rect 15378 27996 15384 28008
rect 14415 27968 15384 27996
rect 14415 27965 14427 27968
rect 14369 27959 14427 27965
rect 15378 27956 15384 27968
rect 15436 27956 15442 28008
rect 16669 27999 16727 28005
rect 16669 27965 16681 27999
rect 16715 27965 16727 27999
rect 16669 27959 16727 27965
rect 17221 27999 17279 28005
rect 17221 27965 17233 27999
rect 17267 27996 17279 27999
rect 17310 27996 17316 28008
rect 17267 27968 17316 27996
rect 17267 27965 17279 27968
rect 17221 27959 17279 27965
rect 15838 27928 15844 27940
rect 7745 27891 7803 27897
rect 13004 27900 13676 27928
rect 15799 27900 15844 27928
rect 13004 27872 13032 27900
rect 15838 27888 15844 27900
rect 15896 27888 15902 27940
rect 16298 27888 16304 27940
rect 16356 27928 16362 27940
rect 16485 27931 16543 27937
rect 16485 27928 16497 27931
rect 16356 27900 16497 27928
rect 16356 27888 16362 27900
rect 16485 27897 16497 27900
rect 16531 27928 16543 27931
rect 16684 27928 16712 27959
rect 17310 27956 17316 27968
rect 17368 27956 17374 28008
rect 17402 27956 17408 28008
rect 17460 27996 17466 28008
rect 17497 27999 17555 28005
rect 17497 27996 17509 27999
rect 17460 27968 17509 27996
rect 17460 27956 17466 27968
rect 17497 27965 17509 27968
rect 17543 27965 17555 27999
rect 17497 27959 17555 27965
rect 16531 27900 16712 27928
rect 17328 27928 17356 27956
rect 18049 27931 18107 27937
rect 18049 27928 18061 27931
rect 17328 27900 18061 27928
rect 16531 27897 16543 27900
rect 16485 27891 16543 27897
rect 18049 27897 18061 27900
rect 18095 27897 18107 27931
rect 18049 27891 18107 27897
rect 4338 27860 4344 27872
rect 4299 27832 4344 27860
rect 4338 27820 4344 27832
rect 4396 27820 4402 27872
rect 5258 27860 5264 27872
rect 5219 27832 5264 27860
rect 5258 27820 5264 27832
rect 5316 27820 5322 27872
rect 5626 27820 5632 27872
rect 5684 27860 5690 27872
rect 5721 27863 5779 27869
rect 5721 27860 5733 27863
rect 5684 27832 5733 27860
rect 5684 27820 5690 27832
rect 5721 27829 5733 27832
rect 5767 27829 5779 27863
rect 5721 27823 5779 27829
rect 9214 27820 9220 27872
rect 9272 27860 9278 27872
rect 10134 27860 10140 27872
rect 9272 27832 10140 27860
rect 9272 27820 9278 27832
rect 10134 27820 10140 27832
rect 10192 27820 10198 27872
rect 11241 27863 11299 27869
rect 11241 27829 11253 27863
rect 11287 27860 11299 27863
rect 12437 27863 12495 27869
rect 12437 27860 12449 27863
rect 11287 27832 12449 27860
rect 11287 27829 11299 27832
rect 11241 27823 11299 27829
rect 12437 27829 12449 27832
rect 12483 27860 12495 27863
rect 12618 27860 12624 27872
rect 12483 27832 12624 27860
rect 12483 27829 12495 27832
rect 12437 27823 12495 27829
rect 12618 27820 12624 27832
rect 12676 27820 12682 27872
rect 12805 27863 12863 27869
rect 12805 27829 12817 27863
rect 12851 27860 12863 27863
rect 12986 27860 12992 27872
rect 12851 27832 12992 27860
rect 12851 27829 12863 27832
rect 12805 27823 12863 27829
rect 12986 27820 12992 27832
rect 13044 27820 13050 27872
rect 13814 27820 13820 27872
rect 13872 27860 13878 27872
rect 14642 27860 14648 27872
rect 13872 27832 14648 27860
rect 13872 27820 13878 27832
rect 14642 27820 14648 27832
rect 14700 27860 14706 27872
rect 15013 27863 15071 27869
rect 15013 27860 15025 27863
rect 14700 27832 15025 27860
rect 14700 27820 14706 27832
rect 15013 27829 15025 27832
rect 15059 27829 15071 27863
rect 15013 27823 15071 27829
rect 1104 27770 18860 27792
rect 1104 27718 7648 27770
rect 7700 27718 7712 27770
rect 7764 27718 7776 27770
rect 7828 27718 7840 27770
rect 7892 27718 14315 27770
rect 14367 27718 14379 27770
rect 14431 27718 14443 27770
rect 14495 27718 14507 27770
rect 14559 27718 18860 27770
rect 1104 27696 18860 27718
rect 5721 27659 5779 27665
rect 5721 27625 5733 27659
rect 5767 27656 5779 27659
rect 5902 27656 5908 27668
rect 5767 27628 5908 27656
rect 5767 27625 5779 27628
rect 5721 27619 5779 27625
rect 5902 27616 5908 27628
rect 5960 27616 5966 27668
rect 7006 27656 7012 27668
rect 6967 27628 7012 27656
rect 7006 27616 7012 27628
rect 7064 27656 7070 27668
rect 8294 27656 8300 27668
rect 7064 27628 7328 27656
rect 7064 27616 7070 27628
rect 3697 27591 3755 27597
rect 3697 27557 3709 27591
rect 3743 27588 3755 27591
rect 4154 27588 4160 27600
rect 3743 27560 4160 27588
rect 3743 27557 3755 27560
rect 3697 27551 3755 27557
rect 4154 27548 4160 27560
rect 4212 27588 4218 27600
rect 4338 27588 4344 27600
rect 4212 27560 4344 27588
rect 4212 27548 4218 27560
rect 4338 27548 4344 27560
rect 4396 27548 4402 27600
rect 5166 27548 5172 27600
rect 5224 27588 5230 27600
rect 5261 27591 5319 27597
rect 5261 27588 5273 27591
rect 5224 27560 5273 27588
rect 5224 27548 5230 27560
rect 5261 27557 5273 27560
rect 5307 27557 5319 27591
rect 5261 27551 5319 27557
rect 6641 27591 6699 27597
rect 6641 27557 6653 27591
rect 6687 27588 6699 27591
rect 7098 27588 7104 27600
rect 6687 27560 7104 27588
rect 6687 27557 6699 27560
rect 6641 27551 6699 27557
rect 7098 27548 7104 27560
rect 7156 27548 7162 27600
rect 7300 27588 7328 27628
rect 8220 27628 8300 27656
rect 7926 27588 7932 27600
rect 7300 27560 7932 27588
rect 1949 27523 2007 27529
rect 1949 27489 1961 27523
rect 1995 27520 2007 27523
rect 2038 27520 2044 27532
rect 1995 27492 2044 27520
rect 1995 27489 2007 27492
rect 1949 27483 2007 27489
rect 2038 27480 2044 27492
rect 2096 27480 2102 27532
rect 3510 27480 3516 27532
rect 3568 27520 3574 27532
rect 4249 27523 4307 27529
rect 4249 27520 4261 27523
rect 3568 27492 4261 27520
rect 3568 27480 3574 27492
rect 4249 27489 4261 27492
rect 4295 27489 4307 27523
rect 4706 27520 4712 27532
rect 4667 27492 4712 27520
rect 4249 27483 4307 27489
rect 4706 27480 4712 27492
rect 4764 27480 4770 27532
rect 7300 27529 7328 27560
rect 7926 27548 7932 27560
rect 7984 27548 7990 27600
rect 4985 27523 5043 27529
rect 4985 27489 4997 27523
rect 5031 27489 5043 27523
rect 4985 27483 5043 27489
rect 7285 27523 7343 27529
rect 7285 27489 7297 27523
rect 7331 27489 7343 27523
rect 8018 27520 8024 27532
rect 7931 27492 8024 27520
rect 7285 27483 7343 27489
rect 1670 27452 1676 27464
rect 1583 27424 1676 27452
rect 1670 27412 1676 27424
rect 1728 27452 1734 27464
rect 2590 27452 2596 27464
rect 1728 27424 2596 27452
rect 1728 27412 1734 27424
rect 2590 27412 2596 27424
rect 2648 27412 2654 27464
rect 2774 27412 2780 27464
rect 2832 27452 2838 27464
rect 4065 27455 4123 27461
rect 4065 27452 4077 27455
rect 2832 27424 4077 27452
rect 2832 27412 2838 27424
rect 4065 27421 4077 27424
rect 4111 27452 4123 27455
rect 5000 27452 5028 27483
rect 8018 27480 8024 27492
rect 8076 27520 8082 27532
rect 8220 27520 8248 27628
rect 8294 27616 8300 27628
rect 8352 27616 8358 27668
rect 8386 27616 8392 27668
rect 8444 27656 8450 27668
rect 8757 27659 8815 27665
rect 8444 27628 8489 27656
rect 8444 27616 8450 27628
rect 8757 27625 8769 27659
rect 8803 27656 8815 27659
rect 9030 27656 9036 27668
rect 8803 27628 9036 27656
rect 8803 27625 8815 27628
rect 8757 27619 8815 27625
rect 9030 27616 9036 27628
rect 9088 27616 9094 27668
rect 11330 27616 11336 27668
rect 11388 27656 11394 27668
rect 12161 27659 12219 27665
rect 12161 27656 12173 27659
rect 11388 27628 12173 27656
rect 11388 27616 11394 27628
rect 12161 27625 12173 27628
rect 12207 27656 12219 27659
rect 12894 27656 12900 27668
rect 12207 27628 12900 27656
rect 12207 27625 12219 27628
rect 12161 27619 12219 27625
rect 12894 27616 12900 27628
rect 12952 27616 12958 27668
rect 15378 27656 15384 27668
rect 15339 27628 15384 27656
rect 15378 27616 15384 27628
rect 15436 27616 15442 27668
rect 16298 27616 16304 27668
rect 16356 27656 16362 27668
rect 16850 27656 16856 27668
rect 16356 27628 16856 27656
rect 16356 27616 16362 27628
rect 16850 27616 16856 27628
rect 16908 27656 16914 27668
rect 17405 27659 17463 27665
rect 17405 27656 17417 27659
rect 16908 27628 17417 27656
rect 16908 27616 16914 27628
rect 17405 27625 17417 27628
rect 17451 27625 17463 27659
rect 17405 27619 17463 27625
rect 13262 27588 13268 27600
rect 13223 27560 13268 27588
rect 13262 27548 13268 27560
rect 13320 27548 13326 27600
rect 16025 27591 16083 27597
rect 16025 27557 16037 27591
rect 16071 27588 16083 27591
rect 16206 27588 16212 27600
rect 16071 27560 16212 27588
rect 16071 27557 16083 27560
rect 16025 27551 16083 27557
rect 16206 27548 16212 27560
rect 16264 27548 16270 27600
rect 17126 27588 17132 27600
rect 16960 27560 17132 27588
rect 10318 27520 10324 27532
rect 8076 27492 8248 27520
rect 10279 27492 10324 27520
rect 8076 27480 8082 27492
rect 10318 27480 10324 27492
rect 10376 27480 10382 27532
rect 11330 27520 11336 27532
rect 11291 27492 11336 27520
rect 11330 27480 11336 27492
rect 11388 27480 11394 27532
rect 12710 27520 12716 27532
rect 12671 27492 12716 27520
rect 12710 27480 12716 27492
rect 12768 27480 12774 27532
rect 13814 27480 13820 27532
rect 13872 27520 13878 27532
rect 14093 27523 14151 27529
rect 14093 27520 14105 27523
rect 13872 27492 14105 27520
rect 13872 27480 13878 27492
rect 14093 27489 14105 27492
rect 14139 27489 14151 27523
rect 14093 27483 14151 27489
rect 14182 27480 14188 27532
rect 14240 27520 14246 27532
rect 14553 27523 14611 27529
rect 14553 27520 14565 27523
rect 14240 27492 14565 27520
rect 14240 27480 14246 27492
rect 14553 27489 14565 27492
rect 14599 27520 14611 27523
rect 15010 27520 15016 27532
rect 14599 27492 15016 27520
rect 14599 27489 14611 27492
rect 14553 27483 14611 27489
rect 15010 27480 15016 27492
rect 15068 27480 15074 27532
rect 16224 27520 16252 27548
rect 16960 27529 16988 27560
rect 17126 27548 17132 27560
rect 17184 27588 17190 27600
rect 17586 27588 17592 27600
rect 17184 27560 17592 27588
rect 17184 27548 17190 27560
rect 17586 27548 17592 27560
rect 17644 27548 17650 27600
rect 16669 27523 16727 27529
rect 16669 27520 16681 27523
rect 16224 27492 16681 27520
rect 16669 27489 16681 27492
rect 16715 27489 16727 27523
rect 16669 27483 16727 27489
rect 16945 27523 17003 27529
rect 16945 27489 16957 27523
rect 16991 27489 17003 27523
rect 17402 27520 17408 27532
rect 16945 27483 17003 27489
rect 17052 27492 17408 27520
rect 14642 27452 14648 27464
rect 4111 27424 5028 27452
rect 14603 27424 14648 27452
rect 4111 27421 4123 27424
rect 4065 27415 4123 27421
rect 14642 27412 14648 27424
rect 14700 27412 14706 27464
rect 16117 27455 16175 27461
rect 16117 27421 16129 27455
rect 16163 27452 16175 27455
rect 17052 27452 17080 27492
rect 17402 27480 17408 27492
rect 17460 27480 17466 27532
rect 16163 27424 17080 27452
rect 17129 27455 17187 27461
rect 16163 27421 16175 27424
rect 16117 27415 16175 27421
rect 17129 27421 17141 27455
rect 17175 27452 17187 27455
rect 17310 27452 17316 27464
rect 17175 27424 17316 27452
rect 17175 27421 17187 27424
rect 17129 27415 17187 27421
rect 17310 27412 17316 27424
rect 17368 27412 17374 27464
rect 11517 27387 11575 27393
rect 11517 27353 11529 27387
rect 11563 27384 11575 27387
rect 12710 27384 12716 27396
rect 11563 27356 12716 27384
rect 11563 27353 11575 27356
rect 11517 27347 11575 27353
rect 12710 27344 12716 27356
rect 12768 27344 12774 27396
rect 16022 27344 16028 27396
rect 16080 27384 16086 27396
rect 16482 27384 16488 27396
rect 16080 27356 16488 27384
rect 16080 27344 16086 27356
rect 16482 27344 16488 27356
rect 16540 27344 16546 27396
rect 16574 27344 16580 27396
rect 16632 27384 16638 27396
rect 17773 27387 17831 27393
rect 17773 27384 17785 27387
rect 16632 27356 17785 27384
rect 16632 27344 16638 27356
rect 17773 27353 17785 27356
rect 17819 27353 17831 27387
rect 17773 27347 17831 27353
rect 3237 27319 3295 27325
rect 3237 27285 3249 27319
rect 3283 27316 3295 27319
rect 3418 27316 3424 27328
rect 3283 27288 3424 27316
rect 3283 27285 3295 27288
rect 3237 27279 3295 27285
rect 3418 27276 3424 27288
rect 3476 27276 3482 27328
rect 6086 27316 6092 27328
rect 6047 27288 6092 27316
rect 6086 27276 6092 27288
rect 6144 27276 6150 27328
rect 7374 27316 7380 27328
rect 7335 27288 7380 27316
rect 7374 27276 7380 27288
rect 7432 27276 7438 27328
rect 8294 27276 8300 27328
rect 8352 27316 8358 27328
rect 8754 27316 8760 27328
rect 8352 27288 8760 27316
rect 8352 27276 8358 27288
rect 8754 27276 8760 27288
rect 8812 27276 8818 27328
rect 10502 27316 10508 27328
rect 10463 27288 10508 27316
rect 10502 27276 10508 27288
rect 10560 27276 10566 27328
rect 11882 27316 11888 27328
rect 11843 27288 11888 27316
rect 11882 27276 11888 27288
rect 11940 27276 11946 27328
rect 13354 27276 13360 27328
rect 13412 27316 13418 27328
rect 13541 27319 13599 27325
rect 13541 27316 13553 27319
rect 13412 27288 13553 27316
rect 13412 27276 13418 27288
rect 13541 27285 13553 27288
rect 13587 27285 13599 27319
rect 13906 27316 13912 27328
rect 13867 27288 13912 27316
rect 13541 27279 13599 27285
rect 13906 27276 13912 27288
rect 13964 27276 13970 27328
rect 1104 27226 18860 27248
rect 1104 27174 4315 27226
rect 4367 27174 4379 27226
rect 4431 27174 4443 27226
rect 4495 27174 4507 27226
rect 4559 27174 10982 27226
rect 11034 27174 11046 27226
rect 11098 27174 11110 27226
rect 11162 27174 11174 27226
rect 11226 27174 17648 27226
rect 17700 27174 17712 27226
rect 17764 27174 17776 27226
rect 17828 27174 17840 27226
rect 17892 27174 18860 27226
rect 1104 27152 18860 27174
rect 1765 27115 1823 27121
rect 1765 27081 1777 27115
rect 1811 27112 1823 27115
rect 2038 27112 2044 27124
rect 1811 27084 2044 27112
rect 1811 27081 1823 27084
rect 1765 27075 1823 27081
rect 2038 27072 2044 27084
rect 2096 27072 2102 27124
rect 3510 27112 3516 27124
rect 3471 27084 3516 27112
rect 3510 27072 3516 27084
rect 3568 27072 3574 27124
rect 3881 27115 3939 27121
rect 3881 27081 3893 27115
rect 3927 27112 3939 27115
rect 4706 27112 4712 27124
rect 3927 27084 4712 27112
rect 3927 27081 3939 27084
rect 3881 27075 3939 27081
rect 4706 27072 4712 27084
rect 4764 27072 4770 27124
rect 6457 27115 6515 27121
rect 6457 27081 6469 27115
rect 6503 27112 6515 27115
rect 8018 27112 8024 27124
rect 6503 27084 8024 27112
rect 6503 27081 6515 27084
rect 6457 27075 6515 27081
rect 8018 27072 8024 27084
rect 8076 27072 8082 27124
rect 10318 27072 10324 27124
rect 10376 27112 10382 27124
rect 10413 27115 10471 27121
rect 10413 27112 10425 27115
rect 10376 27084 10425 27112
rect 10376 27072 10382 27084
rect 10413 27081 10425 27084
rect 10459 27112 10471 27115
rect 12161 27115 12219 27121
rect 12161 27112 12173 27115
rect 10459 27084 12173 27112
rect 10459 27081 10471 27084
rect 10413 27075 10471 27081
rect 12161 27081 12173 27084
rect 12207 27081 12219 27115
rect 12710 27112 12716 27124
rect 12671 27084 12716 27112
rect 12161 27075 12219 27081
rect 12710 27072 12716 27084
rect 12768 27072 12774 27124
rect 13538 27112 13544 27124
rect 13451 27084 13544 27112
rect 13538 27072 13544 27084
rect 13596 27112 13602 27124
rect 14182 27112 14188 27124
rect 13596 27084 14188 27112
rect 13596 27072 13602 27084
rect 14182 27072 14188 27084
rect 14240 27072 14246 27124
rect 15565 27115 15623 27121
rect 15565 27081 15577 27115
rect 15611 27112 15623 27115
rect 17126 27112 17132 27124
rect 15611 27084 17132 27112
rect 15611 27081 15623 27084
rect 15565 27075 15623 27081
rect 17126 27072 17132 27084
rect 17184 27072 17190 27124
rect 3326 27044 3332 27056
rect 2700 27016 3332 27044
rect 2700 26917 2728 27016
rect 3326 27004 3332 27016
rect 3384 27004 3390 27056
rect 6086 27004 6092 27056
rect 6144 27044 6150 27056
rect 7837 27047 7895 27053
rect 7837 27044 7849 27047
rect 6144 27016 7849 27044
rect 6144 27004 6150 27016
rect 7837 27013 7849 27016
rect 7883 27013 7895 27047
rect 7837 27007 7895 27013
rect 7926 27004 7932 27056
rect 7984 27044 7990 27056
rect 8389 27047 8447 27053
rect 8389 27044 8401 27047
rect 7984 27016 8401 27044
rect 7984 27004 7990 27016
rect 8389 27013 8401 27016
rect 8435 27013 8447 27047
rect 8389 27007 8447 27013
rect 11701 27047 11759 27053
rect 11701 27013 11713 27047
rect 11747 27044 11759 27047
rect 11790 27044 11796 27056
rect 11747 27016 11796 27044
rect 11747 27013 11759 27016
rect 11701 27007 11759 27013
rect 11790 27004 11796 27016
rect 11848 27004 11854 27056
rect 15841 27047 15899 27053
rect 15841 27013 15853 27047
rect 15887 27044 15899 27047
rect 16482 27044 16488 27056
rect 15887 27016 16488 27044
rect 15887 27013 15899 27016
rect 15841 27007 15899 27013
rect 16482 27004 16488 27016
rect 16540 27004 16546 27056
rect 17494 27044 17500 27056
rect 17455 27016 17500 27044
rect 17494 27004 17500 27016
rect 17552 27004 17558 27056
rect 2774 26936 2780 26988
rect 2832 26976 2838 26988
rect 5445 26979 5503 26985
rect 5445 26976 5457 26979
rect 2832 26948 2877 26976
rect 3160 26948 5457 26976
rect 2832 26936 2838 26948
rect 2317 26911 2375 26917
rect 2317 26877 2329 26911
rect 2363 26908 2375 26911
rect 2685 26911 2743 26917
rect 2685 26908 2697 26911
rect 2363 26880 2697 26908
rect 2363 26877 2375 26880
rect 2317 26871 2375 26877
rect 2685 26877 2697 26880
rect 2731 26877 2743 26911
rect 2685 26871 2743 26877
rect 2866 26868 2872 26920
rect 2924 26908 2930 26920
rect 3160 26917 3188 26948
rect 5445 26945 5457 26948
rect 5491 26945 5503 26979
rect 5445 26939 5503 26945
rect 7193 26979 7251 26985
rect 7193 26945 7205 26979
rect 7239 26976 7251 26979
rect 8662 26976 8668 26988
rect 7239 26948 8668 26976
rect 7239 26945 7251 26948
rect 7193 26939 7251 26945
rect 8662 26936 8668 26948
rect 8720 26976 8726 26988
rect 8757 26979 8815 26985
rect 8757 26976 8769 26979
rect 8720 26948 8769 26976
rect 8720 26936 8726 26948
rect 8757 26945 8769 26948
rect 8803 26945 8815 26979
rect 11241 26979 11299 26985
rect 11241 26976 11253 26979
rect 8757 26939 8815 26945
rect 10704 26948 11253 26976
rect 3145 26911 3203 26917
rect 3145 26908 3157 26911
rect 2924 26880 3157 26908
rect 2924 26868 2930 26880
rect 3145 26877 3157 26880
rect 3191 26877 3203 26911
rect 3145 26871 3203 26877
rect 3602 26868 3608 26920
rect 3660 26908 3666 26920
rect 4065 26911 4123 26917
rect 4065 26908 4077 26911
rect 3660 26880 4077 26908
rect 3660 26868 3666 26880
rect 4065 26877 4077 26880
rect 4111 26877 4123 26911
rect 4065 26871 4123 26877
rect 4154 26868 4160 26920
rect 4212 26908 4218 26920
rect 4341 26911 4399 26917
rect 4341 26908 4353 26911
rect 4212 26880 4353 26908
rect 4212 26868 4218 26880
rect 4341 26877 4353 26880
rect 4387 26877 4399 26911
rect 4341 26871 4399 26877
rect 4982 26868 4988 26920
rect 5040 26908 5046 26920
rect 6089 26911 6147 26917
rect 6089 26908 6101 26911
rect 5040 26880 6101 26908
rect 5040 26868 5046 26880
rect 6089 26877 6101 26880
rect 6135 26908 6147 26911
rect 6733 26911 6791 26917
rect 6733 26908 6745 26911
rect 6135 26880 6745 26908
rect 6135 26877 6147 26880
rect 6089 26871 6147 26877
rect 6733 26877 6745 26880
rect 6779 26877 6791 26911
rect 7466 26908 7472 26920
rect 7427 26880 7472 26908
rect 6733 26871 6791 26877
rect 7466 26868 7472 26880
rect 7524 26868 7530 26920
rect 10704 26917 10732 26948
rect 11241 26945 11253 26948
rect 11287 26976 11299 26979
rect 13262 26976 13268 26988
rect 11287 26948 13268 26976
rect 11287 26945 11299 26948
rect 11241 26939 11299 26945
rect 13262 26936 13268 26948
rect 13320 26936 13326 26988
rect 16850 26976 16856 26988
rect 16811 26948 16856 26976
rect 16850 26936 16856 26948
rect 16908 26936 16914 26988
rect 18049 26979 18107 26985
rect 18049 26976 18061 26979
rect 17052 26948 18061 26976
rect 17052 26920 17080 26948
rect 18049 26945 18061 26948
rect 18095 26945 18107 26979
rect 18049 26939 18107 26945
rect 7837 26911 7895 26917
rect 7837 26877 7849 26911
rect 7883 26877 7895 26911
rect 7837 26871 7895 26877
rect 10689 26911 10747 26917
rect 10689 26877 10701 26911
rect 10735 26877 10747 26911
rect 10689 26871 10747 26877
rect 5718 26800 5724 26852
rect 5776 26840 5782 26852
rect 5776 26812 6592 26840
rect 5776 26800 5782 26812
rect 6564 26781 6592 26812
rect 7098 26800 7104 26852
rect 7156 26840 7162 26852
rect 7852 26840 7880 26871
rect 11146 26868 11152 26920
rect 11204 26908 11210 26920
rect 11977 26911 12035 26917
rect 11977 26908 11989 26911
rect 11204 26880 11989 26908
rect 11204 26868 11210 26880
rect 11977 26877 11989 26880
rect 12023 26877 12035 26911
rect 13906 26908 13912 26920
rect 13867 26880 13912 26908
rect 11977 26871 12035 26877
rect 13906 26868 13912 26880
rect 13964 26868 13970 26920
rect 14182 26908 14188 26920
rect 14143 26880 14188 26908
rect 14182 26868 14188 26880
rect 14240 26868 14246 26920
rect 15657 26911 15715 26917
rect 15657 26877 15669 26911
rect 15703 26908 15715 26911
rect 17034 26908 17040 26920
rect 15703 26880 16068 26908
rect 16995 26880 17040 26908
rect 15703 26877 15715 26880
rect 15657 26871 15715 26877
rect 11882 26840 11888 26852
rect 7156 26812 7880 26840
rect 11843 26812 11888 26840
rect 7156 26800 7162 26812
rect 11882 26800 11888 26812
rect 11940 26800 11946 26852
rect 13173 26843 13231 26849
rect 13173 26809 13185 26843
rect 13219 26840 13231 26843
rect 14200 26840 14228 26868
rect 13219 26812 14228 26840
rect 14369 26843 14427 26849
rect 13219 26809 13231 26812
rect 13173 26803 13231 26809
rect 14369 26809 14381 26843
rect 14415 26840 14427 26843
rect 15010 26840 15016 26852
rect 14415 26812 15016 26840
rect 14415 26809 14427 26812
rect 14369 26803 14427 26809
rect 15010 26800 15016 26812
rect 15068 26800 15074 26852
rect 16040 26784 16068 26880
rect 17034 26868 17040 26880
rect 17092 26868 17098 26920
rect 17402 26868 17408 26920
rect 17460 26908 17466 26920
rect 17589 26911 17647 26917
rect 17589 26908 17601 26911
rect 17460 26880 17601 26908
rect 17460 26868 17466 26880
rect 17589 26877 17601 26880
rect 17635 26908 17647 26911
rect 18417 26911 18475 26917
rect 18417 26908 18429 26911
rect 17635 26880 18429 26908
rect 17635 26877 17647 26880
rect 17589 26871 17647 26877
rect 18417 26877 18429 26880
rect 18463 26877 18475 26911
rect 18417 26871 18475 26877
rect 6549 26775 6607 26781
rect 6549 26741 6561 26775
rect 6595 26741 6607 26775
rect 10870 26772 10876 26784
rect 10831 26744 10876 26772
rect 6549 26735 6607 26741
rect 10870 26732 10876 26744
rect 10928 26732 10934 26784
rect 11609 26775 11667 26781
rect 11609 26741 11621 26775
rect 11655 26772 11667 26775
rect 11790 26772 11796 26784
rect 11655 26744 11796 26772
rect 11655 26741 11667 26744
rect 11609 26735 11667 26741
rect 11790 26732 11796 26744
rect 11848 26772 11854 26784
rect 13262 26772 13268 26784
rect 11848 26744 13268 26772
rect 11848 26732 11854 26744
rect 13262 26732 13268 26744
rect 13320 26732 13326 26784
rect 13814 26732 13820 26784
rect 13872 26772 13878 26784
rect 14645 26775 14703 26781
rect 14645 26772 14657 26775
rect 13872 26744 14657 26772
rect 13872 26732 13878 26744
rect 14645 26741 14657 26744
rect 14691 26741 14703 26775
rect 14645 26735 14703 26741
rect 16022 26732 16028 26784
rect 16080 26772 16086 26784
rect 16117 26775 16175 26781
rect 16117 26772 16129 26775
rect 16080 26744 16129 26772
rect 16080 26732 16086 26744
rect 16117 26741 16129 26744
rect 16163 26741 16175 26775
rect 16117 26735 16175 26741
rect 16577 26775 16635 26781
rect 16577 26741 16589 26775
rect 16623 26772 16635 26775
rect 17310 26772 17316 26784
rect 16623 26744 17316 26772
rect 16623 26741 16635 26744
rect 16577 26735 16635 26741
rect 17310 26732 17316 26744
rect 17368 26732 17374 26784
rect 1104 26682 18860 26704
rect 1104 26630 7648 26682
rect 7700 26630 7712 26682
rect 7764 26630 7776 26682
rect 7828 26630 7840 26682
rect 7892 26630 14315 26682
rect 14367 26630 14379 26682
rect 14431 26630 14443 26682
rect 14495 26630 14507 26682
rect 14559 26630 18860 26682
rect 1104 26608 18860 26630
rect 4614 26568 4620 26580
rect 4448 26540 4620 26568
rect 3602 26500 3608 26512
rect 3436 26472 3608 26500
rect 1578 26432 1584 26444
rect 1539 26404 1584 26432
rect 1578 26392 1584 26404
rect 1636 26392 1642 26444
rect 1670 26392 1676 26444
rect 1728 26432 1734 26444
rect 1857 26435 1915 26441
rect 1857 26432 1869 26435
rect 1728 26404 1869 26432
rect 1728 26392 1734 26404
rect 1857 26401 1869 26404
rect 1903 26432 1915 26435
rect 2314 26432 2320 26444
rect 1903 26404 2320 26432
rect 1903 26401 1915 26404
rect 1857 26395 1915 26401
rect 2314 26392 2320 26404
rect 2372 26392 2378 26444
rect 3436 26432 3464 26472
rect 3602 26460 3608 26472
rect 3660 26460 3666 26512
rect 2424 26404 3464 26432
rect 1596 26364 1624 26392
rect 2038 26364 2044 26376
rect 1596 26336 2044 26364
rect 2038 26324 2044 26336
rect 2096 26364 2102 26376
rect 2424 26364 2452 26404
rect 3510 26392 3516 26444
rect 3568 26432 3574 26444
rect 4448 26441 4476 26540
rect 4614 26528 4620 26540
rect 4672 26568 4678 26580
rect 5626 26568 5632 26580
rect 4672 26540 5632 26568
rect 4672 26528 4678 26540
rect 5626 26528 5632 26540
rect 5684 26528 5690 26580
rect 5721 26571 5779 26577
rect 5721 26537 5733 26571
rect 5767 26568 5779 26571
rect 6454 26568 6460 26580
rect 5767 26540 6460 26568
rect 5767 26537 5779 26540
rect 5721 26531 5779 26537
rect 6454 26528 6460 26540
rect 6512 26528 6518 26580
rect 6641 26571 6699 26577
rect 6641 26537 6653 26571
rect 6687 26568 6699 26571
rect 7466 26568 7472 26580
rect 6687 26540 7472 26568
rect 6687 26537 6699 26540
rect 6641 26531 6699 26537
rect 7466 26528 7472 26540
rect 7524 26528 7530 26580
rect 8478 26568 8484 26580
rect 8439 26540 8484 26568
rect 8478 26528 8484 26540
rect 8536 26528 8542 26580
rect 8662 26568 8668 26580
rect 8623 26540 8668 26568
rect 8662 26528 8668 26540
rect 8720 26528 8726 26580
rect 11514 26568 11520 26580
rect 11475 26540 11520 26568
rect 11514 26528 11520 26540
rect 11572 26528 11578 26580
rect 16025 26571 16083 26577
rect 16025 26537 16037 26571
rect 16071 26568 16083 26571
rect 16206 26568 16212 26580
rect 16071 26540 16212 26568
rect 16071 26537 16083 26540
rect 16025 26531 16083 26537
rect 16206 26528 16212 26540
rect 16264 26568 16270 26580
rect 16264 26540 16712 26568
rect 16264 26528 16270 26540
rect 5166 26500 5172 26512
rect 5127 26472 5172 26500
rect 5166 26460 5172 26472
rect 5224 26460 5230 26512
rect 7650 26460 7656 26512
rect 7708 26500 7714 26512
rect 7745 26503 7803 26509
rect 7745 26500 7757 26503
rect 7708 26472 7757 26500
rect 7708 26460 7714 26472
rect 7745 26469 7757 26472
rect 7791 26500 7803 26503
rect 8386 26500 8392 26512
rect 7791 26472 8392 26500
rect 7791 26469 7803 26472
rect 7745 26463 7803 26469
rect 8386 26460 8392 26472
rect 8444 26460 8450 26512
rect 16117 26503 16175 26509
rect 16117 26469 16129 26503
rect 16163 26500 16175 26503
rect 16574 26500 16580 26512
rect 16163 26472 16580 26500
rect 16163 26469 16175 26472
rect 16117 26463 16175 26469
rect 16574 26460 16580 26472
rect 16632 26460 16638 26512
rect 4065 26435 4123 26441
rect 4065 26432 4077 26435
rect 3568 26404 4077 26432
rect 3568 26392 3574 26404
rect 4065 26401 4077 26404
rect 4111 26401 4123 26435
rect 4065 26395 4123 26401
rect 4433 26435 4491 26441
rect 4433 26401 4445 26435
rect 4479 26401 4491 26435
rect 4893 26435 4951 26441
rect 4893 26432 4905 26435
rect 4433 26395 4491 26401
rect 4540 26404 4905 26432
rect 3234 26364 3240 26376
rect 2096 26336 2452 26364
rect 3195 26336 3240 26364
rect 2096 26324 2102 26336
rect 3234 26324 3240 26336
rect 3292 26324 3298 26376
rect 3973 26299 4031 26305
rect 3973 26265 3985 26299
rect 4019 26296 4031 26299
rect 4540 26296 4568 26404
rect 4893 26401 4905 26404
rect 4939 26401 4951 26435
rect 4893 26395 4951 26401
rect 7098 26392 7104 26444
rect 7156 26432 7162 26444
rect 7561 26435 7619 26441
rect 7561 26432 7573 26435
rect 7156 26404 7573 26432
rect 7156 26392 7162 26404
rect 7561 26401 7573 26404
rect 7607 26432 7619 26435
rect 8110 26432 8116 26444
rect 7607 26404 8116 26432
rect 7607 26401 7619 26404
rect 7561 26395 7619 26401
rect 8110 26392 8116 26404
rect 8168 26392 8174 26444
rect 8754 26432 8760 26444
rect 8715 26404 8760 26432
rect 8754 26392 8760 26404
rect 8812 26392 8818 26444
rect 9306 26432 9312 26444
rect 9267 26404 9312 26432
rect 9306 26392 9312 26404
rect 9364 26392 9370 26444
rect 11333 26435 11391 26441
rect 11333 26401 11345 26435
rect 11379 26432 11391 26435
rect 11422 26432 11428 26444
rect 11379 26404 11428 26432
rect 11379 26401 11391 26404
rect 11333 26395 11391 26401
rect 11422 26392 11428 26404
rect 11480 26392 11486 26444
rect 13354 26432 13360 26444
rect 13315 26404 13360 26432
rect 13354 26392 13360 26404
rect 13412 26392 13418 26444
rect 13541 26435 13599 26441
rect 13541 26401 13553 26435
rect 13587 26401 13599 26435
rect 14090 26432 14096 26444
rect 14051 26404 14096 26432
rect 13541 26395 13599 26401
rect 8662 26324 8668 26376
rect 8720 26364 8726 26376
rect 9401 26367 9459 26373
rect 9401 26364 9413 26367
rect 8720 26336 9413 26364
rect 8720 26324 8726 26336
rect 9401 26333 9413 26336
rect 9447 26333 9459 26367
rect 12161 26367 12219 26373
rect 12161 26364 12173 26367
rect 9401 26327 9459 26333
rect 11164 26336 12173 26364
rect 11164 26308 11192 26336
rect 12161 26333 12173 26336
rect 12207 26333 12219 26367
rect 12161 26327 12219 26333
rect 12710 26324 12716 26376
rect 12768 26364 12774 26376
rect 12986 26364 12992 26376
rect 12768 26336 12992 26364
rect 12768 26324 12774 26336
rect 12986 26324 12992 26336
rect 13044 26364 13050 26376
rect 13556 26364 13584 26395
rect 14090 26392 14096 26404
rect 14148 26392 14154 26444
rect 16684 26441 16712 26540
rect 16850 26528 16856 26580
rect 16908 26568 16914 26580
rect 17405 26571 17463 26577
rect 17405 26568 17417 26571
rect 16908 26540 17417 26568
rect 16908 26528 16914 26540
rect 17405 26537 17417 26540
rect 17451 26537 17463 26571
rect 17405 26531 17463 26537
rect 16669 26435 16727 26441
rect 16669 26401 16681 26435
rect 16715 26401 16727 26435
rect 16669 26395 16727 26401
rect 16945 26435 17003 26441
rect 16945 26401 16957 26435
rect 16991 26401 17003 26435
rect 16945 26395 17003 26401
rect 13044 26336 13584 26364
rect 13044 26324 13050 26336
rect 14182 26324 14188 26376
rect 14240 26364 14246 26376
rect 14369 26367 14427 26373
rect 14369 26364 14381 26367
rect 14240 26336 14381 26364
rect 14240 26324 14246 26336
rect 14369 26333 14381 26336
rect 14415 26364 14427 26367
rect 15102 26364 15108 26376
rect 14415 26336 15108 26364
rect 14415 26333 14427 26336
rect 14369 26327 14427 26333
rect 15102 26324 15108 26336
rect 15160 26324 15166 26376
rect 16960 26364 16988 26395
rect 16592 26336 16988 26364
rect 17129 26367 17187 26373
rect 4019 26268 4568 26296
rect 8113 26299 8171 26305
rect 4019 26265 4031 26268
rect 3973 26259 4031 26265
rect 4172 26240 4200 26268
rect 8113 26265 8125 26299
rect 8159 26296 8171 26299
rect 11146 26296 11152 26308
rect 8159 26268 8248 26296
rect 11107 26268 11152 26296
rect 8159 26265 8171 26268
rect 8113 26259 8171 26265
rect 4154 26188 4160 26240
rect 4212 26188 4218 26240
rect 8220 26228 8248 26268
rect 11146 26256 11152 26268
rect 11204 26256 11210 26308
rect 11882 26296 11888 26308
rect 11843 26268 11888 26296
rect 11882 26256 11888 26268
rect 11940 26256 11946 26308
rect 12805 26299 12863 26305
rect 12805 26265 12817 26299
rect 12851 26296 12863 26299
rect 13722 26296 13728 26308
rect 12851 26268 13728 26296
rect 12851 26265 12863 26268
rect 12805 26259 12863 26265
rect 13722 26256 13728 26268
rect 13780 26256 13786 26308
rect 8570 26228 8576 26240
rect 8220 26200 8576 26228
rect 8570 26188 8576 26200
rect 8628 26188 8634 26240
rect 10045 26231 10103 26237
rect 10045 26197 10057 26231
rect 10091 26228 10103 26231
rect 10134 26228 10140 26240
rect 10091 26200 10140 26228
rect 10091 26197 10103 26200
rect 10045 26191 10103 26197
rect 10134 26188 10140 26200
rect 10192 26228 10198 26240
rect 10686 26228 10692 26240
rect 10192 26200 10692 26228
rect 10192 26188 10198 26200
rect 10686 26188 10692 26200
rect 10744 26188 10750 26240
rect 15746 26188 15752 26240
rect 15804 26228 15810 26240
rect 16592 26228 16620 26336
rect 17129 26333 17141 26367
rect 17175 26364 17187 26367
rect 17310 26364 17316 26376
rect 17175 26336 17316 26364
rect 17175 26333 17187 26336
rect 17129 26327 17187 26333
rect 17310 26324 17316 26336
rect 17368 26324 17374 26376
rect 15804 26200 16620 26228
rect 15804 26188 15810 26200
rect 1104 26138 18860 26160
rect 1104 26086 4315 26138
rect 4367 26086 4379 26138
rect 4431 26086 4443 26138
rect 4495 26086 4507 26138
rect 4559 26086 10982 26138
rect 11034 26086 11046 26138
rect 11098 26086 11110 26138
rect 11162 26086 11174 26138
rect 11226 26086 17648 26138
rect 17700 26086 17712 26138
rect 17764 26086 17776 26138
rect 17828 26086 17840 26138
rect 17892 26086 18860 26138
rect 1104 26064 18860 26086
rect 1670 26024 1676 26036
rect 1631 25996 1676 26024
rect 1670 25984 1676 25996
rect 1728 25984 1734 26036
rect 2038 26024 2044 26036
rect 1999 25996 2044 26024
rect 2038 25984 2044 25996
rect 2096 25984 2102 26036
rect 2501 26027 2559 26033
rect 2501 25993 2513 26027
rect 2547 26024 2559 26027
rect 2866 26024 2872 26036
rect 2547 25996 2872 26024
rect 2547 25993 2559 25996
rect 2501 25987 2559 25993
rect 2866 25984 2872 25996
rect 2924 25984 2930 26036
rect 3326 25984 3332 26036
rect 3384 26024 3390 26036
rect 3421 26027 3479 26033
rect 3421 26024 3433 26027
rect 3384 25996 3433 26024
rect 3384 25984 3390 25996
rect 3421 25993 3433 25996
rect 3467 25993 3479 26027
rect 3421 25987 3479 25993
rect 3436 25888 3464 25987
rect 3510 25984 3516 26036
rect 3568 26024 3574 26036
rect 3789 26027 3847 26033
rect 3789 26024 3801 26027
rect 3568 25996 3801 26024
rect 3568 25984 3574 25996
rect 3789 25993 3801 25996
rect 3835 25993 3847 26027
rect 4154 26024 4160 26036
rect 4115 25996 4160 26024
rect 3789 25987 3847 25993
rect 4154 25984 4160 25996
rect 4212 25984 4218 26036
rect 7098 26024 7104 26036
rect 7059 25996 7104 26024
rect 7098 25984 7104 25996
rect 7156 25984 7162 26036
rect 7650 26024 7656 26036
rect 7611 25996 7656 26024
rect 7650 25984 7656 25996
rect 7708 25984 7714 26036
rect 9125 26027 9183 26033
rect 9125 25993 9137 26027
rect 9171 26024 9183 26027
rect 9306 26024 9312 26036
rect 9171 25996 9312 26024
rect 9171 25993 9183 25996
rect 9125 25987 9183 25993
rect 9306 25984 9312 25996
rect 9364 25984 9370 26036
rect 12802 26024 12808 26036
rect 12763 25996 12808 26024
rect 12802 25984 12808 25996
rect 12860 25984 12866 26036
rect 15470 25984 15476 26036
rect 15528 26024 15534 26036
rect 15565 26027 15623 26033
rect 15565 26024 15577 26027
rect 15528 25996 15577 26024
rect 15528 25984 15534 25996
rect 15565 25993 15577 25996
rect 15611 26024 15623 26027
rect 15746 26024 15752 26036
rect 15611 25996 15752 26024
rect 15611 25993 15623 25996
rect 15565 25987 15623 25993
rect 15746 25984 15752 25996
rect 15804 25984 15810 26036
rect 15841 26027 15899 26033
rect 15841 25993 15853 26027
rect 15887 26024 15899 26027
rect 16022 26024 16028 26036
rect 15887 25996 16028 26024
rect 15887 25993 15899 25996
rect 15841 25987 15899 25993
rect 16022 25984 16028 25996
rect 16080 25984 16086 26036
rect 16850 25984 16856 26036
rect 16908 26024 16914 26036
rect 18049 26027 18107 26033
rect 18049 26024 18061 26027
rect 16908 25996 18061 26024
rect 16908 25984 16914 25996
rect 18049 25993 18061 25996
rect 18095 25993 18107 26027
rect 18049 25987 18107 25993
rect 4706 25916 4712 25968
rect 4764 25956 4770 25968
rect 5721 25959 5779 25965
rect 5721 25956 5733 25959
rect 4764 25928 5733 25956
rect 4764 25916 4770 25928
rect 5721 25925 5733 25928
rect 5767 25925 5779 25959
rect 5721 25919 5779 25925
rect 8021 25959 8079 25965
rect 8021 25925 8033 25959
rect 8067 25956 8079 25959
rect 8754 25956 8760 25968
rect 8067 25928 8760 25956
rect 8067 25925 8079 25928
rect 8021 25919 8079 25925
rect 8754 25916 8760 25928
rect 8812 25916 8818 25968
rect 17494 25956 17500 25968
rect 17455 25928 17500 25956
rect 17494 25916 17500 25928
rect 17552 25916 17558 25968
rect 6454 25888 6460 25900
rect 3436 25860 4660 25888
rect 6415 25860 6460 25888
rect 3694 25780 3700 25832
rect 3752 25820 3758 25832
rect 4632 25829 4660 25860
rect 6454 25848 6460 25860
rect 6512 25848 6518 25900
rect 9858 25888 9864 25900
rect 9819 25860 9864 25888
rect 9858 25848 9864 25860
rect 9916 25848 9922 25900
rect 12437 25891 12495 25897
rect 12437 25857 12449 25891
rect 12483 25888 12495 25891
rect 16850 25888 16856 25900
rect 12483 25860 13400 25888
rect 16811 25860 16856 25888
rect 12483 25857 12495 25860
rect 12437 25851 12495 25857
rect 13372 25832 13400 25860
rect 16850 25848 16856 25860
rect 16908 25848 16914 25900
rect 18417 25891 18475 25897
rect 18417 25888 18429 25891
rect 17052 25860 18429 25888
rect 17052 25832 17080 25860
rect 18417 25857 18429 25860
rect 18463 25857 18475 25891
rect 18417 25851 18475 25857
rect 4065 25823 4123 25829
rect 4065 25820 4077 25823
rect 3752 25792 4077 25820
rect 3752 25780 3758 25792
rect 4065 25789 4077 25792
rect 4111 25789 4123 25823
rect 4065 25783 4123 25789
rect 4617 25823 4675 25829
rect 4617 25789 4629 25823
rect 4663 25789 4675 25823
rect 4617 25783 4675 25789
rect 5169 25823 5227 25829
rect 5169 25789 5181 25823
rect 5215 25820 5227 25823
rect 5813 25823 5871 25829
rect 5813 25820 5825 25823
rect 5215 25792 5825 25820
rect 5215 25789 5227 25792
rect 5169 25783 5227 25789
rect 5813 25789 5825 25792
rect 5859 25820 5871 25823
rect 5902 25820 5908 25832
rect 5859 25792 5908 25820
rect 5859 25789 5871 25792
rect 5813 25783 5871 25789
rect 5902 25780 5908 25792
rect 5960 25780 5966 25832
rect 6362 25820 6368 25832
rect 6323 25792 6368 25820
rect 6362 25780 6368 25792
rect 6420 25780 6426 25832
rect 7650 25780 7656 25832
rect 7708 25820 7714 25832
rect 8205 25823 8263 25829
rect 8205 25820 8217 25823
rect 7708 25792 8217 25820
rect 7708 25780 7714 25792
rect 8205 25789 8217 25792
rect 8251 25789 8263 25823
rect 8205 25783 8263 25789
rect 8389 25823 8447 25829
rect 8389 25789 8401 25823
rect 8435 25820 8447 25823
rect 8478 25820 8484 25832
rect 8435 25792 8484 25820
rect 8435 25789 8447 25792
rect 8389 25783 8447 25789
rect 8478 25780 8484 25792
rect 8536 25780 8542 25832
rect 8570 25780 8576 25832
rect 8628 25820 8634 25832
rect 9493 25823 9551 25829
rect 8628 25792 8673 25820
rect 8628 25780 8634 25792
rect 9493 25789 9505 25823
rect 9539 25820 9551 25823
rect 9766 25820 9772 25832
rect 9539 25792 9772 25820
rect 9539 25789 9551 25792
rect 9493 25783 9551 25789
rect 9766 25780 9772 25792
rect 9824 25780 9830 25832
rect 10134 25820 10140 25832
rect 10095 25792 10140 25820
rect 10134 25780 10140 25792
rect 10192 25780 10198 25832
rect 10410 25780 10416 25832
rect 10468 25820 10474 25832
rect 10505 25823 10563 25829
rect 10505 25820 10517 25823
rect 10468 25792 10517 25820
rect 10468 25780 10474 25792
rect 10505 25789 10517 25792
rect 10551 25789 10563 25823
rect 10505 25783 10563 25789
rect 12066 25780 12072 25832
rect 12124 25820 12130 25832
rect 12986 25820 12992 25832
rect 12124 25792 12992 25820
rect 12124 25780 12130 25792
rect 12986 25780 12992 25792
rect 13044 25780 13050 25832
rect 13354 25820 13360 25832
rect 13315 25792 13360 25820
rect 13354 25780 13360 25792
rect 13412 25780 13418 25832
rect 13449 25823 13507 25829
rect 13449 25789 13461 25823
rect 13495 25789 13507 25823
rect 13449 25783 13507 25789
rect 5537 25755 5595 25761
rect 5537 25721 5549 25755
rect 5583 25752 5595 25755
rect 6380 25752 6408 25780
rect 5583 25724 6408 25752
rect 5583 25721 5595 25724
rect 5537 25715 5595 25721
rect 10870 25712 10876 25764
rect 10928 25752 10934 25764
rect 11885 25755 11943 25761
rect 11885 25752 11897 25755
rect 10928 25724 11897 25752
rect 10928 25712 10934 25724
rect 11885 25721 11897 25724
rect 11931 25752 11943 25755
rect 12526 25752 12532 25764
rect 11931 25724 12532 25752
rect 11931 25721 11943 25724
rect 11885 25715 11943 25721
rect 12526 25712 12532 25724
rect 12584 25752 12590 25764
rect 13464 25752 13492 25783
rect 13814 25780 13820 25832
rect 13872 25820 13878 25832
rect 14001 25823 14059 25829
rect 14001 25820 14013 25823
rect 13872 25792 14013 25820
rect 13872 25780 13878 25792
rect 14001 25789 14013 25792
rect 14047 25789 14059 25823
rect 15654 25820 15660 25832
rect 15567 25792 15660 25820
rect 14001 25783 14059 25789
rect 15654 25780 15660 25792
rect 15712 25820 15718 25832
rect 16117 25823 16175 25829
rect 16117 25820 16129 25823
rect 15712 25792 16129 25820
rect 15712 25780 15718 25792
rect 16117 25789 16129 25792
rect 16163 25789 16175 25823
rect 17034 25820 17040 25832
rect 16995 25792 17040 25820
rect 16117 25783 16175 25789
rect 17034 25780 17040 25792
rect 17092 25780 17098 25832
rect 17402 25780 17408 25832
rect 17460 25820 17466 25832
rect 17497 25823 17555 25829
rect 17497 25820 17509 25823
rect 17460 25792 17509 25820
rect 17460 25780 17466 25792
rect 17497 25789 17509 25792
rect 17543 25789 17555 25823
rect 17497 25783 17555 25789
rect 14090 25752 14096 25764
rect 12584 25724 14096 25752
rect 12584 25712 12590 25724
rect 14090 25712 14096 25724
rect 14148 25752 14154 25764
rect 14461 25755 14519 25761
rect 14461 25752 14473 25755
rect 14148 25724 14473 25752
rect 14148 25712 14154 25724
rect 14461 25721 14473 25724
rect 14507 25721 14519 25755
rect 14461 25715 14519 25721
rect 11422 25684 11428 25696
rect 11383 25656 11428 25684
rect 11422 25644 11428 25656
rect 11480 25644 11486 25696
rect 12158 25684 12164 25696
rect 12119 25656 12164 25684
rect 12158 25644 12164 25656
rect 12216 25684 12222 25696
rect 12437 25687 12495 25693
rect 12437 25684 12449 25687
rect 12216 25656 12449 25684
rect 12216 25644 12222 25656
rect 12437 25653 12449 25656
rect 12483 25653 12495 25687
rect 12437 25647 12495 25653
rect 12621 25687 12679 25693
rect 12621 25653 12633 25687
rect 12667 25684 12679 25687
rect 12710 25684 12716 25696
rect 12667 25656 12716 25684
rect 12667 25653 12679 25656
rect 12621 25647 12679 25653
rect 12710 25644 12716 25656
rect 12768 25644 12774 25696
rect 16577 25687 16635 25693
rect 16577 25653 16589 25687
rect 16623 25684 16635 25687
rect 17310 25684 17316 25696
rect 16623 25656 17316 25684
rect 16623 25653 16635 25656
rect 16577 25647 16635 25653
rect 17310 25644 17316 25656
rect 17368 25644 17374 25696
rect 1104 25594 18860 25616
rect 1104 25542 7648 25594
rect 7700 25542 7712 25594
rect 7764 25542 7776 25594
rect 7828 25542 7840 25594
rect 7892 25542 14315 25594
rect 14367 25542 14379 25594
rect 14431 25542 14443 25594
rect 14495 25542 14507 25594
rect 14559 25542 18860 25594
rect 1104 25520 18860 25542
rect 5905 25483 5963 25489
rect 5905 25449 5917 25483
rect 5951 25480 5963 25483
rect 6546 25480 6552 25492
rect 5951 25452 6552 25480
rect 5951 25449 5963 25452
rect 5905 25443 5963 25449
rect 6546 25440 6552 25452
rect 6604 25440 6610 25492
rect 8662 25480 8668 25492
rect 8623 25452 8668 25480
rect 8662 25440 8668 25452
rect 8720 25440 8726 25492
rect 8754 25440 8760 25492
rect 8812 25480 8818 25492
rect 8941 25483 8999 25489
rect 8941 25480 8953 25483
rect 8812 25452 8953 25480
rect 8812 25440 8818 25452
rect 8941 25449 8953 25452
rect 8987 25449 8999 25483
rect 9490 25480 9496 25492
rect 9451 25452 9496 25480
rect 8941 25443 8999 25449
rect 9490 25440 9496 25452
rect 9548 25440 9554 25492
rect 9861 25483 9919 25489
rect 9861 25449 9873 25483
rect 9907 25480 9919 25483
rect 10410 25480 10416 25492
rect 9907 25452 10416 25480
rect 9907 25449 9919 25452
rect 9861 25443 9919 25449
rect 10410 25440 10416 25452
rect 10468 25440 10474 25492
rect 12066 25440 12072 25492
rect 12124 25480 12130 25492
rect 12161 25483 12219 25489
rect 12161 25480 12173 25483
rect 12124 25452 12173 25480
rect 12124 25440 12130 25452
rect 12161 25449 12173 25452
rect 12207 25449 12219 25483
rect 13630 25480 13636 25492
rect 13591 25452 13636 25480
rect 12161 25443 12219 25449
rect 13630 25440 13636 25452
rect 13688 25440 13694 25492
rect 15286 25440 15292 25492
rect 15344 25480 15350 25492
rect 15381 25483 15439 25489
rect 15381 25480 15393 25483
rect 15344 25452 15393 25480
rect 15344 25440 15350 25452
rect 15381 25449 15393 25452
rect 15427 25449 15439 25483
rect 15381 25443 15439 25449
rect 6641 25415 6699 25421
rect 6641 25381 6653 25415
rect 6687 25412 6699 25415
rect 7098 25412 7104 25424
rect 6687 25384 7104 25412
rect 6687 25381 6699 25384
rect 6641 25375 6699 25381
rect 7098 25372 7104 25384
rect 7156 25412 7162 25424
rect 7156 25384 7972 25412
rect 7156 25372 7162 25384
rect 3878 25304 3884 25356
rect 3936 25344 3942 25356
rect 4065 25347 4123 25353
rect 4065 25344 4077 25347
rect 3936 25316 4077 25344
rect 3936 25304 3942 25316
rect 4065 25313 4077 25316
rect 4111 25344 4123 25347
rect 4614 25344 4620 25356
rect 4111 25316 4620 25344
rect 4111 25313 4123 25316
rect 4065 25307 4123 25313
rect 4614 25304 4620 25316
rect 4672 25304 4678 25356
rect 5721 25347 5779 25353
rect 5721 25313 5733 25347
rect 5767 25344 5779 25347
rect 5902 25344 5908 25356
rect 5767 25316 5908 25344
rect 5767 25313 5779 25316
rect 5721 25307 5779 25313
rect 5902 25304 5908 25316
rect 5960 25304 5966 25356
rect 7285 25347 7343 25353
rect 7285 25313 7297 25347
rect 7331 25344 7343 25347
rect 7374 25344 7380 25356
rect 7331 25316 7380 25344
rect 7331 25313 7343 25316
rect 7285 25307 7343 25313
rect 7374 25304 7380 25316
rect 7432 25304 7438 25356
rect 7466 25304 7472 25356
rect 7524 25344 7530 25356
rect 7944 25353 7972 25384
rect 10042 25372 10048 25424
rect 10100 25412 10106 25424
rect 10100 25384 10916 25412
rect 10100 25372 10106 25384
rect 7929 25347 7987 25353
rect 7524 25316 7569 25344
rect 7524 25304 7530 25316
rect 7929 25313 7941 25347
rect 7975 25313 7987 25347
rect 7929 25307 7987 25313
rect 9030 25304 9036 25356
rect 9088 25344 9094 25356
rect 9309 25347 9367 25353
rect 9309 25344 9321 25347
rect 9088 25316 9321 25344
rect 9088 25304 9094 25316
rect 9309 25313 9321 25316
rect 9355 25313 9367 25347
rect 9309 25307 9367 25313
rect 9398 25304 9404 25356
rect 9456 25344 9462 25356
rect 10888 25353 10916 25384
rect 12618 25372 12624 25424
rect 12676 25412 12682 25424
rect 12676 25384 12940 25412
rect 12676 25372 12682 25384
rect 12912 25356 12940 25384
rect 10137 25347 10195 25353
rect 10137 25344 10149 25347
rect 9456 25316 10149 25344
rect 9456 25304 9462 25316
rect 10137 25313 10149 25316
rect 10183 25344 10195 25347
rect 10321 25347 10379 25353
rect 10321 25344 10333 25347
rect 10183 25316 10333 25344
rect 10183 25313 10195 25316
rect 10137 25307 10195 25313
rect 10321 25313 10333 25316
rect 10367 25313 10379 25347
rect 10321 25307 10379 25313
rect 10873 25347 10931 25353
rect 10873 25313 10885 25347
rect 10919 25313 10931 25347
rect 12710 25344 12716 25356
rect 12671 25316 12716 25344
rect 10873 25307 10931 25313
rect 12710 25304 12716 25316
rect 12768 25304 12774 25356
rect 12894 25344 12900 25356
rect 12855 25316 12900 25344
rect 12894 25304 12900 25316
rect 12952 25304 12958 25356
rect 13262 25344 13268 25356
rect 13223 25316 13268 25344
rect 13262 25304 13268 25316
rect 13320 25304 13326 25356
rect 15194 25344 15200 25356
rect 15155 25316 15200 25344
rect 15194 25304 15200 25316
rect 15252 25304 15258 25356
rect 15562 25344 15568 25356
rect 15523 25316 15568 25344
rect 15562 25304 15568 25316
rect 15620 25304 15626 25356
rect 15746 25304 15752 25356
rect 15804 25344 15810 25356
rect 15933 25347 15991 25353
rect 15933 25344 15945 25347
rect 15804 25316 15945 25344
rect 15804 25304 15810 25316
rect 15933 25313 15945 25316
rect 15979 25313 15991 25347
rect 15933 25307 15991 25313
rect 6273 25279 6331 25285
rect 6273 25245 6285 25279
rect 6319 25276 6331 25279
rect 6638 25276 6644 25288
rect 6319 25248 6644 25276
rect 6319 25245 6331 25248
rect 6273 25239 6331 25245
rect 6638 25236 6644 25248
rect 6696 25236 6702 25288
rect 9858 25236 9864 25288
rect 9916 25276 9922 25288
rect 11149 25279 11207 25285
rect 11149 25276 11161 25279
rect 9916 25248 11161 25276
rect 9916 25236 9922 25248
rect 11149 25245 11161 25248
rect 11195 25245 11207 25279
rect 11149 25239 11207 25245
rect 13354 25236 13360 25288
rect 13412 25276 13418 25288
rect 13817 25279 13875 25285
rect 13817 25276 13829 25279
rect 13412 25248 13829 25276
rect 13412 25236 13418 25248
rect 13817 25245 13829 25248
rect 13863 25245 13875 25279
rect 13817 25239 13875 25245
rect 16761 25279 16819 25285
rect 16761 25245 16773 25279
rect 16807 25276 16819 25279
rect 17034 25276 17040 25288
rect 16807 25248 17040 25276
rect 16807 25245 16819 25248
rect 16761 25239 16819 25245
rect 17034 25236 17040 25248
rect 17092 25236 17098 25288
rect 3329 25211 3387 25217
rect 3329 25177 3341 25211
rect 3375 25208 3387 25211
rect 3786 25208 3792 25220
rect 3375 25180 3792 25208
rect 3375 25177 3387 25180
rect 3329 25171 3387 25177
rect 3786 25168 3792 25180
rect 3844 25168 3850 25220
rect 6362 25168 6368 25220
rect 6420 25208 6426 25220
rect 7929 25211 7987 25217
rect 7929 25208 7941 25211
rect 6420 25180 7941 25208
rect 6420 25168 6426 25180
rect 7929 25177 7941 25180
rect 7975 25177 7987 25211
rect 10410 25208 10416 25220
rect 10371 25180 10416 25208
rect 7929 25171 7987 25177
rect 10410 25168 10416 25180
rect 10468 25168 10474 25220
rect 1394 25100 1400 25152
rect 1452 25140 1458 25152
rect 1581 25143 1639 25149
rect 1581 25140 1593 25143
rect 1452 25112 1593 25140
rect 1452 25100 1458 25112
rect 1581 25109 1593 25112
rect 1627 25109 1639 25143
rect 3694 25140 3700 25152
rect 3655 25112 3700 25140
rect 1581 25103 1639 25109
rect 3694 25100 3700 25112
rect 3752 25100 3758 25152
rect 4614 25140 4620 25152
rect 4575 25112 4620 25140
rect 4614 25100 4620 25112
rect 4672 25100 4678 25152
rect 13538 25100 13544 25152
rect 13596 25140 13602 25152
rect 13633 25143 13691 25149
rect 13633 25140 13645 25143
rect 13596 25112 13645 25140
rect 13596 25100 13602 25112
rect 13633 25109 13645 25112
rect 13679 25109 13691 25143
rect 13633 25103 13691 25109
rect 16758 25100 16764 25152
rect 16816 25140 16822 25152
rect 17037 25143 17095 25149
rect 17037 25140 17049 25143
rect 16816 25112 17049 25140
rect 16816 25100 16822 25112
rect 17037 25109 17049 25112
rect 17083 25140 17095 25143
rect 17402 25140 17408 25152
rect 17083 25112 17408 25140
rect 17083 25109 17095 25112
rect 17037 25103 17095 25109
rect 17402 25100 17408 25112
rect 17460 25100 17466 25152
rect 1104 25050 18860 25072
rect 1104 24998 4315 25050
rect 4367 24998 4379 25050
rect 4431 24998 4443 25050
rect 4495 24998 4507 25050
rect 4559 24998 10982 25050
rect 11034 24998 11046 25050
rect 11098 24998 11110 25050
rect 11162 24998 11174 25050
rect 11226 24998 17648 25050
rect 17700 24998 17712 25050
rect 17764 24998 17776 25050
rect 17828 24998 17840 25050
rect 17892 24998 18860 25050
rect 1104 24976 18860 24998
rect 3694 24896 3700 24948
rect 3752 24936 3758 24948
rect 5445 24939 5503 24945
rect 5445 24936 5457 24939
rect 3752 24908 5457 24936
rect 3752 24896 3758 24908
rect 5445 24905 5457 24908
rect 5491 24905 5503 24939
rect 9030 24936 9036 24948
rect 8991 24908 9036 24936
rect 5445 24899 5503 24905
rect 9030 24896 9036 24908
rect 9088 24896 9094 24948
rect 15102 24936 15108 24948
rect 15015 24908 15108 24936
rect 15102 24896 15108 24908
rect 15160 24936 15166 24948
rect 15562 24936 15568 24948
rect 15160 24908 15568 24936
rect 15160 24896 15166 24908
rect 15562 24896 15568 24908
rect 15620 24896 15626 24948
rect 3878 24868 3884 24880
rect 3839 24840 3884 24868
rect 3878 24828 3884 24840
rect 3936 24828 3942 24880
rect 7374 24868 7380 24880
rect 6840 24840 7380 24868
rect 1673 24803 1731 24809
rect 1673 24769 1685 24803
rect 1719 24800 1731 24803
rect 1854 24800 1860 24812
rect 1719 24772 1860 24800
rect 1719 24769 1731 24772
rect 1673 24763 1731 24769
rect 1854 24760 1860 24772
rect 1912 24760 1918 24812
rect 3513 24803 3571 24809
rect 3513 24769 3525 24803
rect 3559 24800 3571 24803
rect 6457 24803 6515 24809
rect 3559 24772 4384 24800
rect 3559 24769 3571 24772
rect 3513 24763 3571 24769
rect 1394 24732 1400 24744
rect 1355 24704 1400 24732
rect 1394 24692 1400 24704
rect 1452 24692 1458 24744
rect 3878 24692 3884 24744
rect 3936 24732 3942 24744
rect 4356 24741 4384 24772
rect 6457 24769 6469 24803
rect 6503 24800 6515 24803
rect 6840 24800 6868 24840
rect 7374 24828 7380 24840
rect 7432 24828 7438 24880
rect 8294 24868 8300 24880
rect 8220 24840 8300 24868
rect 8018 24800 8024 24812
rect 6503 24772 6868 24800
rect 7979 24772 8024 24800
rect 6503 24769 6515 24772
rect 6457 24763 6515 24769
rect 8018 24760 8024 24772
rect 8076 24760 8082 24812
rect 4065 24735 4123 24741
rect 4065 24732 4077 24735
rect 3936 24704 4077 24732
rect 3936 24692 3942 24704
rect 4065 24701 4077 24704
rect 4111 24701 4123 24735
rect 4065 24695 4123 24701
rect 4341 24735 4399 24741
rect 4341 24701 4353 24735
rect 4387 24732 4399 24735
rect 4614 24732 4620 24744
rect 4387 24704 4620 24732
rect 4387 24701 4399 24704
rect 4341 24695 4399 24701
rect 4614 24692 4620 24704
rect 4672 24692 4678 24744
rect 6638 24692 6644 24744
rect 6696 24732 6702 24744
rect 6733 24735 6791 24741
rect 6733 24732 6745 24735
rect 6696 24704 6745 24732
rect 6696 24692 6702 24704
rect 6733 24701 6745 24704
rect 6779 24701 6791 24735
rect 6733 24695 6791 24701
rect 7190 24692 7196 24744
rect 7248 24732 7254 24744
rect 7374 24732 7380 24744
rect 7248 24704 7380 24732
rect 7248 24692 7254 24704
rect 7374 24692 7380 24704
rect 7432 24732 7438 24744
rect 7469 24735 7527 24741
rect 7469 24732 7481 24735
rect 7432 24704 7481 24732
rect 7432 24692 7438 24704
rect 7469 24701 7481 24704
rect 7515 24701 7527 24735
rect 7469 24695 7527 24701
rect 8113 24735 8171 24741
rect 8113 24701 8125 24735
rect 8159 24732 8171 24735
rect 8220 24732 8248 24840
rect 8294 24828 8300 24840
rect 8352 24828 8358 24880
rect 9858 24868 9864 24880
rect 9600 24840 9864 24868
rect 9493 24803 9551 24809
rect 9493 24769 9505 24803
rect 9539 24800 9551 24803
rect 9600 24800 9628 24840
rect 9858 24828 9864 24840
rect 9916 24828 9922 24880
rect 12986 24828 12992 24880
rect 13044 24868 13050 24880
rect 15194 24868 15200 24880
rect 13044 24840 13860 24868
rect 13044 24828 13050 24840
rect 9539 24772 9628 24800
rect 10137 24803 10195 24809
rect 9539 24769 9551 24772
rect 9493 24763 9551 24769
rect 10137 24769 10149 24803
rect 10183 24800 10195 24803
rect 13832 24800 13860 24840
rect 15120 24840 15200 24868
rect 13906 24800 13912 24812
rect 10183 24772 10548 24800
rect 13819 24772 13912 24800
rect 10183 24769 10195 24772
rect 10137 24763 10195 24769
rect 8159 24704 8248 24732
rect 8159 24701 8171 24704
rect 8113 24695 8171 24701
rect 3053 24667 3111 24673
rect 3053 24633 3065 24667
rect 3099 24664 3111 24667
rect 3510 24664 3516 24676
rect 3099 24636 3516 24664
rect 3099 24633 3111 24636
rect 3053 24627 3111 24633
rect 3510 24624 3516 24636
rect 3568 24624 3574 24676
rect 7006 24624 7012 24676
rect 7064 24664 7070 24676
rect 7285 24667 7343 24673
rect 7285 24664 7297 24667
rect 7064 24636 7297 24664
rect 7064 24624 7070 24636
rect 7285 24633 7297 24636
rect 7331 24664 7343 24667
rect 8128 24664 8156 24695
rect 8294 24692 8300 24744
rect 8352 24732 8358 24744
rect 8481 24735 8539 24741
rect 8481 24732 8493 24735
rect 8352 24704 8493 24732
rect 8352 24692 8358 24704
rect 8481 24701 8493 24704
rect 8527 24732 8539 24735
rect 8846 24732 8852 24744
rect 8527 24704 8852 24732
rect 8527 24701 8539 24704
rect 8481 24695 8539 24701
rect 8846 24692 8852 24704
rect 8904 24692 8910 24744
rect 10226 24732 10232 24744
rect 10187 24704 10232 24732
rect 10226 24692 10232 24704
rect 10284 24692 10290 24744
rect 10520 24741 10548 24772
rect 13906 24760 13912 24772
rect 13964 24800 13970 24812
rect 14737 24803 14795 24809
rect 14737 24800 14749 24803
rect 13964 24772 14749 24800
rect 13964 24760 13970 24772
rect 14737 24769 14749 24772
rect 14783 24800 14795 24803
rect 15120 24800 15148 24840
rect 15194 24828 15200 24840
rect 15252 24828 15258 24880
rect 17494 24868 17500 24880
rect 17455 24840 17500 24868
rect 17494 24828 17500 24840
rect 17552 24828 17558 24880
rect 15565 24803 15623 24809
rect 15565 24800 15577 24803
rect 14783 24772 15148 24800
rect 15212 24772 15577 24800
rect 14783 24769 14795 24772
rect 14737 24763 14795 24769
rect 10505 24735 10563 24741
rect 10505 24701 10517 24735
rect 10551 24732 10563 24735
rect 10778 24732 10784 24744
rect 10551 24704 10784 24732
rect 10551 24701 10563 24704
rect 10505 24695 10563 24701
rect 10778 24692 10784 24704
rect 10836 24692 10842 24744
rect 13817 24735 13875 24741
rect 13817 24701 13829 24735
rect 13863 24701 13875 24735
rect 14182 24732 14188 24744
rect 14095 24704 14188 24732
rect 13817 24695 13875 24701
rect 7331 24636 8156 24664
rect 7331 24633 7343 24636
rect 7285 24627 7343 24633
rect 12618 24624 12624 24676
rect 12676 24664 12682 24676
rect 13173 24667 13231 24673
rect 13173 24664 13185 24667
rect 12676 24636 13185 24664
rect 12676 24624 12682 24636
rect 13173 24633 13185 24636
rect 13219 24664 13231 24667
rect 13262 24664 13268 24676
rect 13219 24636 13268 24664
rect 13219 24633 13231 24636
rect 13173 24627 13231 24633
rect 13262 24624 13268 24636
rect 13320 24624 13326 24676
rect 13832 24664 13860 24695
rect 14182 24692 14188 24704
rect 14240 24732 14246 24744
rect 14826 24732 14832 24744
rect 14240 24704 14832 24732
rect 14240 24692 14246 24704
rect 14826 24692 14832 24704
rect 14884 24692 14890 24744
rect 13998 24664 14004 24676
rect 13832 24636 14004 24664
rect 13998 24624 14004 24636
rect 14056 24664 14062 24676
rect 15212 24664 15240 24772
rect 15565 24769 15577 24772
rect 15611 24800 15623 24803
rect 15746 24800 15752 24812
rect 15611 24772 15752 24800
rect 15611 24769 15623 24772
rect 15565 24763 15623 24769
rect 15746 24760 15752 24772
rect 15804 24760 15810 24812
rect 16574 24800 16580 24812
rect 16535 24772 16580 24800
rect 16574 24760 16580 24772
rect 16632 24800 16638 24812
rect 16761 24803 16819 24809
rect 16761 24800 16773 24803
rect 16632 24772 16773 24800
rect 16632 24760 16638 24772
rect 16761 24769 16773 24772
rect 16807 24769 16819 24803
rect 16761 24763 16819 24769
rect 15654 24732 15660 24744
rect 15615 24704 15660 24732
rect 15654 24692 15660 24704
rect 15712 24732 15718 24744
rect 16117 24735 16175 24741
rect 16117 24732 16129 24735
rect 15712 24704 16129 24732
rect 15712 24692 15718 24704
rect 16117 24701 16129 24704
rect 16163 24701 16175 24735
rect 17034 24732 17040 24744
rect 16995 24704 17040 24732
rect 16117 24695 16175 24701
rect 17034 24692 17040 24704
rect 17092 24692 17098 24744
rect 17402 24692 17408 24744
rect 17460 24732 17466 24744
rect 17497 24735 17555 24741
rect 17497 24732 17509 24735
rect 17460 24704 17509 24732
rect 17460 24692 17466 24704
rect 17497 24701 17509 24704
rect 17543 24701 17555 24735
rect 17497 24695 17555 24701
rect 16206 24664 16212 24676
rect 14056 24636 15240 24664
rect 15856 24636 16212 24664
rect 14056 24624 14062 24636
rect 5902 24556 5908 24608
rect 5960 24596 5966 24608
rect 5997 24599 6055 24605
rect 5997 24596 6009 24599
rect 5960 24568 6009 24596
rect 5960 24556 5966 24568
rect 5997 24565 6009 24568
rect 6043 24565 6055 24599
rect 5997 24559 6055 24565
rect 6362 24556 6368 24608
rect 6420 24596 6426 24608
rect 6549 24599 6607 24605
rect 6549 24596 6561 24599
rect 6420 24568 6561 24596
rect 6420 24556 6426 24568
rect 6549 24565 6561 24568
rect 6595 24565 6607 24599
rect 6549 24559 6607 24565
rect 11514 24556 11520 24608
rect 11572 24596 11578 24608
rect 11609 24599 11667 24605
rect 11609 24596 11621 24599
rect 11572 24568 11621 24596
rect 11572 24556 11578 24568
rect 11609 24565 11621 24568
rect 11655 24565 11667 24599
rect 11609 24559 11667 24565
rect 12529 24599 12587 24605
rect 12529 24565 12541 24599
rect 12575 24596 12587 24599
rect 12710 24596 12716 24608
rect 12575 24568 12716 24596
rect 12575 24565 12587 24568
rect 12529 24559 12587 24565
rect 12710 24556 12716 24568
rect 12768 24556 12774 24608
rect 12897 24599 12955 24605
rect 12897 24565 12909 24599
rect 12943 24596 12955 24599
rect 12986 24596 12992 24608
rect 12943 24568 12992 24596
rect 12943 24565 12955 24568
rect 12897 24559 12955 24565
rect 12986 24556 12992 24568
rect 13044 24556 13050 24608
rect 13814 24556 13820 24608
rect 13872 24596 13878 24608
rect 15856 24605 15884 24636
rect 16206 24624 16212 24636
rect 16264 24624 16270 24676
rect 13909 24599 13967 24605
rect 13909 24596 13921 24599
rect 13872 24568 13921 24596
rect 13872 24556 13878 24568
rect 13909 24565 13921 24568
rect 13955 24565 13967 24599
rect 13909 24559 13967 24565
rect 15841 24599 15899 24605
rect 15841 24565 15853 24599
rect 15887 24565 15899 24599
rect 15841 24559 15899 24565
rect 1104 24506 18860 24528
rect 1104 24454 7648 24506
rect 7700 24454 7712 24506
rect 7764 24454 7776 24506
rect 7828 24454 7840 24506
rect 7892 24454 14315 24506
rect 14367 24454 14379 24506
rect 14431 24454 14443 24506
rect 14495 24454 14507 24506
rect 14559 24454 18860 24506
rect 1104 24432 18860 24454
rect 1673 24395 1731 24401
rect 1673 24361 1685 24395
rect 1719 24392 1731 24395
rect 1854 24392 1860 24404
rect 1719 24364 1860 24392
rect 1719 24361 1731 24364
rect 1673 24355 1731 24361
rect 1854 24352 1860 24364
rect 1912 24352 1918 24404
rect 4982 24392 4988 24404
rect 4943 24364 4988 24392
rect 4982 24352 4988 24364
rect 5040 24352 5046 24404
rect 5534 24352 5540 24404
rect 5592 24392 5598 24404
rect 5905 24395 5963 24401
rect 5905 24392 5917 24395
rect 5592 24364 5917 24392
rect 5592 24352 5598 24364
rect 5905 24361 5917 24364
rect 5951 24392 5963 24395
rect 6546 24392 6552 24404
rect 5951 24364 6552 24392
rect 5951 24361 5963 24364
rect 5905 24355 5963 24361
rect 6546 24352 6552 24364
rect 6604 24352 6610 24404
rect 7098 24392 7104 24404
rect 7059 24364 7104 24392
rect 7098 24352 7104 24364
rect 7156 24352 7162 24404
rect 7374 24352 7380 24404
rect 7432 24392 7438 24404
rect 7837 24395 7895 24401
rect 7837 24392 7849 24395
rect 7432 24364 7849 24392
rect 7432 24352 7438 24364
rect 7837 24361 7849 24364
rect 7883 24361 7895 24395
rect 8294 24392 8300 24404
rect 8255 24364 8300 24392
rect 7837 24355 7895 24361
rect 8294 24352 8300 24364
rect 8352 24352 8358 24404
rect 10042 24352 10048 24404
rect 10100 24392 10106 24404
rect 10321 24395 10379 24401
rect 10321 24392 10333 24395
rect 10100 24364 10333 24392
rect 10100 24352 10106 24364
rect 10321 24361 10333 24364
rect 10367 24361 10379 24395
rect 10321 24355 10379 24361
rect 13817 24395 13875 24401
rect 13817 24361 13829 24395
rect 13863 24392 13875 24395
rect 13998 24392 14004 24404
rect 13863 24364 14004 24392
rect 13863 24361 13875 24364
rect 13817 24355 13875 24361
rect 13998 24352 14004 24364
rect 14056 24352 14062 24404
rect 14182 24392 14188 24404
rect 14143 24364 14188 24392
rect 14182 24352 14188 24364
rect 14240 24352 14246 24404
rect 16666 24392 16672 24404
rect 16627 24364 16672 24392
rect 16666 24352 16672 24364
rect 16724 24352 16730 24404
rect 16850 24352 16856 24404
rect 16908 24392 16914 24404
rect 17405 24395 17463 24401
rect 17405 24392 17417 24395
rect 16908 24364 17417 24392
rect 16908 24352 16914 24364
rect 17405 24361 17417 24364
rect 17451 24361 17463 24395
rect 17405 24355 17463 24361
rect 4525 24327 4583 24333
rect 4525 24293 4537 24327
rect 4571 24324 4583 24327
rect 6638 24324 6644 24336
rect 4571 24296 6644 24324
rect 4571 24293 4583 24296
rect 4525 24287 4583 24293
rect 2774 24216 2780 24268
rect 2832 24256 2838 24268
rect 5184 24265 5212 24296
rect 6638 24284 6644 24296
rect 6696 24284 6702 24336
rect 10226 24284 10232 24336
rect 10284 24324 10290 24336
rect 11517 24327 11575 24333
rect 11517 24324 11529 24327
rect 10284 24296 11529 24324
rect 10284 24284 10290 24296
rect 11517 24293 11529 24296
rect 11563 24293 11575 24327
rect 13446 24324 13452 24336
rect 13407 24296 13452 24324
rect 11517 24287 11575 24293
rect 13446 24284 13452 24296
rect 13504 24284 13510 24336
rect 16684 24324 16712 24352
rect 17218 24324 17224 24336
rect 16684 24296 17224 24324
rect 17218 24284 17224 24296
rect 17276 24284 17282 24336
rect 5169 24259 5227 24265
rect 2832 24228 2877 24256
rect 2832 24216 2838 24228
rect 5169 24225 5181 24259
rect 5215 24225 5227 24259
rect 5721 24259 5779 24265
rect 5721 24256 5733 24259
rect 5169 24219 5227 24225
rect 5460 24228 5733 24256
rect 1854 24148 1860 24200
rect 1912 24188 1918 24200
rect 2501 24191 2559 24197
rect 2501 24188 2513 24191
rect 1912 24160 2513 24188
rect 1912 24148 1918 24160
rect 2501 24157 2513 24160
rect 2547 24157 2559 24191
rect 2501 24151 2559 24157
rect 4893 24123 4951 24129
rect 4893 24089 4905 24123
rect 4939 24120 4951 24123
rect 5350 24120 5356 24132
rect 4939 24092 5356 24120
rect 4939 24089 4951 24092
rect 4893 24083 4951 24089
rect 5350 24080 5356 24092
rect 5408 24080 5414 24132
rect 4062 24052 4068 24064
rect 4023 24024 4068 24052
rect 4062 24012 4068 24024
rect 4120 24012 4126 24064
rect 5074 24012 5080 24064
rect 5132 24052 5138 24064
rect 5460 24061 5488 24228
rect 5721 24225 5733 24228
rect 5767 24256 5779 24259
rect 5902 24256 5908 24268
rect 5767 24228 5908 24256
rect 5767 24225 5779 24228
rect 5721 24219 5779 24225
rect 5902 24216 5908 24228
rect 5960 24216 5966 24268
rect 7006 24256 7012 24268
rect 6967 24228 7012 24256
rect 7006 24216 7012 24228
rect 7064 24216 7070 24268
rect 8938 24216 8944 24268
rect 8996 24256 9002 24268
rect 9125 24259 9183 24265
rect 9125 24256 9137 24259
rect 8996 24228 9137 24256
rect 8996 24216 9002 24228
rect 9125 24225 9137 24228
rect 9171 24225 9183 24259
rect 9125 24219 9183 24225
rect 9585 24259 9643 24265
rect 9585 24225 9597 24259
rect 9631 24256 9643 24259
rect 10042 24256 10048 24268
rect 9631 24228 10048 24256
rect 9631 24225 9643 24228
rect 9585 24219 9643 24225
rect 10042 24216 10048 24228
rect 10100 24216 10106 24268
rect 10781 24259 10839 24265
rect 10781 24225 10793 24259
rect 10827 24256 10839 24259
rect 10870 24256 10876 24268
rect 10827 24228 10876 24256
rect 10827 24225 10839 24228
rect 10781 24219 10839 24225
rect 10870 24216 10876 24228
rect 10928 24216 10934 24268
rect 11241 24259 11299 24265
rect 11241 24225 11253 24259
rect 11287 24256 11299 24259
rect 11330 24256 11336 24268
rect 11287 24228 11336 24256
rect 11287 24225 11299 24228
rect 11241 24219 11299 24225
rect 11330 24216 11336 24228
rect 11388 24216 11394 24268
rect 12894 24256 12900 24268
rect 12855 24228 12900 24256
rect 12894 24216 12900 24228
rect 12952 24216 12958 24268
rect 13170 24216 13176 24268
rect 13228 24256 13234 24268
rect 14369 24259 14427 24265
rect 14369 24256 14381 24259
rect 13228 24228 14381 24256
rect 13228 24216 13234 24228
rect 14369 24225 14381 24228
rect 14415 24256 14427 24259
rect 14550 24256 14556 24268
rect 14415 24228 14556 24256
rect 14415 24225 14427 24228
rect 14369 24219 14427 24225
rect 14550 24216 14556 24228
rect 14608 24216 14614 24268
rect 17034 24256 17040 24268
rect 16995 24228 17040 24256
rect 17034 24216 17040 24228
rect 17092 24216 17098 24268
rect 8389 24191 8447 24197
rect 8389 24157 8401 24191
rect 8435 24188 8447 24191
rect 9030 24188 9036 24200
rect 8435 24160 9036 24188
rect 8435 24157 8447 24160
rect 8389 24151 8447 24157
rect 9030 24148 9036 24160
rect 9088 24148 9094 24200
rect 12802 24148 12808 24200
rect 12860 24188 12866 24200
rect 13188 24188 13216 24216
rect 12860 24160 13216 24188
rect 15013 24191 15071 24197
rect 12860 24148 12866 24160
rect 15013 24157 15025 24191
rect 15059 24188 15071 24191
rect 15102 24188 15108 24200
rect 15059 24160 15108 24188
rect 15059 24157 15071 24160
rect 15013 24151 15071 24157
rect 15102 24148 15108 24160
rect 15160 24148 15166 24200
rect 6273 24123 6331 24129
rect 6273 24089 6285 24123
rect 6319 24120 6331 24123
rect 8018 24120 8024 24132
rect 6319 24092 8024 24120
rect 6319 24089 6331 24092
rect 6273 24083 6331 24089
rect 8018 24080 8024 24092
rect 8076 24080 8082 24132
rect 8662 24120 8668 24132
rect 8623 24092 8668 24120
rect 8662 24080 8668 24092
rect 8720 24080 8726 24132
rect 9858 24080 9864 24132
rect 9916 24120 9922 24132
rect 10597 24123 10655 24129
rect 10597 24120 10609 24123
rect 9916 24092 10609 24120
rect 9916 24080 9922 24092
rect 10597 24089 10609 24092
rect 10643 24089 10655 24123
rect 10597 24083 10655 24089
rect 5445 24055 5503 24061
rect 5445 24052 5457 24055
rect 5132 24024 5457 24052
rect 5132 24012 5138 24024
rect 5445 24021 5457 24024
rect 5491 24021 5503 24055
rect 6638 24052 6644 24064
rect 6599 24024 6644 24052
rect 5445 24015 5503 24021
rect 6638 24012 6644 24024
rect 6696 24012 6702 24064
rect 1104 23962 18860 23984
rect 1104 23910 4315 23962
rect 4367 23910 4379 23962
rect 4431 23910 4443 23962
rect 4495 23910 4507 23962
rect 4559 23910 10982 23962
rect 11034 23910 11046 23962
rect 11098 23910 11110 23962
rect 11162 23910 11174 23962
rect 11226 23910 17648 23962
rect 17700 23910 17712 23962
rect 17764 23910 17776 23962
rect 17828 23910 17840 23962
rect 17892 23910 18860 23962
rect 1104 23888 18860 23910
rect 11330 23848 11336 23860
rect 11291 23820 11336 23848
rect 11330 23808 11336 23820
rect 11388 23808 11394 23860
rect 11701 23851 11759 23857
rect 11701 23817 11713 23851
rect 11747 23848 11759 23851
rect 11974 23848 11980 23860
rect 11747 23820 11980 23848
rect 11747 23817 11759 23820
rect 11701 23811 11759 23817
rect 11974 23808 11980 23820
rect 12032 23808 12038 23860
rect 14550 23808 14556 23860
rect 14608 23848 14614 23860
rect 14645 23851 14703 23857
rect 14645 23848 14657 23851
rect 14608 23820 14657 23848
rect 14608 23808 14614 23820
rect 14645 23817 14657 23820
rect 14691 23817 14703 23851
rect 14645 23811 14703 23817
rect 10137 23783 10195 23789
rect 10137 23749 10149 23783
rect 10183 23780 10195 23783
rect 10870 23780 10876 23792
rect 10183 23752 10876 23780
rect 10183 23749 10195 23752
rect 10137 23743 10195 23749
rect 10870 23740 10876 23752
rect 10928 23740 10934 23792
rect 15930 23740 15936 23792
rect 15988 23780 15994 23792
rect 16942 23780 16948 23792
rect 15988 23752 16948 23780
rect 15988 23740 15994 23752
rect 16942 23740 16948 23752
rect 17000 23780 17006 23792
rect 18049 23783 18107 23789
rect 18049 23780 18061 23783
rect 17000 23752 18061 23780
rect 17000 23740 17006 23752
rect 1762 23712 1768 23724
rect 1723 23684 1768 23712
rect 1762 23672 1768 23684
rect 1820 23672 1826 23724
rect 5629 23715 5687 23721
rect 5629 23681 5641 23715
rect 5675 23712 5687 23715
rect 5994 23712 6000 23724
rect 5675 23684 6000 23712
rect 5675 23681 5687 23684
rect 5629 23675 5687 23681
rect 5994 23672 6000 23684
rect 6052 23672 6058 23724
rect 6733 23715 6791 23721
rect 6733 23681 6745 23715
rect 6779 23712 6791 23715
rect 7006 23712 7012 23724
rect 6779 23684 7012 23712
rect 6779 23681 6791 23684
rect 6733 23675 6791 23681
rect 7006 23672 7012 23684
rect 7064 23672 7070 23724
rect 8478 23672 8484 23724
rect 8536 23712 8542 23724
rect 10042 23712 10048 23724
rect 8536 23684 10048 23712
rect 8536 23672 8542 23684
rect 10042 23672 10048 23684
rect 10100 23712 10106 23724
rect 10689 23715 10747 23721
rect 10689 23712 10701 23715
rect 10100 23684 10701 23712
rect 10100 23672 10106 23684
rect 10689 23681 10701 23684
rect 10735 23681 10747 23715
rect 16758 23712 16764 23724
rect 16719 23684 16764 23712
rect 10689 23675 10747 23681
rect 16758 23672 16764 23684
rect 16816 23672 16822 23724
rect 17328 23721 17356 23752
rect 18049 23749 18061 23752
rect 18095 23749 18107 23783
rect 18049 23743 18107 23749
rect 17313 23715 17371 23721
rect 17313 23681 17325 23715
rect 17359 23681 17371 23715
rect 17313 23675 17371 23681
rect 17402 23672 17408 23724
rect 17460 23712 17466 23724
rect 17773 23715 17831 23721
rect 17773 23712 17785 23715
rect 17460 23684 17785 23712
rect 17460 23672 17466 23684
rect 17773 23681 17785 23684
rect 17819 23681 17831 23715
rect 17773 23675 17831 23681
rect 1489 23647 1547 23653
rect 1489 23613 1501 23647
rect 1535 23644 1547 23647
rect 1854 23644 1860 23656
rect 1535 23616 1860 23644
rect 1535 23613 1547 23616
rect 1489 23607 1547 23613
rect 1854 23604 1860 23616
rect 1912 23604 1918 23656
rect 4433 23647 4491 23653
rect 4433 23613 4445 23647
rect 4479 23644 4491 23647
rect 4893 23647 4951 23653
rect 4893 23644 4905 23647
rect 4479 23616 4905 23644
rect 4479 23613 4491 23616
rect 4433 23607 4491 23613
rect 4893 23613 4905 23616
rect 4939 23644 4951 23647
rect 5442 23644 5448 23656
rect 4939 23616 5448 23644
rect 4939 23613 4951 23616
rect 4893 23607 4951 23613
rect 5442 23604 5448 23616
rect 5500 23604 5506 23656
rect 6546 23644 6552 23656
rect 6507 23616 6552 23644
rect 6546 23604 6552 23616
rect 6604 23604 6610 23656
rect 7098 23644 7104 23656
rect 7059 23616 7104 23644
rect 7098 23604 7104 23616
rect 7156 23604 7162 23656
rect 7282 23644 7288 23656
rect 7243 23616 7288 23644
rect 7282 23604 7288 23616
rect 7340 23604 7346 23656
rect 7374 23604 7380 23656
rect 7432 23644 7438 23656
rect 7653 23647 7711 23653
rect 7653 23644 7665 23647
rect 7432 23616 7665 23644
rect 7432 23604 7438 23616
rect 7653 23613 7665 23616
rect 7699 23613 7711 23647
rect 8018 23644 8024 23656
rect 7979 23616 8024 23644
rect 7653 23607 7711 23613
rect 8018 23604 8024 23616
rect 8076 23604 8082 23656
rect 9677 23647 9735 23653
rect 9677 23644 9689 23647
rect 9048 23616 9689 23644
rect 3142 23576 3148 23588
rect 3103 23548 3148 23576
rect 3142 23536 3148 23548
rect 3200 23536 3206 23588
rect 4801 23579 4859 23585
rect 4801 23545 4813 23579
rect 4847 23576 4859 23579
rect 5166 23576 5172 23588
rect 4847 23548 5172 23576
rect 4847 23545 4859 23548
rect 4801 23539 4859 23545
rect 5166 23536 5172 23548
rect 5224 23536 5230 23588
rect 5261 23579 5319 23585
rect 5261 23545 5273 23579
rect 5307 23576 5319 23579
rect 5997 23579 6055 23585
rect 5997 23576 6009 23579
rect 5307 23548 6009 23576
rect 5307 23545 5319 23548
rect 5261 23539 5319 23545
rect 5997 23545 6009 23548
rect 6043 23576 6055 23579
rect 6365 23579 6423 23585
rect 6365 23576 6377 23579
rect 6043 23548 6377 23576
rect 6043 23545 6055 23548
rect 5997 23539 6055 23545
rect 6365 23545 6377 23548
rect 6411 23576 6423 23579
rect 7116 23576 7144 23604
rect 6411 23548 7144 23576
rect 6411 23545 6423 23548
rect 6365 23539 6423 23545
rect 9048 23520 9076 23616
rect 9677 23613 9689 23616
rect 9723 23613 9735 23647
rect 9677 23607 9735 23613
rect 10413 23647 10471 23653
rect 10413 23613 10425 23647
rect 10459 23613 10471 23647
rect 12066 23644 12072 23656
rect 12027 23616 12072 23644
rect 10413 23607 10471 23613
rect 9493 23579 9551 23585
rect 9493 23545 9505 23579
rect 9539 23576 9551 23579
rect 10134 23576 10140 23588
rect 9539 23548 10140 23576
rect 9539 23545 9551 23548
rect 9493 23539 9551 23545
rect 10134 23536 10140 23548
rect 10192 23576 10198 23588
rect 10428 23576 10456 23607
rect 12066 23604 12072 23616
rect 12124 23604 12130 23656
rect 12894 23644 12900 23656
rect 12855 23616 12900 23644
rect 12894 23604 12900 23616
rect 12952 23604 12958 23656
rect 13630 23644 13636 23656
rect 13591 23616 13636 23644
rect 13630 23604 13636 23616
rect 13688 23604 13694 23656
rect 14001 23647 14059 23653
rect 14001 23613 14013 23647
rect 14047 23644 14059 23647
rect 14090 23644 14096 23656
rect 14047 23616 14096 23644
rect 14047 23613 14059 23616
rect 14001 23607 14059 23613
rect 14090 23604 14096 23616
rect 14148 23604 14154 23656
rect 14369 23647 14427 23653
rect 14369 23613 14381 23647
rect 14415 23644 14427 23647
rect 15102 23644 15108 23656
rect 14415 23616 15108 23644
rect 14415 23613 14427 23616
rect 14369 23607 14427 23613
rect 10192 23548 10456 23576
rect 12529 23579 12587 23585
rect 10192 23536 10198 23548
rect 12529 23545 12541 23579
rect 12575 23576 12587 23579
rect 12618 23576 12624 23588
rect 12575 23548 12624 23576
rect 12575 23545 12587 23548
rect 12529 23539 12587 23545
rect 12618 23536 12624 23548
rect 12676 23536 12682 23588
rect 13541 23579 13599 23585
rect 13541 23545 13553 23579
rect 13587 23576 13599 23579
rect 14384 23576 14412 23607
rect 15102 23604 15108 23616
rect 15160 23604 15166 23656
rect 15749 23647 15807 23653
rect 15749 23613 15761 23647
rect 15795 23644 15807 23647
rect 15838 23644 15844 23656
rect 15795 23616 15844 23644
rect 15795 23613 15807 23616
rect 15749 23607 15807 23613
rect 15838 23604 15844 23616
rect 15896 23644 15902 23656
rect 16209 23647 16267 23653
rect 16209 23644 16221 23647
rect 15896 23616 16221 23644
rect 15896 23604 15902 23616
rect 16209 23613 16221 23616
rect 16255 23613 16267 23647
rect 17126 23644 17132 23656
rect 16209 23607 16267 23613
rect 16776 23616 17132 23644
rect 16776 23588 16804 23616
rect 17126 23604 17132 23616
rect 17184 23604 17190 23656
rect 17589 23647 17647 23653
rect 17589 23613 17601 23647
rect 17635 23613 17647 23647
rect 17589 23607 17647 23613
rect 13587 23548 14412 23576
rect 13587 23545 13599 23548
rect 13541 23539 13599 23545
rect 16758 23536 16764 23588
rect 16816 23536 16822 23588
rect 16850 23536 16856 23588
rect 16908 23576 16914 23588
rect 17604 23576 17632 23607
rect 16908 23548 17632 23576
rect 16908 23536 16914 23548
rect 17328 23520 17356 23548
rect 5074 23508 5080 23520
rect 5035 23480 5080 23508
rect 5074 23468 5080 23480
rect 5132 23468 5138 23520
rect 8757 23511 8815 23517
rect 8757 23477 8769 23511
rect 8803 23508 8815 23511
rect 9030 23508 9036 23520
rect 8803 23480 9036 23508
rect 8803 23477 8815 23480
rect 8757 23471 8815 23477
rect 9030 23468 9036 23480
rect 9088 23468 9094 23520
rect 15930 23508 15936 23520
rect 15891 23480 15936 23508
rect 15930 23468 15936 23480
rect 15988 23468 15994 23520
rect 16206 23468 16212 23520
rect 16264 23508 16270 23520
rect 16577 23511 16635 23517
rect 16577 23508 16589 23511
rect 16264 23480 16589 23508
rect 16264 23468 16270 23480
rect 16577 23477 16589 23480
rect 16623 23508 16635 23511
rect 17034 23508 17040 23520
rect 16623 23480 17040 23508
rect 16623 23477 16635 23480
rect 16577 23471 16635 23477
rect 17034 23468 17040 23480
rect 17092 23468 17098 23520
rect 17310 23468 17316 23520
rect 17368 23468 17374 23520
rect 1104 23418 18860 23440
rect 1104 23366 7648 23418
rect 7700 23366 7712 23418
rect 7764 23366 7776 23418
rect 7828 23366 7840 23418
rect 7892 23366 14315 23418
rect 14367 23366 14379 23418
rect 14431 23366 14443 23418
rect 14495 23366 14507 23418
rect 14559 23366 18860 23418
rect 1104 23344 18860 23366
rect 1673 23307 1731 23313
rect 1673 23273 1685 23307
rect 1719 23304 1731 23307
rect 1762 23304 1768 23316
rect 1719 23276 1768 23304
rect 1719 23273 1731 23276
rect 1673 23267 1731 23273
rect 1762 23264 1768 23276
rect 1820 23264 1826 23316
rect 2593 23307 2651 23313
rect 2593 23273 2605 23307
rect 2639 23304 2651 23307
rect 2682 23304 2688 23316
rect 2639 23276 2688 23304
rect 2639 23273 2651 23276
rect 2593 23267 2651 23273
rect 2682 23264 2688 23276
rect 2740 23264 2746 23316
rect 2961 23307 3019 23313
rect 2961 23273 2973 23307
rect 3007 23304 3019 23307
rect 3697 23307 3755 23313
rect 3697 23304 3709 23307
rect 3007 23276 3709 23304
rect 3007 23273 3019 23276
rect 2961 23267 3019 23273
rect 3697 23273 3709 23276
rect 3743 23304 3755 23307
rect 3878 23304 3884 23316
rect 3743 23276 3884 23304
rect 3743 23273 3755 23276
rect 3697 23267 3755 23273
rect 1854 22992 1860 23044
rect 1912 23032 1918 23044
rect 1949 23035 2007 23041
rect 1949 23032 1961 23035
rect 1912 23004 1961 23032
rect 1912 22992 1918 23004
rect 1949 23001 1961 23004
rect 1995 23032 2007 23035
rect 2976 23032 3004 23267
rect 3878 23264 3884 23276
rect 3936 23304 3942 23316
rect 6549 23307 6607 23313
rect 3936 23276 4016 23304
rect 3936 23264 3942 23276
rect 3786 23128 3792 23180
rect 3844 23168 3850 23180
rect 3988 23177 4016 23276
rect 6549 23273 6561 23307
rect 6595 23304 6607 23307
rect 7374 23304 7380 23316
rect 6595 23276 7380 23304
rect 6595 23273 6607 23276
rect 6549 23267 6607 23273
rect 7374 23264 7380 23276
rect 7432 23264 7438 23316
rect 8478 23304 8484 23316
rect 8439 23276 8484 23304
rect 8478 23264 8484 23276
rect 8536 23264 8542 23316
rect 8849 23307 8907 23313
rect 8849 23273 8861 23307
rect 8895 23304 8907 23307
rect 8938 23304 8944 23316
rect 8895 23276 8944 23304
rect 8895 23273 8907 23276
rect 8849 23267 8907 23273
rect 8938 23264 8944 23276
rect 8996 23264 9002 23316
rect 11054 23304 11060 23316
rect 11015 23276 11060 23304
rect 11054 23264 11060 23276
rect 11112 23264 11118 23316
rect 13630 23304 13636 23316
rect 13591 23276 13636 23304
rect 13630 23264 13636 23276
rect 13688 23264 13694 23316
rect 5258 23196 5264 23248
rect 5316 23236 5322 23248
rect 7929 23239 7987 23245
rect 7929 23236 7941 23239
rect 5316 23208 7941 23236
rect 5316 23196 5322 23208
rect 7929 23205 7941 23208
rect 7975 23205 7987 23239
rect 7929 23199 7987 23205
rect 12342 23196 12348 23248
rect 12400 23236 12406 23248
rect 13648 23236 13676 23264
rect 14918 23236 14924 23248
rect 12400 23208 14924 23236
rect 12400 23196 12406 23208
rect 14918 23196 14924 23208
rect 14976 23196 14982 23248
rect 15010 23196 15016 23248
rect 15068 23236 15074 23248
rect 15841 23239 15899 23245
rect 15841 23236 15853 23239
rect 15068 23208 15853 23236
rect 15068 23196 15074 23208
rect 15841 23205 15853 23208
rect 15887 23236 15899 23239
rect 15887 23208 16988 23236
rect 15887 23205 15899 23208
rect 15841 23199 15899 23205
rect 3881 23171 3939 23177
rect 3881 23168 3893 23171
rect 3844 23140 3893 23168
rect 3844 23128 3850 23140
rect 3881 23137 3893 23140
rect 3927 23137 3939 23171
rect 3881 23131 3939 23137
rect 3973 23171 4031 23177
rect 3973 23137 3985 23171
rect 4019 23168 4031 23171
rect 4706 23168 4712 23180
rect 4019 23140 4712 23168
rect 4019 23137 4031 23140
rect 3973 23131 4031 23137
rect 4706 23128 4712 23140
rect 4764 23128 4770 23180
rect 5350 23128 5356 23180
rect 5408 23168 5414 23180
rect 6546 23168 6552 23180
rect 5408 23140 6552 23168
rect 5408 23128 5414 23140
rect 6546 23128 6552 23140
rect 6604 23168 6610 23180
rect 6825 23171 6883 23177
rect 6825 23168 6837 23171
rect 6604 23140 6837 23168
rect 6604 23128 6610 23140
rect 6825 23137 6837 23140
rect 6871 23168 6883 23171
rect 7282 23168 7288 23180
rect 6871 23140 7288 23168
rect 6871 23137 6883 23140
rect 6825 23131 6883 23137
rect 7282 23128 7288 23140
rect 7340 23128 7346 23180
rect 7469 23171 7527 23177
rect 7469 23137 7481 23171
rect 7515 23168 7527 23171
rect 7558 23168 7564 23180
rect 7515 23140 7564 23168
rect 7515 23137 7527 23140
rect 7469 23131 7527 23137
rect 7558 23128 7564 23140
rect 7616 23128 7622 23180
rect 7653 23171 7711 23177
rect 7653 23137 7665 23171
rect 7699 23137 7711 23171
rect 7653 23131 7711 23137
rect 9861 23171 9919 23177
rect 9861 23137 9873 23171
rect 9907 23168 9919 23171
rect 9950 23168 9956 23180
rect 9907 23140 9956 23168
rect 9907 23137 9919 23140
rect 9861 23131 9919 23137
rect 4154 23060 4160 23112
rect 4212 23100 4218 23112
rect 4249 23103 4307 23109
rect 4249 23100 4261 23103
rect 4212 23072 4261 23100
rect 4212 23060 4218 23072
rect 4249 23069 4261 23072
rect 4295 23069 4307 23103
rect 4249 23063 4307 23069
rect 5902 23060 5908 23112
rect 5960 23100 5966 23112
rect 5997 23103 6055 23109
rect 5997 23100 6009 23103
rect 5960 23072 6009 23100
rect 5960 23060 5966 23072
rect 5997 23069 6009 23072
rect 6043 23100 6055 23103
rect 7374 23100 7380 23112
rect 6043 23072 7380 23100
rect 6043 23069 6055 23072
rect 5997 23063 6055 23069
rect 7374 23060 7380 23072
rect 7432 23100 7438 23112
rect 7668 23100 7696 23131
rect 9950 23128 9956 23140
rect 10008 23128 10014 23180
rect 10229 23171 10287 23177
rect 10229 23137 10241 23171
rect 10275 23168 10287 23171
rect 10410 23168 10416 23180
rect 10275 23140 10416 23168
rect 10275 23137 10287 23140
rect 10229 23131 10287 23137
rect 10410 23128 10416 23140
rect 10468 23128 10474 23180
rect 10594 23168 10600 23180
rect 10555 23140 10600 23168
rect 10594 23128 10600 23140
rect 10652 23128 10658 23180
rect 11882 23128 11888 23180
rect 11940 23168 11946 23180
rect 12434 23168 12440 23180
rect 11940 23140 12440 23168
rect 11940 23128 11946 23140
rect 12434 23128 12440 23140
rect 12492 23168 12498 23180
rect 12894 23168 12900 23180
rect 12492 23140 12585 23168
rect 12855 23140 12900 23168
rect 12492 23128 12498 23140
rect 12894 23128 12900 23140
rect 12952 23128 12958 23180
rect 13906 23128 13912 23180
rect 13964 23168 13970 23180
rect 14369 23171 14427 23177
rect 14369 23168 14381 23171
rect 13964 23140 14381 23168
rect 13964 23128 13970 23140
rect 14369 23137 14381 23140
rect 14415 23137 14427 23171
rect 14550 23168 14556 23180
rect 14511 23140 14556 23168
rect 14369 23131 14427 23137
rect 14550 23128 14556 23140
rect 14608 23128 14614 23180
rect 14737 23171 14795 23177
rect 14737 23137 14749 23171
rect 14783 23137 14795 23171
rect 16574 23168 16580 23180
rect 16535 23140 16580 23168
rect 14737 23131 14795 23137
rect 7432 23072 7696 23100
rect 10781 23103 10839 23109
rect 7432 23060 7438 23072
rect 10781 23069 10793 23103
rect 10827 23100 10839 23103
rect 11422 23100 11428 23112
rect 10827 23072 11428 23100
rect 10827 23069 10839 23072
rect 10781 23063 10839 23069
rect 11422 23060 11428 23072
rect 11480 23060 11486 23112
rect 13262 23100 13268 23112
rect 13223 23072 13268 23100
rect 13262 23060 13268 23072
rect 13320 23100 13326 23112
rect 14752 23100 14780 23131
rect 16574 23128 16580 23140
rect 16632 23128 16638 23180
rect 16960 23177 16988 23208
rect 16945 23171 17003 23177
rect 16945 23137 16957 23171
rect 16991 23137 17003 23171
rect 16945 23131 17003 23137
rect 17034 23128 17040 23180
rect 17092 23168 17098 23180
rect 17092 23140 17137 23168
rect 17092 23128 17098 23140
rect 13320 23072 14780 23100
rect 13320 23060 13326 23072
rect 16114 23060 16120 23112
rect 16172 23100 16178 23112
rect 16485 23103 16543 23109
rect 16485 23100 16497 23103
rect 16172 23072 16497 23100
rect 16172 23060 16178 23072
rect 16485 23069 16497 23072
rect 16531 23069 16543 23103
rect 16485 23063 16543 23069
rect 1995 23004 3004 23032
rect 14185 23035 14243 23041
rect 1995 23001 2007 23004
rect 1949 22995 2007 23001
rect 14185 23001 14197 23035
rect 14231 23032 14243 23035
rect 15470 23032 15476 23044
rect 14231 23004 15476 23032
rect 14231 23001 14243 23004
rect 14185 22995 14243 23001
rect 15470 22992 15476 23004
rect 15528 22992 15534 23044
rect 5350 22964 5356 22976
rect 5311 22936 5356 22964
rect 5350 22924 5356 22936
rect 5408 22924 5414 22976
rect 9490 22964 9496 22976
rect 9451 22936 9496 22964
rect 9490 22924 9496 22936
rect 9548 22924 9554 22976
rect 12621 22967 12679 22973
rect 12621 22933 12633 22967
rect 12667 22964 12679 22967
rect 12710 22964 12716 22976
rect 12667 22936 12716 22964
rect 12667 22933 12679 22936
rect 12621 22927 12679 22933
rect 12710 22924 12716 22936
rect 12768 22924 12774 22976
rect 16022 22964 16028 22976
rect 15983 22936 16028 22964
rect 16022 22924 16028 22936
rect 16080 22924 16086 22976
rect 17034 22924 17040 22976
rect 17092 22964 17098 22976
rect 17402 22964 17408 22976
rect 17092 22936 17408 22964
rect 17092 22924 17098 22936
rect 17402 22924 17408 22936
rect 17460 22924 17466 22976
rect 1104 22874 18860 22896
rect 1104 22822 4315 22874
rect 4367 22822 4379 22874
rect 4431 22822 4443 22874
rect 4495 22822 4507 22874
rect 4559 22822 10982 22874
rect 11034 22822 11046 22874
rect 11098 22822 11110 22874
rect 11162 22822 11174 22874
rect 11226 22822 17648 22874
rect 17700 22822 17712 22874
rect 17764 22822 17776 22874
rect 17828 22822 17840 22874
rect 17892 22822 18860 22874
rect 1104 22800 18860 22822
rect 4062 22720 4068 22772
rect 4120 22760 4126 22772
rect 4249 22763 4307 22769
rect 4249 22760 4261 22763
rect 4120 22732 4261 22760
rect 4120 22720 4126 22732
rect 4249 22729 4261 22732
rect 4295 22729 4307 22763
rect 6546 22760 6552 22772
rect 6507 22732 6552 22760
rect 4249 22723 4307 22729
rect 6546 22720 6552 22732
rect 6604 22760 6610 22772
rect 6730 22760 6736 22772
rect 6604 22732 6736 22760
rect 6604 22720 6610 22732
rect 6730 22720 6736 22732
rect 6788 22720 6794 22772
rect 7929 22763 7987 22769
rect 7929 22729 7941 22763
rect 7975 22760 7987 22763
rect 8110 22760 8116 22772
rect 7975 22732 8116 22760
rect 7975 22729 7987 22732
rect 7929 22723 7987 22729
rect 8110 22720 8116 22732
rect 8168 22720 8174 22772
rect 9125 22763 9183 22769
rect 9125 22729 9137 22763
rect 9171 22760 9183 22763
rect 10410 22760 10416 22772
rect 9171 22732 10416 22760
rect 9171 22729 9183 22732
rect 9125 22723 9183 22729
rect 10410 22720 10416 22732
rect 10468 22720 10474 22772
rect 10594 22720 10600 22772
rect 10652 22760 10658 22772
rect 11057 22763 11115 22769
rect 11057 22760 11069 22763
rect 10652 22732 11069 22760
rect 10652 22720 10658 22732
rect 10980 22704 11008 22732
rect 11057 22729 11069 22732
rect 11103 22729 11115 22763
rect 11422 22760 11428 22772
rect 11383 22732 11428 22760
rect 11057 22723 11115 22729
rect 11422 22720 11428 22732
rect 11480 22720 11486 22772
rect 12897 22763 12955 22769
rect 12897 22760 12909 22763
rect 12452 22732 12909 22760
rect 9401 22695 9459 22701
rect 9401 22661 9413 22695
rect 9447 22692 9459 22695
rect 9950 22692 9956 22704
rect 9447 22664 9956 22692
rect 9447 22661 9459 22664
rect 9401 22655 9459 22661
rect 9950 22652 9956 22664
rect 10008 22652 10014 22704
rect 10962 22652 10968 22704
rect 11020 22652 11026 22704
rect 4709 22627 4767 22633
rect 4709 22593 4721 22627
rect 4755 22624 4767 22627
rect 5350 22624 5356 22636
rect 4755 22596 5356 22624
rect 4755 22593 4767 22596
rect 4709 22587 4767 22593
rect 5350 22584 5356 22596
rect 5408 22624 5414 22636
rect 5445 22627 5503 22633
rect 5445 22624 5457 22627
rect 5408 22596 5457 22624
rect 5408 22584 5414 22596
rect 5445 22593 5457 22596
rect 5491 22593 5503 22627
rect 5445 22587 5503 22593
rect 8389 22627 8447 22633
rect 8389 22593 8401 22627
rect 8435 22624 8447 22627
rect 9490 22624 9496 22636
rect 8435 22596 9496 22624
rect 8435 22593 8447 22596
rect 8389 22587 8447 22593
rect 9490 22584 9496 22596
rect 9548 22624 9554 22636
rect 11440 22624 11468 22720
rect 12452 22692 12480 22732
rect 12897 22729 12909 22732
rect 12943 22760 12955 22763
rect 13078 22760 13084 22772
rect 12943 22732 13084 22760
rect 12943 22729 12955 22732
rect 12897 22723 12955 22729
rect 13078 22720 13084 22732
rect 13136 22720 13142 22772
rect 13188 22732 14320 22760
rect 13188 22701 13216 22732
rect 9548 22596 9720 22624
rect 9548 22584 9554 22596
rect 4982 22556 4988 22568
rect 4943 22528 4988 22556
rect 4982 22516 4988 22528
rect 5040 22516 5046 22568
rect 5166 22556 5172 22568
rect 5127 22528 5172 22556
rect 5166 22516 5172 22528
rect 5224 22516 5230 22568
rect 8110 22556 8116 22568
rect 8071 22528 8116 22556
rect 8110 22516 8116 22528
rect 8168 22556 8174 22568
rect 8294 22556 8300 22568
rect 8168 22528 8300 22556
rect 8168 22516 8174 22528
rect 8294 22516 8300 22528
rect 8352 22516 8358 22568
rect 9692 22565 9720 22596
rect 10428 22596 11468 22624
rect 12360 22664 12480 22692
rect 12529 22695 12587 22701
rect 10428 22565 10456 22596
rect 8757 22559 8815 22565
rect 8757 22525 8769 22559
rect 8803 22525 8815 22559
rect 8757 22519 8815 22525
rect 9677 22559 9735 22565
rect 9677 22525 9689 22559
rect 9723 22525 9735 22559
rect 9677 22519 9735 22525
rect 10413 22559 10471 22565
rect 10413 22525 10425 22559
rect 10459 22525 10471 22559
rect 10413 22519 10471 22525
rect 7558 22488 7564 22500
rect 7300 22460 7564 22488
rect 3786 22420 3792 22432
rect 3747 22392 3792 22420
rect 3786 22380 3792 22392
rect 3844 22380 3850 22432
rect 4798 22420 4804 22432
rect 4759 22392 4804 22420
rect 4798 22380 4804 22392
rect 4856 22380 4862 22432
rect 7098 22420 7104 22432
rect 7059 22392 7104 22420
rect 7098 22380 7104 22392
rect 7156 22420 7162 22432
rect 7300 22420 7328 22460
rect 7558 22448 7564 22460
rect 7616 22448 7622 22500
rect 8478 22448 8484 22500
rect 8536 22488 8542 22500
rect 8772 22488 8800 22519
rect 10502 22516 10508 22568
rect 10560 22556 10566 22568
rect 12360 22565 12388 22664
rect 12529 22661 12541 22695
rect 12575 22692 12587 22695
rect 13173 22695 13231 22701
rect 13173 22692 13185 22695
rect 12575 22664 13185 22692
rect 12575 22661 12587 22664
rect 12529 22655 12587 22661
rect 13173 22661 13185 22664
rect 13219 22661 13231 22695
rect 13630 22692 13636 22704
rect 13591 22664 13636 22692
rect 13173 22655 13231 22661
rect 13630 22652 13636 22664
rect 13688 22652 13694 22704
rect 12894 22584 12900 22636
rect 12952 22624 12958 22636
rect 14292 22633 14320 22732
rect 14826 22720 14832 22772
rect 14884 22760 14890 22772
rect 15565 22763 15623 22769
rect 15565 22760 15577 22763
rect 14884 22732 15577 22760
rect 14884 22720 14890 22732
rect 15565 22729 15577 22732
rect 15611 22729 15623 22763
rect 15565 22723 15623 22729
rect 16114 22720 16120 22772
rect 16172 22760 16178 22772
rect 16485 22763 16543 22769
rect 16485 22760 16497 22763
rect 16172 22732 16497 22760
rect 16172 22720 16178 22732
rect 16485 22729 16497 22732
rect 16531 22729 16543 22763
rect 16485 22723 16543 22729
rect 14918 22652 14924 22704
rect 14976 22692 14982 22704
rect 15013 22695 15071 22701
rect 15013 22692 15025 22695
rect 14976 22664 15025 22692
rect 14976 22652 14982 22664
rect 15013 22661 15025 22664
rect 15059 22661 15071 22695
rect 17494 22692 17500 22704
rect 17455 22664 17500 22692
rect 15013 22655 15071 22661
rect 14277 22627 14335 22633
rect 12952 22596 14228 22624
rect 12952 22584 12958 22596
rect 12345 22559 12403 22565
rect 10560 22528 10605 22556
rect 10560 22516 10566 22528
rect 12345 22525 12357 22559
rect 12391 22525 12403 22559
rect 12345 22519 12403 22525
rect 13078 22516 13084 22568
rect 13136 22556 13142 22568
rect 13354 22556 13360 22568
rect 13136 22528 13360 22556
rect 13136 22516 13142 22528
rect 13354 22516 13360 22528
rect 13412 22516 13418 22568
rect 13446 22516 13452 22568
rect 13504 22556 13510 22568
rect 14200 22565 14228 22596
rect 14277 22593 14289 22627
rect 14323 22624 14335 22627
rect 14550 22624 14556 22636
rect 14323 22596 14556 22624
rect 14323 22593 14335 22596
rect 14277 22587 14335 22593
rect 14550 22584 14556 22596
rect 14608 22624 14614 22636
rect 14645 22627 14703 22633
rect 14645 22624 14657 22627
rect 14608 22596 14657 22624
rect 14608 22584 14614 22596
rect 14645 22593 14657 22596
rect 14691 22593 14703 22627
rect 14645 22587 14703 22593
rect 13817 22559 13875 22565
rect 13817 22556 13829 22559
rect 13504 22528 13829 22556
rect 13504 22516 13510 22528
rect 13817 22525 13829 22528
rect 13863 22525 13875 22559
rect 13817 22519 13875 22525
rect 14185 22559 14243 22565
rect 14185 22525 14197 22559
rect 14231 22525 14243 22559
rect 15028 22556 15056 22655
rect 17494 22652 17500 22664
rect 17552 22652 17558 22704
rect 15194 22584 15200 22636
rect 15252 22624 15258 22636
rect 15289 22627 15347 22633
rect 15289 22624 15301 22627
rect 15252 22596 15301 22624
rect 15252 22584 15258 22596
rect 15289 22593 15301 22596
rect 15335 22624 15347 22627
rect 16117 22627 16175 22633
rect 16117 22624 16129 22627
rect 15335 22596 16129 22624
rect 15335 22593 15347 22596
rect 15289 22587 15347 22593
rect 16117 22593 16129 22596
rect 16163 22593 16175 22627
rect 16117 22587 16175 22593
rect 16758 22584 16764 22636
rect 16816 22624 16822 22636
rect 18049 22627 18107 22633
rect 18049 22624 18061 22627
rect 16816 22596 18061 22624
rect 16816 22584 16822 22596
rect 15381 22559 15439 22565
rect 15381 22556 15393 22559
rect 15028 22528 15393 22556
rect 14185 22519 14243 22525
rect 15381 22525 15393 22528
rect 15427 22525 15439 22559
rect 16666 22556 16672 22568
rect 16627 22528 16672 22556
rect 15381 22519 15439 22525
rect 16666 22516 16672 22528
rect 16724 22516 16730 22568
rect 17052 22565 17080 22596
rect 18049 22593 18061 22596
rect 18095 22593 18107 22627
rect 18049 22587 18107 22593
rect 17037 22559 17095 22565
rect 17037 22525 17049 22559
rect 17083 22525 17095 22559
rect 17037 22519 17095 22525
rect 17589 22559 17647 22565
rect 17589 22525 17601 22559
rect 17635 22556 17647 22559
rect 18417 22559 18475 22565
rect 18417 22556 18429 22559
rect 17635 22528 18429 22556
rect 17635 22525 17647 22528
rect 17589 22519 17647 22525
rect 18417 22525 18429 22528
rect 18463 22525 18475 22559
rect 18417 22519 18475 22525
rect 9858 22488 9864 22500
rect 8536 22460 9864 22488
rect 8536 22448 8542 22460
rect 9858 22448 9864 22460
rect 9916 22448 9922 22500
rect 16850 22448 16856 22500
rect 16908 22488 16914 22500
rect 17604 22488 17632 22519
rect 16908 22460 17632 22488
rect 16908 22448 16914 22460
rect 7156 22392 7328 22420
rect 7156 22380 7162 22392
rect 7374 22380 7380 22432
rect 7432 22420 7438 22432
rect 7469 22423 7527 22429
rect 7469 22420 7481 22423
rect 7432 22392 7481 22420
rect 7432 22380 7438 22392
rect 7469 22389 7481 22392
rect 7515 22389 7527 22423
rect 9766 22420 9772 22432
rect 9727 22392 9772 22420
rect 7469 22383 7527 22389
rect 9766 22380 9772 22392
rect 9824 22380 9830 22432
rect 11330 22380 11336 22432
rect 11388 22420 11394 22432
rect 12161 22423 12219 22429
rect 12161 22420 12173 22423
rect 11388 22392 12173 22420
rect 11388 22380 11394 22392
rect 12161 22389 12173 22392
rect 12207 22420 12219 22423
rect 12434 22420 12440 22432
rect 12207 22392 12440 22420
rect 12207 22389 12219 22392
rect 12161 22383 12219 22389
rect 12434 22380 12440 22392
rect 12492 22380 12498 22432
rect 1104 22330 18860 22352
rect 1104 22278 7648 22330
rect 7700 22278 7712 22330
rect 7764 22278 7776 22330
rect 7828 22278 7840 22330
rect 7892 22278 14315 22330
rect 14367 22278 14379 22330
rect 14431 22278 14443 22330
rect 14495 22278 14507 22330
rect 14559 22278 18860 22330
rect 1104 22256 18860 22278
rect 3786 22176 3792 22228
rect 3844 22216 3850 22228
rect 4525 22219 4583 22225
rect 3844 22188 4108 22216
rect 3844 22176 3850 22188
rect 3878 22108 3884 22160
rect 3936 22148 3942 22160
rect 3973 22151 4031 22157
rect 3973 22148 3985 22151
rect 3936 22120 3985 22148
rect 3936 22108 3942 22120
rect 3973 22117 3985 22120
rect 4019 22117 4031 22151
rect 3973 22111 4031 22117
rect 1854 22080 1860 22092
rect 1815 22052 1860 22080
rect 1854 22040 1860 22052
rect 1912 22040 1918 22092
rect 2130 22080 2136 22092
rect 2091 22052 2136 22080
rect 2130 22040 2136 22052
rect 2188 22040 2194 22092
rect 4080 22080 4108 22188
rect 4525 22185 4537 22219
rect 4571 22216 4583 22219
rect 4706 22216 4712 22228
rect 4571 22188 4712 22216
rect 4571 22185 4583 22188
rect 4525 22179 4583 22185
rect 4706 22176 4712 22188
rect 4764 22176 4770 22228
rect 4893 22219 4951 22225
rect 4893 22185 4905 22219
rect 4939 22216 4951 22219
rect 4982 22216 4988 22228
rect 4939 22188 4988 22216
rect 4939 22185 4951 22188
rect 4893 22179 4951 22185
rect 4982 22176 4988 22188
rect 5040 22176 5046 22228
rect 5905 22219 5963 22225
rect 5905 22185 5917 22219
rect 5951 22216 5963 22219
rect 6178 22216 6184 22228
rect 5951 22188 6184 22216
rect 5951 22185 5963 22188
rect 5905 22179 5963 22185
rect 6178 22176 6184 22188
rect 6236 22176 6242 22228
rect 6454 22216 6460 22228
rect 6415 22188 6460 22216
rect 6454 22176 6460 22188
rect 6512 22176 6518 22228
rect 8478 22216 8484 22228
rect 8439 22188 8484 22216
rect 8478 22176 8484 22188
rect 8536 22176 8542 22228
rect 14642 22176 14648 22228
rect 14700 22216 14706 22228
rect 14700 22188 15148 22216
rect 14700 22176 14706 22188
rect 6730 22108 6736 22160
rect 6788 22148 6794 22160
rect 7561 22151 7619 22157
rect 7561 22148 7573 22151
rect 6788 22120 7573 22148
rect 6788 22108 6794 22120
rect 7561 22117 7573 22120
rect 7607 22117 7619 22151
rect 7561 22111 7619 22117
rect 9674 22108 9680 22160
rect 9732 22148 9738 22160
rect 9732 22120 9777 22148
rect 9732 22108 9738 22120
rect 5353 22083 5411 22089
rect 4080 22052 5212 22080
rect 5074 21904 5080 21956
rect 5132 21944 5138 21956
rect 5184 21953 5212 22052
rect 5353 22049 5365 22083
rect 5399 22049 5411 22083
rect 5718 22080 5724 22092
rect 5679 22052 5724 22080
rect 5353 22043 5411 22049
rect 5368 22012 5396 22043
rect 5718 22040 5724 22052
rect 5776 22040 5782 22092
rect 7006 22080 7012 22092
rect 6967 22052 7012 22080
rect 7006 22040 7012 22052
rect 7064 22040 7070 22092
rect 7098 22040 7104 22092
rect 7156 22080 7162 22092
rect 7653 22083 7711 22089
rect 7653 22080 7665 22083
rect 7156 22052 7665 22080
rect 7156 22040 7162 22052
rect 7653 22049 7665 22052
rect 7699 22049 7711 22083
rect 7653 22043 7711 22049
rect 9585 22083 9643 22089
rect 9585 22049 9597 22083
rect 9631 22080 9643 22083
rect 9692 22080 9720 22108
rect 9631 22052 9720 22080
rect 9631 22049 9643 22052
rect 9585 22043 9643 22049
rect 9858 22040 9864 22092
rect 9916 22080 9922 22092
rect 10042 22080 10048 22092
rect 9916 22052 10048 22080
rect 9916 22040 9922 22052
rect 10042 22040 10048 22052
rect 10100 22080 10106 22092
rect 10505 22083 10563 22089
rect 10505 22080 10517 22083
rect 10100 22052 10517 22080
rect 10100 22040 10106 22052
rect 10505 22049 10517 22052
rect 10551 22080 10563 22083
rect 10962 22080 10968 22092
rect 10551 22052 10968 22080
rect 10551 22049 10563 22052
rect 10505 22043 10563 22049
rect 10962 22040 10968 22052
rect 11020 22040 11026 22092
rect 12710 22040 12716 22092
rect 12768 22080 12774 22092
rect 12897 22083 12955 22089
rect 12897 22080 12909 22083
rect 12768 22052 12909 22080
rect 12768 22040 12774 22052
rect 12897 22049 12909 22052
rect 12943 22049 12955 22083
rect 12897 22043 12955 22049
rect 14645 22083 14703 22089
rect 14645 22049 14657 22083
rect 14691 22049 14703 22083
rect 15010 22080 15016 22092
rect 14971 22052 15016 22080
rect 14645 22043 14703 22049
rect 6362 22012 6368 22024
rect 5368 21984 6368 22012
rect 6362 21972 6368 21984
rect 6420 21972 6426 22024
rect 8110 22012 8116 22024
rect 8071 21984 8116 22012
rect 8110 21972 8116 21984
rect 8168 21972 8174 22024
rect 8570 21972 8576 22024
rect 8628 22012 8634 22024
rect 10226 22012 10232 22024
rect 8628 21984 10232 22012
rect 8628 21972 8634 21984
rect 10226 21972 10232 21984
rect 10284 21972 10290 22024
rect 10686 22012 10692 22024
rect 10647 21984 10692 22012
rect 10686 21972 10692 21984
rect 10744 22012 10750 22024
rect 11514 22012 11520 22024
rect 10744 21984 11520 22012
rect 10744 21972 10750 21984
rect 11514 21972 11520 21984
rect 11572 21972 11578 22024
rect 14660 22012 14688 22043
rect 15010 22040 15016 22052
rect 15068 22040 15074 22092
rect 15120 22089 15148 22188
rect 15654 22108 15660 22160
rect 15712 22148 15718 22160
rect 15712 22120 16344 22148
rect 15712 22108 15718 22120
rect 15105 22083 15163 22089
rect 15105 22049 15117 22083
rect 15151 22049 15163 22083
rect 15105 22043 15163 22049
rect 15565 22083 15623 22089
rect 15565 22049 15577 22083
rect 15611 22080 15623 22083
rect 16206 22080 16212 22092
rect 15611 22052 16212 22080
rect 15611 22049 15623 22052
rect 15565 22043 15623 22049
rect 16206 22040 16212 22052
rect 16264 22040 16270 22092
rect 16316 22080 16344 22120
rect 16577 22083 16635 22089
rect 16577 22080 16589 22083
rect 16316 22052 16589 22080
rect 16577 22049 16589 22052
rect 16623 22080 16635 22083
rect 16666 22080 16672 22092
rect 16623 22052 16672 22080
rect 16623 22049 16635 22052
rect 16577 22043 16635 22049
rect 16666 22040 16672 22052
rect 16724 22040 16730 22092
rect 16850 22080 16856 22092
rect 16811 22052 16856 22080
rect 16850 22040 16856 22052
rect 16908 22040 16914 22092
rect 14918 22012 14924 22024
rect 14660 21984 14924 22012
rect 14918 21972 14924 21984
rect 14976 21972 14982 22024
rect 15654 21972 15660 22024
rect 15712 22012 15718 22024
rect 16117 22015 16175 22021
rect 16117 22012 16129 22015
rect 15712 21984 16129 22012
rect 15712 21972 15718 21984
rect 16117 21981 16129 21984
rect 16163 22012 16175 22015
rect 16758 22012 16764 22024
rect 16163 21984 16764 22012
rect 16163 21981 16175 21984
rect 16117 21975 16175 21981
rect 16758 21972 16764 21984
rect 16816 22012 16822 22024
rect 17405 22015 17463 22021
rect 17405 22012 17417 22015
rect 16816 21984 17417 22012
rect 16816 21972 16822 21984
rect 17405 21981 17417 21984
rect 17451 21981 17463 22015
rect 17405 21975 17463 21981
rect 5169 21947 5227 21953
rect 5169 21944 5181 21947
rect 5132 21916 5181 21944
rect 5132 21904 5138 21916
rect 5169 21913 5181 21916
rect 5215 21913 5227 21947
rect 5169 21907 5227 21913
rect 13081 21947 13139 21953
rect 13081 21913 13093 21947
rect 13127 21944 13139 21947
rect 13630 21944 13636 21956
rect 13127 21916 13636 21944
rect 13127 21913 13139 21916
rect 13081 21907 13139 21913
rect 13630 21904 13636 21916
rect 13688 21904 13694 21956
rect 14461 21947 14519 21953
rect 14461 21913 14473 21947
rect 14507 21944 14519 21947
rect 15378 21944 15384 21956
rect 14507 21916 15384 21944
rect 14507 21913 14519 21916
rect 14461 21907 14519 21913
rect 15378 21904 15384 21916
rect 15436 21904 15442 21956
rect 16482 21904 16488 21956
rect 16540 21944 16546 21956
rect 16853 21947 16911 21953
rect 16853 21944 16865 21947
rect 16540 21916 16865 21944
rect 16540 21904 16546 21916
rect 16853 21913 16865 21916
rect 16899 21913 16911 21947
rect 16853 21907 16911 21913
rect 3418 21876 3424 21888
rect 3379 21848 3424 21876
rect 3418 21836 3424 21848
rect 3476 21836 3482 21888
rect 7374 21876 7380 21888
rect 7335 21848 7380 21876
rect 7374 21836 7380 21848
rect 7432 21836 7438 21888
rect 13446 21876 13452 21888
rect 13407 21848 13452 21876
rect 13446 21836 13452 21848
rect 13504 21836 13510 21888
rect 13906 21876 13912 21888
rect 13867 21848 13912 21876
rect 13906 21836 13912 21848
rect 13964 21836 13970 21888
rect 15562 21836 15568 21888
rect 15620 21876 15626 21888
rect 15933 21879 15991 21885
rect 15933 21876 15945 21879
rect 15620 21848 15945 21876
rect 15620 21836 15626 21848
rect 15933 21845 15945 21848
rect 15979 21876 15991 21879
rect 16574 21876 16580 21888
rect 15979 21848 16580 21876
rect 15979 21845 15991 21848
rect 15933 21839 15991 21845
rect 16574 21836 16580 21848
rect 16632 21836 16638 21888
rect 1104 21786 18860 21808
rect 1104 21734 4315 21786
rect 4367 21734 4379 21786
rect 4431 21734 4443 21786
rect 4495 21734 4507 21786
rect 4559 21734 10982 21786
rect 11034 21734 11046 21786
rect 11098 21734 11110 21786
rect 11162 21734 11174 21786
rect 11226 21734 17648 21786
rect 17700 21734 17712 21786
rect 17764 21734 17776 21786
rect 17828 21734 17840 21786
rect 17892 21734 18860 21786
rect 1104 21712 18860 21734
rect 1949 21675 2007 21681
rect 1949 21641 1961 21675
rect 1995 21672 2007 21675
rect 2130 21672 2136 21684
rect 1995 21644 2136 21672
rect 1995 21641 2007 21644
rect 1949 21635 2007 21641
rect 2130 21632 2136 21644
rect 2188 21632 2194 21684
rect 7374 21632 7380 21684
rect 7432 21672 7438 21684
rect 8021 21675 8079 21681
rect 8021 21672 8033 21675
rect 7432 21644 8033 21672
rect 7432 21632 7438 21644
rect 8021 21641 8033 21644
rect 8067 21641 8079 21675
rect 8021 21635 8079 21641
rect 8294 21632 8300 21684
rect 8352 21672 8358 21684
rect 8389 21675 8447 21681
rect 8389 21672 8401 21675
rect 8352 21644 8401 21672
rect 8352 21632 8358 21644
rect 8389 21641 8401 21644
rect 8435 21641 8447 21675
rect 8389 21635 8447 21641
rect 9953 21675 10011 21681
rect 9953 21641 9965 21675
rect 9999 21672 10011 21675
rect 10042 21672 10048 21684
rect 9999 21644 10048 21672
rect 9999 21641 10011 21644
rect 9953 21635 10011 21641
rect 10042 21632 10048 21644
rect 10100 21632 10106 21684
rect 10226 21672 10232 21684
rect 10187 21644 10232 21672
rect 10226 21632 10232 21644
rect 10284 21632 10290 21684
rect 12161 21675 12219 21681
rect 12161 21641 12173 21675
rect 12207 21672 12219 21675
rect 12342 21672 12348 21684
rect 12207 21644 12348 21672
rect 12207 21641 12219 21644
rect 12161 21635 12219 21641
rect 1854 21564 1860 21616
rect 1912 21604 1918 21616
rect 2225 21607 2283 21613
rect 2225 21604 2237 21607
rect 1912 21576 2237 21604
rect 1912 21564 1918 21576
rect 2225 21573 2237 21576
rect 2271 21573 2283 21607
rect 2225 21567 2283 21573
rect 9493 21607 9551 21613
rect 9493 21573 9505 21607
rect 9539 21604 9551 21607
rect 10686 21604 10692 21616
rect 9539 21576 10692 21604
rect 9539 21573 9551 21576
rect 9493 21567 9551 21573
rect 10686 21564 10692 21576
rect 10744 21564 10750 21616
rect 5534 21496 5540 21548
rect 5592 21536 5598 21548
rect 6638 21536 6644 21548
rect 5592 21508 6644 21536
rect 5592 21496 5598 21508
rect 6638 21496 6644 21508
rect 6696 21496 6702 21548
rect 4893 21471 4951 21477
rect 4893 21437 4905 21471
rect 4939 21468 4951 21471
rect 5261 21471 5319 21477
rect 5261 21468 5273 21471
rect 4939 21440 5273 21468
rect 4939 21437 4951 21440
rect 4893 21431 4951 21437
rect 5261 21437 5273 21440
rect 5307 21468 5319 21471
rect 6362 21468 6368 21480
rect 5307 21440 6368 21468
rect 5307 21437 5319 21440
rect 5261 21431 5319 21437
rect 6362 21428 6368 21440
rect 6420 21468 6426 21480
rect 6549 21471 6607 21477
rect 6549 21468 6561 21471
rect 6420 21440 6561 21468
rect 6420 21428 6426 21440
rect 6549 21437 6561 21440
rect 6595 21437 6607 21471
rect 7282 21468 7288 21480
rect 7243 21440 7288 21468
rect 6549 21431 6607 21437
rect 7282 21428 7288 21440
rect 7340 21428 7346 21480
rect 8202 21468 8208 21480
rect 8163 21440 8208 21468
rect 8202 21428 8208 21440
rect 8260 21468 8266 21480
rect 8665 21471 8723 21477
rect 8665 21468 8677 21471
rect 8260 21440 8677 21468
rect 8260 21428 8266 21440
rect 8665 21437 8677 21440
rect 8711 21437 8723 21471
rect 8665 21431 8723 21437
rect 11609 21471 11667 21477
rect 11609 21437 11621 21471
rect 11655 21468 11667 21471
rect 12176 21468 12204 21635
rect 12342 21632 12348 21644
rect 12400 21632 12406 21684
rect 12526 21672 12532 21684
rect 12439 21644 12532 21672
rect 12526 21632 12532 21644
rect 12584 21672 12590 21684
rect 15010 21672 15016 21684
rect 12584 21644 15016 21672
rect 12584 21632 12590 21644
rect 15010 21632 15016 21644
rect 15068 21632 15074 21684
rect 15654 21672 15660 21684
rect 15615 21644 15660 21672
rect 15654 21632 15660 21644
rect 15712 21632 15718 21684
rect 13725 21607 13783 21613
rect 13725 21573 13737 21607
rect 13771 21604 13783 21607
rect 14182 21604 14188 21616
rect 13771 21576 14188 21604
rect 13771 21573 13783 21576
rect 13725 21567 13783 21573
rect 14182 21564 14188 21576
rect 14240 21604 14246 21616
rect 15286 21604 15292 21616
rect 14240 21576 15292 21604
rect 14240 21564 14246 21576
rect 15286 21564 15292 21576
rect 15344 21564 15350 21616
rect 15933 21607 15991 21613
rect 15933 21573 15945 21607
rect 15979 21604 15991 21607
rect 17034 21604 17040 21616
rect 15979 21576 17040 21604
rect 15979 21573 15991 21576
rect 15933 21567 15991 21573
rect 17034 21564 17040 21576
rect 17092 21564 17098 21616
rect 14366 21536 14372 21548
rect 14327 21508 14372 21536
rect 14366 21496 14372 21508
rect 14424 21496 14430 21548
rect 14642 21536 14648 21548
rect 14603 21508 14648 21536
rect 14642 21496 14648 21508
rect 14700 21536 14706 21548
rect 15010 21536 15016 21548
rect 14700 21508 15016 21536
rect 14700 21496 14706 21508
rect 15010 21496 15016 21508
rect 15068 21496 15074 21548
rect 17218 21496 17224 21548
rect 17276 21536 17282 21548
rect 18049 21539 18107 21545
rect 18049 21536 18061 21539
rect 17276 21508 18061 21536
rect 17276 21496 17282 21508
rect 11655 21440 12204 21468
rect 12621 21471 12679 21477
rect 11655 21437 11667 21440
rect 11609 21431 11667 21437
rect 12621 21437 12633 21471
rect 12667 21468 12679 21471
rect 12897 21471 12955 21477
rect 12897 21468 12909 21471
rect 12667 21440 12909 21468
rect 12667 21437 12679 21440
rect 12621 21431 12679 21437
rect 12897 21437 12909 21440
rect 12943 21437 12955 21471
rect 12897 21431 12955 21437
rect 13633 21471 13691 21477
rect 13633 21437 13645 21471
rect 13679 21437 13691 21471
rect 13633 21431 13691 21437
rect 5718 21360 5724 21412
rect 5776 21400 5782 21412
rect 5813 21403 5871 21409
rect 5813 21400 5825 21403
rect 5776 21372 5825 21400
rect 5776 21360 5782 21372
rect 5813 21369 5825 21372
rect 5859 21400 5871 21403
rect 6822 21400 6828 21412
rect 5859 21372 6828 21400
rect 5859 21369 5871 21372
rect 5813 21363 5871 21369
rect 6822 21360 6828 21372
rect 6880 21360 6886 21412
rect 12526 21360 12532 21412
rect 12584 21400 12590 21412
rect 12710 21400 12716 21412
rect 12584 21372 12716 21400
rect 12584 21360 12590 21372
rect 12710 21360 12716 21372
rect 12768 21400 12774 21412
rect 13081 21403 13139 21409
rect 13081 21400 13093 21403
rect 12768 21372 13093 21400
rect 12768 21360 12774 21372
rect 13081 21369 13093 21372
rect 13127 21369 13139 21403
rect 13081 21363 13139 21369
rect 13170 21360 13176 21412
rect 13228 21400 13234 21412
rect 13648 21400 13676 21431
rect 13814 21428 13820 21480
rect 13872 21468 13878 21480
rect 13909 21471 13967 21477
rect 13909 21468 13921 21471
rect 13872 21440 13921 21468
rect 13872 21428 13878 21440
rect 13909 21437 13921 21440
rect 13955 21437 13967 21471
rect 13909 21431 13967 21437
rect 14734 21428 14740 21480
rect 14792 21468 14798 21480
rect 17604 21477 17632 21508
rect 18049 21505 18061 21508
rect 18095 21505 18107 21539
rect 18049 21499 18107 21505
rect 15749 21471 15807 21477
rect 15749 21468 15761 21471
rect 14792 21440 15761 21468
rect 14792 21428 14798 21440
rect 15749 21437 15761 21440
rect 15795 21468 15807 21471
rect 16209 21471 16267 21477
rect 16209 21468 16221 21471
rect 15795 21440 16221 21468
rect 15795 21437 15807 21440
rect 15749 21431 15807 21437
rect 16209 21437 16221 21440
rect 16255 21437 16267 21471
rect 17313 21471 17371 21477
rect 17313 21468 17325 21471
rect 16209 21431 16267 21437
rect 16592 21440 17325 21468
rect 15562 21400 15568 21412
rect 13228 21372 15568 21400
rect 13228 21360 13234 21372
rect 15562 21360 15568 21372
rect 15620 21360 15626 21412
rect 16592 21344 16620 21440
rect 17313 21437 17325 21440
rect 17359 21437 17371 21471
rect 17313 21431 17371 21437
rect 17589 21471 17647 21477
rect 17589 21437 17601 21471
rect 17635 21437 17647 21471
rect 17589 21431 17647 21437
rect 17773 21471 17831 21477
rect 17773 21437 17785 21471
rect 17819 21437 17831 21471
rect 17773 21431 17831 21437
rect 16758 21400 16764 21412
rect 16719 21372 16764 21400
rect 16758 21360 16764 21372
rect 16816 21360 16822 21412
rect 17034 21360 17040 21412
rect 17092 21400 17098 21412
rect 17218 21400 17224 21412
rect 17092 21372 17224 21400
rect 17092 21360 17098 21372
rect 17218 21360 17224 21372
rect 17276 21400 17282 21412
rect 17788 21400 17816 21431
rect 17276 21372 17816 21400
rect 17276 21360 17282 21372
rect 6178 21332 6184 21344
rect 6139 21304 6184 21332
rect 6178 21292 6184 21304
rect 6236 21292 6242 21344
rect 6362 21332 6368 21344
rect 6323 21304 6368 21332
rect 6362 21292 6368 21304
rect 6420 21292 6426 21344
rect 7098 21292 7104 21344
rect 7156 21332 7162 21344
rect 7745 21335 7803 21341
rect 7745 21332 7757 21335
rect 7156 21304 7757 21332
rect 7156 21292 7162 21304
rect 7745 21301 7757 21304
rect 7791 21332 7803 21335
rect 8754 21332 8760 21344
rect 7791 21304 8760 21332
rect 7791 21301 7803 21304
rect 7745 21295 7803 21301
rect 8754 21292 8760 21304
rect 8812 21292 8818 21344
rect 11793 21335 11851 21341
rect 11793 21301 11805 21335
rect 11839 21332 11851 21335
rect 12066 21332 12072 21344
rect 11839 21304 12072 21332
rect 11839 21301 11851 21304
rect 11793 21295 11851 21301
rect 12066 21292 12072 21304
rect 12124 21292 12130 21344
rect 12802 21332 12808 21344
rect 12763 21304 12808 21332
rect 12802 21292 12808 21304
rect 12860 21292 12866 21344
rect 12897 21335 12955 21341
rect 12897 21301 12909 21335
rect 12943 21332 12955 21335
rect 13541 21335 13599 21341
rect 13541 21332 13553 21335
rect 12943 21304 13553 21332
rect 12943 21301 12955 21304
rect 12897 21295 12955 21301
rect 13541 21301 13553 21304
rect 13587 21332 13599 21335
rect 13722 21332 13728 21344
rect 13587 21304 13728 21332
rect 13587 21301 13599 21304
rect 13541 21295 13599 21301
rect 13722 21292 13728 21304
rect 13780 21292 13786 21344
rect 14918 21292 14924 21344
rect 14976 21332 14982 21344
rect 15013 21335 15071 21341
rect 15013 21332 15025 21335
rect 14976 21304 15025 21332
rect 14976 21292 14982 21304
rect 15013 21301 15025 21304
rect 15059 21301 15071 21335
rect 16574 21332 16580 21344
rect 16535 21304 16580 21332
rect 15013 21295 15071 21301
rect 16574 21292 16580 21304
rect 16632 21292 16638 21344
rect 1104 21242 18860 21264
rect 1104 21190 7648 21242
rect 7700 21190 7712 21242
rect 7764 21190 7776 21242
rect 7828 21190 7840 21242
rect 7892 21190 14315 21242
rect 14367 21190 14379 21242
rect 14431 21190 14443 21242
rect 14495 21190 14507 21242
rect 14559 21190 18860 21242
rect 1104 21168 18860 21190
rect 1394 21088 1400 21140
rect 1452 21128 1458 21140
rect 3881 21131 3939 21137
rect 3881 21128 3893 21131
rect 1452 21100 3893 21128
rect 1452 21088 1458 21100
rect 3881 21097 3893 21100
rect 3927 21097 3939 21131
rect 3881 21091 3939 21097
rect 6178 21088 6184 21140
rect 6236 21128 6242 21140
rect 6273 21131 6331 21137
rect 6273 21128 6285 21131
rect 6236 21100 6285 21128
rect 6236 21088 6242 21100
rect 6273 21097 6285 21100
rect 6319 21128 6331 21131
rect 6730 21128 6736 21140
rect 6319 21100 6736 21128
rect 6319 21097 6331 21100
rect 6273 21091 6331 21097
rect 6730 21088 6736 21100
rect 6788 21128 6794 21140
rect 7282 21128 7288 21140
rect 6788 21100 7288 21128
rect 6788 21088 6794 21100
rect 7282 21088 7288 21100
rect 7340 21128 7346 21140
rect 8205 21131 8263 21137
rect 8205 21128 8217 21131
rect 7340 21100 8217 21128
rect 7340 21088 7346 21100
rect 8205 21097 8217 21100
rect 8251 21097 8263 21131
rect 8205 21091 8263 21097
rect 12434 21088 12440 21140
rect 12492 21128 12498 21140
rect 12710 21128 12716 21140
rect 12492 21100 12716 21128
rect 12492 21088 12498 21100
rect 12710 21088 12716 21100
rect 12768 21088 12774 21140
rect 13170 21128 13176 21140
rect 13131 21100 13176 21128
rect 13170 21088 13176 21100
rect 13228 21088 13234 21140
rect 13814 21128 13820 21140
rect 13775 21100 13820 21128
rect 13814 21088 13820 21100
rect 13872 21088 13878 21140
rect 14182 21128 14188 21140
rect 14143 21100 14188 21128
rect 14182 21088 14188 21100
rect 14240 21088 14246 21140
rect 16666 21088 16672 21140
rect 16724 21128 16730 21140
rect 17773 21131 17831 21137
rect 17773 21128 17785 21131
rect 16724 21100 17785 21128
rect 16724 21088 16730 21100
rect 17773 21097 17785 21100
rect 17819 21097 17831 21131
rect 17773 21091 17831 21097
rect 5902 21060 5908 21072
rect 5863 21032 5908 21060
rect 5902 21020 5908 21032
rect 5960 21020 5966 21072
rect 6638 21060 6644 21072
rect 6599 21032 6644 21060
rect 6638 21020 6644 21032
rect 6696 21060 6702 21072
rect 6696 21032 7696 21060
rect 6696 21020 6702 21032
rect 1394 20992 1400 21004
rect 1355 20964 1400 20992
rect 1394 20952 1400 20964
rect 1452 20952 1458 21004
rect 1670 20992 1676 21004
rect 1631 20964 1676 20992
rect 1670 20952 1676 20964
rect 1728 20952 1734 21004
rect 3789 20995 3847 21001
rect 3789 20961 3801 20995
rect 3835 20992 3847 20995
rect 3878 20992 3884 21004
rect 3835 20964 3884 20992
rect 3835 20961 3847 20964
rect 3789 20955 3847 20961
rect 3878 20952 3884 20964
rect 3936 20992 3942 21004
rect 4065 20995 4123 21001
rect 4065 20992 4077 20995
rect 3936 20964 4077 20992
rect 3936 20952 3942 20964
rect 4065 20961 4077 20964
rect 4111 20992 4123 20995
rect 4798 20992 4804 21004
rect 4111 20964 4804 20992
rect 4111 20961 4123 20964
rect 4065 20955 4123 20961
rect 4798 20952 4804 20964
rect 4856 20952 4862 21004
rect 5810 20992 5816 21004
rect 5771 20964 5816 20992
rect 5810 20952 5816 20964
rect 5868 20952 5874 21004
rect 7098 20992 7104 21004
rect 7059 20964 7104 20992
rect 7098 20952 7104 20964
rect 7156 20952 7162 21004
rect 7466 20992 7472 21004
rect 7427 20964 7472 20992
rect 7466 20952 7472 20964
rect 7524 20952 7530 21004
rect 7668 21001 7696 21032
rect 8570 21020 8576 21072
rect 8628 21060 8634 21072
rect 8757 21063 8815 21069
rect 8757 21060 8769 21063
rect 8628 21032 8769 21060
rect 8628 21020 8634 21032
rect 8757 21029 8769 21032
rect 8803 21029 8815 21063
rect 8757 21023 8815 21029
rect 15197 21063 15255 21069
rect 15197 21029 15209 21063
rect 15243 21060 15255 21063
rect 15562 21060 15568 21072
rect 15243 21032 15568 21060
rect 15243 21029 15255 21032
rect 15197 21023 15255 21029
rect 15562 21020 15568 21032
rect 15620 21020 15626 21072
rect 15933 21063 15991 21069
rect 15933 21029 15945 21063
rect 15979 21060 15991 21063
rect 16758 21060 16764 21072
rect 15979 21032 16764 21060
rect 15979 21029 15991 21032
rect 15933 21023 15991 21029
rect 16758 21020 16764 21032
rect 16816 21060 16822 21072
rect 17126 21060 17132 21072
rect 16816 21032 16896 21060
rect 17087 21032 17132 21060
rect 16816 21020 16822 21032
rect 7653 20995 7711 21001
rect 7653 20961 7665 20995
rect 7699 20961 7711 20995
rect 7653 20955 7711 20961
rect 7929 20995 7987 21001
rect 7929 20961 7941 20995
rect 7975 20992 7987 20995
rect 8849 20995 8907 21001
rect 8849 20992 8861 20995
rect 7975 20964 8861 20992
rect 7975 20961 7987 20964
rect 7929 20955 7987 20961
rect 8849 20961 8861 20964
rect 8895 20992 8907 20995
rect 9030 20992 9036 21004
rect 8895 20964 9036 20992
rect 8895 20961 8907 20964
rect 8849 20955 8907 20961
rect 9030 20952 9036 20964
rect 9088 20952 9094 21004
rect 13265 20995 13323 21001
rect 13265 20961 13277 20995
rect 13311 20992 13323 20995
rect 13354 20992 13360 21004
rect 13311 20964 13360 20992
rect 13311 20961 13323 20964
rect 13265 20955 13323 20961
rect 13354 20952 13360 20964
rect 13412 20952 13418 21004
rect 15102 20992 15108 21004
rect 15063 20964 15108 20992
rect 15102 20952 15108 20964
rect 15160 20952 15166 21004
rect 15654 20952 15660 21004
rect 15712 20992 15718 21004
rect 16022 20992 16028 21004
rect 15712 20964 16028 20992
rect 15712 20952 15718 20964
rect 16022 20952 16028 20964
rect 16080 20952 16086 21004
rect 16298 20952 16304 21004
rect 16356 20992 16362 21004
rect 16868 21001 16896 21032
rect 17126 21020 17132 21032
rect 17184 21020 17190 21072
rect 16393 20995 16451 21001
rect 16393 20992 16405 20995
rect 16356 20964 16405 20992
rect 16356 20952 16362 20964
rect 16393 20961 16405 20964
rect 16439 20961 16451 20995
rect 16393 20955 16451 20961
rect 16853 20995 16911 21001
rect 16853 20961 16865 20995
rect 16899 20992 16911 20995
rect 17494 20992 17500 21004
rect 16899 20964 17500 20992
rect 16899 20961 16911 20964
rect 16853 20955 16911 20961
rect 17494 20952 17500 20964
rect 17552 20952 17558 21004
rect 2958 20788 2964 20800
rect 2919 20760 2964 20788
rect 2958 20748 2964 20760
rect 3016 20748 3022 20800
rect 4154 20748 4160 20800
rect 4212 20788 4218 20800
rect 4341 20791 4399 20797
rect 4341 20788 4353 20791
rect 4212 20760 4353 20788
rect 4212 20748 4218 20760
rect 4341 20757 4353 20760
rect 4387 20757 4399 20791
rect 4341 20751 4399 20757
rect 12434 20748 12440 20800
rect 12492 20788 12498 20800
rect 12621 20791 12679 20797
rect 12621 20788 12633 20791
rect 12492 20760 12633 20788
rect 12492 20748 12498 20760
rect 12621 20757 12633 20760
rect 12667 20757 12679 20791
rect 12621 20751 12679 20757
rect 13170 20748 13176 20800
rect 13228 20788 13234 20800
rect 13449 20791 13507 20797
rect 13449 20788 13461 20791
rect 13228 20760 13461 20788
rect 13228 20748 13234 20760
rect 13449 20757 13461 20760
rect 13495 20788 13507 20791
rect 13722 20788 13728 20800
rect 13495 20760 13728 20788
rect 13495 20757 13507 20760
rect 13449 20751 13507 20757
rect 13722 20748 13728 20760
rect 13780 20748 13786 20800
rect 15565 20791 15623 20797
rect 15565 20757 15577 20791
rect 15611 20788 15623 20791
rect 16758 20788 16764 20800
rect 15611 20760 16764 20788
rect 15611 20757 15623 20760
rect 15565 20751 15623 20757
rect 16758 20748 16764 20760
rect 16816 20748 16822 20800
rect 17218 20748 17224 20800
rect 17276 20788 17282 20800
rect 17405 20791 17463 20797
rect 17405 20788 17417 20791
rect 17276 20760 17417 20788
rect 17276 20748 17282 20760
rect 17405 20757 17417 20760
rect 17451 20757 17463 20791
rect 17405 20751 17463 20757
rect 1104 20698 18860 20720
rect 1104 20646 4315 20698
rect 4367 20646 4379 20698
rect 4431 20646 4443 20698
rect 4495 20646 4507 20698
rect 4559 20646 10982 20698
rect 11034 20646 11046 20698
rect 11098 20646 11110 20698
rect 11162 20646 11174 20698
rect 11226 20646 17648 20698
rect 17700 20646 17712 20698
rect 17764 20646 17776 20698
rect 17828 20646 17840 20698
rect 17892 20646 18860 20698
rect 1104 20624 18860 20646
rect 1670 20584 1676 20596
rect 1631 20556 1676 20584
rect 1670 20544 1676 20556
rect 1728 20544 1734 20596
rect 3602 20584 3608 20596
rect 3563 20556 3608 20584
rect 3602 20544 3608 20556
rect 3660 20544 3666 20596
rect 6089 20587 6147 20593
rect 6089 20553 6101 20587
rect 6135 20584 6147 20587
rect 7098 20584 7104 20596
rect 6135 20556 7104 20584
rect 6135 20553 6147 20556
rect 6089 20547 6147 20553
rect 7098 20544 7104 20556
rect 7156 20544 7162 20596
rect 8754 20584 8760 20596
rect 8715 20556 8760 20584
rect 8754 20544 8760 20556
rect 8812 20544 8818 20596
rect 9030 20584 9036 20596
rect 8991 20556 9036 20584
rect 9030 20544 9036 20556
rect 9088 20544 9094 20596
rect 13354 20584 13360 20596
rect 13315 20556 13360 20584
rect 13354 20544 13360 20556
rect 13412 20544 13418 20596
rect 14737 20587 14795 20593
rect 14737 20553 14749 20587
rect 14783 20584 14795 20587
rect 14826 20584 14832 20596
rect 14783 20556 14832 20584
rect 14783 20553 14795 20556
rect 14737 20547 14795 20553
rect 1394 20476 1400 20528
rect 1452 20516 1458 20528
rect 1949 20519 2007 20525
rect 1949 20516 1961 20519
rect 1452 20488 1961 20516
rect 1452 20476 1458 20488
rect 1949 20485 1961 20488
rect 1995 20485 2007 20519
rect 1949 20479 2007 20485
rect 3620 20448 3648 20544
rect 6457 20519 6515 20525
rect 6457 20485 6469 20519
rect 6503 20516 6515 20519
rect 6638 20516 6644 20528
rect 6503 20488 6644 20516
rect 6503 20485 6515 20488
rect 6457 20479 6515 20485
rect 6638 20476 6644 20488
rect 6696 20516 6702 20528
rect 9398 20516 9404 20528
rect 6696 20488 7604 20516
rect 9359 20488 9404 20516
rect 6696 20476 6702 20488
rect 4341 20451 4399 20457
rect 4341 20448 4353 20451
rect 3620 20420 4353 20448
rect 4341 20417 4353 20420
rect 4387 20417 4399 20451
rect 7466 20448 7472 20460
rect 4341 20411 4399 20417
rect 6840 20420 7472 20448
rect 3237 20383 3295 20389
rect 3237 20349 3249 20383
rect 3283 20380 3295 20383
rect 3878 20380 3884 20392
rect 3283 20352 3884 20380
rect 3283 20349 3295 20352
rect 3237 20343 3295 20349
rect 3878 20340 3884 20352
rect 3936 20340 3942 20392
rect 4062 20380 4068 20392
rect 4023 20352 4068 20380
rect 4062 20340 4068 20352
rect 4120 20340 4126 20392
rect 6840 20389 6868 20420
rect 7466 20408 7472 20420
rect 7524 20408 7530 20460
rect 7576 20389 7604 20488
rect 9398 20476 9404 20488
rect 9456 20476 9462 20528
rect 7745 20451 7803 20457
rect 7745 20417 7757 20451
rect 7791 20448 7803 20451
rect 8202 20448 8208 20460
rect 7791 20420 8208 20448
rect 7791 20417 7803 20420
rect 7745 20411 7803 20417
rect 8202 20408 8208 20420
rect 8260 20408 8266 20460
rect 9416 20448 9444 20476
rect 10137 20451 10195 20457
rect 10137 20448 10149 20451
rect 9416 20420 10149 20448
rect 10137 20417 10149 20420
rect 10183 20417 10195 20451
rect 12342 20448 12348 20460
rect 12303 20420 12348 20448
rect 10137 20411 10195 20417
rect 12342 20408 12348 20420
rect 12400 20408 12406 20460
rect 6825 20383 6883 20389
rect 6825 20349 6837 20383
rect 6871 20349 6883 20383
rect 6825 20343 6883 20349
rect 7193 20383 7251 20389
rect 7193 20349 7205 20383
rect 7239 20349 7251 20383
rect 7193 20343 7251 20349
rect 7561 20383 7619 20389
rect 7561 20349 7573 20383
rect 7607 20349 7619 20383
rect 8573 20383 8631 20389
rect 8573 20380 8585 20383
rect 7561 20343 7619 20349
rect 8404 20352 8585 20380
rect 3694 20244 3700 20256
rect 3655 20216 3700 20244
rect 3694 20204 3700 20216
rect 3752 20204 3758 20256
rect 5442 20244 5448 20256
rect 5403 20216 5448 20244
rect 5442 20204 5448 20216
rect 5500 20204 5506 20256
rect 6914 20204 6920 20256
rect 6972 20244 6978 20256
rect 7208 20244 7236 20343
rect 8018 20244 8024 20256
rect 6972 20216 8024 20244
rect 6972 20204 6978 20216
rect 8018 20204 8024 20216
rect 8076 20244 8082 20256
rect 8404 20253 8432 20352
rect 8573 20349 8585 20352
rect 8619 20349 8631 20383
rect 9858 20380 9864 20392
rect 9819 20352 9864 20380
rect 8573 20343 8631 20349
rect 9858 20340 9864 20352
rect 9916 20340 9922 20392
rect 12253 20383 12311 20389
rect 12253 20349 12265 20383
rect 12299 20380 12311 20383
rect 12526 20380 12532 20392
rect 12299 20352 12532 20380
rect 12299 20349 12311 20352
rect 12253 20343 12311 20349
rect 12526 20340 12532 20352
rect 12584 20340 12590 20392
rect 12621 20383 12679 20389
rect 12621 20349 12633 20383
rect 12667 20380 12679 20383
rect 12986 20380 12992 20392
rect 12667 20352 12992 20380
rect 12667 20349 12679 20352
rect 12621 20343 12679 20349
rect 11882 20312 11888 20324
rect 11795 20284 11888 20312
rect 11882 20272 11888 20284
rect 11940 20312 11946 20324
rect 12636 20312 12664 20343
rect 12986 20340 12992 20352
rect 13044 20340 13050 20392
rect 14185 20383 14243 20389
rect 14185 20349 14197 20383
rect 14231 20380 14243 20383
rect 14752 20380 14780 20547
rect 14826 20544 14832 20556
rect 14884 20544 14890 20596
rect 15102 20584 15108 20596
rect 15063 20556 15108 20584
rect 15102 20544 15108 20556
rect 15160 20544 15166 20596
rect 15565 20587 15623 20593
rect 15565 20553 15577 20587
rect 15611 20584 15623 20587
rect 16022 20584 16028 20596
rect 15611 20556 16028 20584
rect 15611 20553 15623 20556
rect 15565 20547 15623 20553
rect 16022 20544 16028 20556
rect 16080 20584 16086 20596
rect 16485 20587 16543 20593
rect 16485 20584 16497 20587
rect 16080 20556 16497 20584
rect 16080 20544 16086 20556
rect 16485 20553 16497 20556
rect 16531 20553 16543 20587
rect 16485 20547 16543 20553
rect 16500 20448 16528 20547
rect 16574 20476 16580 20528
rect 16632 20516 16638 20528
rect 17497 20519 17555 20525
rect 17497 20516 17509 20519
rect 16632 20488 17509 20516
rect 16632 20476 16638 20488
rect 17497 20485 17509 20488
rect 17543 20485 17555 20519
rect 17497 20479 17555 20485
rect 16761 20451 16819 20457
rect 16761 20448 16773 20451
rect 16500 20420 16773 20448
rect 16761 20417 16773 20420
rect 16807 20417 16819 20451
rect 16761 20411 16819 20417
rect 14231 20352 14780 20380
rect 14231 20349 14243 20352
rect 14185 20343 14243 20349
rect 15194 20340 15200 20392
rect 15252 20380 15258 20392
rect 15657 20383 15715 20389
rect 15657 20380 15669 20383
rect 15252 20352 15669 20380
rect 15252 20340 15258 20352
rect 15657 20349 15669 20352
rect 15703 20380 15715 20383
rect 15838 20380 15844 20392
rect 15703 20352 15844 20380
rect 15703 20349 15715 20352
rect 15657 20343 15715 20349
rect 15838 20340 15844 20352
rect 15896 20380 15902 20392
rect 16117 20383 16175 20389
rect 16117 20380 16129 20383
rect 15896 20352 16129 20380
rect 15896 20340 15902 20352
rect 16117 20349 16129 20352
rect 16163 20349 16175 20383
rect 16117 20343 16175 20349
rect 17221 20383 17279 20389
rect 17221 20349 17233 20383
rect 17267 20380 17279 20383
rect 17402 20380 17408 20392
rect 17267 20352 17408 20380
rect 17267 20349 17279 20352
rect 17221 20343 17279 20349
rect 17402 20340 17408 20352
rect 17460 20340 17466 20392
rect 17494 20340 17500 20392
rect 17552 20380 17558 20392
rect 17552 20352 17597 20380
rect 17552 20340 17558 20352
rect 11940 20284 12664 20312
rect 12713 20315 12771 20321
rect 11940 20272 11946 20284
rect 12713 20281 12725 20315
rect 12759 20281 12771 20315
rect 13078 20312 13084 20324
rect 13039 20284 13084 20312
rect 12713 20275 12771 20281
rect 8389 20247 8447 20253
rect 8389 20244 8401 20247
rect 8076 20216 8401 20244
rect 8076 20204 8082 20216
rect 8389 20213 8401 20216
rect 8435 20213 8447 20247
rect 8389 20207 8447 20213
rect 11425 20247 11483 20253
rect 11425 20213 11437 20247
rect 11471 20244 11483 20247
rect 12158 20244 12164 20256
rect 11471 20216 12164 20244
rect 11471 20213 11483 20216
rect 11425 20207 11483 20213
rect 12158 20204 12164 20216
rect 12216 20204 12222 20256
rect 12728 20244 12756 20275
rect 13078 20272 13084 20284
rect 13136 20272 13142 20324
rect 13814 20244 13820 20256
rect 12728 20216 13820 20244
rect 13814 20204 13820 20216
rect 13872 20204 13878 20256
rect 14369 20247 14427 20253
rect 14369 20213 14381 20247
rect 14415 20244 14427 20247
rect 14918 20244 14924 20256
rect 14415 20216 14924 20244
rect 14415 20213 14427 20216
rect 14369 20207 14427 20213
rect 14918 20204 14924 20216
rect 14976 20204 14982 20256
rect 15562 20204 15568 20256
rect 15620 20244 15626 20256
rect 15841 20247 15899 20253
rect 15841 20244 15853 20247
rect 15620 20216 15853 20244
rect 15620 20204 15626 20216
rect 15841 20213 15853 20216
rect 15887 20213 15899 20247
rect 15841 20207 15899 20213
rect 1104 20154 18860 20176
rect 1104 20102 7648 20154
rect 7700 20102 7712 20154
rect 7764 20102 7776 20154
rect 7828 20102 7840 20154
rect 7892 20102 14315 20154
rect 14367 20102 14379 20154
rect 14431 20102 14443 20154
rect 14495 20102 14507 20154
rect 14559 20102 18860 20154
rect 1104 20080 18860 20102
rect 1394 20000 1400 20052
rect 1452 20040 1458 20052
rect 1581 20043 1639 20049
rect 1581 20040 1593 20043
rect 1452 20012 1593 20040
rect 1452 20000 1458 20012
rect 1581 20009 1593 20012
rect 1627 20009 1639 20043
rect 1581 20003 1639 20009
rect 5261 20043 5319 20049
rect 5261 20009 5273 20043
rect 5307 20040 5319 20043
rect 5810 20040 5816 20052
rect 5307 20012 5816 20040
rect 5307 20009 5319 20012
rect 5261 20003 5319 20009
rect 5810 20000 5816 20012
rect 5868 20040 5874 20052
rect 6365 20043 6423 20049
rect 6365 20040 6377 20043
rect 5868 20012 6377 20040
rect 5868 20000 5874 20012
rect 6365 20009 6377 20012
rect 6411 20040 6423 20043
rect 6546 20040 6552 20052
rect 6411 20012 6552 20040
rect 6411 20009 6423 20012
rect 6365 20003 6423 20009
rect 6546 20000 6552 20012
rect 6604 20040 6610 20052
rect 7466 20040 7472 20052
rect 6604 20012 7472 20040
rect 6604 20000 6610 20012
rect 7466 20000 7472 20012
rect 7524 20040 7530 20052
rect 7653 20043 7711 20049
rect 7653 20040 7665 20043
rect 7524 20012 7665 20040
rect 7524 20000 7530 20012
rect 7653 20009 7665 20012
rect 7699 20009 7711 20043
rect 12158 20040 12164 20052
rect 12119 20012 12164 20040
rect 7653 20003 7711 20009
rect 12158 20000 12164 20012
rect 12216 20000 12222 20052
rect 16298 20040 16304 20052
rect 16259 20012 16304 20040
rect 16298 20000 16304 20012
rect 16356 20000 16362 20052
rect 17402 20000 17408 20052
rect 17460 20040 17466 20052
rect 17497 20043 17555 20049
rect 17497 20040 17509 20043
rect 17460 20012 17509 20040
rect 17460 20000 17466 20012
rect 17497 20009 17509 20012
rect 17543 20009 17555 20043
rect 17497 20003 17555 20009
rect 12176 19972 12204 20000
rect 12176 19944 13492 19972
rect 3418 19904 3424 19916
rect 3379 19876 3424 19904
rect 3418 19864 3424 19876
rect 3476 19864 3482 19916
rect 6362 19864 6368 19916
rect 6420 19904 6426 19916
rect 6641 19907 6699 19913
rect 6641 19904 6653 19907
rect 6420 19876 6653 19904
rect 6420 19864 6426 19876
rect 6641 19873 6653 19876
rect 6687 19873 6699 19907
rect 6914 19904 6920 19916
rect 6875 19876 6920 19904
rect 6641 19867 6699 19873
rect 6914 19864 6920 19876
rect 6972 19864 6978 19916
rect 13365 19907 13423 19913
rect 13365 19873 13377 19907
rect 13411 19904 13423 19907
rect 13464 19904 13492 19944
rect 13411 19876 13492 19904
rect 13411 19873 13423 19876
rect 13365 19867 13423 19873
rect 15286 19864 15292 19916
rect 15344 19904 15350 19916
rect 15381 19907 15439 19913
rect 15381 19904 15393 19907
rect 15344 19876 15393 19904
rect 15344 19864 15350 19876
rect 15381 19873 15393 19876
rect 15427 19873 15439 19907
rect 15381 19867 15439 19873
rect 15749 19907 15807 19913
rect 15749 19873 15761 19907
rect 15795 19873 15807 19907
rect 15749 19867 15807 19873
rect 3145 19839 3203 19845
rect 3145 19805 3157 19839
rect 3191 19836 3203 19839
rect 3602 19836 3608 19848
rect 3191 19808 3608 19836
rect 3191 19805 3203 19808
rect 3145 19799 3203 19805
rect 3602 19796 3608 19808
rect 3660 19796 3666 19848
rect 6730 19796 6736 19848
rect 6788 19836 6794 19848
rect 6825 19839 6883 19845
rect 6825 19836 6837 19839
rect 6788 19808 6837 19836
rect 6788 19796 6794 19808
rect 6825 19805 6837 19808
rect 6871 19805 6883 19839
rect 6825 19799 6883 19805
rect 12529 19839 12587 19845
rect 12529 19805 12541 19839
rect 12575 19805 12587 19839
rect 12529 19799 12587 19805
rect 12544 19768 12572 19799
rect 12618 19796 12624 19848
rect 12676 19836 12682 19848
rect 12676 19808 12721 19836
rect 12676 19796 12682 19808
rect 12802 19796 12808 19848
rect 12860 19836 12866 19848
rect 13449 19839 13507 19845
rect 13449 19836 13461 19839
rect 12860 19808 13461 19836
rect 12860 19796 12866 19808
rect 13449 19805 13461 19808
rect 13495 19836 13507 19839
rect 13722 19836 13728 19848
rect 13495 19808 13728 19836
rect 13495 19805 13507 19808
rect 13449 19799 13507 19805
rect 13722 19796 13728 19808
rect 13780 19796 13786 19848
rect 15764 19836 15792 19867
rect 15838 19864 15844 19916
rect 15896 19904 15902 19916
rect 17221 19907 17279 19913
rect 15896 19876 15941 19904
rect 15896 19864 15902 19876
rect 17221 19873 17233 19907
rect 17267 19904 17279 19907
rect 17494 19904 17500 19916
rect 17267 19876 17500 19904
rect 17267 19873 17279 19876
rect 17221 19867 17279 19873
rect 17494 19864 17500 19876
rect 17552 19864 17558 19916
rect 14752 19808 15792 19836
rect 14752 19780 14780 19808
rect 12986 19768 12992 19780
rect 12544 19740 12992 19768
rect 12986 19728 12992 19740
rect 13044 19728 13050 19780
rect 14734 19768 14740 19780
rect 14695 19740 14740 19768
rect 14734 19728 14740 19740
rect 14792 19728 14798 19780
rect 15194 19768 15200 19780
rect 15155 19740 15200 19768
rect 15194 19728 15200 19740
rect 15252 19728 15258 19780
rect 4706 19700 4712 19712
rect 4667 19672 4712 19700
rect 4706 19660 4712 19672
rect 4764 19660 4770 19712
rect 6457 19703 6515 19709
rect 6457 19669 6469 19703
rect 6503 19700 6515 19703
rect 6822 19700 6828 19712
rect 6503 19672 6828 19700
rect 6503 19669 6515 19672
rect 6457 19663 6515 19669
rect 6822 19660 6828 19672
rect 6880 19660 6886 19712
rect 7006 19660 7012 19712
rect 7064 19700 7070 19712
rect 7101 19703 7159 19709
rect 7101 19700 7113 19703
rect 7064 19672 7113 19700
rect 7064 19660 7070 19672
rect 7101 19669 7113 19672
rect 7147 19669 7159 19703
rect 9858 19700 9864 19712
rect 9819 19672 9864 19700
rect 7101 19663 7159 19669
rect 9858 19660 9864 19672
rect 9916 19660 9922 19712
rect 13814 19700 13820 19712
rect 13775 19672 13820 19700
rect 13814 19660 13820 19672
rect 13872 19660 13878 19712
rect 14182 19700 14188 19712
rect 14143 19672 14188 19700
rect 14182 19660 14188 19672
rect 14240 19660 14246 19712
rect 16853 19703 16911 19709
rect 16853 19669 16865 19703
rect 16899 19700 16911 19703
rect 17218 19700 17224 19712
rect 16899 19672 17224 19700
rect 16899 19669 16911 19672
rect 16853 19663 16911 19669
rect 17218 19660 17224 19672
rect 17276 19700 17282 19712
rect 17494 19700 17500 19712
rect 17276 19672 17500 19700
rect 17276 19660 17282 19672
rect 17494 19660 17500 19672
rect 17552 19660 17558 19712
rect 1104 19610 18860 19632
rect 1104 19558 4315 19610
rect 4367 19558 4379 19610
rect 4431 19558 4443 19610
rect 4495 19558 4507 19610
rect 4559 19558 10982 19610
rect 11034 19558 11046 19610
rect 11098 19558 11110 19610
rect 11162 19558 11174 19610
rect 11226 19558 17648 19610
rect 17700 19558 17712 19610
rect 17764 19558 17776 19610
rect 17828 19558 17840 19610
rect 17892 19558 18860 19610
rect 1104 19536 18860 19558
rect 3418 19496 3424 19508
rect 3379 19468 3424 19496
rect 3418 19456 3424 19468
rect 3476 19456 3482 19508
rect 3694 19496 3700 19508
rect 3655 19468 3700 19496
rect 3694 19456 3700 19468
rect 3752 19456 3758 19508
rect 6546 19496 6552 19508
rect 6507 19468 6552 19496
rect 6546 19456 6552 19468
rect 6604 19456 6610 19508
rect 6730 19456 6736 19508
rect 6788 19496 6794 19508
rect 7101 19499 7159 19505
rect 7101 19496 7113 19499
rect 6788 19468 7113 19496
rect 6788 19456 6794 19468
rect 7101 19465 7113 19468
rect 7147 19465 7159 19499
rect 7101 19459 7159 19465
rect 12158 19456 12164 19508
rect 12216 19496 12222 19508
rect 13722 19496 13728 19508
rect 12216 19468 13584 19496
rect 13683 19468 13728 19496
rect 12216 19456 12222 19468
rect 12342 19388 12348 19440
rect 12400 19428 12406 19440
rect 12802 19428 12808 19440
rect 12400 19400 12808 19428
rect 12400 19388 12406 19400
rect 12802 19388 12808 19400
rect 12860 19388 12866 19440
rect 13170 19388 13176 19440
rect 13228 19428 13234 19440
rect 13556 19428 13584 19468
rect 13722 19456 13728 19468
rect 13780 19456 13786 19508
rect 13814 19428 13820 19440
rect 13228 19400 13492 19428
rect 13556 19400 13820 19428
rect 13228 19388 13234 19400
rect 1394 19360 1400 19372
rect 1355 19332 1400 19360
rect 1394 19320 1400 19332
rect 1452 19320 1458 19372
rect 12989 19363 13047 19369
rect 4908 19332 5304 19360
rect 1486 19252 1492 19304
rect 1544 19292 1550 19304
rect 1673 19295 1731 19301
rect 1673 19292 1685 19295
rect 1544 19264 1685 19292
rect 1544 19252 1550 19264
rect 1673 19261 1685 19264
rect 1719 19261 1731 19295
rect 1673 19255 1731 19261
rect 4801 19295 4859 19301
rect 4801 19261 4813 19295
rect 4847 19292 4859 19295
rect 4908 19292 4936 19332
rect 5074 19292 5080 19304
rect 4847 19264 4936 19292
rect 5035 19264 5080 19292
rect 4847 19261 4859 19264
rect 4801 19255 4859 19261
rect 5074 19252 5080 19264
rect 5132 19252 5138 19304
rect 5176 19295 5234 19301
rect 5176 19261 5188 19295
rect 5222 19261 5234 19295
rect 5276 19292 5304 19332
rect 12989 19329 13001 19363
rect 13035 19360 13047 19363
rect 13078 19360 13084 19372
rect 13035 19332 13084 19360
rect 13035 19329 13047 19332
rect 12989 19323 13047 19329
rect 13078 19320 13084 19332
rect 13136 19320 13142 19372
rect 13464 19360 13492 19400
rect 13814 19388 13820 19400
rect 13872 19388 13878 19440
rect 16298 19388 16304 19440
rect 16356 19428 16362 19440
rect 16577 19431 16635 19437
rect 16577 19428 16589 19431
rect 16356 19400 16589 19428
rect 16356 19388 16362 19400
rect 16577 19397 16589 19400
rect 16623 19428 16635 19431
rect 16623 19400 17448 19428
rect 16623 19397 16635 19400
rect 16577 19391 16635 19397
rect 13464 19332 15148 19360
rect 5442 19292 5448 19304
rect 5276 19264 5448 19292
rect 5176 19255 5234 19261
rect 3053 19227 3111 19233
rect 3053 19193 3065 19227
rect 3099 19224 3111 19227
rect 4062 19224 4068 19236
rect 3099 19196 4068 19224
rect 3099 19193 3111 19196
rect 3053 19187 3111 19193
rect 4062 19184 4068 19196
rect 4120 19184 4126 19236
rect 4154 19116 4160 19168
rect 4212 19156 4218 19168
rect 4893 19159 4951 19165
rect 4893 19156 4905 19159
rect 4212 19128 4905 19156
rect 4212 19116 4218 19128
rect 4893 19125 4905 19128
rect 4939 19156 4951 19159
rect 5184 19156 5212 19255
rect 5442 19252 5448 19264
rect 5500 19252 5506 19304
rect 6362 19252 6368 19304
rect 6420 19292 6426 19304
rect 7837 19295 7895 19301
rect 7837 19292 7849 19295
rect 6420 19264 7849 19292
rect 6420 19252 6426 19264
rect 7837 19261 7849 19264
rect 7883 19292 7895 19295
rect 8113 19295 8171 19301
rect 8113 19292 8125 19295
rect 7883 19264 8125 19292
rect 7883 19261 7895 19264
rect 7837 19255 7895 19261
rect 8113 19261 8125 19264
rect 8159 19261 8171 19295
rect 8113 19255 8171 19261
rect 10597 19295 10655 19301
rect 10597 19261 10609 19295
rect 10643 19292 10655 19295
rect 11333 19295 11391 19301
rect 11333 19292 11345 19295
rect 10643 19264 11345 19292
rect 10643 19261 10655 19264
rect 10597 19255 10655 19261
rect 11333 19261 11345 19264
rect 11379 19292 11391 19295
rect 12897 19295 12955 19301
rect 12897 19292 12909 19295
rect 11379 19264 12909 19292
rect 11379 19261 11391 19264
rect 11333 19255 11391 19261
rect 7561 19227 7619 19233
rect 7561 19193 7573 19227
rect 7607 19224 7619 19227
rect 8018 19224 8024 19236
rect 7607 19196 8024 19224
rect 7607 19193 7619 19196
rect 7561 19187 7619 19193
rect 8018 19184 8024 19196
rect 8076 19184 8082 19236
rect 11425 19227 11483 19233
rect 11425 19193 11437 19227
rect 11471 19224 11483 19227
rect 11606 19224 11612 19236
rect 11471 19196 11612 19224
rect 11471 19193 11483 19196
rect 11425 19187 11483 19193
rect 11606 19184 11612 19196
rect 11664 19184 11670 19236
rect 12176 19168 12204 19264
rect 12897 19261 12909 19264
rect 12943 19261 12955 19295
rect 12897 19255 12955 19261
rect 13170 19252 13176 19304
rect 13228 19292 13234 19304
rect 13265 19295 13323 19301
rect 13265 19292 13277 19295
rect 13228 19264 13277 19292
rect 13228 19252 13234 19264
rect 13265 19261 13277 19264
rect 13311 19261 13323 19295
rect 13265 19255 13323 19261
rect 13449 19295 13507 19301
rect 13449 19261 13461 19295
rect 13495 19292 13507 19295
rect 13538 19292 13544 19304
rect 13495 19264 13544 19292
rect 13495 19261 13507 19264
rect 13449 19255 13507 19261
rect 13538 19252 13544 19264
rect 13596 19252 13602 19304
rect 15010 19292 15016 19304
rect 14971 19264 15016 19292
rect 15010 19252 15016 19264
rect 15068 19252 15074 19304
rect 15120 19292 15148 19332
rect 15289 19295 15347 19301
rect 15289 19292 15301 19295
rect 15120 19264 15301 19292
rect 15289 19261 15301 19264
rect 15335 19292 15347 19295
rect 15838 19292 15844 19304
rect 15335 19264 15844 19292
rect 15335 19261 15347 19264
rect 15289 19255 15347 19261
rect 15838 19252 15844 19264
rect 15896 19252 15902 19304
rect 16301 19295 16359 19301
rect 16301 19261 16313 19295
rect 16347 19292 16359 19295
rect 17310 19292 17316 19304
rect 16347 19264 17316 19292
rect 16347 19261 16359 19264
rect 16301 19255 16359 19261
rect 17310 19252 17316 19264
rect 17368 19252 17374 19304
rect 17420 19292 17448 19400
rect 17494 19320 17500 19372
rect 17552 19360 17558 19372
rect 17773 19363 17831 19369
rect 17773 19360 17785 19363
rect 17552 19332 17785 19360
rect 17552 19320 17558 19332
rect 17773 19329 17785 19332
rect 17819 19329 17831 19363
rect 17773 19323 17831 19329
rect 17589 19295 17647 19301
rect 17589 19292 17601 19295
rect 17420 19264 17601 19292
rect 17589 19261 17601 19264
rect 17635 19261 17647 19295
rect 17589 19255 17647 19261
rect 12253 19227 12311 19233
rect 12253 19193 12265 19227
rect 12299 19224 12311 19227
rect 13354 19224 13360 19236
rect 12299 19196 13360 19224
rect 12299 19193 12311 19196
rect 12253 19187 12311 19193
rect 13354 19184 13360 19196
rect 13412 19184 13418 19236
rect 14185 19227 14243 19233
rect 14185 19193 14197 19227
rect 14231 19224 14243 19227
rect 14734 19224 14740 19236
rect 14231 19196 14740 19224
rect 14231 19193 14243 19196
rect 14185 19187 14243 19193
rect 14734 19184 14740 19196
rect 14792 19224 14798 19236
rect 16758 19224 16764 19236
rect 14792 19196 15516 19224
rect 16719 19196 16764 19224
rect 14792 19184 14798 19196
rect 5718 19156 5724 19168
rect 4939 19128 5724 19156
rect 4939 19125 4951 19128
rect 4893 19119 4951 19125
rect 5718 19116 5724 19128
rect 5776 19116 5782 19168
rect 7374 19116 7380 19168
rect 7432 19156 7438 19168
rect 7653 19159 7711 19165
rect 7653 19156 7665 19159
rect 7432 19128 7665 19156
rect 7432 19116 7438 19128
rect 7653 19125 7665 19128
rect 7699 19125 7711 19159
rect 11790 19156 11796 19168
rect 11751 19128 11796 19156
rect 7653 19119 7711 19125
rect 11790 19116 11796 19128
rect 11848 19116 11854 19168
rect 12158 19156 12164 19168
rect 12119 19128 12164 19156
rect 12158 19116 12164 19128
rect 12216 19116 12222 19168
rect 14645 19159 14703 19165
rect 14645 19125 14657 19159
rect 14691 19156 14703 19159
rect 15286 19156 15292 19168
rect 14691 19128 15292 19156
rect 14691 19125 14703 19128
rect 14645 19119 14703 19125
rect 15286 19116 15292 19128
rect 15344 19116 15350 19168
rect 15488 19165 15516 19196
rect 16758 19184 16764 19196
rect 16816 19184 16822 19236
rect 15473 19159 15531 19165
rect 15473 19125 15485 19159
rect 15519 19125 15531 19159
rect 15473 19119 15531 19125
rect 1104 19066 18860 19088
rect 1104 19014 7648 19066
rect 7700 19014 7712 19066
rect 7764 19014 7776 19066
rect 7828 19014 7840 19066
rect 7892 19014 14315 19066
rect 14367 19014 14379 19066
rect 14431 19014 14443 19066
rect 14495 19014 14507 19066
rect 14559 19014 18860 19066
rect 1104 18992 18860 19014
rect 1486 18912 1492 18964
rect 1544 18952 1550 18964
rect 1581 18955 1639 18961
rect 1581 18952 1593 18955
rect 1544 18924 1593 18952
rect 1544 18912 1550 18924
rect 1581 18921 1593 18924
rect 1627 18921 1639 18955
rect 1581 18915 1639 18921
rect 4985 18955 5043 18961
rect 4985 18921 4997 18955
rect 5031 18952 5043 18955
rect 5074 18952 5080 18964
rect 5031 18924 5080 18952
rect 5031 18921 5043 18924
rect 4985 18915 5043 18921
rect 5074 18912 5080 18924
rect 5132 18912 5138 18964
rect 6362 18912 6368 18964
rect 6420 18952 6426 18964
rect 6457 18955 6515 18961
rect 6457 18952 6469 18955
rect 6420 18924 6469 18952
rect 6420 18912 6426 18924
rect 6457 18921 6469 18924
rect 6503 18921 6515 18955
rect 6457 18915 6515 18921
rect 12434 18912 12440 18964
rect 12492 18952 12498 18964
rect 12621 18955 12679 18961
rect 12621 18952 12633 18955
rect 12492 18924 12633 18952
rect 12492 18912 12498 18924
rect 12621 18921 12633 18924
rect 12667 18921 12679 18955
rect 12621 18915 12679 18921
rect 12989 18955 13047 18961
rect 12989 18921 13001 18955
rect 13035 18952 13047 18955
rect 13078 18952 13084 18964
rect 13035 18924 13084 18952
rect 13035 18921 13047 18924
rect 12989 18915 13047 18921
rect 13078 18912 13084 18924
rect 13136 18912 13142 18964
rect 10778 18816 10784 18828
rect 10739 18788 10784 18816
rect 10778 18776 10784 18788
rect 10836 18776 10842 18828
rect 10870 18776 10876 18828
rect 10928 18816 10934 18828
rect 11330 18816 11336 18828
rect 10928 18788 11336 18816
rect 10928 18776 10934 18788
rect 11330 18776 11336 18788
rect 11388 18816 11394 18828
rect 11882 18816 11888 18828
rect 11388 18788 11888 18816
rect 11388 18776 11394 18788
rect 11882 18776 11888 18788
rect 11940 18776 11946 18828
rect 12437 18819 12495 18825
rect 12437 18785 12449 18819
rect 12483 18816 12495 18819
rect 12526 18816 12532 18828
rect 12483 18788 12532 18816
rect 12483 18785 12495 18788
rect 12437 18779 12495 18785
rect 12526 18776 12532 18788
rect 12584 18776 12590 18828
rect 13998 18776 14004 18828
rect 14056 18816 14062 18828
rect 14185 18819 14243 18825
rect 14185 18816 14197 18819
rect 14056 18788 14197 18816
rect 14056 18776 14062 18788
rect 14185 18785 14197 18788
rect 14231 18785 14243 18819
rect 14185 18779 14243 18785
rect 14274 18776 14280 18828
rect 14332 18816 14338 18828
rect 14553 18819 14611 18825
rect 14553 18816 14565 18819
rect 14332 18788 14565 18816
rect 14332 18776 14338 18788
rect 14553 18785 14565 18788
rect 14599 18785 14611 18819
rect 14553 18779 14611 18785
rect 14918 18776 14924 18828
rect 14976 18816 14982 18828
rect 15746 18816 15752 18828
rect 14976 18788 15752 18816
rect 14976 18776 14982 18788
rect 15746 18776 15752 18788
rect 15804 18816 15810 18828
rect 16025 18819 16083 18825
rect 16025 18816 16037 18819
rect 15804 18788 16037 18816
rect 15804 18776 15810 18788
rect 16025 18785 16037 18788
rect 16071 18785 16083 18819
rect 16482 18816 16488 18828
rect 16443 18788 16488 18816
rect 16025 18779 16083 18785
rect 16482 18776 16488 18788
rect 16540 18776 16546 18828
rect 11514 18748 11520 18760
rect 11427 18720 11520 18748
rect 11514 18708 11520 18720
rect 11572 18748 11578 18760
rect 11793 18751 11851 18757
rect 11793 18748 11805 18751
rect 11572 18720 11805 18748
rect 11572 18708 11578 18720
rect 11793 18717 11805 18720
rect 11839 18717 11851 18751
rect 11793 18711 11851 18717
rect 14645 18751 14703 18757
rect 14645 18717 14657 18751
rect 14691 18748 14703 18751
rect 14734 18748 14740 18760
rect 14691 18720 14740 18748
rect 14691 18717 14703 18720
rect 14645 18711 14703 18717
rect 11808 18680 11836 18711
rect 14734 18708 14740 18720
rect 14792 18708 14798 18760
rect 15381 18751 15439 18757
rect 15381 18717 15393 18751
rect 15427 18748 15439 18751
rect 15841 18751 15899 18757
rect 15841 18748 15853 18751
rect 15427 18720 15853 18748
rect 15427 18717 15439 18720
rect 15381 18711 15439 18717
rect 15841 18717 15853 18720
rect 15887 18748 15899 18751
rect 16114 18748 16120 18760
rect 15887 18720 16120 18748
rect 15887 18717 15899 18720
rect 15841 18711 15899 18717
rect 16114 18708 16120 18720
rect 16172 18708 16178 18760
rect 11882 18680 11888 18692
rect 11808 18652 11888 18680
rect 11882 18640 11888 18652
rect 11940 18640 11946 18692
rect 13170 18680 13176 18692
rect 12636 18652 13176 18680
rect 12636 18624 12664 18652
rect 13170 18640 13176 18652
rect 13228 18640 13234 18692
rect 14001 18683 14059 18689
rect 14001 18649 14013 18683
rect 14047 18680 14059 18683
rect 15102 18680 15108 18692
rect 14047 18652 15108 18680
rect 14047 18649 14059 18652
rect 14001 18643 14059 18649
rect 15102 18640 15108 18652
rect 15160 18640 15166 18692
rect 16574 18680 16580 18692
rect 16535 18652 16580 18680
rect 16574 18640 16580 18652
rect 16632 18640 16638 18692
rect 5353 18615 5411 18621
rect 5353 18581 5365 18615
rect 5399 18612 5411 18615
rect 5718 18612 5724 18624
rect 5399 18584 5724 18612
rect 5399 18581 5411 18584
rect 5353 18575 5411 18581
rect 5718 18572 5724 18584
rect 5776 18572 5782 18624
rect 12253 18615 12311 18621
rect 12253 18581 12265 18615
rect 12299 18612 12311 18615
rect 12618 18612 12624 18624
rect 12299 18584 12624 18612
rect 12299 18581 12311 18584
rect 12253 18575 12311 18581
rect 12618 18572 12624 18584
rect 12676 18572 12682 18624
rect 12986 18572 12992 18624
rect 13044 18612 13050 18624
rect 13265 18615 13323 18621
rect 13265 18612 13277 18615
rect 13044 18584 13277 18612
rect 13044 18572 13050 18584
rect 13265 18581 13277 18584
rect 13311 18581 13323 18615
rect 13265 18575 13323 18581
rect 1104 18522 18860 18544
rect 1104 18470 4315 18522
rect 4367 18470 4379 18522
rect 4431 18470 4443 18522
rect 4495 18470 4507 18522
rect 4559 18470 10982 18522
rect 11034 18470 11046 18522
rect 11098 18470 11110 18522
rect 11162 18470 11174 18522
rect 11226 18470 17648 18522
rect 17700 18470 17712 18522
rect 17764 18470 17776 18522
rect 17828 18470 17840 18522
rect 17892 18470 18860 18522
rect 1104 18448 18860 18470
rect 3786 18408 3792 18420
rect 3747 18380 3792 18408
rect 3786 18368 3792 18380
rect 3844 18368 3850 18420
rect 8018 18408 8024 18420
rect 7979 18380 8024 18408
rect 8018 18368 8024 18380
rect 8076 18368 8082 18420
rect 10870 18408 10876 18420
rect 10831 18380 10876 18408
rect 10870 18368 10876 18380
rect 10928 18368 10934 18420
rect 14642 18408 14648 18420
rect 14603 18380 14648 18408
rect 14642 18368 14648 18380
rect 14700 18368 14706 18420
rect 12158 18340 12164 18352
rect 12119 18312 12164 18340
rect 12158 18300 12164 18312
rect 12216 18300 12222 18352
rect 12526 18300 12532 18352
rect 12584 18340 12590 18352
rect 12621 18343 12679 18349
rect 12621 18340 12633 18343
rect 12584 18312 12633 18340
rect 12584 18300 12590 18312
rect 12621 18309 12633 18312
rect 12667 18309 12679 18343
rect 13630 18340 13636 18352
rect 13591 18312 13636 18340
rect 12621 18303 12679 18309
rect 13630 18300 13636 18312
rect 13688 18300 13694 18352
rect 13814 18300 13820 18352
rect 13872 18300 13878 18352
rect 3694 18232 3700 18284
rect 3752 18272 3758 18284
rect 4154 18272 4160 18284
rect 3752 18244 4160 18272
rect 3752 18232 3758 18244
rect 4154 18232 4160 18244
rect 4212 18232 4218 18284
rect 13832 18272 13860 18300
rect 15933 18275 15991 18281
rect 13832 18244 14228 18272
rect 3786 18164 3792 18216
rect 3844 18204 3850 18216
rect 4433 18207 4491 18213
rect 4433 18204 4445 18207
rect 3844 18176 4445 18204
rect 3844 18164 3850 18176
rect 4433 18173 4445 18176
rect 4479 18173 4491 18207
rect 4433 18167 4491 18173
rect 6365 18207 6423 18213
rect 6365 18173 6377 18207
rect 6411 18204 6423 18207
rect 6641 18207 6699 18213
rect 6641 18204 6653 18207
rect 6411 18176 6653 18204
rect 6411 18173 6423 18176
rect 6365 18167 6423 18173
rect 6641 18173 6653 18176
rect 6687 18173 6699 18207
rect 6917 18207 6975 18213
rect 6917 18204 6929 18207
rect 6641 18167 6699 18173
rect 6748 18176 6929 18204
rect 5813 18139 5871 18145
rect 5813 18105 5825 18139
rect 5859 18136 5871 18139
rect 6457 18139 6515 18145
rect 6457 18136 6469 18139
rect 5859 18108 6469 18136
rect 5859 18105 5871 18108
rect 5813 18099 5871 18105
rect 6457 18105 6469 18108
rect 6503 18136 6515 18139
rect 6748 18136 6776 18176
rect 6917 18173 6929 18176
rect 6963 18173 6975 18207
rect 6917 18167 6975 18173
rect 10505 18207 10563 18213
rect 10505 18173 10517 18207
rect 10551 18204 10563 18207
rect 11425 18207 11483 18213
rect 11425 18204 11437 18207
rect 10551 18176 11437 18204
rect 10551 18173 10563 18176
rect 10505 18167 10563 18173
rect 11425 18173 11437 18176
rect 11471 18173 11483 18207
rect 11790 18204 11796 18216
rect 11751 18176 11796 18204
rect 11425 18167 11483 18173
rect 6503 18108 6776 18136
rect 11440 18136 11468 18167
rect 11790 18164 11796 18176
rect 11848 18164 11854 18216
rect 11882 18164 11888 18216
rect 11940 18204 11946 18216
rect 14200 18213 14228 18244
rect 15933 18241 15945 18275
rect 15979 18272 15991 18275
rect 16390 18272 16396 18284
rect 15979 18244 16396 18272
rect 15979 18241 15991 18244
rect 15933 18235 15991 18241
rect 16390 18232 16396 18244
rect 16448 18232 16454 18284
rect 12069 18207 12127 18213
rect 12069 18204 12081 18207
rect 11940 18176 12081 18204
rect 11940 18164 11946 18176
rect 12069 18173 12081 18176
rect 12115 18173 12127 18207
rect 12069 18167 12127 18173
rect 13817 18207 13875 18213
rect 13817 18173 13829 18207
rect 13863 18173 13875 18207
rect 13817 18167 13875 18173
rect 14185 18207 14243 18213
rect 14185 18173 14197 18207
rect 14231 18173 14243 18207
rect 14185 18167 14243 18173
rect 14277 18207 14335 18213
rect 14277 18173 14289 18207
rect 14323 18204 14335 18207
rect 14734 18204 14740 18216
rect 14323 18176 14740 18204
rect 14323 18173 14335 18176
rect 14277 18167 14335 18173
rect 12526 18136 12532 18148
rect 11440 18108 12532 18136
rect 6503 18105 6515 18108
rect 6457 18099 6515 18105
rect 12526 18096 12532 18108
rect 12584 18096 12590 18148
rect 13265 18139 13323 18145
rect 13265 18105 13277 18139
rect 13311 18136 13323 18139
rect 13832 18136 13860 18167
rect 14734 18164 14740 18176
rect 14792 18164 14798 18216
rect 14918 18164 14924 18216
rect 14976 18204 14982 18216
rect 15657 18207 15715 18213
rect 15657 18204 15669 18207
rect 14976 18176 15669 18204
rect 14976 18164 14982 18176
rect 15657 18173 15669 18176
rect 15703 18173 15715 18207
rect 15657 18167 15715 18173
rect 16114 18164 16120 18216
rect 16172 18204 16178 18216
rect 16485 18207 16543 18213
rect 16485 18204 16497 18207
rect 16172 18176 16497 18204
rect 16172 18164 16178 18176
rect 16485 18173 16497 18176
rect 16531 18173 16543 18207
rect 16850 18204 16856 18216
rect 16811 18176 16856 18204
rect 16485 18167 16543 18173
rect 16850 18164 16856 18176
rect 16908 18164 16914 18216
rect 14550 18136 14556 18148
rect 13311 18108 14556 18136
rect 13311 18105 13323 18108
rect 13265 18099 13323 18105
rect 14550 18096 14556 18108
rect 14608 18096 14614 18148
rect 1670 18068 1676 18080
rect 1631 18040 1676 18068
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 5718 18028 5724 18080
rect 5776 18068 5782 18080
rect 6089 18071 6147 18077
rect 6089 18068 6101 18071
rect 5776 18040 6101 18068
rect 5776 18028 5782 18040
rect 6089 18037 6101 18040
rect 6135 18068 6147 18071
rect 6365 18071 6423 18077
rect 6365 18068 6377 18071
rect 6135 18040 6377 18068
rect 6135 18037 6147 18040
rect 6089 18031 6147 18037
rect 6365 18037 6377 18040
rect 6411 18037 6423 18071
rect 6365 18031 6423 18037
rect 11606 18028 11612 18080
rect 11664 18068 11670 18080
rect 12066 18068 12072 18080
rect 11664 18040 12072 18068
rect 11664 18028 11670 18040
rect 12066 18028 12072 18040
rect 12124 18028 12130 18080
rect 15105 18071 15163 18077
rect 15105 18037 15117 18071
rect 15151 18068 15163 18071
rect 15746 18068 15752 18080
rect 15151 18040 15752 18068
rect 15151 18037 15163 18040
rect 15105 18031 15163 18037
rect 15746 18028 15752 18040
rect 15804 18028 15810 18080
rect 16206 18068 16212 18080
rect 16167 18040 16212 18068
rect 16206 18028 16212 18040
rect 16264 18028 16270 18080
rect 1104 17978 18860 18000
rect 1104 17926 7648 17978
rect 7700 17926 7712 17978
rect 7764 17926 7776 17978
rect 7828 17926 7840 17978
rect 7892 17926 14315 17978
rect 14367 17926 14379 17978
rect 14431 17926 14443 17978
rect 14495 17926 14507 17978
rect 14559 17926 18860 17978
rect 1104 17904 18860 17926
rect 4154 17864 4160 17876
rect 4115 17836 4160 17864
rect 4154 17824 4160 17836
rect 4212 17824 4218 17876
rect 10778 17864 10784 17876
rect 10739 17836 10784 17864
rect 10778 17824 10784 17836
rect 10836 17824 10842 17876
rect 11790 17864 11796 17876
rect 11751 17836 11796 17864
rect 11790 17824 11796 17836
rect 11848 17824 11854 17876
rect 12253 17867 12311 17873
rect 12253 17833 12265 17867
rect 12299 17864 12311 17867
rect 12434 17864 12440 17876
rect 12299 17836 12440 17864
rect 12299 17833 12311 17836
rect 12253 17827 12311 17833
rect 12434 17824 12440 17836
rect 12492 17824 12498 17876
rect 16482 17864 16488 17876
rect 15764 17836 16488 17864
rect 8941 17799 8999 17805
rect 8941 17765 8953 17799
rect 8987 17796 8999 17799
rect 9306 17796 9312 17808
rect 8987 17768 9312 17796
rect 8987 17765 8999 17768
rect 8941 17759 8999 17765
rect 9306 17756 9312 17768
rect 9364 17756 9370 17808
rect 15764 17805 15792 17836
rect 16482 17824 16488 17836
rect 16540 17824 16546 17876
rect 15749 17799 15807 17805
rect 15749 17765 15761 17799
rect 15795 17765 15807 17799
rect 15749 17759 15807 17765
rect 1489 17731 1547 17737
rect 1489 17697 1501 17731
rect 1535 17728 1547 17731
rect 1578 17728 1584 17740
rect 1535 17700 1584 17728
rect 1535 17697 1547 17700
rect 1489 17691 1547 17697
rect 1578 17688 1584 17700
rect 1636 17688 1642 17740
rect 1762 17728 1768 17740
rect 1723 17700 1768 17728
rect 1762 17688 1768 17700
rect 1820 17688 1826 17740
rect 7285 17731 7343 17737
rect 7285 17697 7297 17731
rect 7331 17728 7343 17731
rect 7374 17728 7380 17740
rect 7331 17700 7380 17728
rect 7331 17697 7343 17700
rect 7285 17691 7343 17697
rect 7374 17688 7380 17700
rect 7432 17728 7438 17740
rect 8018 17728 8024 17740
rect 7432 17700 8024 17728
rect 7432 17688 7438 17700
rect 8018 17688 8024 17700
rect 8076 17688 8082 17740
rect 11330 17728 11336 17740
rect 11291 17700 11336 17728
rect 11330 17688 11336 17700
rect 11388 17688 11394 17740
rect 13354 17688 13360 17740
rect 13412 17728 13418 17740
rect 13633 17731 13691 17737
rect 13633 17728 13645 17731
rect 13412 17700 13645 17728
rect 13412 17688 13418 17700
rect 13633 17697 13645 17700
rect 13679 17697 13691 17731
rect 13633 17691 13691 17697
rect 14001 17731 14059 17737
rect 14001 17697 14013 17731
rect 14047 17728 14059 17731
rect 14366 17728 14372 17740
rect 14047 17700 14372 17728
rect 14047 17697 14059 17700
rect 14001 17691 14059 17697
rect 14366 17688 14372 17700
rect 14424 17688 14430 17740
rect 15102 17728 15108 17740
rect 15063 17700 15108 17728
rect 15102 17688 15108 17700
rect 15160 17688 15166 17740
rect 3142 17660 3148 17672
rect 3103 17632 3148 17660
rect 3142 17620 3148 17632
rect 3200 17620 3206 17672
rect 7558 17660 7564 17672
rect 7519 17632 7564 17660
rect 7558 17620 7564 17632
rect 7616 17620 7622 17672
rect 13722 17660 13728 17672
rect 13683 17632 13728 17660
rect 13722 17620 13728 17632
rect 13780 17620 13786 17672
rect 14093 17663 14151 17669
rect 14093 17629 14105 17663
rect 14139 17660 14151 17663
rect 14139 17632 14964 17660
rect 14139 17629 14151 17632
rect 14093 17623 14151 17629
rect 12897 17595 12955 17601
rect 12897 17561 12909 17595
rect 12943 17592 12955 17595
rect 14734 17592 14740 17604
rect 12943 17564 14740 17592
rect 12943 17561 12955 17564
rect 12897 17555 12955 17561
rect 14734 17552 14740 17564
rect 14792 17552 14798 17604
rect 14936 17536 14964 17632
rect 11517 17527 11575 17533
rect 11517 17493 11529 17527
rect 11563 17524 11575 17527
rect 11882 17524 11888 17536
rect 11563 17496 11888 17524
rect 11563 17493 11575 17496
rect 11517 17487 11575 17493
rect 11882 17484 11888 17496
rect 11940 17484 11946 17536
rect 13081 17527 13139 17533
rect 13081 17493 13093 17527
rect 13127 17524 13139 17527
rect 13446 17524 13452 17536
rect 13127 17496 13452 17524
rect 13127 17493 13139 17496
rect 13081 17487 13139 17493
rect 13446 17484 13452 17496
rect 13504 17524 13510 17536
rect 13630 17524 13636 17536
rect 13504 17496 13636 17524
rect 13504 17484 13510 17496
rect 13630 17484 13636 17496
rect 13688 17484 13694 17536
rect 13998 17484 14004 17536
rect 14056 17524 14062 17536
rect 14461 17527 14519 17533
rect 14461 17524 14473 17527
rect 14056 17496 14473 17524
rect 14056 17484 14062 17496
rect 14461 17493 14473 17496
rect 14507 17493 14519 17527
rect 14918 17524 14924 17536
rect 14879 17496 14924 17524
rect 14461 17487 14519 17493
rect 14918 17484 14924 17496
rect 14976 17484 14982 17536
rect 16114 17524 16120 17536
rect 16075 17496 16120 17524
rect 16114 17484 16120 17496
rect 16172 17484 16178 17536
rect 16390 17484 16396 17536
rect 16448 17524 16454 17536
rect 16761 17527 16819 17533
rect 16761 17524 16773 17527
rect 16448 17496 16773 17524
rect 16448 17484 16454 17496
rect 16761 17493 16773 17496
rect 16807 17493 16819 17527
rect 16761 17487 16819 17493
rect 1104 17434 18860 17456
rect 1104 17382 4315 17434
rect 4367 17382 4379 17434
rect 4431 17382 4443 17434
rect 4495 17382 4507 17434
rect 4559 17382 10982 17434
rect 11034 17382 11046 17434
rect 11098 17382 11110 17434
rect 11162 17382 11174 17434
rect 11226 17382 17648 17434
rect 17700 17382 17712 17434
rect 17764 17382 17776 17434
rect 17828 17382 17840 17434
rect 17892 17382 18860 17434
rect 1104 17360 18860 17382
rect 1670 17320 1676 17332
rect 1504 17292 1676 17320
rect 1504 17193 1532 17292
rect 1670 17280 1676 17292
rect 1728 17320 1734 17332
rect 1854 17320 1860 17332
rect 1728 17292 1860 17320
rect 1728 17280 1734 17292
rect 1854 17280 1860 17292
rect 1912 17280 1918 17332
rect 9398 17320 9404 17332
rect 9359 17292 9404 17320
rect 9398 17280 9404 17292
rect 9456 17280 9462 17332
rect 11330 17280 11336 17332
rect 11388 17320 11394 17332
rect 11609 17323 11667 17329
rect 11609 17320 11621 17323
rect 11388 17292 11621 17320
rect 11388 17280 11394 17292
rect 11609 17289 11621 17292
rect 11655 17289 11667 17323
rect 11609 17283 11667 17289
rect 1489 17187 1547 17193
rect 1489 17153 1501 17187
rect 1535 17153 1547 17187
rect 1489 17147 1547 17153
rect 1670 17144 1676 17196
rect 1728 17184 1734 17196
rect 1765 17187 1823 17193
rect 1765 17184 1777 17187
rect 1728 17156 1777 17184
rect 1728 17144 1734 17156
rect 1765 17153 1777 17156
rect 1811 17153 1823 17187
rect 1765 17147 1823 17153
rect 4154 17144 4160 17196
rect 4212 17184 4218 17196
rect 4706 17184 4712 17196
rect 4212 17156 4712 17184
rect 4212 17144 4218 17156
rect 4706 17144 4712 17156
rect 4764 17144 4770 17196
rect 6365 17187 6423 17193
rect 6365 17153 6377 17187
rect 6411 17184 6423 17187
rect 7285 17187 7343 17193
rect 7285 17184 7297 17187
rect 6411 17156 7297 17184
rect 6411 17153 6423 17156
rect 6365 17147 6423 17153
rect 7285 17153 7297 17156
rect 7331 17184 7343 17187
rect 7558 17184 7564 17196
rect 7331 17156 7564 17184
rect 7331 17153 7343 17156
rect 7285 17147 7343 17153
rect 7558 17144 7564 17156
rect 7616 17144 7622 17196
rect 9416 17184 9444 17280
rect 12158 17212 12164 17264
rect 12216 17252 12222 17264
rect 12434 17252 12440 17264
rect 12216 17224 12440 17252
rect 12216 17212 12222 17224
rect 12434 17212 12440 17224
rect 12492 17252 12498 17264
rect 12492 17224 12940 17252
rect 12492 17212 12498 17224
rect 9953 17187 10011 17193
rect 9953 17184 9965 17187
rect 9416 17156 9965 17184
rect 9953 17153 9965 17156
rect 9999 17153 10011 17187
rect 12802 17184 12808 17196
rect 9953 17147 10011 17153
rect 11992 17156 12664 17184
rect 12763 17156 12808 17184
rect 4985 17119 5043 17125
rect 4985 17116 4997 17119
rect 4816 17088 4997 17116
rect 3145 17051 3203 17057
rect 3145 17017 3157 17051
rect 3191 17048 3203 17051
rect 4525 17051 4583 17057
rect 4525 17048 4537 17051
rect 3191 17020 4537 17048
rect 3191 17017 3203 17020
rect 3145 17011 3203 17017
rect 4525 17017 4537 17020
rect 4571 17048 4583 17051
rect 4816 17048 4844 17088
rect 4985 17085 4997 17088
rect 5031 17085 5043 17119
rect 9674 17116 9680 17128
rect 9635 17088 9680 17116
rect 4985 17079 5043 17085
rect 9674 17076 9680 17088
rect 9732 17076 9738 17128
rect 4571 17020 4844 17048
rect 4571 17017 4583 17020
rect 4525 17011 4583 17017
rect 7745 16983 7803 16989
rect 7745 16949 7757 16983
rect 7791 16980 7803 16983
rect 8018 16980 8024 16992
rect 7791 16952 8024 16980
rect 7791 16949 7803 16952
rect 7745 16943 7803 16949
rect 8018 16940 8024 16952
rect 8076 16940 8082 16992
rect 11054 16980 11060 16992
rect 11015 16952 11060 16980
rect 11054 16940 11060 16952
rect 11112 16940 11118 16992
rect 11882 16940 11888 16992
rect 11940 16980 11946 16992
rect 11992 16989 12020 17156
rect 12434 17076 12440 17128
rect 12492 17116 12498 17128
rect 12636 17125 12664 17156
rect 12802 17144 12808 17156
rect 12860 17144 12866 17196
rect 12912 17125 12940 17224
rect 13354 17212 13360 17264
rect 13412 17252 13418 17264
rect 15013 17255 15071 17261
rect 15013 17252 15025 17255
rect 13412 17224 15025 17252
rect 13412 17212 13418 17224
rect 15013 17221 15025 17224
rect 15059 17252 15071 17255
rect 15102 17252 15108 17264
rect 15059 17224 15108 17252
rect 15059 17221 15071 17224
rect 15013 17215 15071 17221
rect 15102 17212 15108 17224
rect 15160 17212 15166 17264
rect 15562 17252 15568 17264
rect 15523 17224 15568 17252
rect 15562 17212 15568 17224
rect 15620 17212 15626 17264
rect 14734 17184 14740 17196
rect 14647 17156 14740 17184
rect 14734 17144 14740 17156
rect 14792 17184 14798 17196
rect 14792 17156 16252 17184
rect 14792 17144 14798 17156
rect 12621 17119 12679 17125
rect 12492 17088 12537 17116
rect 12492 17076 12498 17088
rect 12621 17085 12633 17119
rect 12667 17085 12679 17119
rect 12621 17079 12679 17085
rect 12897 17119 12955 17125
rect 12897 17085 12909 17119
rect 12943 17085 12955 17119
rect 12897 17079 12955 17085
rect 13449 17119 13507 17125
rect 13449 17085 13461 17119
rect 13495 17085 13507 17119
rect 13449 17079 13507 17085
rect 13464 17048 13492 17079
rect 15286 17076 15292 17128
rect 15344 17116 15350 17128
rect 16224 17125 16252 17156
rect 15749 17119 15807 17125
rect 15749 17116 15761 17119
rect 15344 17088 15761 17116
rect 15344 17076 15350 17088
rect 15749 17085 15761 17088
rect 15795 17085 15807 17119
rect 15749 17079 15807 17085
rect 16117 17119 16175 17125
rect 16117 17085 16129 17119
rect 16163 17085 16175 17119
rect 16117 17079 16175 17085
rect 16209 17119 16267 17125
rect 16209 17085 16221 17119
rect 16255 17116 16267 17119
rect 16298 17116 16304 17128
rect 16255 17088 16304 17116
rect 16255 17085 16267 17088
rect 16209 17079 16267 17085
rect 14366 17048 14372 17060
rect 12452 17020 13492 17048
rect 14279 17020 14372 17048
rect 12452 16992 12480 17020
rect 14366 17008 14372 17020
rect 14424 17048 14430 17060
rect 14734 17048 14740 17060
rect 14424 17020 14740 17048
rect 14424 17008 14430 17020
rect 14734 17008 14740 17020
rect 14792 17008 14798 17060
rect 15654 17008 15660 17060
rect 15712 17048 15718 17060
rect 16132 17048 16160 17079
rect 16298 17076 16304 17088
rect 16356 17076 16362 17128
rect 15712 17020 16160 17048
rect 15712 17008 15718 17020
rect 11977 16983 12035 16989
rect 11977 16980 11989 16983
rect 11940 16952 11989 16980
rect 11940 16940 11946 16952
rect 11977 16949 11989 16952
rect 12023 16949 12035 16983
rect 11977 16943 12035 16949
rect 12250 16940 12256 16992
rect 12308 16980 12314 16992
rect 12434 16980 12440 16992
rect 12308 16952 12440 16980
rect 12308 16940 12314 16952
rect 12434 16940 12440 16952
rect 12492 16940 12498 16992
rect 13722 16940 13728 16992
rect 13780 16980 13786 16992
rect 13909 16983 13967 16989
rect 13909 16980 13921 16983
rect 13780 16952 13921 16980
rect 13780 16940 13786 16952
rect 13909 16949 13921 16952
rect 13955 16949 13967 16983
rect 13909 16943 13967 16949
rect 1104 16890 18860 16912
rect 1104 16838 7648 16890
rect 7700 16838 7712 16890
rect 7764 16838 7776 16890
rect 7828 16838 7840 16890
rect 7892 16838 14315 16890
rect 14367 16838 14379 16890
rect 14431 16838 14443 16890
rect 14495 16838 14507 16890
rect 14559 16838 18860 16890
rect 1104 16816 18860 16838
rect 1670 16776 1676 16788
rect 1631 16748 1676 16776
rect 1670 16736 1676 16748
rect 1728 16736 1734 16788
rect 1762 16736 1768 16788
rect 1820 16776 1826 16788
rect 1949 16779 2007 16785
rect 1949 16776 1961 16779
rect 1820 16748 1961 16776
rect 1820 16736 1826 16748
rect 1949 16745 1961 16748
rect 1995 16745 2007 16779
rect 4706 16776 4712 16788
rect 4667 16748 4712 16776
rect 1949 16739 2007 16745
rect 4706 16736 4712 16748
rect 4764 16736 4770 16788
rect 12253 16779 12311 16785
rect 12253 16745 12265 16779
rect 12299 16776 12311 16779
rect 12434 16776 12440 16788
rect 12299 16748 12440 16776
rect 12299 16745 12311 16748
rect 12253 16739 12311 16745
rect 12434 16736 12440 16748
rect 12492 16736 12498 16788
rect 12526 16736 12532 16788
rect 12584 16776 12590 16788
rect 12621 16779 12679 16785
rect 12621 16776 12633 16779
rect 12584 16748 12633 16776
rect 12584 16736 12590 16748
rect 12621 16745 12633 16748
rect 12667 16745 12679 16779
rect 12621 16739 12679 16745
rect 13081 16779 13139 16785
rect 13081 16745 13093 16779
rect 13127 16776 13139 16779
rect 13354 16776 13360 16788
rect 13127 16748 13360 16776
rect 13127 16745 13139 16748
rect 13081 16739 13139 16745
rect 1578 16668 1584 16720
rect 1636 16708 1642 16720
rect 2314 16708 2320 16720
rect 1636 16680 2320 16708
rect 1636 16668 1642 16680
rect 2314 16668 2320 16680
rect 2372 16668 2378 16720
rect 12636 16708 12664 16739
rect 13354 16736 13360 16748
rect 13412 16736 13418 16788
rect 16114 16776 16120 16788
rect 16075 16748 16120 16776
rect 16114 16736 16120 16748
rect 16172 16736 16178 16788
rect 12636 16680 14504 16708
rect 3050 16640 3056 16652
rect 3011 16612 3056 16640
rect 3050 16600 3056 16612
rect 3108 16600 3114 16652
rect 4433 16643 4491 16649
rect 4433 16609 4445 16643
rect 4479 16640 4491 16643
rect 4706 16640 4712 16652
rect 4479 16612 4712 16640
rect 4479 16609 4491 16612
rect 4433 16603 4491 16609
rect 4706 16600 4712 16612
rect 4764 16600 4770 16652
rect 9674 16640 9680 16652
rect 9635 16612 9680 16640
rect 9674 16600 9680 16612
rect 9732 16600 9738 16652
rect 13354 16600 13360 16652
rect 13412 16640 13418 16652
rect 14093 16643 14151 16649
rect 14093 16640 14105 16643
rect 13412 16612 14105 16640
rect 13412 16600 13418 16612
rect 14093 16609 14105 16612
rect 14139 16609 14151 16643
rect 14093 16603 14151 16609
rect 14182 16600 14188 16652
rect 14240 16640 14246 16652
rect 14476 16649 14504 16680
rect 14277 16643 14335 16649
rect 14277 16640 14289 16643
rect 14240 16612 14289 16640
rect 14240 16600 14246 16612
rect 14277 16609 14289 16612
rect 14323 16609 14335 16643
rect 14277 16603 14335 16609
rect 14461 16643 14519 16649
rect 14461 16609 14473 16643
rect 14507 16609 14519 16643
rect 14461 16603 14519 16609
rect 16114 16600 16120 16652
rect 16172 16640 16178 16652
rect 16172 16612 16217 16640
rect 16172 16600 16178 16612
rect 1854 16532 1860 16584
rect 1912 16572 1918 16584
rect 2682 16572 2688 16584
rect 1912 16544 2688 16572
rect 1912 16532 1918 16544
rect 2682 16532 2688 16544
rect 2740 16572 2746 16584
rect 2777 16575 2835 16581
rect 2777 16572 2789 16575
rect 2740 16544 2789 16572
rect 2740 16532 2746 16544
rect 2777 16541 2789 16544
rect 2823 16541 2835 16575
rect 2777 16535 2835 16541
rect 11790 16532 11796 16584
rect 11848 16572 11854 16584
rect 15654 16572 15660 16584
rect 11848 16544 15660 16572
rect 11848 16532 11854 16544
rect 15654 16532 15660 16544
rect 15712 16532 15718 16584
rect 13814 16464 13820 16516
rect 13872 16504 13878 16516
rect 13909 16507 13967 16513
rect 13909 16504 13921 16507
rect 13872 16476 13921 16504
rect 13872 16464 13878 16476
rect 13909 16473 13921 16476
rect 13955 16504 13967 16507
rect 15286 16504 15292 16516
rect 13955 16476 15292 16504
rect 13955 16473 13967 16476
rect 13909 16467 13967 16473
rect 15286 16464 15292 16476
rect 15344 16464 15350 16516
rect 11149 16439 11207 16445
rect 11149 16405 11161 16439
rect 11195 16436 11207 16439
rect 11606 16436 11612 16448
rect 11195 16408 11612 16436
rect 11195 16405 11207 16408
rect 11149 16399 11207 16405
rect 11606 16396 11612 16408
rect 11664 16396 11670 16448
rect 13446 16436 13452 16448
rect 13407 16408 13452 16436
rect 13446 16396 13452 16408
rect 13504 16436 13510 16448
rect 14918 16436 14924 16448
rect 13504 16408 14924 16436
rect 13504 16396 13510 16408
rect 14918 16396 14924 16408
rect 14976 16396 14982 16448
rect 1104 16346 18860 16368
rect 1104 16294 4315 16346
rect 4367 16294 4379 16346
rect 4431 16294 4443 16346
rect 4495 16294 4507 16346
rect 4559 16294 10982 16346
rect 11034 16294 11046 16346
rect 11098 16294 11110 16346
rect 11162 16294 11174 16346
rect 11226 16294 17648 16346
rect 17700 16294 17712 16346
rect 17764 16294 17776 16346
rect 17828 16294 17840 16346
rect 17892 16294 18860 16346
rect 1104 16272 18860 16294
rect 3050 16192 3056 16244
rect 3108 16232 3114 16244
rect 3421 16235 3479 16241
rect 3421 16232 3433 16235
rect 3108 16204 3433 16232
rect 3108 16192 3114 16204
rect 3421 16201 3433 16204
rect 3467 16201 3479 16235
rect 3421 16195 3479 16201
rect 3881 16235 3939 16241
rect 3881 16201 3893 16235
rect 3927 16232 3939 16235
rect 3970 16232 3976 16244
rect 3927 16204 3976 16232
rect 3927 16201 3939 16204
rect 3881 16195 3939 16201
rect 3970 16192 3976 16204
rect 4028 16192 4034 16244
rect 10597 16235 10655 16241
rect 10597 16201 10609 16235
rect 10643 16232 10655 16235
rect 10870 16232 10876 16244
rect 10643 16204 10876 16232
rect 10643 16201 10655 16204
rect 10597 16195 10655 16201
rect 10870 16192 10876 16204
rect 10928 16192 10934 16244
rect 12802 16232 12808 16244
rect 12763 16204 12808 16232
rect 12802 16192 12808 16204
rect 12860 16192 12866 16244
rect 13354 16192 13360 16244
rect 13412 16232 13418 16244
rect 14001 16235 14059 16241
rect 14001 16232 14013 16235
rect 13412 16204 14013 16232
rect 13412 16192 13418 16204
rect 14001 16201 14013 16204
rect 14047 16201 14059 16235
rect 14001 16195 14059 16201
rect 14182 16192 14188 16244
rect 14240 16232 14246 16244
rect 14369 16235 14427 16241
rect 14369 16232 14381 16235
rect 14240 16204 14381 16232
rect 14240 16192 14246 16204
rect 14369 16201 14381 16204
rect 14415 16201 14427 16235
rect 14369 16195 14427 16201
rect 1394 16056 1400 16108
rect 1452 16096 1458 16108
rect 1765 16099 1823 16105
rect 1765 16096 1777 16099
rect 1452 16068 1777 16096
rect 1452 16056 1458 16068
rect 1765 16065 1777 16068
rect 1811 16065 1823 16099
rect 3988 16096 4016 16192
rect 10888 16164 10916 16192
rect 15565 16167 15623 16173
rect 10888 16136 12020 16164
rect 4341 16099 4399 16105
rect 4341 16096 4353 16099
rect 3988 16068 4353 16096
rect 1765 16059 1823 16065
rect 4341 16065 4353 16068
rect 4387 16065 4399 16099
rect 4341 16059 4399 16065
rect 11241 16099 11299 16105
rect 11241 16065 11253 16099
rect 11287 16096 11299 16099
rect 11330 16096 11336 16108
rect 11287 16068 11336 16096
rect 11287 16065 11299 16068
rect 11241 16059 11299 16065
rect 11330 16056 11336 16068
rect 11388 16056 11394 16108
rect 1486 16028 1492 16040
rect 1447 16000 1492 16028
rect 1486 15988 1492 16000
rect 1544 15988 1550 16040
rect 3142 16028 3148 16040
rect 3103 16000 3148 16028
rect 3142 15988 3148 16000
rect 3200 15988 3206 16040
rect 4062 16028 4068 16040
rect 4023 16000 4068 16028
rect 4062 15988 4068 16000
rect 4120 15988 4126 16040
rect 11149 16031 11207 16037
rect 11149 15997 11161 16031
rect 11195 16028 11207 16031
rect 11606 16028 11612 16040
rect 11195 16000 11612 16028
rect 11195 15997 11207 16000
rect 11149 15991 11207 15997
rect 11606 15988 11612 16000
rect 11664 15988 11670 16040
rect 11992 16037 12020 16136
rect 15565 16133 15577 16167
rect 15611 16164 15623 16167
rect 15930 16164 15936 16176
rect 15611 16136 15936 16164
rect 15611 16133 15623 16136
rect 15565 16127 15623 16133
rect 15930 16124 15936 16136
rect 15988 16124 15994 16176
rect 12069 16099 12127 16105
rect 12069 16065 12081 16099
rect 12115 16096 12127 16099
rect 12342 16096 12348 16108
rect 12115 16068 12348 16096
rect 12115 16065 12127 16068
rect 12069 16059 12127 16065
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 15997 12035 16031
rect 11977 15991 12035 15997
rect 10870 15920 10876 15972
rect 10928 15960 10934 15972
rect 10965 15963 11023 15969
rect 10965 15960 10977 15963
rect 10928 15932 10977 15960
rect 10928 15920 10934 15932
rect 10965 15929 10977 15932
rect 11011 15960 11023 15963
rect 12084 15960 12112 16059
rect 12342 16056 12348 16068
rect 12400 16056 12406 16108
rect 13722 16096 13728 16108
rect 13683 16068 13728 16096
rect 13722 16056 13728 16068
rect 13780 16056 13786 16108
rect 15654 16056 15660 16108
rect 15712 16096 15718 16108
rect 16390 16096 16396 16108
rect 15712 16068 16396 16096
rect 15712 16056 15718 16068
rect 12802 15988 12808 16040
rect 12860 16028 12866 16040
rect 13081 16031 13139 16037
rect 13081 16028 13093 16031
rect 12860 16000 13093 16028
rect 12860 15988 12866 16000
rect 13081 15997 13093 16000
rect 13127 15997 13139 16031
rect 13081 15991 13139 15997
rect 15378 15988 15384 16040
rect 15436 16028 15442 16040
rect 16132 16037 16160 16068
rect 16390 16056 16396 16068
rect 16448 16056 16454 16108
rect 15749 16031 15807 16037
rect 15749 16028 15761 16031
rect 15436 16000 15761 16028
rect 15436 15988 15442 16000
rect 15749 15997 15761 16000
rect 15795 15997 15807 16031
rect 15749 15991 15807 15997
rect 15933 16031 15991 16037
rect 15933 15997 15945 16031
rect 15979 15997 15991 16031
rect 15933 15991 15991 15997
rect 16117 16031 16175 16037
rect 16117 15997 16129 16031
rect 16163 15997 16175 16031
rect 16117 15991 16175 15997
rect 11011 15932 12112 15960
rect 11011 15929 11023 15932
rect 10965 15923 11023 15929
rect 5626 15892 5632 15904
rect 5587 15864 5632 15892
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 14918 15852 14924 15904
rect 14976 15892 14982 15904
rect 15013 15895 15071 15901
rect 15013 15892 15025 15895
rect 14976 15864 15025 15892
rect 14976 15852 14982 15864
rect 15013 15861 15025 15864
rect 15059 15892 15071 15895
rect 15948 15892 15976 15991
rect 15059 15864 15976 15892
rect 15059 15861 15071 15864
rect 15013 15855 15071 15861
rect 16114 15852 16120 15904
rect 16172 15892 16178 15904
rect 16669 15895 16727 15901
rect 16669 15892 16681 15895
rect 16172 15864 16681 15892
rect 16172 15852 16178 15864
rect 16669 15861 16681 15864
rect 16715 15892 16727 15895
rect 17034 15892 17040 15904
rect 16715 15864 17040 15892
rect 16715 15861 16727 15864
rect 16669 15855 16727 15861
rect 17034 15852 17040 15864
rect 17092 15852 17098 15904
rect 1104 15802 18860 15824
rect 1104 15750 7648 15802
rect 7700 15750 7712 15802
rect 7764 15750 7776 15802
rect 7828 15750 7840 15802
rect 7892 15750 14315 15802
rect 14367 15750 14379 15802
rect 14431 15750 14443 15802
rect 14495 15750 14507 15802
rect 14559 15750 18860 15802
rect 1104 15728 18860 15750
rect 1394 15648 1400 15700
rect 1452 15688 1458 15700
rect 1581 15691 1639 15697
rect 1581 15688 1593 15691
rect 1452 15660 1593 15688
rect 1452 15648 1458 15660
rect 1581 15657 1593 15660
rect 1627 15657 1639 15691
rect 1581 15651 1639 15657
rect 2869 15691 2927 15697
rect 2869 15657 2881 15691
rect 2915 15688 2927 15691
rect 3421 15691 3479 15697
rect 3421 15688 3433 15691
rect 2915 15660 3433 15688
rect 2915 15657 2927 15660
rect 2869 15651 2927 15657
rect 3421 15657 3433 15660
rect 3467 15688 3479 15691
rect 4062 15688 4068 15700
rect 3467 15660 4068 15688
rect 3467 15657 3479 15660
rect 3421 15651 3479 15657
rect 1486 15308 1492 15360
rect 1544 15348 1550 15360
rect 2041 15351 2099 15357
rect 2041 15348 2053 15351
rect 1544 15320 2053 15348
rect 1544 15308 1550 15320
rect 2041 15317 2053 15320
rect 2087 15348 2099 15351
rect 2682 15348 2688 15360
rect 2087 15320 2688 15348
rect 2087 15317 2099 15320
rect 2041 15311 2099 15317
rect 2682 15308 2688 15320
rect 2740 15348 2746 15360
rect 2884 15348 2912 15651
rect 3528 15561 3556 15660
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 8849 15691 8907 15697
rect 8849 15657 8861 15691
rect 8895 15688 8907 15691
rect 10134 15688 10140 15700
rect 8895 15660 10140 15688
rect 8895 15657 8907 15660
rect 8849 15651 8907 15657
rect 10134 15648 10140 15660
rect 10192 15648 10198 15700
rect 12526 15648 12532 15700
rect 12584 15688 12590 15700
rect 13449 15691 13507 15697
rect 13449 15688 13461 15691
rect 12584 15660 13461 15688
rect 12584 15648 12590 15660
rect 13449 15657 13461 15660
rect 13495 15688 13507 15691
rect 13817 15691 13875 15697
rect 13817 15688 13829 15691
rect 13495 15660 13829 15688
rect 13495 15657 13507 15660
rect 13449 15651 13507 15657
rect 13817 15657 13829 15660
rect 13863 15688 13875 15691
rect 15378 15688 15384 15700
rect 13863 15660 14872 15688
rect 15339 15660 15384 15688
rect 13863 15657 13875 15660
rect 13817 15651 13875 15657
rect 11422 15620 11428 15632
rect 11383 15592 11428 15620
rect 11422 15580 11428 15592
rect 11480 15580 11486 15632
rect 3513 15555 3571 15561
rect 3513 15521 3525 15555
rect 3559 15521 3571 15555
rect 3786 15552 3792 15564
rect 3747 15524 3792 15552
rect 3513 15515 3571 15521
rect 3786 15512 3792 15524
rect 3844 15512 3850 15564
rect 6914 15512 6920 15564
rect 6972 15552 6978 15564
rect 7285 15555 7343 15561
rect 7285 15552 7297 15555
rect 6972 15524 7297 15552
rect 6972 15512 6978 15524
rect 7285 15521 7297 15524
rect 7331 15552 7343 15555
rect 7650 15552 7656 15564
rect 7331 15524 7656 15552
rect 7331 15521 7343 15524
rect 7285 15515 7343 15521
rect 7650 15512 7656 15524
rect 7708 15512 7714 15564
rect 9858 15512 9864 15564
rect 9916 15552 9922 15564
rect 10045 15555 10103 15561
rect 10045 15552 10057 15555
rect 9916 15524 10057 15552
rect 9916 15512 9922 15524
rect 10045 15521 10057 15524
rect 10091 15521 10103 15555
rect 10045 15515 10103 15521
rect 12894 15512 12900 15564
rect 12952 15552 12958 15564
rect 12989 15555 13047 15561
rect 12989 15552 13001 15555
rect 12952 15524 13001 15552
rect 12952 15512 12958 15524
rect 12989 15521 13001 15524
rect 13035 15521 13047 15555
rect 12989 15515 13047 15521
rect 13814 15512 13820 15564
rect 13872 15552 13878 15564
rect 14844 15561 14872 15660
rect 15378 15648 15384 15660
rect 15436 15648 15442 15700
rect 14461 15555 14519 15561
rect 14461 15552 14473 15555
rect 13872 15524 14473 15552
rect 13872 15512 13878 15524
rect 14461 15521 14473 15524
rect 14507 15521 14519 15555
rect 14461 15515 14519 15521
rect 14829 15555 14887 15561
rect 14829 15521 14841 15555
rect 14875 15521 14887 15555
rect 14829 15515 14887 15521
rect 15102 15512 15108 15564
rect 15160 15552 15166 15564
rect 16117 15555 16175 15561
rect 16117 15552 16129 15555
rect 15160 15524 16129 15552
rect 15160 15512 15166 15524
rect 16117 15521 16129 15524
rect 16163 15552 16175 15555
rect 16206 15552 16212 15564
rect 16163 15524 16212 15552
rect 16163 15521 16175 15524
rect 16117 15515 16175 15521
rect 16206 15512 16212 15524
rect 16264 15512 16270 15564
rect 16482 15552 16488 15564
rect 16443 15524 16488 15552
rect 16482 15512 16488 15524
rect 16540 15512 16546 15564
rect 7558 15484 7564 15496
rect 7519 15456 7564 15484
rect 7558 15444 7564 15456
rect 7616 15444 7622 15496
rect 9766 15484 9772 15496
rect 9679 15456 9772 15484
rect 9766 15444 9772 15456
rect 9824 15484 9830 15496
rect 10226 15484 10232 15496
rect 9824 15456 10232 15484
rect 9824 15444 9830 15456
rect 10226 15444 10232 15456
rect 10284 15444 10290 15496
rect 14918 15484 14924 15496
rect 14879 15456 14924 15484
rect 14918 15444 14924 15456
rect 14976 15444 14982 15496
rect 14274 15416 14280 15428
rect 14235 15388 14280 15416
rect 14274 15376 14280 15388
rect 14332 15376 14338 15428
rect 15378 15376 15384 15428
rect 15436 15416 15442 15428
rect 15933 15419 15991 15425
rect 15933 15416 15945 15419
rect 15436 15388 15945 15416
rect 15436 15376 15442 15388
rect 15933 15385 15945 15388
rect 15979 15385 15991 15419
rect 15933 15379 15991 15385
rect 5074 15348 5080 15360
rect 2740 15320 2912 15348
rect 5035 15320 5080 15348
rect 2740 15308 2746 15320
rect 5074 15308 5080 15320
rect 5132 15308 5138 15360
rect 11790 15348 11796 15360
rect 11751 15320 11796 15348
rect 11790 15308 11796 15320
rect 11848 15308 11854 15360
rect 13173 15351 13231 15357
rect 13173 15317 13185 15351
rect 13219 15348 13231 15351
rect 13446 15348 13452 15360
rect 13219 15320 13452 15348
rect 13219 15317 13231 15320
rect 13173 15311 13231 15317
rect 13446 15308 13452 15320
rect 13504 15308 13510 15360
rect 15654 15348 15660 15360
rect 15615 15320 15660 15348
rect 15654 15308 15660 15320
rect 15712 15308 15718 15360
rect 16298 15308 16304 15360
rect 16356 15348 16362 15360
rect 16850 15348 16856 15360
rect 16356 15320 16856 15348
rect 16356 15308 16362 15320
rect 16850 15308 16856 15320
rect 16908 15308 16914 15360
rect 1104 15258 18860 15280
rect 1104 15206 4315 15258
rect 4367 15206 4379 15258
rect 4431 15206 4443 15258
rect 4495 15206 4507 15258
rect 4559 15206 10982 15258
rect 11034 15206 11046 15258
rect 11098 15206 11110 15258
rect 11162 15206 11174 15258
rect 11226 15206 17648 15258
rect 17700 15206 17712 15258
rect 17764 15206 17776 15258
rect 17828 15206 17840 15258
rect 17892 15206 18860 15258
rect 1104 15184 18860 15206
rect 3605 15147 3663 15153
rect 3605 15113 3617 15147
rect 3651 15144 3663 15147
rect 3786 15144 3792 15156
rect 3651 15116 3792 15144
rect 3651 15113 3663 15116
rect 3605 15107 3663 15113
rect 3786 15104 3792 15116
rect 3844 15104 3850 15156
rect 4154 15104 4160 15156
rect 4212 15144 4218 15156
rect 4249 15147 4307 15153
rect 4249 15144 4261 15147
rect 4212 15116 4261 15144
rect 4212 15104 4218 15116
rect 4249 15113 4261 15116
rect 4295 15113 4307 15147
rect 4706 15144 4712 15156
rect 4667 15116 4712 15144
rect 4249 15107 4307 15113
rect 4264 14940 4292 15107
rect 4706 15104 4712 15116
rect 4764 15104 4770 15156
rect 6457 15147 6515 15153
rect 6457 15113 6469 15147
rect 6503 15144 6515 15147
rect 7377 15147 7435 15153
rect 7377 15144 7389 15147
rect 6503 15116 7389 15144
rect 6503 15113 6515 15116
rect 6457 15107 6515 15113
rect 7377 15113 7389 15116
rect 7423 15144 7435 15147
rect 7558 15144 7564 15156
rect 7423 15116 7564 15144
rect 7423 15113 7435 15116
rect 7377 15107 7435 15113
rect 7558 15104 7564 15116
rect 7616 15104 7622 15156
rect 7650 15104 7656 15156
rect 7708 15144 7714 15156
rect 10870 15144 10876 15156
rect 7708 15116 7753 15144
rect 10831 15116 10876 15144
rect 7708 15104 7714 15116
rect 10870 15104 10876 15116
rect 10928 15104 10934 15156
rect 12894 15104 12900 15156
rect 12952 15144 12958 15156
rect 12989 15147 13047 15153
rect 12989 15144 13001 15147
rect 12952 15116 13001 15144
rect 12952 15104 12958 15116
rect 12989 15113 13001 15116
rect 13035 15113 13047 15147
rect 13722 15144 13728 15156
rect 13683 15116 13728 15144
rect 12989 15107 13047 15113
rect 4724 15008 4752 15104
rect 11241 15079 11299 15085
rect 11241 15045 11253 15079
rect 11287 15076 11299 15079
rect 11698 15076 11704 15088
rect 11287 15048 11704 15076
rect 11287 15045 11299 15048
rect 11241 15039 11299 15045
rect 11532 15017 11560 15048
rect 11698 15036 11704 15048
rect 11756 15036 11762 15088
rect 5169 15011 5227 15017
rect 5169 15008 5181 15011
rect 4724 14980 5181 15008
rect 5169 14977 5181 14980
rect 5215 14977 5227 15011
rect 5169 14971 5227 14977
rect 11517 15011 11575 15017
rect 11517 14977 11529 15011
rect 11563 14977 11575 15011
rect 12342 15008 12348 15020
rect 12303 14980 12348 15008
rect 11517 14971 11575 14977
rect 12342 14968 12348 14980
rect 12400 14968 12406 15020
rect 4890 14940 4896 14952
rect 4264 14912 4896 14940
rect 4890 14900 4896 14912
rect 4948 14900 4954 14952
rect 10870 14900 10876 14952
rect 10928 14940 10934 14952
rect 11701 14943 11759 14949
rect 11701 14940 11713 14943
rect 10928 14912 11713 14940
rect 10928 14900 10934 14912
rect 11701 14909 11713 14912
rect 11747 14909 11759 14943
rect 11701 14903 11759 14909
rect 11790 14900 11796 14952
rect 11848 14940 11854 14952
rect 12161 14943 12219 14949
rect 12161 14940 12173 14943
rect 11848 14912 12173 14940
rect 11848 14900 11854 14912
rect 12161 14909 12173 14912
rect 12207 14909 12219 14943
rect 13004 14940 13032 15107
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 15102 15144 15108 15156
rect 15063 15116 15108 15144
rect 15102 15104 15108 15116
rect 15160 15104 15166 15156
rect 15933 15147 15991 15153
rect 15933 15113 15945 15147
rect 15979 15144 15991 15147
rect 16482 15144 16488 15156
rect 15979 15116 16488 15144
rect 15979 15113 15991 15116
rect 15933 15107 15991 15113
rect 16482 15104 16488 15116
rect 16540 15104 16546 15156
rect 16390 15076 16396 15088
rect 16351 15048 16396 15076
rect 16390 15036 16396 15048
rect 16448 15036 16454 15088
rect 13722 14940 13728 14952
rect 13004 14912 13728 14940
rect 12161 14903 12219 14909
rect 13722 14900 13728 14912
rect 13780 14900 13786 14952
rect 14185 14943 14243 14949
rect 14185 14909 14197 14943
rect 14231 14940 14243 14943
rect 14461 14943 14519 14949
rect 14461 14940 14473 14943
rect 14231 14912 14473 14940
rect 14231 14909 14243 14912
rect 14185 14903 14243 14909
rect 14461 14909 14473 14912
rect 14507 14909 14519 14943
rect 14461 14903 14519 14909
rect 15565 14943 15623 14949
rect 15565 14909 15577 14943
rect 15611 14940 15623 14943
rect 16577 14943 16635 14949
rect 16577 14940 16589 14943
rect 15611 14912 16589 14940
rect 15611 14909 15623 14912
rect 15565 14903 15623 14909
rect 16577 14909 16589 14912
rect 16623 14940 16635 14943
rect 16666 14940 16672 14952
rect 16623 14912 16672 14940
rect 16623 14909 16635 14912
rect 16577 14903 16635 14909
rect 16666 14900 16672 14912
rect 16724 14900 16730 14952
rect 16761 14943 16819 14949
rect 16761 14909 16773 14943
rect 16807 14909 16819 14943
rect 16942 14940 16948 14952
rect 16903 14912 16948 14940
rect 16761 14903 16819 14909
rect 14093 14875 14151 14881
rect 14093 14841 14105 14875
rect 14139 14872 14151 14875
rect 14918 14872 14924 14884
rect 14139 14844 14924 14872
rect 14139 14841 14151 14844
rect 14093 14835 14151 14841
rect 9858 14804 9864 14816
rect 9819 14776 9864 14804
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 10226 14804 10232 14816
rect 10187 14776 10232 14804
rect 10226 14764 10232 14776
rect 10284 14764 10290 14816
rect 14384 14813 14412 14844
rect 14918 14832 14924 14844
rect 14976 14872 14982 14884
rect 15102 14872 15108 14884
rect 14976 14844 15108 14872
rect 14976 14832 14982 14844
rect 15102 14832 15108 14844
rect 15160 14832 15166 14884
rect 16776 14872 16804 14903
rect 16942 14900 16948 14912
rect 17000 14940 17006 14952
rect 17405 14943 17463 14949
rect 17405 14940 17417 14943
rect 17000 14912 17417 14940
rect 17000 14900 17006 14912
rect 17405 14909 17417 14912
rect 17451 14909 17463 14943
rect 17405 14903 17463 14909
rect 16850 14872 16856 14884
rect 16776 14844 16856 14872
rect 16850 14832 16856 14844
rect 16908 14832 16914 14884
rect 14369 14807 14427 14813
rect 14369 14773 14381 14807
rect 14415 14773 14427 14807
rect 14369 14767 14427 14773
rect 14461 14807 14519 14813
rect 14461 14773 14473 14807
rect 14507 14804 14519 14807
rect 14737 14807 14795 14813
rect 14737 14804 14749 14807
rect 14507 14776 14749 14804
rect 14507 14773 14519 14776
rect 14461 14767 14519 14773
rect 14737 14773 14749 14776
rect 14783 14804 14795 14807
rect 15286 14804 15292 14816
rect 14783 14776 15292 14804
rect 14783 14773 14795 14776
rect 14737 14767 14795 14773
rect 15286 14764 15292 14776
rect 15344 14804 15350 14816
rect 15838 14804 15844 14816
rect 15344 14776 15844 14804
rect 15344 14764 15350 14776
rect 15838 14764 15844 14776
rect 15896 14764 15902 14816
rect 1104 14714 18860 14736
rect 1104 14662 7648 14714
rect 7700 14662 7712 14714
rect 7764 14662 7776 14714
rect 7828 14662 7840 14714
rect 7892 14662 14315 14714
rect 14367 14662 14379 14714
rect 14431 14662 14443 14714
rect 14495 14662 14507 14714
rect 14559 14662 18860 14714
rect 1104 14640 18860 14662
rect 4890 14600 4896 14612
rect 4851 14572 4896 14600
rect 4890 14560 4896 14572
rect 4948 14560 4954 14612
rect 12253 14603 12311 14609
rect 12253 14569 12265 14603
rect 12299 14600 12311 14603
rect 12434 14600 12440 14612
rect 12299 14572 12440 14600
rect 12299 14569 12311 14572
rect 12253 14563 12311 14569
rect 12434 14560 12440 14572
rect 12492 14600 12498 14612
rect 13354 14600 13360 14612
rect 12492 14572 13360 14600
rect 12492 14560 12498 14572
rect 13354 14560 13360 14572
rect 13412 14560 13418 14612
rect 15378 14600 15384 14612
rect 15339 14572 15384 14600
rect 15378 14560 15384 14572
rect 15436 14600 15442 14612
rect 15436 14572 16804 14600
rect 15436 14560 15442 14572
rect 11517 14535 11575 14541
rect 11517 14501 11529 14535
rect 11563 14532 11575 14535
rect 11698 14532 11704 14544
rect 11563 14504 11704 14532
rect 11563 14501 11575 14504
rect 11517 14495 11575 14501
rect 11698 14492 11704 14504
rect 11756 14492 11762 14544
rect 12710 14532 12716 14544
rect 12671 14504 12716 14532
rect 12710 14492 12716 14504
rect 12768 14492 12774 14544
rect 2314 14464 2320 14476
rect 2275 14436 2320 14464
rect 2314 14424 2320 14436
rect 2372 14424 2378 14476
rect 2590 14464 2596 14476
rect 2551 14436 2596 14464
rect 2590 14424 2596 14436
rect 2648 14424 2654 14476
rect 10686 14424 10692 14476
rect 10744 14464 10750 14476
rect 10873 14467 10931 14473
rect 10873 14464 10885 14467
rect 10744 14436 10885 14464
rect 10744 14424 10750 14436
rect 10873 14433 10885 14436
rect 10919 14433 10931 14467
rect 10873 14427 10931 14433
rect 13814 14424 13820 14476
rect 13872 14464 13878 14476
rect 14458 14464 14464 14476
rect 13872 14436 14464 14464
rect 13872 14424 13878 14436
rect 14458 14424 14464 14436
rect 14516 14424 14522 14476
rect 14550 14424 14556 14476
rect 14608 14464 14614 14476
rect 14645 14467 14703 14473
rect 14645 14464 14657 14467
rect 14608 14436 14657 14464
rect 14608 14424 14614 14436
rect 14645 14433 14657 14436
rect 14691 14433 14703 14467
rect 14645 14427 14703 14433
rect 14829 14467 14887 14473
rect 14829 14433 14841 14467
rect 14875 14433 14887 14467
rect 14829 14427 14887 14433
rect 16393 14467 16451 14473
rect 16393 14433 16405 14467
rect 16439 14464 16451 14467
rect 16482 14464 16488 14476
rect 16439 14436 16488 14464
rect 16439 14433 16451 14436
rect 16393 14427 16451 14433
rect 3970 14396 3976 14408
rect 3931 14368 3976 14396
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 14734 14396 14740 14408
rect 13832 14368 14740 14396
rect 13832 14272 13860 14368
rect 14734 14356 14740 14368
rect 14792 14396 14798 14408
rect 14844 14396 14872 14427
rect 16482 14424 16488 14436
rect 16540 14424 16546 14476
rect 16776 14473 16804 14572
rect 16761 14467 16819 14473
rect 16761 14433 16773 14467
rect 16807 14433 16819 14467
rect 16761 14427 16819 14433
rect 16850 14424 16856 14476
rect 16908 14464 16914 14476
rect 16908 14436 16953 14464
rect 16908 14424 16914 14436
rect 14792 14368 14872 14396
rect 15841 14399 15899 14405
rect 14792 14356 14798 14368
rect 15841 14365 15853 14399
rect 15887 14396 15899 14399
rect 16868 14396 16896 14424
rect 15887 14368 16896 14396
rect 15887 14365 15899 14368
rect 15841 14359 15899 14365
rect 14277 14331 14335 14337
rect 14277 14297 14289 14331
rect 14323 14328 14335 14331
rect 15010 14328 15016 14340
rect 14323 14300 15016 14328
rect 14323 14297 14335 14300
rect 14277 14291 14335 14297
rect 15010 14288 15016 14300
rect 15068 14288 15074 14340
rect 16206 14328 16212 14340
rect 16167 14300 16212 14328
rect 16206 14288 16212 14300
rect 16264 14288 16270 14340
rect 11698 14220 11704 14272
rect 11756 14260 11762 14272
rect 12069 14263 12127 14269
rect 12069 14260 12081 14263
rect 11756 14232 12081 14260
rect 11756 14220 11762 14232
rect 12069 14229 12081 14232
rect 12115 14260 12127 14263
rect 12253 14263 12311 14269
rect 12253 14260 12265 14263
rect 12115 14232 12265 14260
rect 12115 14229 12127 14232
rect 12069 14223 12127 14229
rect 12253 14229 12265 14232
rect 12299 14229 12311 14263
rect 12253 14223 12311 14229
rect 12894 14220 12900 14272
rect 12952 14260 12958 14272
rect 12989 14263 13047 14269
rect 12989 14260 13001 14263
rect 12952 14232 13001 14260
rect 12952 14220 12958 14232
rect 12989 14229 13001 14232
rect 13035 14229 13047 14263
rect 13814 14260 13820 14272
rect 13775 14232 13820 14260
rect 12989 14223 13047 14229
rect 13814 14220 13820 14232
rect 13872 14220 13878 14272
rect 1104 14170 18860 14192
rect 1104 14118 4315 14170
rect 4367 14118 4379 14170
rect 4431 14118 4443 14170
rect 4495 14118 4507 14170
rect 4559 14118 10982 14170
rect 11034 14118 11046 14170
rect 11098 14118 11110 14170
rect 11162 14118 11174 14170
rect 11226 14118 17648 14170
rect 17700 14118 17712 14170
rect 17764 14118 17776 14170
rect 17828 14118 17840 14170
rect 17892 14118 18860 14170
rect 1104 14096 18860 14118
rect 2409 14059 2467 14065
rect 2409 14025 2421 14059
rect 2455 14056 2467 14059
rect 2590 14056 2596 14068
rect 2455 14028 2596 14056
rect 2455 14025 2467 14028
rect 2409 14019 2467 14025
rect 2590 14016 2596 14028
rect 2648 14016 2654 14068
rect 5626 14056 5632 14068
rect 5587 14028 5632 14056
rect 5626 14016 5632 14028
rect 5684 14016 5690 14068
rect 7282 14056 7288 14068
rect 7243 14028 7288 14056
rect 7282 14016 7288 14028
rect 7340 14016 7346 14068
rect 11333 14059 11391 14065
rect 11333 14025 11345 14059
rect 11379 14056 11391 14059
rect 11609 14059 11667 14065
rect 11609 14056 11621 14059
rect 11379 14028 11621 14056
rect 11379 14025 11391 14028
rect 11333 14019 11391 14025
rect 11609 14025 11621 14028
rect 11655 14056 11667 14059
rect 12158 14056 12164 14068
rect 11655 14028 12164 14056
rect 11655 14025 11667 14028
rect 11609 14019 11667 14025
rect 12158 14016 12164 14028
rect 12216 14016 12222 14068
rect 14093 14059 14151 14065
rect 14093 14025 14105 14059
rect 14139 14056 14151 14059
rect 14550 14056 14556 14068
rect 14139 14028 14556 14056
rect 14139 14025 14151 14028
rect 14093 14019 14151 14025
rect 14550 14016 14556 14028
rect 14608 14056 14614 14068
rect 15473 14059 15531 14065
rect 15473 14056 15485 14059
rect 14608 14028 15485 14056
rect 14608 14016 14614 14028
rect 15473 14025 15485 14028
rect 15519 14056 15531 14059
rect 16298 14056 16304 14068
rect 15519 14028 16304 14056
rect 15519 14025 15531 14028
rect 15473 14019 15531 14025
rect 16298 14016 16304 14028
rect 16356 14016 16362 14068
rect 16393 14059 16451 14065
rect 16393 14025 16405 14059
rect 16439 14056 16451 14059
rect 16574 14056 16580 14068
rect 16439 14028 16580 14056
rect 16439 14025 16451 14028
rect 16393 14019 16451 14025
rect 16574 14016 16580 14028
rect 16632 14016 16638 14068
rect 2314 13948 2320 14000
rect 2372 13988 2378 14000
rect 2685 13991 2743 13997
rect 2685 13988 2697 13991
rect 2372 13960 2697 13988
rect 2372 13948 2378 13960
rect 2685 13957 2697 13960
rect 2731 13957 2743 13991
rect 2685 13951 2743 13957
rect 5644 13920 5672 14016
rect 12434 13948 12440 14000
rect 12492 13988 12498 14000
rect 12710 13988 12716 14000
rect 12492 13960 12716 13988
rect 12492 13948 12498 13960
rect 12710 13948 12716 13960
rect 12768 13948 12774 14000
rect 14458 13988 14464 14000
rect 14419 13960 14464 13988
rect 14458 13948 14464 13960
rect 14516 13948 14522 14000
rect 16758 13988 16764 14000
rect 16719 13960 16764 13988
rect 16758 13948 16764 13960
rect 16816 13948 16822 14000
rect 5997 13923 6055 13929
rect 5997 13920 6009 13923
rect 5644 13892 6009 13920
rect 5997 13889 6009 13892
rect 6043 13889 6055 13923
rect 11885 13923 11943 13929
rect 11885 13920 11897 13923
rect 5997 13883 6055 13889
rect 10796 13892 11897 13920
rect 5718 13852 5724 13864
rect 5679 13824 5724 13852
rect 5718 13812 5724 13824
rect 5776 13812 5782 13864
rect 10686 13812 10692 13864
rect 10744 13852 10750 13864
rect 10796 13861 10824 13892
rect 11885 13889 11897 13892
rect 11931 13889 11943 13923
rect 17402 13920 17408 13932
rect 11885 13883 11943 13889
rect 16960 13892 17408 13920
rect 10781 13855 10839 13861
rect 10781 13852 10793 13855
rect 10744 13824 10793 13852
rect 10744 13812 10750 13824
rect 10781 13821 10793 13824
rect 10827 13821 10839 13855
rect 10781 13815 10839 13821
rect 11057 13855 11115 13861
rect 11057 13821 11069 13855
rect 11103 13852 11115 13855
rect 11333 13855 11391 13861
rect 11333 13852 11345 13855
rect 11103 13824 11345 13852
rect 11103 13821 11115 13824
rect 11057 13815 11115 13821
rect 11333 13821 11345 13824
rect 11379 13821 11391 13855
rect 11900 13852 11928 13883
rect 12069 13855 12127 13861
rect 12069 13852 12081 13855
rect 11900 13824 12081 13852
rect 11333 13815 11391 13821
rect 12069 13821 12081 13824
rect 12115 13821 12127 13855
rect 12069 13815 12127 13821
rect 12529 13855 12587 13861
rect 12529 13821 12541 13855
rect 12575 13821 12587 13855
rect 12529 13815 12587 13821
rect 12544 13784 12572 13815
rect 12710 13812 12716 13864
rect 12768 13852 12774 13864
rect 12805 13855 12863 13861
rect 12805 13852 12817 13855
rect 12768 13824 12817 13852
rect 12768 13812 12774 13824
rect 12805 13821 12817 13824
rect 12851 13821 12863 13855
rect 13262 13852 13268 13864
rect 13223 13824 13268 13852
rect 12805 13815 12863 13821
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 13354 13812 13360 13864
rect 13412 13852 13418 13864
rect 15013 13855 15071 13861
rect 15013 13852 15025 13855
rect 13412 13824 13457 13852
rect 13740 13824 15025 13852
rect 13412 13812 13418 13824
rect 12618 13784 12624 13796
rect 12544 13756 12624 13784
rect 12618 13744 12624 13756
rect 12676 13744 12682 13796
rect 13740 13784 13768 13824
rect 15013 13821 15025 13824
rect 15059 13852 15071 13855
rect 15286 13852 15292 13864
rect 15059 13824 15292 13852
rect 15059 13821 15071 13824
rect 15013 13815 15071 13821
rect 15286 13812 15292 13824
rect 15344 13812 15350 13864
rect 16025 13855 16083 13861
rect 16025 13821 16037 13855
rect 16071 13852 16083 13855
rect 16482 13852 16488 13864
rect 16071 13824 16488 13852
rect 16071 13821 16083 13824
rect 16025 13815 16083 13821
rect 16482 13812 16488 13824
rect 16540 13812 16546 13864
rect 16574 13812 16580 13864
rect 16632 13852 16638 13864
rect 16960 13861 16988 13892
rect 17402 13880 17408 13892
rect 17460 13880 17466 13932
rect 16945 13855 17003 13861
rect 16945 13852 16957 13855
rect 16632 13824 16957 13852
rect 16632 13812 16638 13824
rect 16945 13821 16957 13824
rect 16991 13821 17003 13855
rect 17126 13852 17132 13864
rect 17087 13824 17132 13852
rect 16945 13815 17003 13821
rect 17126 13812 17132 13824
rect 17184 13812 17190 13864
rect 17313 13855 17371 13861
rect 17313 13821 17325 13855
rect 17359 13821 17371 13855
rect 17313 13815 17371 13821
rect 12728 13756 13768 13784
rect 12728 13728 12756 13756
rect 16850 13744 16856 13796
rect 16908 13784 16914 13796
rect 17328 13784 17356 13815
rect 16908 13756 17356 13784
rect 16908 13744 16914 13756
rect 10318 13716 10324 13728
rect 10279 13688 10324 13716
rect 10318 13676 10324 13688
rect 10376 13676 10382 13728
rect 10870 13676 10876 13728
rect 10928 13716 10934 13728
rect 11241 13719 11299 13725
rect 11241 13716 11253 13719
rect 10928 13688 11253 13716
rect 10928 13676 10934 13688
rect 11241 13685 11253 13688
rect 11287 13685 11299 13719
rect 11241 13679 11299 13685
rect 12710 13676 12716 13728
rect 12768 13676 12774 13728
rect 1104 13626 18860 13648
rect 1104 13574 7648 13626
rect 7700 13574 7712 13626
rect 7764 13574 7776 13626
rect 7828 13574 7840 13626
rect 7892 13574 14315 13626
rect 14367 13574 14379 13626
rect 14431 13574 14443 13626
rect 14495 13574 14507 13626
rect 14559 13574 18860 13626
rect 1104 13552 18860 13574
rect 1486 13472 1492 13524
rect 1544 13512 1550 13524
rect 1673 13515 1731 13521
rect 1673 13512 1685 13515
rect 1544 13484 1685 13512
rect 1544 13472 1550 13484
rect 1673 13481 1685 13484
rect 1719 13512 1731 13515
rect 2314 13512 2320 13524
rect 1719 13484 2320 13512
rect 1719 13481 1731 13484
rect 1673 13475 1731 13481
rect 2314 13472 2320 13484
rect 2372 13472 2378 13524
rect 4890 13512 4896 13524
rect 4851 13484 4896 13512
rect 4890 13472 4896 13484
rect 4948 13472 4954 13524
rect 5718 13512 5724 13524
rect 5679 13484 5724 13512
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 11330 13472 11336 13524
rect 11388 13512 11394 13524
rect 12161 13515 12219 13521
rect 12161 13512 12173 13515
rect 11388 13484 12173 13512
rect 11388 13472 11394 13484
rect 12161 13481 12173 13484
rect 12207 13512 12219 13515
rect 12618 13512 12624 13524
rect 12207 13484 12624 13512
rect 12207 13481 12219 13484
rect 12161 13475 12219 13481
rect 12618 13472 12624 13484
rect 12676 13512 12682 13524
rect 13170 13512 13176 13524
rect 12676 13484 13176 13512
rect 12676 13472 12682 13484
rect 13170 13472 13176 13484
rect 13228 13472 13234 13524
rect 16298 13472 16304 13524
rect 16356 13512 16362 13524
rect 16485 13515 16543 13521
rect 16485 13512 16497 13515
rect 16356 13484 16497 13512
rect 16356 13472 16362 13484
rect 16485 13481 16497 13484
rect 16531 13481 16543 13515
rect 16850 13512 16856 13524
rect 16811 13484 16856 13512
rect 16485 13475 16543 13481
rect 16850 13472 16856 13484
rect 16908 13472 16914 13524
rect 2332 13376 2360 13472
rect 11517 13447 11575 13453
rect 11517 13413 11529 13447
rect 11563 13444 11575 13447
rect 12894 13444 12900 13456
rect 11563 13416 12900 13444
rect 11563 13413 11575 13416
rect 11517 13407 11575 13413
rect 12894 13404 12900 13416
rect 12952 13404 12958 13456
rect 14918 13404 14924 13456
rect 14976 13444 14982 13456
rect 14976 13416 15700 13444
rect 14976 13404 14982 13416
rect 2958 13376 2964 13388
rect 2332 13348 2964 13376
rect 2958 13336 2964 13348
rect 3016 13336 3022 13388
rect 3234 13376 3240 13388
rect 3195 13348 3240 13376
rect 3234 13336 3240 13348
rect 3292 13336 3298 13388
rect 7466 13336 7472 13388
rect 7524 13376 7530 13388
rect 7561 13379 7619 13385
rect 7561 13376 7573 13379
rect 7524 13348 7573 13376
rect 7524 13336 7530 13348
rect 7561 13345 7573 13348
rect 7607 13345 7619 13379
rect 7561 13339 7619 13345
rect 9217 13379 9275 13385
rect 9217 13345 9229 13379
rect 9263 13376 9275 13379
rect 9490 13376 9496 13388
rect 9263 13348 9496 13376
rect 9263 13345 9275 13348
rect 9217 13339 9275 13345
rect 9490 13336 9496 13348
rect 9548 13336 9554 13388
rect 10318 13376 10324 13388
rect 10279 13348 10324 13376
rect 10318 13336 10324 13348
rect 10376 13336 10382 13388
rect 10870 13376 10876 13388
rect 10831 13348 10876 13376
rect 10870 13336 10876 13348
rect 10928 13336 10934 13388
rect 11333 13379 11391 13385
rect 11333 13345 11345 13379
rect 11379 13376 11391 13379
rect 11422 13376 11428 13388
rect 11379 13348 11428 13376
rect 11379 13345 11391 13348
rect 11333 13339 11391 13345
rect 11422 13336 11428 13348
rect 11480 13336 11486 13388
rect 12529 13379 12587 13385
rect 12529 13345 12541 13379
rect 12575 13345 12587 13379
rect 12802 13376 12808 13388
rect 12763 13348 12808 13376
rect 12529 13339 12587 13345
rect 4614 13308 4620 13320
rect 4575 13280 4620 13308
rect 4614 13268 4620 13280
rect 4672 13268 4678 13320
rect 7834 13308 7840 13320
rect 7795 13280 7840 13308
rect 7834 13268 7840 13280
rect 7892 13268 7898 13320
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13308 10287 13311
rect 10888 13308 10916 13336
rect 10275 13280 10916 13308
rect 12544 13308 12572 13339
rect 12802 13336 12808 13348
rect 12860 13336 12866 13388
rect 13814 13336 13820 13388
rect 13872 13376 13878 13388
rect 14366 13376 14372 13388
rect 13872 13348 14372 13376
rect 13872 13336 13878 13348
rect 14366 13336 14372 13348
rect 14424 13376 14430 13388
rect 15672 13385 15700 13416
rect 14461 13379 14519 13385
rect 14461 13376 14473 13379
rect 14424 13348 14473 13376
rect 14424 13336 14430 13348
rect 14461 13345 14473 13348
rect 14507 13345 14519 13379
rect 14461 13339 14519 13345
rect 15473 13379 15531 13385
rect 15473 13345 15485 13379
rect 15519 13345 15531 13379
rect 15473 13339 15531 13345
rect 15657 13379 15715 13385
rect 15657 13345 15669 13379
rect 15703 13376 15715 13379
rect 15838 13376 15844 13388
rect 15703 13348 15844 13376
rect 15703 13345 15715 13348
rect 15657 13339 15715 13345
rect 12710 13308 12716 13320
rect 12544 13280 12716 13308
rect 10275 13277 10287 13280
rect 10229 13271 10287 13277
rect 12710 13268 12716 13280
rect 12768 13268 12774 13320
rect 13265 13311 13323 13317
rect 13265 13277 13277 13311
rect 13311 13308 13323 13311
rect 13446 13308 13452 13320
rect 13311 13280 13452 13308
rect 13311 13277 13323 13280
rect 13265 13271 13323 13277
rect 13446 13268 13452 13280
rect 13504 13308 13510 13320
rect 13909 13311 13967 13317
rect 13909 13308 13921 13311
rect 13504 13280 13921 13308
rect 13504 13268 13510 13280
rect 13909 13277 13921 13280
rect 13955 13277 13967 13311
rect 14734 13308 14740 13320
rect 14695 13280 14740 13308
rect 13909 13271 13967 13277
rect 14734 13268 14740 13280
rect 14792 13268 14798 13320
rect 15488 13308 15516 13339
rect 15838 13336 15844 13348
rect 15896 13336 15902 13388
rect 15488 13280 15700 13308
rect 15672 13252 15700 13280
rect 12618 13240 12624 13252
rect 12579 13212 12624 13240
rect 12618 13200 12624 13212
rect 12676 13200 12682 13252
rect 14182 13200 14188 13252
rect 14240 13240 14246 13252
rect 15013 13243 15071 13249
rect 15013 13240 15025 13243
rect 14240 13212 15025 13240
rect 14240 13200 14246 13212
rect 15013 13209 15025 13212
rect 15059 13209 15071 13243
rect 15013 13203 15071 13209
rect 15654 13200 15660 13252
rect 15712 13200 15718 13252
rect 9766 13172 9772 13184
rect 9727 13144 9772 13172
rect 9766 13132 9772 13144
rect 9824 13132 9830 13184
rect 13633 13175 13691 13181
rect 13633 13141 13645 13175
rect 13679 13172 13691 13175
rect 13722 13172 13728 13184
rect 13679 13144 13728 13172
rect 13679 13141 13691 13144
rect 13633 13135 13691 13141
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 1104 13082 18860 13104
rect 1104 13030 4315 13082
rect 4367 13030 4379 13082
rect 4431 13030 4443 13082
rect 4495 13030 4507 13082
rect 4559 13030 10982 13082
rect 11034 13030 11046 13082
rect 11098 13030 11110 13082
rect 11162 13030 11174 13082
rect 11226 13030 17648 13082
rect 17700 13030 17712 13082
rect 17764 13030 17776 13082
rect 17828 13030 17840 13082
rect 17892 13030 18860 13082
rect 1104 13008 18860 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 1670 12928 1676 12980
rect 1728 12968 1734 12980
rect 2041 12971 2099 12977
rect 2041 12968 2053 12971
rect 1728 12940 2053 12968
rect 1728 12928 1734 12940
rect 2041 12937 2053 12940
rect 2087 12968 2099 12971
rect 2682 12968 2688 12980
rect 2087 12940 2688 12968
rect 2087 12937 2099 12940
rect 2041 12931 2099 12937
rect 2682 12928 2688 12940
rect 2740 12928 2746 12980
rect 2958 12928 2964 12980
rect 3016 12968 3022 12980
rect 3326 12968 3332 12980
rect 3016 12940 3332 12968
rect 3016 12928 3022 12940
rect 3326 12928 3332 12940
rect 3384 12928 3390 12980
rect 3786 12968 3792 12980
rect 3747 12940 3792 12968
rect 3786 12928 3792 12940
rect 3844 12928 3850 12980
rect 5626 12968 5632 12980
rect 5587 12940 5632 12968
rect 5626 12928 5632 12940
rect 5684 12928 5690 12980
rect 7466 12928 7472 12980
rect 7524 12968 7530 12980
rect 7653 12971 7711 12977
rect 7653 12968 7665 12971
rect 7524 12940 7665 12968
rect 7524 12928 7530 12940
rect 7653 12937 7665 12940
rect 7699 12968 7711 12971
rect 7834 12968 7840 12980
rect 7699 12940 7840 12968
rect 7699 12937 7711 12940
rect 7653 12931 7711 12937
rect 7834 12928 7840 12940
rect 7892 12928 7898 12980
rect 14185 12971 14243 12977
rect 14185 12937 14197 12971
rect 14231 12968 14243 12971
rect 14366 12968 14372 12980
rect 14231 12940 14372 12968
rect 14231 12937 14243 12940
rect 14185 12931 14243 12937
rect 14366 12928 14372 12940
rect 14424 12928 14430 12980
rect 15286 12928 15292 12980
rect 15344 12968 15350 12980
rect 16298 12968 16304 12980
rect 15344 12940 16304 12968
rect 15344 12928 15350 12940
rect 3053 12903 3111 12909
rect 3053 12869 3065 12903
rect 3099 12900 3111 12903
rect 3234 12900 3240 12912
rect 3099 12872 3240 12900
rect 3099 12869 3111 12872
rect 3053 12863 3111 12869
rect 3234 12860 3240 12872
rect 3292 12860 3298 12912
rect 3804 12832 3832 12928
rect 7098 12860 7104 12912
rect 7156 12900 7162 12912
rect 7558 12900 7564 12912
rect 7156 12872 7564 12900
rect 7156 12860 7162 12872
rect 7558 12860 7564 12872
rect 7616 12900 7622 12912
rect 7929 12903 7987 12909
rect 7929 12900 7941 12903
rect 7616 12872 7941 12900
rect 7616 12860 7622 12872
rect 7929 12869 7941 12872
rect 7975 12869 7987 12903
rect 7929 12863 7987 12869
rect 10045 12903 10103 12909
rect 10045 12869 10057 12903
rect 10091 12900 10103 12903
rect 10413 12903 10471 12909
rect 10413 12900 10425 12903
rect 10091 12872 10425 12900
rect 10091 12869 10103 12872
rect 10045 12863 10103 12869
rect 10413 12869 10425 12872
rect 10459 12900 10471 12903
rect 10459 12872 11560 12900
rect 10459 12869 10471 12872
rect 10413 12863 10471 12869
rect 11532 12844 11560 12872
rect 12066 12860 12072 12912
rect 12124 12900 12130 12912
rect 12250 12900 12256 12912
rect 12124 12872 12256 12900
rect 12124 12860 12130 12872
rect 12250 12860 12256 12872
rect 12308 12860 12314 12912
rect 15562 12900 15568 12912
rect 15523 12872 15568 12900
rect 15562 12860 15568 12872
rect 15620 12860 15626 12912
rect 4341 12835 4399 12841
rect 4341 12832 4353 12835
rect 3804 12804 4353 12832
rect 4341 12801 4353 12804
rect 4387 12801 4399 12835
rect 4341 12795 4399 12801
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12832 9551 12835
rect 9539 12804 10916 12832
rect 9539 12801 9551 12804
rect 9493 12795 9551 12801
rect 10888 12776 10916 12804
rect 11514 12792 11520 12844
rect 11572 12792 11578 12844
rect 11790 12832 11796 12844
rect 11751 12804 11796 12832
rect 11790 12792 11796 12804
rect 11848 12792 11854 12844
rect 12529 12835 12587 12841
rect 12529 12801 12541 12835
rect 12575 12832 12587 12835
rect 12802 12832 12808 12844
rect 12575 12804 12808 12832
rect 12575 12801 12587 12804
rect 12529 12795 12587 12801
rect 12802 12792 12808 12804
rect 12860 12792 12866 12844
rect 14553 12835 14611 12841
rect 14553 12801 14565 12835
rect 14599 12832 14611 12835
rect 15654 12832 15660 12844
rect 14599 12804 15660 12832
rect 14599 12801 14611 12804
rect 14553 12795 14611 12801
rect 15654 12792 15660 12804
rect 15712 12792 15718 12844
rect 16224 12841 16252 12940
rect 16298 12928 16304 12940
rect 16356 12968 16362 12980
rect 16577 12971 16635 12977
rect 16577 12968 16589 12971
rect 16356 12940 16589 12968
rect 16356 12928 16362 12940
rect 16577 12937 16589 12940
rect 16623 12968 16635 12971
rect 16758 12968 16764 12980
rect 16623 12940 16764 12968
rect 16623 12937 16635 12940
rect 16577 12931 16635 12937
rect 16758 12928 16764 12940
rect 16816 12968 16822 12980
rect 17126 12968 17132 12980
rect 16816 12940 17132 12968
rect 16816 12928 16822 12940
rect 17126 12928 17132 12940
rect 17184 12928 17190 12980
rect 16209 12835 16267 12841
rect 16209 12801 16221 12835
rect 16255 12801 16267 12835
rect 16209 12795 16267 12801
rect 4062 12764 4068 12776
rect 3975 12736 4068 12764
rect 4062 12724 4068 12736
rect 4120 12764 4126 12776
rect 4798 12764 4804 12776
rect 4120 12736 4804 12764
rect 4120 12724 4126 12736
rect 4798 12724 4804 12736
rect 4856 12724 4862 12776
rect 9766 12724 9772 12776
rect 9824 12764 9830 12776
rect 10597 12767 10655 12773
rect 10597 12764 10609 12767
rect 9824 12736 10609 12764
rect 9824 12724 9830 12736
rect 10597 12733 10609 12736
rect 10643 12733 10655 12767
rect 10597 12727 10655 12733
rect 10870 12724 10876 12776
rect 10928 12764 10934 12776
rect 11241 12767 11299 12773
rect 11241 12764 11253 12767
rect 10928 12736 11253 12764
rect 10928 12724 10934 12736
rect 11241 12733 11253 12736
rect 11287 12733 11299 12767
rect 11241 12727 11299 12733
rect 11425 12767 11483 12773
rect 11425 12733 11437 12767
rect 11471 12764 11483 12767
rect 11532 12764 11560 12792
rect 12894 12764 12900 12776
rect 11471 12736 11560 12764
rect 12855 12736 12900 12764
rect 11471 12733 11483 12736
rect 11425 12727 11483 12733
rect 11256 12696 11284 12727
rect 12894 12724 12900 12736
rect 12952 12724 12958 12776
rect 13078 12764 13084 12776
rect 13039 12736 13084 12764
rect 13078 12724 13084 12736
rect 13136 12724 13142 12776
rect 13446 12764 13452 12776
rect 13407 12736 13452 12764
rect 13446 12724 13452 12736
rect 13504 12724 13510 12776
rect 15105 12767 15163 12773
rect 15105 12733 15117 12767
rect 15151 12764 15163 12767
rect 15378 12764 15384 12776
rect 15151 12736 15384 12764
rect 15151 12733 15163 12736
rect 15105 12727 15163 12733
rect 15378 12724 15384 12736
rect 15436 12764 15442 12776
rect 15749 12767 15807 12773
rect 15749 12764 15761 12767
rect 15436 12736 15761 12764
rect 15436 12724 15442 12736
rect 15749 12733 15761 12736
rect 15795 12733 15807 12767
rect 16114 12764 16120 12776
rect 16075 12736 16120 12764
rect 15749 12727 15807 12733
rect 16114 12724 16120 12736
rect 16172 12764 16178 12776
rect 17313 12767 17371 12773
rect 17313 12764 17325 12767
rect 16172 12736 17325 12764
rect 16172 12724 16178 12736
rect 17313 12733 17325 12736
rect 17359 12733 17371 12767
rect 17313 12727 17371 12733
rect 11514 12696 11520 12708
rect 11256 12668 11520 12696
rect 11514 12656 11520 12668
rect 11572 12656 11578 12708
rect 13722 12696 13728 12708
rect 13683 12668 13728 12696
rect 13722 12656 13728 12668
rect 13780 12656 13786 12708
rect 1946 12588 1952 12640
rect 2004 12628 2010 12640
rect 2317 12631 2375 12637
rect 2317 12628 2329 12631
rect 2004 12600 2329 12628
rect 2004 12588 2010 12600
rect 2317 12597 2329 12600
rect 2363 12597 2375 12631
rect 2317 12591 2375 12597
rect 10502 12588 10508 12640
rect 10560 12628 10566 12640
rect 12161 12631 12219 12637
rect 12161 12628 12173 12631
rect 10560 12600 12173 12628
rect 10560 12588 10566 12600
rect 12161 12597 12173 12600
rect 12207 12628 12219 12631
rect 12618 12628 12624 12640
rect 12207 12600 12624 12628
rect 12207 12597 12219 12600
rect 12161 12591 12219 12597
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 16942 12628 16948 12640
rect 16903 12600 16948 12628
rect 16942 12588 16948 12600
rect 17000 12588 17006 12640
rect 1104 12538 18860 12560
rect 1104 12486 7648 12538
rect 7700 12486 7712 12538
rect 7764 12486 7776 12538
rect 7828 12486 7840 12538
rect 7892 12486 14315 12538
rect 14367 12486 14379 12538
rect 14431 12486 14443 12538
rect 14495 12486 14507 12538
rect 14559 12486 18860 12538
rect 1104 12464 18860 12486
rect 11330 12384 11336 12436
rect 11388 12424 11394 12436
rect 11388 12396 11560 12424
rect 11388 12384 11394 12396
rect 3050 12356 3056 12368
rect 3011 12328 3056 12356
rect 3050 12316 3056 12328
rect 3108 12316 3114 12368
rect 8481 12359 8539 12365
rect 8481 12325 8493 12359
rect 8527 12356 8539 12359
rect 9214 12356 9220 12368
rect 8527 12328 9220 12356
rect 8527 12325 8539 12328
rect 8481 12319 8539 12325
rect 9214 12316 9220 12328
rect 9272 12316 9278 12368
rect 10502 12356 10508 12368
rect 10463 12328 10508 12356
rect 10502 12316 10508 12328
rect 10560 12316 10566 12368
rect 11532 12356 11560 12396
rect 11698 12384 11704 12436
rect 11756 12424 11762 12436
rect 11790 12424 11796 12436
rect 11756 12396 11796 12424
rect 11756 12384 11762 12396
rect 11790 12384 11796 12396
rect 11848 12384 11854 12436
rect 11974 12384 11980 12436
rect 12032 12384 12038 12436
rect 12710 12384 12716 12436
rect 12768 12424 12774 12436
rect 12989 12427 13047 12433
rect 12989 12424 13001 12427
rect 12768 12396 13001 12424
rect 12768 12384 12774 12396
rect 12989 12393 13001 12396
rect 13035 12393 13047 12427
rect 14918 12424 14924 12436
rect 14879 12396 14924 12424
rect 12989 12387 13047 12393
rect 14918 12384 14924 12396
rect 14976 12384 14982 12436
rect 11992 12356 12020 12384
rect 12250 12356 12256 12368
rect 11532 12328 12020 12356
rect 12211 12328 12256 12356
rect 12250 12316 12256 12328
rect 12308 12316 12314 12368
rect 15930 12316 15936 12368
rect 15988 12356 15994 12368
rect 15988 12328 16068 12356
rect 15988 12316 15994 12328
rect 1670 12288 1676 12300
rect 1631 12260 1676 12288
rect 1670 12248 1676 12260
rect 1728 12248 1734 12300
rect 3786 12248 3792 12300
rect 3844 12288 3850 12300
rect 4525 12291 4583 12297
rect 4525 12288 4537 12291
rect 3844 12260 4537 12288
rect 3844 12248 3850 12260
rect 4525 12257 4537 12260
rect 4571 12257 4583 12291
rect 4525 12251 4583 12257
rect 6546 12248 6552 12300
rect 6604 12288 6610 12300
rect 7101 12291 7159 12297
rect 7101 12288 7113 12291
rect 6604 12260 7113 12288
rect 6604 12248 6610 12260
rect 7101 12257 7113 12260
rect 7147 12257 7159 12291
rect 7101 12251 7159 12257
rect 10134 12248 10140 12300
rect 10192 12288 10198 12300
rect 10413 12291 10471 12297
rect 10413 12288 10425 12291
rect 10192 12260 10425 12288
rect 10192 12248 10198 12260
rect 10413 12257 10425 12260
rect 10459 12288 10471 12291
rect 11333 12291 11391 12297
rect 11333 12288 11345 12291
rect 10459 12260 11345 12288
rect 10459 12257 10471 12260
rect 10413 12251 10471 12257
rect 11333 12257 11345 12260
rect 11379 12288 11391 12291
rect 11882 12288 11888 12300
rect 11379 12260 11888 12288
rect 11379 12257 11391 12260
rect 11333 12251 11391 12257
rect 11882 12248 11888 12260
rect 11940 12248 11946 12300
rect 13262 12288 13268 12300
rect 13223 12260 13268 12288
rect 13262 12248 13268 12260
rect 13320 12248 13326 12300
rect 13722 12288 13728 12300
rect 13683 12260 13728 12288
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 14182 12288 14188 12300
rect 14143 12260 14188 12288
rect 14182 12248 14188 12260
rect 14240 12248 14246 12300
rect 14461 12291 14519 12297
rect 14461 12257 14473 12291
rect 14507 12257 14519 12291
rect 14461 12251 14519 12257
rect 1397 12223 1455 12229
rect 1397 12189 1409 12223
rect 1443 12220 1455 12223
rect 1854 12220 1860 12232
rect 1443 12192 1860 12220
rect 1443 12189 1455 12192
rect 1397 12183 1455 12189
rect 1854 12180 1860 12192
rect 1912 12180 1918 12232
rect 4249 12223 4307 12229
rect 4249 12220 4261 12223
rect 4080 12192 4261 12220
rect 4080 12096 4108 12192
rect 4249 12189 4261 12192
rect 4295 12189 4307 12223
rect 4249 12183 4307 12189
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12220 6883 12223
rect 7006 12220 7012 12232
rect 6871 12192 7012 12220
rect 6871 12189 6883 12192
rect 6825 12183 6883 12189
rect 7006 12180 7012 12192
rect 7064 12180 7070 12232
rect 10045 12223 10103 12229
rect 10045 12189 10057 12223
rect 10091 12220 10103 12223
rect 11057 12223 11115 12229
rect 11057 12220 11069 12223
rect 10091 12192 11069 12220
rect 10091 12189 10103 12192
rect 10045 12183 10103 12189
rect 11057 12189 11069 12192
rect 11103 12220 11115 12223
rect 11238 12220 11244 12232
rect 11103 12192 11244 12220
rect 11103 12189 11115 12192
rect 11057 12183 11115 12189
rect 11238 12180 11244 12192
rect 11296 12180 11302 12232
rect 11517 12223 11575 12229
rect 11517 12189 11529 12223
rect 11563 12220 11575 12223
rect 13538 12220 13544 12232
rect 11563 12192 13544 12220
rect 11563 12189 11575 12192
rect 11517 12183 11575 12189
rect 10502 12112 10508 12164
rect 10560 12152 10566 12164
rect 11532 12152 11560 12183
rect 13538 12180 13544 12192
rect 13596 12180 13602 12232
rect 13814 12220 13820 12232
rect 13775 12192 13820 12220
rect 13814 12180 13820 12192
rect 13872 12180 13878 12232
rect 13998 12180 14004 12232
rect 14056 12220 14062 12232
rect 14476 12220 14504 12251
rect 15746 12248 15752 12300
rect 15804 12248 15810 12300
rect 14056 12192 14504 12220
rect 15657 12223 15715 12229
rect 14056 12180 14062 12192
rect 15657 12189 15669 12223
rect 15703 12220 15715 12223
rect 15764 12220 15792 12248
rect 16040 12232 16068 12328
rect 16574 12288 16580 12300
rect 16535 12260 16580 12288
rect 16574 12248 16580 12260
rect 16632 12248 16638 12300
rect 16758 12288 16764 12300
rect 16719 12260 16764 12288
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 16945 12291 17003 12297
rect 16945 12257 16957 12291
rect 16991 12288 17003 12291
rect 17310 12288 17316 12300
rect 16991 12260 17316 12288
rect 16991 12257 17003 12260
rect 16945 12251 17003 12257
rect 17310 12248 17316 12260
rect 17368 12248 17374 12300
rect 15930 12220 15936 12232
rect 15703 12192 15936 12220
rect 15703 12189 15715 12192
rect 15657 12183 15715 12189
rect 15930 12180 15936 12192
rect 15988 12180 15994 12232
rect 16022 12180 16028 12232
rect 16080 12180 16086 12232
rect 16390 12152 16396 12164
rect 10560 12124 11560 12152
rect 16351 12124 16396 12152
rect 10560 12112 10566 12124
rect 16390 12112 16396 12124
rect 16448 12112 16454 12164
rect 4062 12084 4068 12096
rect 4023 12056 4068 12084
rect 4062 12044 4068 12056
rect 4120 12044 4126 12096
rect 5810 12084 5816 12096
rect 5771 12056 5816 12084
rect 5810 12044 5816 12056
rect 5868 12044 5874 12096
rect 11422 12044 11428 12096
rect 11480 12084 11486 12096
rect 11606 12084 11612 12096
rect 11480 12056 11612 12084
rect 11480 12044 11486 12056
rect 11606 12044 11612 12056
rect 11664 12084 11670 12096
rect 11793 12087 11851 12093
rect 11793 12084 11805 12087
rect 11664 12056 11805 12084
rect 11664 12044 11670 12056
rect 11793 12053 11805 12056
rect 11839 12053 11851 12087
rect 12710 12084 12716 12096
rect 12671 12056 12716 12084
rect 11793 12047 11851 12053
rect 12710 12044 12716 12056
rect 12768 12084 12774 12096
rect 13078 12084 13084 12096
rect 12768 12056 13084 12084
rect 12768 12044 12774 12056
rect 13078 12044 13084 12056
rect 13136 12044 13142 12096
rect 14182 12044 14188 12096
rect 14240 12084 14246 12096
rect 14734 12084 14740 12096
rect 14240 12056 14740 12084
rect 14240 12044 14246 12056
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 14826 12044 14832 12096
rect 14884 12084 14890 12096
rect 15286 12084 15292 12096
rect 14884 12056 15292 12084
rect 14884 12044 14890 12056
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 15746 12044 15752 12096
rect 15804 12084 15810 12096
rect 15933 12087 15991 12093
rect 15933 12084 15945 12087
rect 15804 12056 15945 12084
rect 15804 12044 15810 12056
rect 15933 12053 15945 12056
rect 15979 12053 15991 12087
rect 15933 12047 15991 12053
rect 1104 11994 18860 12016
rect 1104 11942 4315 11994
rect 4367 11942 4379 11994
rect 4431 11942 4443 11994
rect 4495 11942 4507 11994
rect 4559 11942 10982 11994
rect 11034 11942 11046 11994
rect 11098 11942 11110 11994
rect 11162 11942 11174 11994
rect 11226 11942 17648 11994
rect 17700 11942 17712 11994
rect 17764 11942 17776 11994
rect 17828 11942 17840 11994
rect 17892 11942 18860 11994
rect 1104 11920 18860 11942
rect 2958 11880 2964 11892
rect 2919 11852 2964 11880
rect 2958 11840 2964 11852
rect 3016 11840 3022 11892
rect 3786 11880 3792 11892
rect 3747 11852 3792 11880
rect 3786 11840 3792 11852
rect 3844 11840 3850 11892
rect 5902 11880 5908 11892
rect 5863 11852 5908 11880
rect 5902 11840 5908 11852
rect 5960 11840 5966 11892
rect 8478 11880 8484 11892
rect 8439 11852 8484 11880
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 10502 11880 10508 11892
rect 10463 11852 10508 11880
rect 10502 11840 10508 11852
rect 10560 11840 10566 11892
rect 13262 11840 13268 11892
rect 13320 11880 13326 11892
rect 14645 11883 14703 11889
rect 14645 11880 14657 11883
rect 13320 11852 14657 11880
rect 13320 11840 13326 11852
rect 14645 11849 14657 11852
rect 14691 11880 14703 11883
rect 14734 11880 14740 11892
rect 14691 11852 14740 11880
rect 14691 11849 14703 11852
rect 14645 11843 14703 11849
rect 14734 11840 14740 11852
rect 14792 11840 14798 11892
rect 16574 11840 16580 11892
rect 16632 11880 16638 11892
rect 16945 11883 17003 11889
rect 16945 11880 16957 11883
rect 16632 11852 16957 11880
rect 16632 11840 16638 11852
rect 16945 11849 16957 11852
rect 16991 11849 17003 11883
rect 16945 11843 17003 11849
rect 13630 11812 13636 11824
rect 13591 11784 13636 11812
rect 13630 11772 13636 11784
rect 13688 11772 13694 11824
rect 16485 11815 16543 11821
rect 16485 11781 16497 11815
rect 16531 11812 16543 11815
rect 16666 11812 16672 11824
rect 16531 11784 16672 11812
rect 16531 11781 16543 11784
rect 16485 11775 16543 11781
rect 16666 11772 16672 11784
rect 16724 11772 16730 11824
rect 1578 11704 1584 11756
rect 1636 11744 1642 11756
rect 1673 11747 1731 11753
rect 1673 11744 1685 11747
rect 1636 11716 1685 11744
rect 1636 11704 1642 11716
rect 1673 11713 1685 11716
rect 1719 11713 1731 11747
rect 1673 11707 1731 11713
rect 9306 11704 9312 11756
rect 9364 11744 9370 11756
rect 9582 11744 9588 11756
rect 9364 11716 9588 11744
rect 9364 11704 9370 11716
rect 9582 11704 9588 11716
rect 9640 11704 9646 11756
rect 11054 11744 11060 11756
rect 11015 11716 11060 11744
rect 11054 11704 11060 11716
rect 11112 11704 11118 11756
rect 12897 11747 12955 11753
rect 12897 11713 12909 11747
rect 12943 11744 12955 11747
rect 13722 11744 13728 11756
rect 12943 11716 13728 11744
rect 12943 11713 12955 11716
rect 12897 11707 12955 11713
rect 13722 11704 13728 11716
rect 13780 11704 13786 11756
rect 15102 11704 15108 11756
rect 15160 11744 15166 11756
rect 15654 11744 15660 11756
rect 15160 11716 15660 11744
rect 15160 11704 15166 11716
rect 15654 11704 15660 11716
rect 15712 11704 15718 11756
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 1486 11676 1492 11688
rect 1443 11648 1492 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 1486 11636 1492 11648
rect 1544 11636 1550 11688
rect 4062 11636 4068 11688
rect 4120 11676 4126 11688
rect 4341 11679 4399 11685
rect 4341 11676 4353 11679
rect 4120 11648 4353 11676
rect 4120 11636 4126 11648
rect 4341 11645 4353 11648
rect 4387 11645 4399 11679
rect 4617 11679 4675 11685
rect 4617 11676 4629 11679
rect 4341 11639 4399 11645
rect 4448 11648 4629 11676
rect 3418 11540 3424 11552
rect 3379 11512 3424 11540
rect 3418 11500 3424 11512
rect 3476 11540 3482 11552
rect 4448 11540 4476 11648
rect 4617 11645 4629 11648
rect 4663 11645 4675 11679
rect 7098 11676 7104 11688
rect 7059 11648 7104 11676
rect 4617 11639 4675 11645
rect 7098 11636 7104 11648
rect 7156 11636 7162 11688
rect 7377 11679 7435 11685
rect 7377 11676 7389 11679
rect 7208 11648 7389 11676
rect 6546 11540 6552 11552
rect 3476 11512 4476 11540
rect 6507 11512 6552 11540
rect 3476 11500 3482 11512
rect 6546 11500 6552 11512
rect 6604 11500 6610 11552
rect 6914 11540 6920 11552
rect 6875 11512 6920 11540
rect 6914 11500 6920 11512
rect 6972 11540 6978 11552
rect 7208 11540 7236 11648
rect 7377 11645 7389 11648
rect 7423 11645 7435 11679
rect 10134 11676 10140 11688
rect 10095 11648 10140 11676
rect 7377 11639 7435 11645
rect 10134 11636 10140 11648
rect 10192 11636 10198 11688
rect 11241 11679 11299 11685
rect 11241 11645 11253 11679
rect 11287 11645 11299 11679
rect 11241 11639 11299 11645
rect 11333 11679 11391 11685
rect 11333 11645 11345 11679
rect 11379 11645 11391 11679
rect 11333 11639 11391 11645
rect 6972 11512 7236 11540
rect 6972 11500 6978 11512
rect 10686 11500 10692 11552
rect 10744 11540 10750 11552
rect 10873 11543 10931 11549
rect 10873 11540 10885 11543
rect 10744 11512 10885 11540
rect 10744 11500 10750 11512
rect 10873 11509 10885 11512
rect 10919 11540 10931 11543
rect 11256 11540 11284 11639
rect 11348 11608 11376 11639
rect 11422 11636 11428 11688
rect 11480 11676 11486 11688
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 11480 11648 11713 11676
rect 11480 11636 11486 11648
rect 11701 11645 11713 11648
rect 11747 11645 11759 11679
rect 11701 11639 11759 11645
rect 11790 11636 11796 11688
rect 11848 11676 11854 11688
rect 12253 11679 12311 11685
rect 12253 11676 12265 11679
rect 11848 11648 12265 11676
rect 11848 11636 11854 11648
rect 12253 11645 12265 11648
rect 12299 11645 12311 11679
rect 13814 11676 13820 11688
rect 13775 11648 13820 11676
rect 12253 11639 12311 11645
rect 13814 11636 13820 11648
rect 13872 11636 13878 11688
rect 14182 11676 14188 11688
rect 14143 11648 14188 11676
rect 14182 11636 14188 11648
rect 14240 11636 14246 11688
rect 14274 11636 14280 11688
rect 14332 11676 14338 11688
rect 14826 11676 14832 11688
rect 14332 11648 14832 11676
rect 14332 11636 14338 11648
rect 14826 11636 14832 11648
rect 14884 11636 14890 11688
rect 15746 11676 15752 11688
rect 15707 11648 15752 11676
rect 15746 11636 15752 11648
rect 15804 11636 15810 11688
rect 15930 11676 15936 11688
rect 15891 11648 15936 11676
rect 15930 11636 15936 11648
rect 15988 11636 15994 11688
rect 16298 11636 16304 11688
rect 16356 11676 16362 11688
rect 16393 11679 16451 11685
rect 16393 11676 16405 11679
rect 16356 11648 16405 11676
rect 16356 11636 16362 11648
rect 16393 11645 16405 11648
rect 16439 11645 16451 11679
rect 16393 11639 16451 11645
rect 11882 11608 11888 11620
rect 11348 11580 11888 11608
rect 11882 11568 11888 11580
rect 11940 11568 11946 11620
rect 11698 11540 11704 11552
rect 10919 11512 11704 11540
rect 10919 11509 10931 11512
rect 10873 11503 10931 11509
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 12710 11500 12716 11552
rect 12768 11540 12774 11552
rect 13265 11543 13323 11549
rect 13265 11540 13277 11543
rect 12768 11512 13277 11540
rect 12768 11500 12774 11512
rect 13265 11509 13277 11512
rect 13311 11540 13323 11543
rect 13998 11540 14004 11552
rect 13311 11512 14004 11540
rect 13311 11509 13323 11512
rect 13265 11503 13323 11509
rect 13998 11500 14004 11512
rect 14056 11500 14062 11552
rect 15102 11540 15108 11552
rect 15063 11512 15108 11540
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 17310 11540 17316 11552
rect 17271 11512 17316 11540
rect 17310 11500 17316 11512
rect 17368 11500 17374 11552
rect 1104 11450 18860 11472
rect 1104 11398 7648 11450
rect 7700 11398 7712 11450
rect 7764 11398 7776 11450
rect 7828 11398 7840 11450
rect 7892 11398 14315 11450
rect 14367 11398 14379 11450
rect 14431 11398 14443 11450
rect 14495 11398 14507 11450
rect 14559 11398 18860 11450
rect 1104 11376 18860 11398
rect 8110 11336 8116 11348
rect 8071 11308 8116 11336
rect 8110 11296 8116 11308
rect 8168 11296 8174 11348
rect 12250 11336 12256 11348
rect 12211 11308 12256 11336
rect 12250 11296 12256 11308
rect 12308 11296 12314 11348
rect 14090 11296 14096 11348
rect 14148 11336 14154 11348
rect 14553 11339 14611 11345
rect 14553 11336 14565 11339
rect 14148 11308 14565 11336
rect 14148 11296 14154 11308
rect 14553 11305 14565 11308
rect 14599 11305 14611 11339
rect 14553 11299 14611 11305
rect 5813 11271 5871 11277
rect 5813 11237 5825 11271
rect 5859 11268 5871 11271
rect 6546 11268 6552 11280
rect 5859 11240 6552 11268
rect 5859 11237 5871 11240
rect 5813 11231 5871 11237
rect 6546 11228 6552 11240
rect 6604 11228 6610 11280
rect 9953 11271 10011 11277
rect 9953 11237 9965 11271
rect 9999 11268 10011 11271
rect 11790 11268 11796 11280
rect 9999 11240 11796 11268
rect 9999 11237 10011 11240
rect 9953 11231 10011 11237
rect 1762 11200 1768 11212
rect 1675 11172 1768 11200
rect 1762 11160 1768 11172
rect 1820 11200 1826 11212
rect 2222 11200 2228 11212
rect 1820 11172 2228 11200
rect 1820 11160 1826 11172
rect 2222 11160 2228 11172
rect 2280 11160 2286 11212
rect 3786 11160 3792 11212
rect 3844 11200 3850 11212
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 3844 11172 4445 11200
rect 3844 11160 3850 11172
rect 4433 11169 4445 11172
rect 4479 11169 4491 11203
rect 10042 11200 10048 11212
rect 10003 11172 10048 11200
rect 4433 11163 4491 11169
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 10134 11160 10140 11212
rect 10192 11200 10198 11212
rect 11348 11209 11376 11240
rect 11790 11228 11796 11240
rect 11848 11228 11854 11280
rect 11882 11228 11888 11280
rect 11940 11268 11946 11280
rect 14568 11268 14596 11299
rect 14826 11296 14832 11348
rect 14884 11336 14890 11348
rect 16117 11339 16175 11345
rect 16117 11336 16129 11339
rect 14884 11308 16129 11336
rect 14884 11296 14890 11308
rect 16117 11305 16129 11308
rect 16163 11305 16175 11339
rect 16117 11299 16175 11305
rect 16577 11339 16635 11345
rect 16577 11305 16589 11339
rect 16623 11336 16635 11339
rect 16758 11336 16764 11348
rect 16623 11308 16764 11336
rect 16623 11305 16635 11308
rect 16577 11299 16635 11305
rect 16758 11296 16764 11308
rect 16816 11296 16822 11348
rect 11940 11240 12848 11268
rect 14568 11240 15792 11268
rect 11940 11228 11946 11240
rect 10689 11203 10747 11209
rect 10689 11200 10701 11203
rect 10192 11172 10701 11200
rect 10192 11160 10198 11172
rect 10689 11169 10701 11172
rect 10735 11169 10747 11203
rect 10689 11163 10747 11169
rect 10781 11203 10839 11209
rect 10781 11169 10793 11203
rect 10827 11169 10839 11203
rect 10781 11163 10839 11169
rect 11333 11203 11391 11209
rect 11333 11169 11345 11203
rect 11379 11169 11391 11203
rect 11333 11163 11391 11169
rect 1489 11135 1547 11141
rect 1489 11101 1501 11135
rect 1535 11132 1547 11135
rect 1946 11132 1952 11144
rect 1535 11104 1952 11132
rect 1535 11101 1547 11104
rect 1489 11095 1547 11101
rect 1946 11092 1952 11104
rect 2004 11132 2010 11144
rect 4157 11135 4215 11141
rect 4157 11132 4169 11135
rect 2004 11104 4169 11132
rect 2004 11092 2010 11104
rect 4080 11008 4108 11104
rect 4157 11101 4169 11104
rect 4203 11101 4215 11135
rect 4157 11095 4215 11101
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 10796 11132 10824 11163
rect 11974 11160 11980 11212
rect 12032 11200 12038 11212
rect 12820 11209 12848 11240
rect 12437 11203 12495 11209
rect 12437 11200 12449 11203
rect 12032 11172 12449 11200
rect 12032 11160 12038 11172
rect 12437 11169 12449 11172
rect 12483 11169 12495 11203
rect 12437 11163 12495 11169
rect 12805 11203 12863 11209
rect 12805 11169 12817 11203
rect 12851 11169 12863 11203
rect 12805 11163 12863 11169
rect 13173 11203 13231 11209
rect 13173 11169 13185 11203
rect 13219 11169 13231 11203
rect 13173 11163 13231 11169
rect 9732 11104 10824 11132
rect 9732 11092 9738 11104
rect 7098 11024 7104 11076
rect 7156 11064 7162 11076
rect 7193 11067 7251 11073
rect 7193 11064 7205 11067
rect 7156 11036 7205 11064
rect 7156 11024 7162 11036
rect 7193 11033 7205 11036
rect 7239 11064 7251 11067
rect 7561 11067 7619 11073
rect 7561 11064 7573 11067
rect 7239 11036 7573 11064
rect 7239 11033 7251 11036
rect 7193 11027 7251 11033
rect 7561 11033 7573 11036
rect 7607 11064 7619 11067
rect 9585 11067 9643 11073
rect 9585 11064 9597 11067
rect 7607 11036 9597 11064
rect 7607 11033 7619 11036
rect 7561 11027 7619 11033
rect 9585 11033 9597 11036
rect 9631 11033 9643 11067
rect 9585 11027 9643 11033
rect 3053 10999 3111 11005
rect 3053 10965 3065 10999
rect 3099 10996 3111 10999
rect 3786 10996 3792 11008
rect 3099 10968 3792 10996
rect 3099 10965 3111 10968
rect 3053 10959 3111 10965
rect 3786 10956 3792 10968
rect 3844 10956 3850 11008
rect 4062 10996 4068 11008
rect 4023 10968 4068 10996
rect 4062 10956 4068 10968
rect 4120 10956 4126 11008
rect 9600 10996 9628 11027
rect 10042 11024 10048 11076
rect 10100 11064 10106 11076
rect 10796 11064 10824 11104
rect 11238 11092 11244 11144
rect 11296 11132 11302 11144
rect 11422 11132 11428 11144
rect 11296 11104 11428 11132
rect 11296 11092 11302 11104
rect 11422 11092 11428 11104
rect 11480 11092 11486 11144
rect 12066 11092 12072 11144
rect 12124 11132 12130 11144
rect 12710 11132 12716 11144
rect 12124 11104 12716 11132
rect 12124 11092 12130 11104
rect 12710 11092 12716 11104
rect 12768 11132 12774 11144
rect 13188 11132 13216 11163
rect 13538 11160 13544 11212
rect 13596 11200 13602 11212
rect 13817 11203 13875 11209
rect 13817 11200 13829 11203
rect 13596 11172 13829 11200
rect 13596 11160 13602 11172
rect 13817 11169 13829 11172
rect 13863 11169 13875 11203
rect 13817 11163 13875 11169
rect 14921 11203 14979 11209
rect 14921 11169 14933 11203
rect 14967 11200 14979 11203
rect 15286 11200 15292 11212
rect 14967 11172 15292 11200
rect 14967 11169 14979 11172
rect 14921 11163 14979 11169
rect 15286 11160 15292 11172
rect 15344 11200 15350 11212
rect 15764 11209 15792 11240
rect 15657 11203 15715 11209
rect 15657 11200 15669 11203
rect 15344 11172 15516 11200
rect 15344 11160 15350 11172
rect 15488 11144 15516 11172
rect 15580 11172 15669 11200
rect 14182 11132 14188 11144
rect 12768 11104 13216 11132
rect 14143 11104 14188 11132
rect 12768 11092 12774 11104
rect 14182 11092 14188 11104
rect 14240 11132 14246 11144
rect 14829 11135 14887 11141
rect 14829 11132 14841 11135
rect 14240 11104 14841 11132
rect 14240 11092 14246 11104
rect 14829 11101 14841 11104
rect 14875 11101 14887 11135
rect 14829 11095 14887 11101
rect 15470 11092 15476 11144
rect 15528 11092 15534 11144
rect 11330 11064 11336 11076
rect 10100 11036 10732 11064
rect 10796 11036 11336 11064
rect 10100 11024 10106 11036
rect 9766 10996 9772 11008
rect 9600 10968 9772 10996
rect 9766 10956 9772 10968
rect 9824 10956 9830 11008
rect 10134 10996 10140 11008
rect 10095 10968 10140 10996
rect 10134 10956 10140 10968
rect 10192 10956 10198 11008
rect 10704 10996 10732 11036
rect 11330 11024 11336 11036
rect 11388 11024 11394 11076
rect 12268 11036 14872 11064
rect 12268 10996 12296 11036
rect 10704 10968 12296 10996
rect 13633 10999 13691 11005
rect 13633 10965 13645 10999
rect 13679 10996 13691 10999
rect 13722 10996 13728 11008
rect 13679 10968 13728 10996
rect 13679 10965 13691 10968
rect 13633 10959 13691 10965
rect 13722 10956 13728 10968
rect 13780 10956 13786 11008
rect 14844 10996 14872 11036
rect 15580 10996 15608 11172
rect 15657 11169 15669 11172
rect 15703 11169 15715 11203
rect 15657 11163 15715 11169
rect 15749 11203 15807 11209
rect 15749 11169 15761 11203
rect 15795 11169 15807 11203
rect 15749 11163 15807 11169
rect 16390 10996 16396 11008
rect 14844 10968 16396 10996
rect 16390 10956 16396 10968
rect 16448 10956 16454 11008
rect 1104 10906 18860 10928
rect 1104 10854 4315 10906
rect 4367 10854 4379 10906
rect 4431 10854 4443 10906
rect 4495 10854 4507 10906
rect 4559 10854 10982 10906
rect 11034 10854 11046 10906
rect 11098 10854 11110 10906
rect 11162 10854 11174 10906
rect 11226 10854 17648 10906
rect 17700 10854 17712 10906
rect 17764 10854 17776 10906
rect 17828 10854 17840 10906
rect 17892 10854 18860 10906
rect 1104 10832 18860 10854
rect 3326 10792 3332 10804
rect 3287 10764 3332 10792
rect 3326 10752 3332 10764
rect 3384 10752 3390 10804
rect 3786 10792 3792 10804
rect 3747 10764 3792 10792
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 5905 10795 5963 10801
rect 5905 10761 5917 10795
rect 5951 10792 5963 10795
rect 6914 10792 6920 10804
rect 5951 10764 6920 10792
rect 5951 10761 5963 10764
rect 5905 10755 5963 10761
rect 6914 10752 6920 10764
rect 6972 10752 6978 10804
rect 9125 10795 9183 10801
rect 9125 10761 9137 10795
rect 9171 10792 9183 10795
rect 9674 10792 9680 10804
rect 9171 10764 9680 10792
rect 9171 10761 9183 10764
rect 9125 10755 9183 10761
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 11609 10795 11667 10801
rect 11609 10761 11621 10795
rect 11655 10792 11667 10795
rect 11882 10792 11888 10804
rect 11655 10764 11888 10792
rect 11655 10761 11667 10764
rect 11609 10755 11667 10761
rect 11882 10752 11888 10764
rect 11940 10792 11946 10804
rect 12069 10795 12127 10801
rect 12069 10792 12081 10795
rect 11940 10764 12081 10792
rect 11940 10752 11946 10764
rect 12069 10761 12081 10764
rect 12115 10761 12127 10795
rect 12069 10755 12127 10761
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 12529 10795 12587 10801
rect 12529 10792 12541 10795
rect 12492 10764 12541 10792
rect 12492 10752 12498 10764
rect 12529 10761 12541 10764
rect 12575 10792 12587 10795
rect 13538 10792 13544 10804
rect 12575 10764 13544 10792
rect 12575 10761 12587 10764
rect 12529 10755 12587 10761
rect 13538 10752 13544 10764
rect 13596 10752 13602 10804
rect 14734 10792 14740 10804
rect 14695 10764 14740 10792
rect 14734 10752 14740 10764
rect 14792 10752 14798 10804
rect 16574 10724 16580 10736
rect 16535 10696 16580 10724
rect 16574 10684 16580 10696
rect 16632 10684 16638 10736
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 2038 10656 2044 10668
rect 1719 10628 2044 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 2038 10616 2044 10628
rect 2096 10656 2102 10668
rect 2406 10656 2412 10668
rect 2096 10628 2412 10656
rect 2096 10616 2102 10628
rect 2406 10616 2412 10628
rect 2464 10616 2470 10668
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 4246 10656 4252 10668
rect 3099 10628 4252 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 4246 10616 4252 10628
rect 4304 10656 4310 10668
rect 4617 10659 4675 10665
rect 4617 10656 4629 10659
rect 4304 10628 4629 10656
rect 4304 10616 4310 10628
rect 4617 10625 4629 10628
rect 4663 10625 4675 10659
rect 8754 10656 8760 10668
rect 8715 10628 8760 10656
rect 4617 10619 4675 10625
rect 8754 10616 8760 10628
rect 8812 10616 8818 10668
rect 13906 10656 13912 10668
rect 13867 10628 13912 10656
rect 13906 10616 13912 10628
rect 13964 10616 13970 10668
rect 15565 10659 15623 10665
rect 15565 10625 15577 10659
rect 15611 10656 15623 10659
rect 15841 10659 15899 10665
rect 15841 10656 15853 10659
rect 15611 10628 15853 10656
rect 15611 10625 15623 10628
rect 15565 10619 15623 10625
rect 15841 10625 15853 10628
rect 15887 10656 15899 10659
rect 16206 10656 16212 10668
rect 15887 10628 16212 10656
rect 15887 10625 15899 10628
rect 15841 10619 15899 10625
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 1486 10588 1492 10600
rect 1443 10560 1492 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 1486 10548 1492 10560
rect 1544 10548 1550 10600
rect 4062 10548 4068 10600
rect 4120 10588 4126 10600
rect 4341 10591 4399 10597
rect 4341 10588 4353 10591
rect 4120 10560 4353 10588
rect 4120 10548 4126 10560
rect 4341 10557 4353 10560
rect 4387 10588 4399 10591
rect 4430 10588 4436 10600
rect 4387 10560 4436 10588
rect 4387 10557 4399 10560
rect 4341 10551 4399 10557
rect 4430 10548 4436 10560
rect 4488 10548 4494 10600
rect 8018 10588 8024 10600
rect 7979 10560 8024 10588
rect 8018 10548 8024 10560
rect 8076 10548 8082 10600
rect 8110 10548 8116 10600
rect 8168 10588 8174 10600
rect 8386 10597 8392 10600
rect 8205 10591 8263 10597
rect 8205 10588 8217 10591
rect 8168 10560 8217 10588
rect 8168 10548 8174 10560
rect 8205 10557 8217 10560
rect 8251 10557 8263 10591
rect 8205 10551 8263 10557
rect 8338 10591 8392 10597
rect 8338 10557 8350 10591
rect 8384 10557 8392 10591
rect 8338 10551 8392 10557
rect 8386 10548 8392 10551
rect 8444 10548 8450 10600
rect 9674 10588 9680 10600
rect 9635 10560 9680 10588
rect 9674 10548 9680 10560
rect 9732 10548 9738 10600
rect 9953 10591 10011 10597
rect 9953 10588 9965 10591
rect 9784 10560 9965 10588
rect 7561 10523 7619 10529
rect 7561 10489 7573 10523
rect 7607 10520 7619 10523
rect 8404 10520 8432 10548
rect 9398 10520 9404 10532
rect 7607 10492 8432 10520
rect 9359 10492 9404 10520
rect 7607 10489 7619 10492
rect 7561 10483 7619 10489
rect 9398 10480 9404 10492
rect 9456 10520 9462 10532
rect 9784 10520 9812 10560
rect 9953 10557 9965 10560
rect 9999 10557 10011 10591
rect 9953 10551 10011 10557
rect 11333 10591 11391 10597
rect 11333 10557 11345 10591
rect 11379 10588 11391 10591
rect 11606 10588 11612 10600
rect 11379 10560 11612 10588
rect 11379 10557 11391 10560
rect 11333 10551 11391 10557
rect 11606 10548 11612 10560
rect 11664 10548 11670 10600
rect 13173 10591 13231 10597
rect 13173 10557 13185 10591
rect 13219 10588 13231 10591
rect 13262 10588 13268 10600
rect 13219 10560 13268 10588
rect 13219 10557 13231 10560
rect 13173 10551 13231 10557
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 13541 10591 13599 10597
rect 13541 10557 13553 10591
rect 13587 10557 13599 10591
rect 13814 10588 13820 10600
rect 13775 10560 13820 10588
rect 13541 10551 13599 10557
rect 9456 10492 9812 10520
rect 13556 10520 13584 10551
rect 13814 10548 13820 10560
rect 13872 10548 13878 10600
rect 14090 10548 14096 10600
rect 14148 10588 14154 10600
rect 14185 10591 14243 10597
rect 14185 10588 14197 10591
rect 14148 10560 14197 10588
rect 14148 10548 14154 10560
rect 14185 10557 14197 10560
rect 14231 10557 14243 10591
rect 15930 10588 15936 10600
rect 14185 10551 14243 10557
rect 15028 10560 15936 10588
rect 13722 10520 13728 10532
rect 13556 10492 13728 10520
rect 9456 10480 9462 10492
rect 13722 10480 13728 10492
rect 13780 10480 13786 10532
rect 7929 10455 7987 10461
rect 7929 10421 7941 10455
rect 7975 10452 7987 10455
rect 8018 10452 8024 10464
rect 7975 10424 8024 10452
rect 7975 10421 7987 10424
rect 7929 10415 7987 10421
rect 8018 10412 8024 10424
rect 8076 10412 8082 10464
rect 14918 10412 14924 10464
rect 14976 10452 14982 10464
rect 15028 10461 15056 10560
rect 15930 10548 15936 10560
rect 15988 10588 15994 10600
rect 16025 10591 16083 10597
rect 16025 10588 16037 10591
rect 15988 10560 16037 10588
rect 15988 10548 15994 10560
rect 16025 10557 16037 10560
rect 16071 10557 16083 10591
rect 16025 10551 16083 10557
rect 16298 10548 16304 10600
rect 16356 10588 16362 10600
rect 16485 10591 16543 10597
rect 16485 10588 16497 10591
rect 16356 10560 16497 10588
rect 16356 10548 16362 10560
rect 16485 10557 16497 10560
rect 16531 10557 16543 10591
rect 16485 10551 16543 10557
rect 15013 10455 15071 10461
rect 15013 10452 15025 10455
rect 14976 10424 15025 10452
rect 14976 10412 14982 10424
rect 15013 10421 15025 10424
rect 15059 10421 15071 10455
rect 15013 10415 15071 10421
rect 1104 10362 18860 10384
rect 1104 10310 7648 10362
rect 7700 10310 7712 10362
rect 7764 10310 7776 10362
rect 7828 10310 7840 10362
rect 7892 10310 14315 10362
rect 14367 10310 14379 10362
rect 14431 10310 14443 10362
rect 14495 10310 14507 10362
rect 14559 10310 18860 10362
rect 1104 10288 18860 10310
rect 4246 10208 4252 10260
rect 4304 10248 4310 10260
rect 4341 10251 4399 10257
rect 4341 10248 4353 10251
rect 4304 10220 4353 10248
rect 4304 10208 4310 10220
rect 4341 10217 4353 10220
rect 4387 10217 4399 10251
rect 11330 10248 11336 10260
rect 11291 10220 11336 10248
rect 4341 10211 4399 10217
rect 11330 10208 11336 10220
rect 11388 10248 11394 10260
rect 11514 10248 11520 10260
rect 11388 10220 11520 10248
rect 11388 10208 11394 10220
rect 11514 10208 11520 10220
rect 11572 10208 11578 10260
rect 12250 10248 12256 10260
rect 12211 10220 12256 10248
rect 12250 10208 12256 10220
rect 12308 10208 12314 10260
rect 12710 10248 12716 10260
rect 12671 10220 12716 10248
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 14829 10251 14887 10257
rect 14829 10248 14841 10251
rect 13872 10220 14841 10248
rect 13872 10208 13878 10220
rect 14829 10217 14841 10220
rect 14875 10217 14887 10251
rect 16390 10248 16396 10260
rect 16351 10220 16396 10248
rect 14829 10211 14887 10217
rect 16390 10208 16396 10220
rect 16448 10208 16454 10260
rect 16574 10208 16580 10260
rect 16632 10248 16638 10260
rect 16761 10251 16819 10257
rect 16761 10248 16773 10251
rect 16632 10220 16773 10248
rect 16632 10208 16638 10220
rect 16761 10217 16773 10220
rect 16807 10217 16819 10251
rect 16761 10211 16819 10217
rect 3142 10180 3148 10192
rect 3103 10152 3148 10180
rect 3142 10140 3148 10152
rect 3200 10140 3206 10192
rect 4065 10183 4123 10189
rect 4065 10149 4077 10183
rect 4111 10180 4123 10183
rect 4430 10180 4436 10192
rect 4111 10152 4436 10180
rect 4111 10149 4123 10152
rect 4065 10143 4123 10149
rect 4430 10140 4436 10152
rect 4488 10180 4494 10192
rect 4709 10183 4767 10189
rect 4709 10180 4721 10183
rect 4488 10152 4721 10180
rect 4488 10140 4494 10152
rect 4709 10149 4721 10152
rect 4755 10149 4767 10183
rect 4709 10143 4767 10149
rect 7929 10183 7987 10189
rect 7929 10149 7941 10183
rect 7975 10180 7987 10183
rect 8110 10180 8116 10192
rect 7975 10152 8116 10180
rect 7975 10149 7987 10152
rect 7929 10143 7987 10149
rect 8110 10140 8116 10152
rect 8168 10140 8174 10192
rect 8478 10180 8484 10192
rect 8439 10152 8484 10180
rect 8478 10140 8484 10152
rect 8536 10140 8542 10192
rect 13354 10140 13360 10192
rect 13412 10180 13418 10192
rect 16206 10180 16212 10192
rect 13412 10152 14504 10180
rect 13412 10140 13418 10152
rect 1210 10072 1216 10124
rect 1268 10112 1274 10124
rect 1765 10115 1823 10121
rect 1765 10112 1777 10115
rect 1268 10084 1777 10112
rect 1268 10072 1274 10084
rect 1765 10081 1777 10084
rect 1811 10112 1823 10115
rect 2222 10112 2228 10124
rect 1811 10084 2228 10112
rect 1811 10081 1823 10084
rect 1765 10075 1823 10081
rect 2222 10072 2228 10084
rect 2280 10072 2286 10124
rect 8021 10115 8079 10121
rect 8021 10081 8033 10115
rect 8067 10112 8079 10115
rect 8202 10112 8208 10124
rect 8067 10084 8208 10112
rect 8067 10081 8079 10084
rect 8021 10075 8079 10081
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 9582 10112 9588 10124
rect 9543 10084 9588 10112
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 12158 10072 12164 10124
rect 12216 10112 12222 10124
rect 12894 10112 12900 10124
rect 12216 10084 12900 10112
rect 12216 10072 12222 10084
rect 12894 10072 12900 10084
rect 12952 10072 12958 10124
rect 13998 10112 14004 10124
rect 13959 10084 14004 10112
rect 13998 10072 14004 10084
rect 14056 10072 14062 10124
rect 14476 10121 14504 10152
rect 15304 10152 16212 10180
rect 15304 10124 15332 10152
rect 16206 10140 16212 10152
rect 16264 10140 16270 10192
rect 14461 10115 14519 10121
rect 14461 10081 14473 10115
rect 14507 10112 14519 10115
rect 15010 10112 15016 10124
rect 14507 10084 15016 10112
rect 14507 10081 14519 10084
rect 14461 10075 14519 10081
rect 15010 10072 15016 10084
rect 15068 10072 15074 10124
rect 15286 10112 15292 10124
rect 15199 10084 15292 10112
rect 15286 10072 15292 10084
rect 15344 10072 15350 10124
rect 15565 10115 15623 10121
rect 15565 10081 15577 10115
rect 15611 10112 15623 10115
rect 15838 10112 15844 10124
rect 15611 10084 15844 10112
rect 15611 10081 15623 10084
rect 15565 10075 15623 10081
rect 1486 10044 1492 10056
rect 1447 10016 1492 10044
rect 1486 10004 1492 10016
rect 1544 10004 1550 10056
rect 9309 10047 9367 10053
rect 9309 10013 9321 10047
rect 9355 10044 9367 10047
rect 9490 10044 9496 10056
rect 9355 10016 9496 10044
rect 9355 10013 9367 10016
rect 9309 10007 9367 10013
rect 9490 10004 9496 10016
rect 9548 10004 9554 10056
rect 14734 10004 14740 10056
rect 14792 10044 14798 10056
rect 15580 10044 15608 10075
rect 15838 10072 15844 10084
rect 15896 10072 15902 10124
rect 14792 10016 15608 10044
rect 14792 10004 14798 10016
rect 14090 9976 14096 9988
rect 13372 9948 14096 9976
rect 7745 9911 7803 9917
rect 7745 9877 7757 9911
rect 7791 9908 7803 9911
rect 7834 9908 7840 9920
rect 7791 9880 7840 9908
rect 7791 9877 7803 9880
rect 7745 9871 7803 9877
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 10870 9908 10876 9920
rect 10831 9880 10876 9908
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 11882 9908 11888 9920
rect 11843 9880 11888 9908
rect 11882 9868 11888 9880
rect 11940 9868 11946 9920
rect 12710 9868 12716 9920
rect 12768 9908 12774 9920
rect 13372 9917 13400 9948
rect 14090 9936 14096 9948
rect 14148 9936 14154 9988
rect 13081 9911 13139 9917
rect 13081 9908 13093 9911
rect 12768 9880 13093 9908
rect 12768 9868 12774 9880
rect 13081 9877 13093 9880
rect 13127 9908 13139 9911
rect 13357 9911 13415 9917
rect 13357 9908 13369 9911
rect 13127 9880 13369 9908
rect 13127 9877 13139 9880
rect 13081 9871 13139 9877
rect 13357 9877 13369 9880
rect 13403 9877 13415 9911
rect 13814 9908 13820 9920
rect 13775 9880 13820 9908
rect 13357 9871 13415 9877
rect 13814 9868 13820 9880
rect 13872 9868 13878 9920
rect 15194 9868 15200 9920
rect 15252 9908 15258 9920
rect 16025 9911 16083 9917
rect 16025 9908 16037 9911
rect 15252 9880 16037 9908
rect 15252 9868 15258 9880
rect 16025 9877 16037 9880
rect 16071 9908 16083 9911
rect 16298 9908 16304 9920
rect 16071 9880 16304 9908
rect 16071 9877 16083 9880
rect 16025 9871 16083 9877
rect 16298 9868 16304 9880
rect 16356 9868 16362 9920
rect 1104 9818 18860 9840
rect 1104 9766 4315 9818
rect 4367 9766 4379 9818
rect 4431 9766 4443 9818
rect 4495 9766 4507 9818
rect 4559 9766 10982 9818
rect 11034 9766 11046 9818
rect 11098 9766 11110 9818
rect 11162 9766 11174 9818
rect 11226 9766 17648 9818
rect 17700 9766 17712 9818
rect 17764 9766 17776 9818
rect 17828 9766 17840 9818
rect 17892 9766 18860 9818
rect 1104 9744 18860 9766
rect 2038 9704 2044 9716
rect 1999 9676 2044 9704
rect 2038 9664 2044 9676
rect 2096 9664 2102 9716
rect 2222 9664 2228 9716
rect 2280 9704 2286 9716
rect 2317 9707 2375 9713
rect 2317 9704 2329 9707
rect 2280 9676 2329 9704
rect 2280 9664 2286 9676
rect 2317 9673 2329 9676
rect 2363 9673 2375 9707
rect 8110 9704 8116 9716
rect 8071 9676 8116 9704
rect 2317 9667 2375 9673
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 8386 9664 8392 9716
rect 8444 9704 8450 9716
rect 11241 9707 11299 9713
rect 11241 9704 11253 9707
rect 8444 9676 11253 9704
rect 8444 9664 8450 9676
rect 11241 9673 11253 9676
rect 11287 9673 11299 9707
rect 11241 9667 11299 9673
rect 11422 9664 11428 9716
rect 11480 9704 11486 9716
rect 11974 9704 11980 9716
rect 11480 9676 11980 9704
rect 11480 9664 11486 9676
rect 11974 9664 11980 9676
rect 12032 9664 12038 9716
rect 12894 9704 12900 9716
rect 12855 9676 12900 9704
rect 12894 9664 12900 9676
rect 12952 9704 12958 9716
rect 13265 9707 13323 9713
rect 13265 9704 13277 9707
rect 12952 9676 13277 9704
rect 12952 9664 12958 9676
rect 13265 9673 13277 9676
rect 13311 9704 13323 9707
rect 13449 9707 13507 9713
rect 13449 9704 13461 9707
rect 13311 9676 13461 9704
rect 13311 9673 13323 9676
rect 13265 9667 13323 9673
rect 13449 9673 13461 9676
rect 13495 9673 13507 9707
rect 15286 9704 15292 9716
rect 13449 9667 13507 9673
rect 15120 9676 15292 9704
rect 1673 9639 1731 9645
rect 1673 9605 1685 9639
rect 1719 9636 1731 9639
rect 1762 9636 1768 9648
rect 1719 9608 1768 9636
rect 1719 9605 1731 9608
rect 1673 9599 1731 9605
rect 1762 9596 1768 9608
rect 1820 9596 1826 9648
rect 9401 9639 9459 9645
rect 9401 9605 9413 9639
rect 9447 9636 9459 9639
rect 9582 9636 9588 9648
rect 9447 9608 9588 9636
rect 9447 9605 9459 9608
rect 9401 9599 9459 9605
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 11330 9596 11336 9648
rect 11388 9636 11394 9648
rect 12434 9636 12440 9648
rect 11388 9608 12440 9636
rect 11388 9596 11394 9608
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 14553 9639 14611 9645
rect 14553 9605 14565 9639
rect 14599 9636 14611 9639
rect 15120 9636 15148 9676
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 14599 9608 15148 9636
rect 14599 9605 14611 9608
rect 14553 9599 14611 9605
rect 15562 9596 15568 9648
rect 15620 9636 15626 9648
rect 16577 9639 16635 9645
rect 16577 9636 16589 9639
rect 15620 9608 16589 9636
rect 15620 9596 15626 9608
rect 16577 9605 16589 9608
rect 16623 9636 16635 9639
rect 17034 9636 17040 9648
rect 16623 9608 17040 9636
rect 16623 9605 16635 9608
rect 16577 9599 16635 9605
rect 17034 9596 17040 9608
rect 17092 9636 17098 9648
rect 17092 9608 17724 9636
rect 17092 9596 17098 9608
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9568 9091 9571
rect 9490 9568 9496 9580
rect 9079 9540 9496 9568
rect 9079 9537 9091 9540
rect 9033 9531 9091 9537
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 10689 9571 10747 9577
rect 10689 9537 10701 9571
rect 10735 9568 10747 9571
rect 10735 9540 12204 9568
rect 10735 9537 10747 9540
rect 10689 9531 10747 9537
rect 7834 9500 7840 9512
rect 7795 9472 7840 9500
rect 7834 9460 7840 9472
rect 7892 9460 7898 9512
rect 11422 9500 11428 9512
rect 11383 9472 11428 9500
rect 11422 9460 11428 9472
rect 11480 9460 11486 9512
rect 11514 9460 11520 9512
rect 11572 9500 11578 9512
rect 12176 9509 12204 9540
rect 12161 9503 12219 9509
rect 11572 9472 11617 9500
rect 11572 9460 11578 9472
rect 12161 9469 12173 9503
rect 12207 9500 12219 9503
rect 12342 9500 12348 9512
rect 12207 9472 12348 9500
rect 12207 9469 12219 9472
rect 12161 9463 12219 9469
rect 12342 9460 12348 9472
rect 12400 9460 12406 9512
rect 12452 9509 12480 9596
rect 14185 9571 14243 9577
rect 14185 9537 14197 9571
rect 14231 9568 14243 9571
rect 15102 9568 15108 9580
rect 14231 9540 15108 9568
rect 14231 9537 14243 9540
rect 14185 9531 14243 9537
rect 15102 9528 15108 9540
rect 15160 9528 15166 9580
rect 16298 9528 16304 9580
rect 16356 9568 16362 9580
rect 17696 9577 17724 9608
rect 17681 9571 17739 9577
rect 16356 9540 17632 9568
rect 16356 9528 16362 9540
rect 12437 9503 12495 9509
rect 12437 9469 12449 9503
rect 12483 9469 12495 9503
rect 12437 9463 12495 9469
rect 13262 9460 13268 9512
rect 13320 9500 13326 9512
rect 13725 9503 13783 9509
rect 13725 9500 13737 9503
rect 13320 9472 13737 9500
rect 13320 9460 13326 9472
rect 13725 9469 13737 9472
rect 13771 9500 13783 9503
rect 14090 9500 14096 9512
rect 13771 9472 14096 9500
rect 13771 9469 13783 9472
rect 13725 9463 13783 9469
rect 14090 9460 14096 9472
rect 14148 9460 14154 9512
rect 14734 9460 14740 9512
rect 14792 9500 14798 9512
rect 14829 9503 14887 9509
rect 14829 9500 14841 9503
rect 14792 9472 14841 9500
rect 14792 9460 14798 9472
rect 14829 9469 14841 9472
rect 14875 9469 14887 9503
rect 14829 9463 14887 9469
rect 15010 9460 15016 9512
rect 15068 9500 15074 9512
rect 15473 9503 15531 9509
rect 15473 9500 15485 9503
rect 15068 9472 15485 9500
rect 15068 9460 15074 9472
rect 15473 9469 15485 9472
rect 15519 9469 15531 9503
rect 15473 9463 15531 9469
rect 16574 9460 16580 9512
rect 16632 9500 16638 9512
rect 17604 9509 17632 9540
rect 17681 9537 17693 9571
rect 17727 9537 17739 9571
rect 17681 9531 17739 9537
rect 17221 9503 17279 9509
rect 17221 9500 17233 9503
rect 16632 9472 17233 9500
rect 16632 9460 16638 9472
rect 17221 9469 17233 9472
rect 17267 9469 17279 9503
rect 17221 9463 17279 9469
rect 17589 9503 17647 9509
rect 17589 9469 17601 9503
rect 17635 9469 17647 9503
rect 17589 9463 17647 9469
rect 13633 9435 13691 9441
rect 13633 9401 13645 9435
rect 13679 9432 13691 9435
rect 13814 9432 13820 9444
rect 13679 9404 13820 9432
rect 13679 9401 13691 9404
rect 13633 9395 13691 9401
rect 13814 9392 13820 9404
rect 13872 9392 13878 9444
rect 15194 9392 15200 9444
rect 15252 9432 15258 9444
rect 15841 9435 15899 9441
rect 15841 9432 15853 9435
rect 15252 9404 15853 9432
rect 15252 9392 15258 9404
rect 15841 9401 15853 9404
rect 15887 9432 15899 9435
rect 16390 9432 16396 9444
rect 15887 9404 16396 9432
rect 15887 9401 15899 9404
rect 15841 9395 15899 9401
rect 16390 9392 16396 9404
rect 16448 9392 16454 9444
rect 16666 9392 16672 9444
rect 16724 9432 16730 9444
rect 16761 9435 16819 9441
rect 16761 9432 16773 9435
rect 16724 9404 16773 9432
rect 16724 9392 16730 9404
rect 16761 9401 16773 9404
rect 16807 9401 16819 9435
rect 16761 9395 16819 9401
rect 8202 9324 8208 9376
rect 8260 9364 8266 9376
rect 8570 9364 8576 9376
rect 8260 9336 8576 9364
rect 8260 9324 8266 9336
rect 8570 9324 8576 9336
rect 8628 9324 8634 9376
rect 10042 9364 10048 9376
rect 10003 9336 10048 9364
rect 10042 9324 10048 9336
rect 10100 9324 10106 9376
rect 11057 9367 11115 9373
rect 11057 9333 11069 9367
rect 11103 9364 11115 9367
rect 11330 9364 11336 9376
rect 11103 9336 11336 9364
rect 11103 9333 11115 9336
rect 11057 9327 11115 9333
rect 11330 9324 11336 9336
rect 11388 9324 11394 9376
rect 16298 9364 16304 9376
rect 16259 9336 16304 9364
rect 16298 9324 16304 9336
rect 16356 9324 16362 9376
rect 1104 9274 18860 9296
rect 1104 9222 7648 9274
rect 7700 9222 7712 9274
rect 7764 9222 7776 9274
rect 7828 9222 7840 9274
rect 7892 9222 14315 9274
rect 14367 9222 14379 9274
rect 14431 9222 14443 9274
rect 14495 9222 14507 9274
rect 14559 9222 18860 9274
rect 1104 9200 18860 9222
rect 1486 9120 1492 9172
rect 1544 9160 1550 9172
rect 1581 9163 1639 9169
rect 1581 9160 1593 9163
rect 1544 9132 1593 9160
rect 1544 9120 1550 9132
rect 1581 9129 1593 9132
rect 1627 9160 1639 9163
rect 1670 9160 1676 9172
rect 1627 9132 1676 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 1946 9160 1952 9172
rect 1907 9132 1952 9160
rect 1946 9120 1952 9132
rect 2004 9120 2010 9172
rect 11422 9120 11428 9172
rect 11480 9160 11486 9172
rect 11793 9163 11851 9169
rect 11793 9160 11805 9163
rect 11480 9132 11805 9160
rect 11480 9120 11486 9132
rect 11793 9129 11805 9132
rect 11839 9129 11851 9163
rect 13814 9160 13820 9172
rect 13775 9132 13820 9160
rect 11793 9123 11851 9129
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 14090 9120 14096 9172
rect 14148 9160 14154 9172
rect 14185 9163 14243 9169
rect 14185 9160 14197 9163
rect 14148 9132 14197 9160
rect 14148 9120 14154 9132
rect 14185 9129 14197 9132
rect 14231 9129 14243 9163
rect 14185 9123 14243 9129
rect 11146 9092 11152 9104
rect 11107 9064 11152 9092
rect 11146 9052 11152 9064
rect 11204 9052 11210 9104
rect 11517 9095 11575 9101
rect 11517 9061 11529 9095
rect 11563 9092 11575 9095
rect 12342 9092 12348 9104
rect 11563 9064 12348 9092
rect 11563 9061 11575 9064
rect 11517 9055 11575 9061
rect 12342 9052 12348 9064
rect 12400 9052 12406 9104
rect 15657 9095 15715 9101
rect 15657 9092 15669 9095
rect 14844 9064 15669 9092
rect 9490 9024 9496 9036
rect 9451 8996 9496 9024
rect 9490 8984 9496 8996
rect 9548 8984 9554 9036
rect 9766 9024 9772 9036
rect 9727 8996 9772 9024
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 12618 9024 12624 9036
rect 12579 8996 12624 9024
rect 12618 8984 12624 8996
rect 12676 8984 12682 9036
rect 12986 9024 12992 9036
rect 12947 8996 12992 9024
rect 12986 8984 12992 8996
rect 13044 8984 13050 9036
rect 13262 9024 13268 9036
rect 13223 8996 13268 9024
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 13906 8984 13912 9036
rect 13964 9024 13970 9036
rect 14844 9033 14872 9064
rect 15657 9061 15669 9064
rect 15703 9061 15715 9095
rect 16206 9092 16212 9104
rect 16167 9064 16212 9092
rect 15657 9055 15715 9061
rect 16206 9052 16212 9064
rect 16264 9052 16270 9104
rect 14829 9027 14887 9033
rect 14829 9024 14841 9027
rect 13964 8996 14841 9024
rect 13964 8984 13970 8996
rect 14829 8993 14841 8996
rect 14875 8993 14887 9027
rect 15194 9024 15200 9036
rect 15155 8996 15200 9024
rect 14829 8987 14887 8993
rect 15194 8984 15200 8996
rect 15252 8984 15258 9036
rect 16298 9024 16304 9036
rect 16259 8996 16304 9024
rect 16298 8984 16304 8996
rect 16356 8984 16362 9036
rect 15102 8916 15108 8968
rect 15160 8956 15166 8968
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 15160 8928 15301 8956
rect 15160 8916 15166 8928
rect 15289 8925 15301 8928
rect 15335 8956 15347 8959
rect 15654 8956 15660 8968
rect 15335 8928 15660 8956
rect 15335 8925 15347 8928
rect 15289 8919 15347 8925
rect 15654 8916 15660 8928
rect 15712 8916 15718 8968
rect 13170 8848 13176 8900
rect 13228 8888 13234 8900
rect 13265 8891 13323 8897
rect 13265 8888 13277 8891
rect 13228 8860 13277 8888
rect 13228 8848 13234 8860
rect 13265 8857 13277 8860
rect 13311 8857 13323 8891
rect 13265 8851 13323 8857
rect 14645 8891 14703 8897
rect 14645 8857 14657 8891
rect 14691 8888 14703 8891
rect 15194 8888 15200 8900
rect 14691 8860 15200 8888
rect 14691 8857 14703 8860
rect 14645 8851 14703 8857
rect 15194 8848 15200 8860
rect 15252 8848 15258 8900
rect 15838 8780 15844 8832
rect 15896 8820 15902 8832
rect 16025 8823 16083 8829
rect 16025 8820 16037 8823
rect 15896 8792 16037 8820
rect 15896 8780 15902 8792
rect 16025 8789 16037 8792
rect 16071 8789 16083 8823
rect 16025 8783 16083 8789
rect 1104 8730 18860 8752
rect 1104 8678 4315 8730
rect 4367 8678 4379 8730
rect 4431 8678 4443 8730
rect 4495 8678 4507 8730
rect 4559 8678 10982 8730
rect 11034 8678 11046 8730
rect 11098 8678 11110 8730
rect 11162 8678 11174 8730
rect 11226 8678 17648 8730
rect 17700 8678 17712 8730
rect 17764 8678 17776 8730
rect 17828 8678 17840 8730
rect 17892 8678 18860 8730
rect 1104 8656 18860 8678
rect 9493 8619 9551 8625
rect 9493 8585 9505 8619
rect 9539 8616 9551 8619
rect 9766 8616 9772 8628
rect 9539 8588 9772 8616
rect 9539 8585 9551 8588
rect 9493 8579 9551 8585
rect 9766 8576 9772 8588
rect 9824 8576 9830 8628
rect 11330 8616 11336 8628
rect 11291 8588 11336 8616
rect 11330 8576 11336 8588
rect 11388 8576 11394 8628
rect 11514 8616 11520 8628
rect 11475 8588 11520 8616
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 12434 8576 12440 8628
rect 12492 8616 12498 8628
rect 13173 8619 13231 8625
rect 13173 8616 13185 8619
rect 12492 8588 13185 8616
rect 12492 8576 12498 8588
rect 13173 8585 13185 8588
rect 13219 8616 13231 8619
rect 13262 8616 13268 8628
rect 13219 8588 13268 8616
rect 13219 8585 13231 8588
rect 13173 8579 13231 8585
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 14461 8619 14519 8625
rect 14461 8616 14473 8619
rect 14056 8588 14473 8616
rect 14056 8576 14062 8588
rect 14461 8585 14473 8588
rect 14507 8616 14519 8619
rect 15102 8616 15108 8628
rect 14507 8588 15108 8616
rect 14507 8585 14519 8588
rect 14461 8579 14519 8585
rect 15102 8576 15108 8588
rect 15160 8576 15166 8628
rect 16390 8576 16396 8628
rect 16448 8616 16454 8628
rect 16577 8619 16635 8625
rect 16577 8616 16589 8619
rect 16448 8588 16589 8616
rect 16448 8576 16454 8588
rect 16577 8585 16589 8588
rect 16623 8585 16635 8619
rect 16577 8579 16635 8585
rect 11348 8548 11376 8576
rect 11348 8520 12756 8548
rect 8754 8480 8760 8492
rect 8667 8452 8760 8480
rect 8754 8440 8760 8452
rect 8812 8480 8818 8492
rect 9490 8480 9496 8492
rect 8812 8452 9496 8480
rect 8812 8440 8818 8452
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 10594 8480 10600 8492
rect 10555 8452 10600 8480
rect 10594 8440 10600 8452
rect 10652 8440 10658 8492
rect 10965 8483 11023 8489
rect 10965 8449 10977 8483
rect 11011 8480 11023 8483
rect 11606 8480 11612 8492
rect 11011 8452 11612 8480
rect 11011 8449 11023 8452
rect 10965 8443 11023 8449
rect 9125 8415 9183 8421
rect 9125 8381 9137 8415
rect 9171 8412 9183 8415
rect 10502 8412 10508 8424
rect 9171 8384 10508 8412
rect 9171 8381 9183 8384
rect 9125 8375 9183 8381
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 11532 8421 11560 8452
rect 11606 8440 11612 8452
rect 11664 8440 11670 8492
rect 11517 8415 11575 8421
rect 11517 8381 11529 8415
rect 11563 8412 11575 8415
rect 12066 8412 12072 8424
rect 11563 8384 11597 8412
rect 12027 8384 12072 8412
rect 11563 8381 11575 8384
rect 11517 8375 11575 8381
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 12342 8412 12348 8424
rect 12303 8384 12348 8412
rect 12342 8372 12348 8384
rect 12400 8372 12406 8424
rect 12728 8421 12756 8520
rect 12986 8508 12992 8560
rect 13044 8548 13050 8560
rect 13909 8551 13967 8557
rect 13909 8548 13921 8551
rect 13044 8520 13921 8548
rect 13044 8508 13050 8520
rect 13909 8517 13921 8520
rect 13955 8517 13967 8551
rect 15562 8548 15568 8560
rect 15523 8520 15568 8548
rect 13909 8511 13967 8517
rect 15562 8508 15568 8520
rect 15620 8508 15626 8560
rect 15654 8440 15660 8492
rect 15712 8480 15718 8492
rect 15712 8452 15976 8480
rect 15712 8440 15718 8452
rect 12713 8415 12771 8421
rect 12713 8381 12725 8415
rect 12759 8381 12771 8415
rect 12713 8375 12771 8381
rect 14826 8372 14832 8424
rect 14884 8412 14890 8424
rect 15749 8415 15807 8421
rect 15749 8412 15761 8415
rect 14884 8384 15761 8412
rect 14884 8372 14890 8384
rect 15749 8381 15761 8384
rect 15795 8412 15807 8415
rect 15838 8412 15844 8424
rect 15795 8384 15844 8412
rect 15795 8381 15807 8384
rect 15749 8375 15807 8381
rect 15838 8372 15844 8384
rect 15896 8372 15902 8424
rect 15948 8421 15976 8452
rect 15933 8415 15991 8421
rect 15933 8381 15945 8415
rect 15979 8381 15991 8415
rect 15933 8375 15991 8381
rect 16117 8415 16175 8421
rect 16117 8381 16129 8415
rect 16163 8381 16175 8415
rect 16117 8375 16175 8381
rect 12618 8304 12624 8356
rect 12676 8344 12682 8356
rect 13354 8344 13360 8356
rect 12676 8316 13360 8344
rect 12676 8304 12682 8316
rect 13354 8304 13360 8316
rect 13412 8344 13418 8356
rect 13541 8347 13599 8353
rect 13541 8344 13553 8347
rect 13412 8316 13553 8344
rect 13412 8304 13418 8316
rect 13541 8313 13553 8316
rect 13587 8313 13599 8347
rect 13541 8307 13599 8313
rect 15654 8304 15660 8356
rect 15712 8344 15718 8356
rect 16132 8344 16160 8375
rect 16945 8347 17003 8353
rect 16945 8344 16957 8347
rect 15712 8316 16957 8344
rect 15712 8304 15718 8316
rect 16945 8313 16957 8316
rect 16991 8313 17003 8347
rect 16945 8307 17003 8313
rect 1104 8186 18860 8208
rect 1104 8134 7648 8186
rect 7700 8134 7712 8186
rect 7764 8134 7776 8186
rect 7828 8134 7840 8186
rect 7892 8134 14315 8186
rect 14367 8134 14379 8186
rect 14431 8134 14443 8186
rect 14495 8134 14507 8186
rect 14559 8134 18860 8186
rect 1104 8112 18860 8134
rect 11517 8075 11575 8081
rect 11517 8041 11529 8075
rect 11563 8072 11575 8075
rect 12066 8072 12072 8084
rect 11563 8044 12072 8072
rect 11563 8041 11575 8044
rect 11517 8035 11575 8041
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 14185 8075 14243 8081
rect 14185 8041 14197 8075
rect 14231 8072 14243 8075
rect 14734 8072 14740 8084
rect 14231 8044 14740 8072
rect 14231 8041 14243 8044
rect 14185 8035 14243 8041
rect 14734 8032 14740 8044
rect 14792 8072 14798 8084
rect 15378 8072 15384 8084
rect 14792 8044 15384 8072
rect 14792 8032 14798 8044
rect 15378 8032 15384 8044
rect 15436 8072 15442 8084
rect 15436 8044 15608 8072
rect 15436 8032 15442 8044
rect 11149 8007 11207 8013
rect 11149 7973 11161 8007
rect 11195 8004 11207 8007
rect 11330 8004 11336 8016
rect 11195 7976 11336 8004
rect 11195 7973 11207 7976
rect 11149 7967 11207 7973
rect 11330 7964 11336 7976
rect 11388 8004 11394 8016
rect 11790 8004 11796 8016
rect 11388 7976 11796 8004
rect 11388 7964 11394 7976
rect 11790 7964 11796 7976
rect 11848 7964 11854 8016
rect 12802 7964 12808 8016
rect 12860 8004 12866 8016
rect 15010 8004 15016 8016
rect 12860 7976 13492 8004
rect 12860 7964 12866 7976
rect 8754 7936 8760 7948
rect 8715 7908 8760 7936
rect 8754 7896 8760 7908
rect 8812 7896 8818 7948
rect 8846 7896 8852 7948
rect 8904 7936 8910 7948
rect 9033 7939 9091 7945
rect 9033 7936 9045 7939
rect 8904 7908 9045 7936
rect 8904 7896 8910 7908
rect 9033 7905 9045 7908
rect 9079 7905 9091 7939
rect 9033 7899 9091 7905
rect 11974 7896 11980 7948
rect 12032 7936 12038 7948
rect 13464 7945 13492 7976
rect 14844 7976 15016 8004
rect 13265 7939 13323 7945
rect 13265 7936 13277 7939
rect 12032 7908 13277 7936
rect 12032 7896 12038 7908
rect 13265 7905 13277 7908
rect 13311 7905 13323 7939
rect 13265 7899 13323 7905
rect 13449 7939 13507 7945
rect 13449 7905 13461 7939
rect 13495 7905 13507 7939
rect 13449 7899 13507 7905
rect 14182 7896 14188 7948
rect 14240 7936 14246 7948
rect 14277 7939 14335 7945
rect 14277 7936 14289 7939
rect 14240 7908 14289 7936
rect 14240 7896 14246 7908
rect 14277 7905 14289 7908
rect 14323 7905 14335 7939
rect 14277 7899 14335 7905
rect 14734 7896 14740 7948
rect 14792 7936 14798 7948
rect 14844 7945 14872 7976
rect 15010 7964 15016 7976
rect 15068 7964 15074 8016
rect 14829 7939 14887 7945
rect 14829 7936 14841 7939
rect 14792 7908 14841 7936
rect 14792 7896 14798 7908
rect 14829 7905 14841 7908
rect 14875 7905 14887 7939
rect 14829 7899 14887 7905
rect 15286 7896 15292 7948
rect 15344 7936 15350 7948
rect 15473 7939 15531 7945
rect 15473 7936 15485 7939
rect 15344 7908 15485 7936
rect 15344 7896 15350 7908
rect 15473 7905 15485 7908
rect 15519 7905 15531 7939
rect 15580 7936 15608 8044
rect 15841 7939 15899 7945
rect 15841 7936 15853 7939
rect 15580 7908 15853 7936
rect 15473 7899 15531 7905
rect 15841 7905 15853 7908
rect 15887 7905 15899 7939
rect 15841 7899 15899 7905
rect 12434 7828 12440 7880
rect 12492 7868 12498 7880
rect 12492 7840 12537 7868
rect 12492 7828 12498 7840
rect 12710 7828 12716 7880
rect 12768 7868 12774 7880
rect 12989 7871 13047 7877
rect 12989 7868 13001 7871
rect 12768 7840 13001 7868
rect 12768 7828 12774 7840
rect 12989 7837 13001 7840
rect 13035 7837 13047 7871
rect 12989 7831 13047 7837
rect 13004 7800 13032 7831
rect 15010 7828 15016 7880
rect 15068 7868 15074 7880
rect 15068 7840 15113 7868
rect 15068 7828 15074 7840
rect 15654 7828 15660 7880
rect 15712 7868 15718 7880
rect 16298 7868 16304 7880
rect 15712 7840 16304 7868
rect 15712 7828 15718 7840
rect 16298 7828 16304 7840
rect 16356 7868 16362 7880
rect 16393 7871 16451 7877
rect 16393 7868 16405 7871
rect 16356 7840 16405 7868
rect 16356 7828 16362 7840
rect 16393 7837 16405 7840
rect 16439 7837 16451 7871
rect 16393 7831 16451 7837
rect 13725 7803 13783 7809
rect 13725 7800 13737 7803
rect 13004 7772 13737 7800
rect 13725 7769 13737 7772
rect 13771 7800 13783 7803
rect 13814 7800 13820 7812
rect 13771 7772 13820 7800
rect 13771 7769 13783 7772
rect 13725 7763 13783 7769
rect 13814 7760 13820 7772
rect 13872 7760 13878 7812
rect 10318 7732 10324 7744
rect 10279 7704 10324 7732
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 1104 7642 18860 7664
rect 1104 7590 4315 7642
rect 4367 7590 4379 7642
rect 4431 7590 4443 7642
rect 4495 7590 4507 7642
rect 4559 7590 10982 7642
rect 11034 7590 11046 7642
rect 11098 7590 11110 7642
rect 11162 7590 11174 7642
rect 11226 7590 17648 7642
rect 17700 7590 17712 7642
rect 17764 7590 17776 7642
rect 17828 7590 17840 7642
rect 17892 7590 18860 7642
rect 1104 7568 18860 7590
rect 8662 7488 8668 7540
rect 8720 7528 8726 7540
rect 9125 7531 9183 7537
rect 9125 7528 9137 7531
rect 8720 7500 9137 7528
rect 8720 7488 8726 7500
rect 9125 7497 9137 7500
rect 9171 7528 9183 7531
rect 9582 7528 9588 7540
rect 9171 7500 9588 7528
rect 9171 7497 9183 7500
rect 9125 7491 9183 7497
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 10686 7488 10692 7540
rect 10744 7528 10750 7540
rect 10873 7531 10931 7537
rect 10873 7528 10885 7531
rect 10744 7500 10885 7528
rect 10744 7488 10750 7500
rect 10873 7497 10885 7500
rect 10919 7497 10931 7531
rect 10873 7491 10931 7497
rect 12529 7531 12587 7537
rect 12529 7497 12541 7531
rect 12575 7528 12587 7531
rect 12802 7528 12808 7540
rect 12575 7500 12808 7528
rect 12575 7497 12587 7500
rect 12529 7491 12587 7497
rect 8754 7460 8760 7472
rect 8715 7432 8760 7460
rect 8754 7420 8760 7432
rect 8812 7420 8818 7472
rect 10888 7460 10916 7491
rect 12802 7488 12808 7500
rect 12860 7488 12866 7540
rect 11514 7460 11520 7472
rect 10888 7432 11520 7460
rect 11514 7420 11520 7432
rect 11572 7460 11578 7472
rect 11572 7432 12112 7460
rect 11572 7420 11578 7432
rect 10318 7352 10324 7404
rect 10376 7392 10382 7404
rect 12084 7401 12112 7432
rect 10597 7395 10655 7401
rect 10597 7392 10609 7395
rect 10376 7364 10609 7392
rect 10376 7352 10382 7364
rect 10597 7361 10609 7364
rect 10643 7392 10655 7395
rect 12069 7395 12127 7401
rect 10643 7364 11468 7392
rect 10643 7361 10655 7364
rect 10597 7355 10655 7361
rect 11440 7336 11468 7364
rect 12069 7361 12081 7395
rect 12115 7361 12127 7395
rect 12820 7392 12848 7488
rect 13081 7395 13139 7401
rect 13081 7392 13093 7395
rect 12820 7364 13093 7392
rect 12069 7355 12127 7361
rect 13081 7361 13093 7364
rect 13127 7392 13139 7395
rect 13170 7392 13176 7404
rect 13127 7364 13176 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 13170 7352 13176 7364
rect 13228 7352 13234 7404
rect 14918 7352 14924 7404
rect 14976 7392 14982 7404
rect 15013 7395 15071 7401
rect 15013 7392 15025 7395
rect 14976 7364 15025 7392
rect 14976 7352 14982 7364
rect 15013 7361 15025 7364
rect 15059 7392 15071 7395
rect 16482 7392 16488 7404
rect 15059 7364 15792 7392
rect 16443 7364 16488 7392
rect 15059 7361 15071 7364
rect 15013 7355 15071 7361
rect 5626 7324 5632 7336
rect 5587 7296 5632 7324
rect 5626 7284 5632 7296
rect 5684 7284 5690 7336
rect 5905 7327 5963 7333
rect 5905 7324 5917 7327
rect 5736 7296 5917 7324
rect 5534 7188 5540 7200
rect 5495 7160 5540 7188
rect 5534 7148 5540 7160
rect 5592 7188 5598 7200
rect 5736 7188 5764 7296
rect 5905 7293 5917 7296
rect 5951 7293 5963 7327
rect 5905 7287 5963 7293
rect 11149 7327 11207 7333
rect 11149 7293 11161 7327
rect 11195 7324 11207 7327
rect 11330 7324 11336 7336
rect 11195 7296 11336 7324
rect 11195 7293 11207 7296
rect 11149 7287 11207 7293
rect 11330 7284 11336 7296
rect 11388 7284 11394 7336
rect 11422 7284 11428 7336
rect 11480 7324 11486 7336
rect 11977 7327 12035 7333
rect 11977 7324 11989 7327
rect 11480 7296 11989 7324
rect 11480 7284 11486 7296
rect 11977 7293 11989 7296
rect 12023 7293 12035 7327
rect 13354 7324 13360 7336
rect 13315 7296 13360 7324
rect 11977 7287 12035 7293
rect 13354 7284 13360 7296
rect 13412 7284 13418 7336
rect 13814 7324 13820 7336
rect 13775 7296 13820 7324
rect 13814 7284 13820 7296
rect 13872 7284 13878 7336
rect 14093 7327 14151 7333
rect 14093 7293 14105 7327
rect 14139 7324 14151 7327
rect 15102 7324 15108 7336
rect 14139 7296 15108 7324
rect 14139 7293 14151 7296
rect 14093 7287 14151 7293
rect 15102 7284 15108 7296
rect 15160 7284 15166 7336
rect 15764 7333 15792 7364
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 15381 7327 15439 7333
rect 15381 7293 15393 7327
rect 15427 7293 15439 7327
rect 15381 7287 15439 7293
rect 15749 7327 15807 7333
rect 15749 7293 15761 7327
rect 15795 7293 15807 7327
rect 16206 7324 16212 7336
rect 16167 7296 16212 7324
rect 15749 7287 15807 7293
rect 7282 7256 7288 7268
rect 7243 7228 7288 7256
rect 7282 7216 7288 7228
rect 7340 7216 7346 7268
rect 11241 7259 11299 7265
rect 11241 7225 11253 7259
rect 11287 7256 11299 7259
rect 11790 7256 11796 7268
rect 11287 7228 11796 7256
rect 11287 7225 11299 7228
rect 11241 7219 11299 7225
rect 11790 7216 11796 7228
rect 11848 7216 11854 7268
rect 14461 7259 14519 7265
rect 14461 7225 14473 7259
rect 14507 7256 14519 7259
rect 15286 7256 15292 7268
rect 14507 7228 15292 7256
rect 14507 7225 14519 7228
rect 14461 7219 14519 7225
rect 15286 7216 15292 7228
rect 15344 7256 15350 7268
rect 15396 7256 15424 7287
rect 16206 7284 16212 7296
rect 16264 7284 16270 7336
rect 15344 7228 15424 7256
rect 15344 7216 15350 7228
rect 5592 7160 5764 7188
rect 5592 7148 5598 7160
rect 1104 7098 18860 7120
rect 1104 7046 7648 7098
rect 7700 7046 7712 7098
rect 7764 7046 7776 7098
rect 7828 7046 7840 7098
rect 7892 7046 14315 7098
rect 14367 7046 14379 7098
rect 14431 7046 14443 7098
rect 14495 7046 14507 7098
rect 14559 7046 18860 7098
rect 1104 7024 18860 7046
rect 5718 6984 5724 6996
rect 5679 6956 5724 6984
rect 5718 6944 5724 6956
rect 5776 6944 5782 6996
rect 12710 6984 12716 6996
rect 12671 6956 12716 6984
rect 12710 6944 12716 6956
rect 12768 6944 12774 6996
rect 13081 6987 13139 6993
rect 13081 6953 13093 6987
rect 13127 6984 13139 6987
rect 13354 6984 13360 6996
rect 13127 6956 13360 6984
rect 13127 6953 13139 6956
rect 13081 6947 13139 6953
rect 13354 6944 13360 6956
rect 13412 6944 13418 6996
rect 13262 6876 13268 6928
rect 13320 6916 13326 6928
rect 14918 6916 14924 6928
rect 13320 6888 13860 6916
rect 14831 6888 14924 6916
rect 13320 6876 13326 6888
rect 10134 6848 10140 6860
rect 10095 6820 10140 6848
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 11517 6851 11575 6857
rect 11517 6817 11529 6851
rect 11563 6848 11575 6851
rect 12158 6848 12164 6860
rect 11563 6820 12164 6848
rect 11563 6817 11575 6820
rect 11517 6811 11575 6817
rect 12158 6808 12164 6820
rect 12216 6848 12222 6860
rect 13173 6851 13231 6857
rect 13173 6848 13185 6851
rect 12216 6820 13185 6848
rect 12216 6808 12222 6820
rect 13173 6817 13185 6820
rect 13219 6817 13231 6851
rect 13173 6811 13231 6817
rect 13725 6851 13783 6857
rect 13725 6817 13737 6851
rect 13771 6817 13783 6851
rect 13832 6848 13860 6888
rect 14844 6857 14872 6888
rect 14918 6876 14924 6888
rect 14976 6916 14982 6928
rect 15378 6916 15384 6928
rect 14976 6888 15384 6916
rect 14976 6876 14982 6888
rect 15378 6876 15384 6888
rect 15436 6876 15442 6928
rect 16776 6888 17080 6916
rect 14369 6851 14427 6857
rect 14369 6848 14381 6851
rect 13832 6820 14381 6848
rect 13725 6811 13783 6817
rect 14369 6817 14381 6820
rect 14415 6817 14427 6851
rect 14369 6811 14427 6817
rect 14829 6851 14887 6857
rect 14829 6817 14841 6851
rect 14875 6817 14887 6851
rect 14829 6811 14887 6817
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 9861 6783 9919 6789
rect 9861 6780 9873 6783
rect 9732 6752 9873 6780
rect 9732 6740 9738 6752
rect 9861 6749 9873 6752
rect 9907 6780 9919 6783
rect 10226 6780 10232 6792
rect 9907 6752 10232 6780
rect 9907 6749 9919 6752
rect 9861 6743 9919 6749
rect 10226 6740 10232 6752
rect 10284 6740 10290 6792
rect 11974 6672 11980 6724
rect 12032 6712 12038 6724
rect 12161 6715 12219 6721
rect 12161 6712 12173 6715
rect 12032 6684 12173 6712
rect 12032 6672 12038 6684
rect 12161 6681 12173 6684
rect 12207 6681 12219 6715
rect 13740 6712 13768 6811
rect 15838 6808 15844 6860
rect 15896 6848 15902 6860
rect 16577 6851 16635 6857
rect 16577 6848 16589 6851
rect 15896 6820 16589 6848
rect 15896 6808 15902 6820
rect 16577 6817 16589 6820
rect 16623 6848 16635 6851
rect 16776 6848 16804 6888
rect 16942 6848 16948 6860
rect 16623 6820 16804 6848
rect 16903 6820 16948 6848
rect 16623 6817 16635 6820
rect 16577 6811 16635 6817
rect 16942 6808 16948 6820
rect 17000 6808 17006 6860
rect 17052 6848 17080 6888
rect 17402 6848 17408 6860
rect 17052 6820 17408 6848
rect 17402 6808 17408 6820
rect 17460 6808 17466 6860
rect 13906 6780 13912 6792
rect 13867 6752 13912 6780
rect 13906 6740 13912 6752
rect 13964 6740 13970 6792
rect 17034 6780 17040 6792
rect 16995 6752 17040 6780
rect 17034 6740 17040 6752
rect 17092 6740 17098 6792
rect 13814 6712 13820 6724
rect 13727 6684 13820 6712
rect 12161 6675 12219 6681
rect 13814 6672 13820 6684
rect 13872 6712 13878 6724
rect 14734 6712 14740 6724
rect 13872 6684 14740 6712
rect 13872 6672 13878 6684
rect 14734 6672 14740 6684
rect 14792 6672 14798 6724
rect 15194 6672 15200 6724
rect 15252 6712 15258 6724
rect 15749 6715 15807 6721
rect 15749 6712 15761 6715
rect 15252 6684 15761 6712
rect 15252 6672 15258 6684
rect 15749 6681 15761 6684
rect 15795 6712 15807 6715
rect 16206 6712 16212 6724
rect 15795 6684 16212 6712
rect 15795 6681 15807 6684
rect 15749 6675 15807 6681
rect 16206 6672 16212 6684
rect 16264 6672 16270 6724
rect 16393 6715 16451 6721
rect 16393 6681 16405 6715
rect 16439 6712 16451 6715
rect 16482 6712 16488 6724
rect 16439 6684 16488 6712
rect 16439 6681 16451 6684
rect 16393 6675 16451 6681
rect 16482 6672 16488 6684
rect 16540 6672 16546 6724
rect 17402 6712 17408 6724
rect 17363 6684 17408 6712
rect 17402 6672 17408 6684
rect 17460 6672 17466 6724
rect 15286 6604 15292 6656
rect 15344 6644 15350 6656
rect 15381 6647 15439 6653
rect 15381 6644 15393 6647
rect 15344 6616 15393 6644
rect 15344 6604 15350 6616
rect 15381 6613 15393 6616
rect 15427 6613 15439 6647
rect 15381 6607 15439 6613
rect 1104 6554 18860 6576
rect 1104 6502 4315 6554
rect 4367 6502 4379 6554
rect 4431 6502 4443 6554
rect 4495 6502 4507 6554
rect 4559 6502 10982 6554
rect 11034 6502 11046 6554
rect 11098 6502 11110 6554
rect 11162 6502 11174 6554
rect 11226 6502 17648 6554
rect 17700 6502 17712 6554
rect 17764 6502 17776 6554
rect 17828 6502 17840 6554
rect 17892 6502 18860 6554
rect 1104 6480 18860 6502
rect 9953 6443 10011 6449
rect 9953 6409 9965 6443
rect 9999 6440 10011 6443
rect 10134 6440 10140 6452
rect 9999 6412 10140 6440
rect 9999 6409 10011 6412
rect 9953 6403 10011 6409
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 10226 6400 10232 6452
rect 10284 6440 10290 6452
rect 10284 6412 10329 6440
rect 10284 6400 10290 6412
rect 10778 6400 10784 6452
rect 10836 6440 10842 6452
rect 10873 6443 10931 6449
rect 10873 6440 10885 6443
rect 10836 6412 10885 6440
rect 10836 6400 10842 6412
rect 10873 6409 10885 6412
rect 10919 6409 10931 6443
rect 10873 6403 10931 6409
rect 11333 6443 11391 6449
rect 11333 6409 11345 6443
rect 11379 6440 11391 6443
rect 11514 6440 11520 6452
rect 11379 6412 11520 6440
rect 11379 6409 11391 6412
rect 11333 6403 11391 6409
rect 10888 6236 10916 6403
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 13170 6440 13176 6452
rect 13131 6412 13176 6440
rect 13170 6400 13176 6412
rect 13228 6400 13234 6452
rect 14182 6400 14188 6452
rect 14240 6440 14246 6452
rect 15013 6443 15071 6449
rect 15013 6440 15025 6443
rect 14240 6412 15025 6440
rect 14240 6400 14246 6412
rect 15013 6409 15025 6412
rect 15059 6409 15071 6443
rect 15838 6440 15844 6452
rect 15799 6412 15844 6440
rect 15013 6403 15071 6409
rect 15838 6400 15844 6412
rect 15896 6400 15902 6452
rect 16209 6443 16267 6449
rect 16209 6409 16221 6443
rect 16255 6440 16267 6443
rect 16577 6443 16635 6449
rect 16577 6440 16589 6443
rect 16255 6412 16589 6440
rect 16255 6409 16267 6412
rect 16209 6403 16267 6409
rect 16577 6409 16589 6412
rect 16623 6440 16635 6443
rect 16942 6440 16948 6452
rect 16623 6412 16948 6440
rect 16623 6409 16635 6412
rect 16577 6403 16635 6409
rect 16942 6400 16948 6412
rect 17000 6440 17006 6452
rect 17000 6412 17172 6440
rect 17000 6400 17006 6412
rect 11532 6372 11560 6400
rect 13630 6372 13636 6384
rect 11532 6344 11744 6372
rect 13591 6344 13636 6372
rect 11606 6304 11612 6316
rect 11567 6276 11612 6304
rect 11606 6264 11612 6276
rect 11664 6264 11670 6316
rect 11716 6304 11744 6344
rect 13630 6332 13636 6344
rect 13688 6332 13694 6384
rect 14734 6372 14740 6384
rect 14695 6344 14740 6372
rect 14734 6332 14740 6344
rect 14792 6332 14798 6384
rect 17034 6372 17040 6384
rect 16995 6344 17040 6372
rect 17034 6332 17040 6344
rect 17092 6332 17098 6384
rect 17144 6316 17172 6412
rect 12437 6307 12495 6313
rect 12437 6304 12449 6307
rect 11716 6276 12449 6304
rect 12437 6273 12449 6276
rect 12483 6273 12495 6307
rect 14642 6304 14648 6316
rect 12437 6267 12495 6273
rect 13832 6276 14648 6304
rect 11517 6239 11575 6245
rect 11517 6236 11529 6239
rect 10888 6208 11529 6236
rect 11517 6205 11529 6208
rect 11563 6205 11575 6239
rect 11517 6199 11575 6205
rect 11698 6196 11704 6248
rect 11756 6236 11762 6248
rect 13832 6245 13860 6276
rect 14642 6264 14648 6276
rect 14700 6264 14706 6316
rect 17126 6304 17132 6316
rect 17039 6276 17132 6304
rect 17126 6264 17132 6276
rect 17184 6304 17190 6316
rect 17184 6276 17448 6304
rect 17184 6264 17190 6276
rect 12345 6239 12403 6245
rect 12345 6236 12357 6239
rect 11756 6208 12357 6236
rect 11756 6196 11762 6208
rect 12345 6205 12357 6208
rect 12391 6205 12403 6239
rect 12345 6199 12403 6205
rect 13817 6239 13875 6245
rect 13817 6205 13829 6239
rect 13863 6205 13875 6239
rect 13998 6236 14004 6248
rect 13959 6208 14004 6236
rect 13817 6199 13875 6205
rect 13998 6196 14004 6208
rect 14056 6196 14062 6248
rect 14185 6239 14243 6245
rect 14185 6205 14197 6239
rect 14231 6205 14243 6239
rect 14185 6199 14243 6205
rect 13262 6128 13268 6180
rect 13320 6168 13326 6180
rect 14200 6168 14228 6199
rect 16758 6196 16764 6248
rect 16816 6236 16822 6248
rect 17221 6239 17279 6245
rect 17221 6236 17233 6239
rect 16816 6208 17233 6236
rect 16816 6196 16822 6208
rect 17221 6205 17233 6208
rect 17267 6236 17279 6239
rect 17310 6236 17316 6248
rect 17267 6208 17316 6236
rect 17267 6205 17279 6208
rect 17221 6199 17279 6205
rect 17310 6196 17316 6208
rect 17368 6196 17374 6248
rect 17420 6245 17448 6276
rect 17405 6239 17463 6245
rect 17405 6205 17417 6239
rect 17451 6205 17463 6239
rect 17405 6199 17463 6205
rect 17494 6196 17500 6248
rect 17552 6236 17558 6248
rect 17589 6239 17647 6245
rect 17589 6236 17601 6239
rect 17552 6208 17601 6236
rect 17552 6196 17558 6208
rect 17589 6205 17601 6208
rect 17635 6205 17647 6239
rect 17589 6199 17647 6205
rect 13320 6140 14228 6168
rect 13320 6128 13326 6140
rect 12897 6103 12955 6109
rect 12897 6069 12909 6103
rect 12943 6100 12955 6103
rect 13998 6100 14004 6112
rect 12943 6072 14004 6100
rect 12943 6069 12955 6072
rect 12897 6063 12955 6069
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 1104 6010 18860 6032
rect 1104 5958 7648 6010
rect 7700 5958 7712 6010
rect 7764 5958 7776 6010
rect 7828 5958 7840 6010
rect 7892 5958 14315 6010
rect 14367 5958 14379 6010
rect 14431 5958 14443 6010
rect 14495 5958 14507 6010
rect 14559 5958 18860 6010
rect 1104 5936 18860 5958
rect 11698 5896 11704 5908
rect 11659 5868 11704 5896
rect 11698 5856 11704 5868
rect 11756 5856 11762 5908
rect 12158 5896 12164 5908
rect 12119 5868 12164 5896
rect 12158 5856 12164 5868
rect 12216 5896 12222 5908
rect 13262 5896 13268 5908
rect 12216 5868 13268 5896
rect 12216 5856 12222 5868
rect 13262 5856 13268 5868
rect 13320 5856 13326 5908
rect 13814 5896 13820 5908
rect 13775 5868 13820 5896
rect 13814 5856 13820 5868
rect 13872 5856 13878 5908
rect 13998 5856 14004 5908
rect 14056 5896 14062 5908
rect 14277 5899 14335 5905
rect 14277 5896 14289 5899
rect 14056 5868 14289 5896
rect 14056 5856 14062 5868
rect 14277 5865 14289 5868
rect 14323 5896 14335 5899
rect 14642 5896 14648 5908
rect 14323 5868 14648 5896
rect 14323 5865 14335 5868
rect 14277 5859 14335 5865
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 16022 5896 16028 5908
rect 15935 5868 16028 5896
rect 16022 5856 16028 5868
rect 16080 5896 16086 5908
rect 16850 5896 16856 5908
rect 16080 5868 16856 5896
rect 16080 5856 16086 5868
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 17310 5856 17316 5908
rect 17368 5896 17374 5908
rect 17405 5899 17463 5905
rect 17405 5896 17417 5899
rect 17368 5868 17417 5896
rect 17368 5856 17374 5868
rect 17405 5865 17417 5868
rect 17451 5865 17463 5899
rect 17405 5859 17463 5865
rect 8938 5828 8944 5840
rect 8899 5800 8944 5828
rect 8938 5788 8944 5800
rect 8996 5788 9002 5840
rect 13170 5828 13176 5840
rect 13131 5800 13176 5828
rect 13170 5788 13176 5800
rect 13228 5788 13234 5840
rect 13541 5831 13599 5837
rect 13541 5797 13553 5831
rect 13587 5828 13599 5831
rect 14918 5828 14924 5840
rect 13587 5800 14924 5828
rect 13587 5797 13599 5800
rect 13541 5791 13599 5797
rect 14918 5788 14924 5800
rect 14976 5788 14982 5840
rect 15286 5828 15292 5840
rect 15247 5800 15292 5828
rect 15286 5788 15292 5800
rect 15344 5788 15350 5840
rect 1670 5720 1676 5772
rect 1728 5760 1734 5772
rect 2133 5763 2191 5769
rect 2133 5760 2145 5763
rect 1728 5732 2145 5760
rect 1728 5720 1734 5732
rect 2133 5729 2145 5732
rect 2179 5729 2191 5763
rect 2133 5723 2191 5729
rect 2222 5720 2228 5772
rect 2280 5760 2286 5772
rect 2409 5763 2467 5769
rect 2409 5760 2421 5763
rect 2280 5732 2421 5760
rect 2280 5720 2286 5732
rect 2409 5729 2421 5732
rect 2455 5729 2467 5763
rect 3786 5760 3792 5772
rect 3747 5732 3792 5760
rect 2409 5723 2467 5729
rect 3786 5720 3792 5732
rect 3844 5720 3850 5772
rect 7374 5720 7380 5772
rect 7432 5760 7438 5772
rect 7561 5763 7619 5769
rect 7561 5760 7573 5763
rect 7432 5732 7573 5760
rect 7432 5720 7438 5732
rect 7561 5729 7573 5732
rect 7607 5729 7619 5763
rect 7561 5723 7619 5729
rect 9674 5720 9680 5772
rect 9732 5760 9738 5772
rect 9769 5763 9827 5769
rect 9769 5760 9781 5763
rect 9732 5732 9781 5760
rect 9732 5720 9738 5732
rect 9769 5729 9781 5732
rect 9815 5729 9827 5763
rect 9769 5723 9827 5729
rect 9858 5720 9864 5772
rect 9916 5760 9922 5772
rect 10045 5763 10103 5769
rect 10045 5760 10057 5763
rect 9916 5732 10057 5760
rect 9916 5720 9922 5732
rect 10045 5729 10057 5732
rect 10091 5729 10103 5763
rect 12526 5760 12532 5772
rect 12487 5732 12532 5760
rect 10045 5723 10103 5729
rect 12526 5720 12532 5732
rect 12584 5720 12590 5772
rect 14642 5760 14648 5772
rect 14603 5732 14648 5760
rect 14642 5720 14648 5732
rect 14700 5720 14706 5772
rect 16574 5760 16580 5772
rect 16535 5732 16580 5760
rect 16574 5720 16580 5732
rect 16632 5720 16638 5772
rect 16942 5760 16948 5772
rect 16903 5732 16948 5760
rect 16942 5720 16948 5732
rect 17000 5720 17006 5772
rect 17037 5763 17095 5769
rect 17037 5729 17049 5763
rect 17083 5760 17095 5763
rect 17126 5760 17132 5772
rect 17083 5732 17132 5760
rect 17083 5729 17095 5732
rect 17037 5723 17095 5729
rect 17126 5720 17132 5732
rect 17184 5720 17190 5772
rect 7285 5695 7343 5701
rect 7285 5661 7297 5695
rect 7331 5692 7343 5695
rect 7742 5692 7748 5704
rect 7331 5664 7748 5692
rect 7331 5661 7343 5664
rect 7285 5655 7343 5661
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 11422 5692 11428 5704
rect 11383 5664 11428 5692
rect 11422 5652 11428 5664
rect 11480 5652 11486 5704
rect 16390 5624 16396 5636
rect 16351 5596 16396 5624
rect 16390 5584 16396 5596
rect 16448 5584 16454 5636
rect 1104 5466 18860 5488
rect 1104 5414 4315 5466
rect 4367 5414 4379 5466
rect 4431 5414 4443 5466
rect 4495 5414 4507 5466
rect 4559 5414 10982 5466
rect 11034 5414 11046 5466
rect 11098 5414 11110 5466
rect 11162 5414 11174 5466
rect 11226 5414 17648 5466
rect 17700 5414 17712 5466
rect 17764 5414 17776 5466
rect 17828 5414 17840 5466
rect 17892 5414 18860 5466
rect 1104 5392 18860 5414
rect 1670 5312 1676 5364
rect 1728 5352 1734 5364
rect 2501 5355 2559 5361
rect 2501 5352 2513 5355
rect 1728 5324 2513 5352
rect 1728 5312 1734 5324
rect 2501 5321 2513 5324
rect 2547 5321 2559 5355
rect 7742 5352 7748 5364
rect 7655 5324 7748 5352
rect 2501 5315 2559 5321
rect 7742 5312 7748 5324
rect 7800 5352 7806 5364
rect 9674 5352 9680 5364
rect 7800 5324 9680 5352
rect 7800 5312 7806 5324
rect 9674 5312 9680 5324
rect 9732 5352 9738 5364
rect 10226 5352 10232 5364
rect 9732 5324 10232 5352
rect 9732 5312 9738 5324
rect 10226 5312 10232 5324
rect 10284 5312 10290 5364
rect 12526 5352 12532 5364
rect 12487 5324 12532 5352
rect 12526 5312 12532 5324
rect 12584 5312 12590 5364
rect 13173 5355 13231 5361
rect 13173 5321 13185 5355
rect 13219 5352 13231 5355
rect 13262 5352 13268 5364
rect 13219 5324 13268 5352
rect 13219 5321 13231 5324
rect 13173 5315 13231 5321
rect 13262 5312 13268 5324
rect 13320 5312 13326 5364
rect 16574 5312 16580 5364
rect 16632 5352 16638 5364
rect 16945 5355 17003 5361
rect 16945 5352 16957 5355
rect 16632 5324 16957 5352
rect 16632 5312 16638 5324
rect 16945 5321 16957 5324
rect 16991 5321 17003 5355
rect 16945 5315 17003 5321
rect 12434 5244 12440 5296
rect 12492 5284 12498 5296
rect 13449 5287 13507 5293
rect 13449 5284 13461 5287
rect 12492 5256 13461 5284
rect 12492 5244 12498 5256
rect 13449 5253 13461 5256
rect 13495 5284 13507 5287
rect 15562 5284 15568 5296
rect 13495 5256 14136 5284
rect 15523 5256 15568 5284
rect 13495 5253 13507 5256
rect 13449 5247 13507 5253
rect 13998 5216 14004 5228
rect 13959 5188 14004 5216
rect 13998 5176 14004 5188
rect 14056 5176 14062 5228
rect 2130 5148 2136 5160
rect 2091 5120 2136 5148
rect 2130 5108 2136 5120
rect 2188 5108 2194 5160
rect 13906 5148 13912 5160
rect 13867 5120 13912 5148
rect 13906 5108 13912 5120
rect 13964 5108 13970 5160
rect 14108 5148 14136 5256
rect 15562 5244 15568 5256
rect 15620 5244 15626 5296
rect 16669 5287 16727 5293
rect 16669 5284 16681 5287
rect 16224 5256 16681 5284
rect 16224 5225 16252 5256
rect 16669 5253 16681 5256
rect 16715 5284 16727 5287
rect 17126 5284 17132 5296
rect 16715 5256 17132 5284
rect 16715 5253 16727 5256
rect 16669 5247 16727 5253
rect 17126 5244 17132 5256
rect 17184 5244 17190 5296
rect 15105 5219 15163 5225
rect 15105 5185 15117 5219
rect 15151 5216 15163 5219
rect 16209 5219 16267 5225
rect 16209 5216 16221 5219
rect 15151 5188 16221 5216
rect 15151 5185 15163 5188
rect 15105 5179 15163 5185
rect 16209 5185 16221 5188
rect 16255 5185 16267 5219
rect 16209 5179 16267 5185
rect 14182 5148 14188 5160
rect 14095 5120 14188 5148
rect 14182 5108 14188 5120
rect 14240 5108 14246 5160
rect 15470 5108 15476 5160
rect 15528 5148 15534 5160
rect 15749 5151 15807 5157
rect 15749 5148 15761 5151
rect 15528 5120 15761 5148
rect 15528 5108 15534 5120
rect 15749 5117 15761 5120
rect 15795 5117 15807 5151
rect 15749 5111 15807 5117
rect 16117 5151 16175 5157
rect 16117 5117 16129 5151
rect 16163 5117 16175 5151
rect 16117 5111 16175 5117
rect 7282 5012 7288 5024
rect 7243 4984 7288 5012
rect 7282 4972 7288 4984
rect 7340 4972 7346 5024
rect 9858 5012 9864 5024
rect 9819 4984 9864 5012
rect 9858 4972 9864 4984
rect 9916 4972 9922 5024
rect 14642 5012 14648 5024
rect 14603 4984 14648 5012
rect 14642 4972 14648 4984
rect 14700 5012 14706 5024
rect 16132 5012 16160 5111
rect 14700 4984 16160 5012
rect 14700 4972 14706 4984
rect 1104 4922 18860 4944
rect 1104 4870 7648 4922
rect 7700 4870 7712 4922
rect 7764 4870 7776 4922
rect 7828 4870 7840 4922
rect 7892 4870 14315 4922
rect 14367 4870 14379 4922
rect 14431 4870 14443 4922
rect 14495 4870 14507 4922
rect 14559 4870 18860 4922
rect 1104 4848 18860 4870
rect 1394 4768 1400 4820
rect 1452 4808 1458 4820
rect 1670 4808 1676 4820
rect 1452 4780 1676 4808
rect 1452 4768 1458 4780
rect 1670 4768 1676 4780
rect 1728 4768 1734 4820
rect 13725 4811 13783 4817
rect 13725 4777 13737 4811
rect 13771 4808 13783 4811
rect 13906 4808 13912 4820
rect 13771 4780 13912 4808
rect 13771 4777 13783 4780
rect 13725 4771 13783 4777
rect 13906 4768 13912 4780
rect 13964 4768 13970 4820
rect 14090 4808 14096 4820
rect 14051 4780 14096 4808
rect 14090 4768 14096 4780
rect 14148 4808 14154 4820
rect 16761 4811 16819 4817
rect 16761 4808 16773 4811
rect 14148 4780 16773 4808
rect 14148 4768 14154 4780
rect 16761 4777 16773 4780
rect 16807 4808 16819 4811
rect 16942 4808 16948 4820
rect 16807 4780 16948 4808
rect 16807 4777 16819 4780
rect 16761 4771 16819 4777
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 14550 4740 14556 4752
rect 14463 4712 14556 4740
rect 14476 4681 14504 4712
rect 14550 4700 14556 4712
rect 14608 4740 14614 4752
rect 15010 4740 15016 4752
rect 14608 4712 15016 4740
rect 14608 4700 14614 4712
rect 15010 4700 15016 4712
rect 15068 4700 15074 4752
rect 15381 4743 15439 4749
rect 15381 4709 15393 4743
rect 15427 4740 15439 4743
rect 15470 4740 15476 4752
rect 15427 4712 15476 4740
rect 15427 4709 15439 4712
rect 15381 4703 15439 4709
rect 15470 4700 15476 4712
rect 15528 4700 15534 4752
rect 15746 4740 15752 4752
rect 15707 4712 15752 4740
rect 15746 4700 15752 4712
rect 15804 4700 15810 4752
rect 14461 4675 14519 4681
rect 14461 4641 14473 4675
rect 14507 4641 14519 4675
rect 14461 4635 14519 4641
rect 14737 4675 14795 4681
rect 14737 4641 14749 4675
rect 14783 4672 14795 4675
rect 15194 4672 15200 4684
rect 14783 4644 15200 4672
rect 14783 4641 14795 4644
rect 14737 4635 14795 4641
rect 14182 4564 14188 4616
rect 14240 4604 14246 4616
rect 14752 4604 14780 4635
rect 15194 4632 15200 4644
rect 15252 4632 15258 4684
rect 15930 4672 15936 4684
rect 15891 4644 15936 4672
rect 15930 4632 15936 4644
rect 15988 4632 15994 4684
rect 14240 4576 14780 4604
rect 14240 4564 14246 4576
rect 14277 4539 14335 4545
rect 14277 4505 14289 4539
rect 14323 4536 14335 4539
rect 14826 4536 14832 4548
rect 14323 4508 14832 4536
rect 14323 4505 14335 4508
rect 14277 4499 14335 4505
rect 14826 4496 14832 4508
rect 14884 4496 14890 4548
rect 1104 4378 18860 4400
rect 1104 4326 4315 4378
rect 4367 4326 4379 4378
rect 4431 4326 4443 4378
rect 4495 4326 4507 4378
rect 4559 4326 10982 4378
rect 11034 4326 11046 4378
rect 11098 4326 11110 4378
rect 11162 4326 11174 4378
rect 11226 4326 17648 4378
rect 17700 4326 17712 4378
rect 17764 4326 17776 4378
rect 17828 4326 17840 4378
rect 17892 4326 18860 4378
rect 1104 4304 18860 4326
rect 14182 4264 14188 4276
rect 14143 4236 14188 4264
rect 14182 4224 14188 4236
rect 14240 4224 14246 4276
rect 14550 4264 14556 4276
rect 14511 4236 14556 4264
rect 14550 4224 14556 4236
rect 14608 4224 14614 4276
rect 15841 4267 15899 4273
rect 15841 4233 15853 4267
rect 15887 4264 15899 4267
rect 15930 4264 15936 4276
rect 15887 4236 15936 4264
rect 15887 4233 15899 4236
rect 15841 4227 15899 4233
rect 15930 4224 15936 4236
rect 15988 4224 15994 4276
rect 1394 4128 1400 4140
rect 1355 4100 1400 4128
rect 1394 4088 1400 4100
rect 1452 4088 1458 4140
rect 1670 4128 1676 4140
rect 1631 4100 1676 4128
rect 1670 4088 1676 4100
rect 1728 4088 1734 4140
rect 3050 4128 3056 4140
rect 3011 4100 3056 4128
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 10226 4128 10232 4140
rect 10187 4100 10232 4128
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 11885 4131 11943 4137
rect 11885 4097 11897 4131
rect 11931 4128 11943 4131
rect 12342 4128 12348 4140
rect 11931 4100 12348 4128
rect 11931 4097 11943 4100
rect 11885 4091 11943 4097
rect 12342 4088 12348 4100
rect 12400 4088 12406 4140
rect 10505 4063 10563 4069
rect 10505 4060 10517 4063
rect 10336 4032 10517 4060
rect 10042 3924 10048 3936
rect 10003 3896 10048 3924
rect 10042 3884 10048 3896
rect 10100 3924 10106 3936
rect 10336 3924 10364 4032
rect 10505 4029 10517 4032
rect 10551 4029 10563 4063
rect 10505 4023 10563 4029
rect 10100 3896 10364 3924
rect 10100 3884 10106 3896
rect 1104 3834 18860 3856
rect 1104 3782 7648 3834
rect 7700 3782 7712 3834
rect 7764 3782 7776 3834
rect 7828 3782 7840 3834
rect 7892 3782 14315 3834
rect 14367 3782 14379 3834
rect 14431 3782 14443 3834
rect 14495 3782 14507 3834
rect 14559 3782 18860 3834
rect 1104 3760 18860 3782
rect 1670 3720 1676 3732
rect 1631 3692 1676 3720
rect 1670 3680 1676 3692
rect 1728 3680 1734 3732
rect 10226 3720 10232 3732
rect 10187 3692 10232 3720
rect 10226 3680 10232 3692
rect 10284 3680 10290 3732
rect 1104 3290 18860 3312
rect 1104 3238 4315 3290
rect 4367 3238 4379 3290
rect 4431 3238 4443 3290
rect 4495 3238 4507 3290
rect 4559 3238 10982 3290
rect 11034 3238 11046 3290
rect 11098 3238 11110 3290
rect 11162 3238 11174 3290
rect 11226 3238 17648 3290
rect 17700 3238 17712 3290
rect 17764 3238 17776 3290
rect 17828 3238 17840 3290
rect 17892 3238 18860 3290
rect 1104 3216 18860 3238
rect 1104 2746 18860 2768
rect 1104 2694 7648 2746
rect 7700 2694 7712 2746
rect 7764 2694 7776 2746
rect 7828 2694 7840 2746
rect 7892 2694 14315 2746
rect 14367 2694 14379 2746
rect 14431 2694 14443 2746
rect 14495 2694 14507 2746
rect 14559 2694 18860 2746
rect 1104 2672 18860 2694
rect 9217 2635 9275 2641
rect 9217 2601 9229 2635
rect 9263 2632 9275 2635
rect 9766 2632 9772 2644
rect 9263 2604 9772 2632
rect 9263 2601 9275 2604
rect 9217 2595 9275 2601
rect 9766 2592 9772 2604
rect 9824 2632 9830 2644
rect 10134 2632 10140 2644
rect 9824 2604 10140 2632
rect 9824 2592 9830 2604
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 9490 2456 9496 2508
rect 9548 2496 9554 2508
rect 10045 2499 10103 2505
rect 10045 2496 10057 2499
rect 9548 2468 10057 2496
rect 9548 2456 9554 2468
rect 10045 2465 10057 2468
rect 10091 2465 10103 2499
rect 10045 2459 10103 2465
rect 9766 2428 9772 2440
rect 9727 2400 9772 2428
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 9490 2292 9496 2304
rect 9451 2264 9496 2292
rect 9490 2252 9496 2264
rect 9548 2252 9554 2304
rect 11330 2292 11336 2304
rect 11291 2264 11336 2292
rect 11330 2252 11336 2264
rect 11388 2292 11394 2304
rect 12250 2292 12256 2304
rect 11388 2264 12256 2292
rect 11388 2252 11394 2264
rect 12250 2252 12256 2264
rect 12308 2252 12314 2304
rect 1104 2202 18860 2224
rect 1104 2150 4315 2202
rect 4367 2150 4379 2202
rect 4431 2150 4443 2202
rect 4495 2150 4507 2202
rect 4559 2150 10982 2202
rect 11034 2150 11046 2202
rect 11098 2150 11110 2202
rect 11162 2150 11174 2202
rect 11226 2150 17648 2202
rect 17700 2150 17712 2202
rect 17764 2150 17776 2202
rect 17828 2150 17840 2202
rect 17892 2150 18860 2202
rect 1104 2128 18860 2150
<< via1 >>
rect 3792 78616 3844 78668
rect 4804 78616 4856 78668
rect 7648 77766 7700 77818
rect 7712 77766 7764 77818
rect 7776 77766 7828 77818
rect 7840 77766 7892 77818
rect 14315 77766 14367 77818
rect 14379 77766 14431 77818
rect 14443 77766 14495 77818
rect 14507 77766 14559 77818
rect 3240 77460 3292 77512
rect 15936 77460 15988 77512
rect 3332 77392 3384 77444
rect 16028 77392 16080 77444
rect 4315 77222 4367 77274
rect 4379 77222 4431 77274
rect 4443 77222 4495 77274
rect 4507 77222 4559 77274
rect 10982 77222 11034 77274
rect 11046 77222 11098 77274
rect 11110 77222 11162 77274
rect 11174 77222 11226 77274
rect 17648 77222 17700 77274
rect 17712 77222 17764 77274
rect 17776 77222 17828 77274
rect 17840 77222 17892 77274
rect 7648 76678 7700 76730
rect 7712 76678 7764 76730
rect 7776 76678 7828 76730
rect 7840 76678 7892 76730
rect 14315 76678 14367 76730
rect 14379 76678 14431 76730
rect 14443 76678 14495 76730
rect 14507 76678 14559 76730
rect 4315 76134 4367 76186
rect 4379 76134 4431 76186
rect 4443 76134 4495 76186
rect 4507 76134 4559 76186
rect 10982 76134 11034 76186
rect 11046 76134 11098 76186
rect 11110 76134 11162 76186
rect 11174 76134 11226 76186
rect 17648 76134 17700 76186
rect 17712 76134 17764 76186
rect 17776 76134 17828 76186
rect 17840 76134 17892 76186
rect 7648 75590 7700 75642
rect 7712 75590 7764 75642
rect 7776 75590 7828 75642
rect 7840 75590 7892 75642
rect 14315 75590 14367 75642
rect 14379 75590 14431 75642
rect 14443 75590 14495 75642
rect 14507 75590 14559 75642
rect 4160 75420 4212 75472
rect 5172 75395 5224 75404
rect 5172 75361 5181 75395
rect 5181 75361 5215 75395
rect 5215 75361 5224 75395
rect 5172 75352 5224 75361
rect 7104 75395 7156 75404
rect 7104 75361 7113 75395
rect 7113 75361 7147 75395
rect 7147 75361 7156 75395
rect 7104 75352 7156 75361
rect 4896 75327 4948 75336
rect 4896 75293 4905 75327
rect 4905 75293 4939 75327
rect 4939 75293 4948 75327
rect 4896 75284 4948 75293
rect 3976 75216 4028 75268
rect 2964 75148 3016 75200
rect 4160 75191 4212 75200
rect 4160 75157 4169 75191
rect 4169 75157 4203 75191
rect 4203 75157 4212 75191
rect 4160 75148 4212 75157
rect 7288 75191 7340 75200
rect 7288 75157 7297 75191
rect 7297 75157 7331 75191
rect 7331 75157 7340 75191
rect 7288 75148 7340 75157
rect 4315 75046 4367 75098
rect 4379 75046 4431 75098
rect 4443 75046 4495 75098
rect 4507 75046 4559 75098
rect 10982 75046 11034 75098
rect 11046 75046 11098 75098
rect 11110 75046 11162 75098
rect 11174 75046 11226 75098
rect 17648 75046 17700 75098
rect 17712 75046 17764 75098
rect 17776 75046 17828 75098
rect 17840 75046 17892 75098
rect 5172 74944 5224 74996
rect 7012 74987 7064 74996
rect 7012 74953 7021 74987
rect 7021 74953 7055 74987
rect 7055 74953 7064 74987
rect 7012 74944 7064 74953
rect 2136 74851 2188 74860
rect 2136 74817 2145 74851
rect 2145 74817 2179 74851
rect 2179 74817 2188 74851
rect 2136 74808 2188 74817
rect 2228 74740 2280 74792
rect 2964 74783 3016 74792
rect 2964 74749 2973 74783
rect 2973 74749 3007 74783
rect 3007 74749 3016 74783
rect 2964 74740 3016 74749
rect 4896 74808 4948 74860
rect 3976 74740 4028 74792
rect 4160 74740 4212 74792
rect 4068 74672 4120 74724
rect 3976 74604 4028 74656
rect 4988 74740 5040 74792
rect 6736 74740 6788 74792
rect 7380 74672 7432 74724
rect 5448 74604 5500 74656
rect 7648 74502 7700 74554
rect 7712 74502 7764 74554
rect 7776 74502 7828 74554
rect 7840 74502 7892 74554
rect 14315 74502 14367 74554
rect 14379 74502 14431 74554
rect 14443 74502 14495 74554
rect 14507 74502 14559 74554
rect 4160 74400 4212 74452
rect 5540 74400 5592 74452
rect 6092 74400 6144 74452
rect 5908 74332 5960 74384
rect 7380 74332 7432 74384
rect 8300 74332 8352 74384
rect 2780 74264 2832 74316
rect 5356 74307 5408 74316
rect 5356 74273 5365 74307
rect 5365 74273 5399 74307
rect 5399 74273 5408 74307
rect 5356 74264 5408 74273
rect 7748 74307 7800 74316
rect 7748 74273 7757 74307
rect 7757 74273 7791 74307
rect 7791 74273 7800 74307
rect 7748 74264 7800 74273
rect 2136 74196 2188 74248
rect 2688 74239 2740 74248
rect 2688 74205 2697 74239
rect 2697 74205 2731 74239
rect 2731 74205 2740 74239
rect 2688 74196 2740 74205
rect 4988 74239 5040 74248
rect 4988 74205 4997 74239
rect 4997 74205 5031 74239
rect 5031 74205 5040 74239
rect 4988 74196 5040 74205
rect 5080 74128 5132 74180
rect 6460 74128 6512 74180
rect 7104 74128 7156 74180
rect 2228 74103 2280 74112
rect 2228 74069 2237 74103
rect 2237 74069 2271 74103
rect 2271 74069 2280 74103
rect 2228 74060 2280 74069
rect 5448 74103 5500 74112
rect 5448 74069 5457 74103
rect 5457 74069 5491 74103
rect 5491 74069 5500 74103
rect 5448 74060 5500 74069
rect 6552 74060 6604 74112
rect 10600 74060 10652 74112
rect 4315 73958 4367 74010
rect 4379 73958 4431 74010
rect 4443 73958 4495 74010
rect 4507 73958 4559 74010
rect 10982 73958 11034 74010
rect 11046 73958 11098 74010
rect 11110 73958 11162 74010
rect 11174 73958 11226 74010
rect 17648 73958 17700 74010
rect 17712 73958 17764 74010
rect 17776 73958 17828 74010
rect 17840 73958 17892 74010
rect 2136 73899 2188 73908
rect 2136 73865 2145 73899
rect 2145 73865 2179 73899
rect 2179 73865 2188 73899
rect 2136 73856 2188 73865
rect 2228 73856 2280 73908
rect 2780 73695 2832 73704
rect 2780 73661 2789 73695
rect 2789 73661 2823 73695
rect 2823 73661 2832 73695
rect 2780 73652 2832 73661
rect 5908 73788 5960 73840
rect 6092 73763 6144 73772
rect 6092 73729 6101 73763
rect 6101 73729 6135 73763
rect 6135 73729 6144 73763
rect 6092 73720 6144 73729
rect 6552 73720 6604 73772
rect 10692 73763 10744 73772
rect 10692 73729 10701 73763
rect 10701 73729 10735 73763
rect 10735 73729 10744 73763
rect 10692 73720 10744 73729
rect 4344 73652 4396 73704
rect 5080 73695 5132 73704
rect 5080 73661 5089 73695
rect 5089 73661 5123 73695
rect 5123 73661 5132 73695
rect 5080 73652 5132 73661
rect 5264 73695 5316 73704
rect 5264 73661 5273 73695
rect 5273 73661 5307 73695
rect 5307 73661 5316 73695
rect 5264 73652 5316 73661
rect 5356 73652 5408 73704
rect 7196 73652 7248 73704
rect 9312 73652 9364 73704
rect 10600 73695 10652 73704
rect 10600 73661 10609 73695
rect 10609 73661 10643 73695
rect 10643 73661 10652 73695
rect 10600 73652 10652 73661
rect 4252 73627 4304 73636
rect 4252 73593 4261 73627
rect 4261 73593 4295 73627
rect 4295 73593 4304 73627
rect 4252 73584 4304 73593
rect 7380 73584 7432 73636
rect 7748 73584 7800 73636
rect 11336 73652 11388 73704
rect 5908 73559 5960 73568
rect 5908 73525 5917 73559
rect 5917 73525 5951 73559
rect 5951 73525 5960 73559
rect 5908 73516 5960 73525
rect 6000 73516 6052 73568
rect 7648 73414 7700 73466
rect 7712 73414 7764 73466
rect 7776 73414 7828 73466
rect 7840 73414 7892 73466
rect 14315 73414 14367 73466
rect 14379 73414 14431 73466
rect 14443 73414 14495 73466
rect 14507 73414 14559 73466
rect 2780 73312 2832 73364
rect 9312 73355 9364 73364
rect 2872 73244 2924 73296
rect 4804 73287 4856 73296
rect 4804 73253 4813 73287
rect 4813 73253 4847 73287
rect 4847 73253 4856 73287
rect 4804 73244 4856 73253
rect 6184 73244 6236 73296
rect 7288 73244 7340 73296
rect 4344 73219 4396 73228
rect 2688 73108 2740 73160
rect 3516 73151 3568 73160
rect 3516 73117 3525 73151
rect 3525 73117 3559 73151
rect 3559 73117 3568 73151
rect 3516 73108 3568 73117
rect 3976 73151 4028 73160
rect 3976 73117 3985 73151
rect 3985 73117 4019 73151
rect 4019 73117 4028 73151
rect 3976 73108 4028 73117
rect 4344 73185 4353 73219
rect 4353 73185 4387 73219
rect 4387 73185 4396 73219
rect 4344 73176 4396 73185
rect 5448 73176 5500 73228
rect 6000 73176 6052 73228
rect 4988 73108 5040 73160
rect 5264 73108 5316 73160
rect 5816 73151 5868 73160
rect 5816 73117 5825 73151
rect 5825 73117 5859 73151
rect 5859 73117 5868 73151
rect 5816 73108 5868 73117
rect 6736 73108 6788 73160
rect 9312 73321 9321 73355
rect 9321 73321 9355 73355
rect 9355 73321 9364 73355
rect 9312 73312 9364 73321
rect 9220 73176 9272 73228
rect 9496 73176 9548 73228
rect 10048 73219 10100 73228
rect 10048 73185 10057 73219
rect 10057 73185 10091 73219
rect 10091 73185 10100 73219
rect 10048 73176 10100 73185
rect 3056 73040 3108 73092
rect 5080 73040 5132 73092
rect 6920 73083 6972 73092
rect 6920 73049 6929 73083
rect 6929 73049 6963 73083
rect 6963 73049 6972 73083
rect 6920 73040 6972 73049
rect 8300 73040 8352 73092
rect 9312 73040 9364 73092
rect 11612 73108 11664 73160
rect 4712 73015 4764 73024
rect 4712 72981 4721 73015
rect 4721 72981 4755 73015
rect 4755 72981 4764 73015
rect 4712 72972 4764 72981
rect 6460 73015 6512 73024
rect 6460 72981 6469 73015
rect 6469 72981 6503 73015
rect 6503 72981 6512 73015
rect 6460 72972 6512 72981
rect 8576 72972 8628 73024
rect 10876 72972 10928 73024
rect 4315 72870 4367 72922
rect 4379 72870 4431 72922
rect 4443 72870 4495 72922
rect 4507 72870 4559 72922
rect 10982 72870 11034 72922
rect 11046 72870 11098 72922
rect 11110 72870 11162 72922
rect 11174 72870 11226 72922
rect 17648 72870 17700 72922
rect 17712 72870 17764 72922
rect 17776 72870 17828 72922
rect 17840 72870 17892 72922
rect 2688 72811 2740 72820
rect 2688 72777 2697 72811
rect 2697 72777 2731 72811
rect 2731 72777 2740 72811
rect 2688 72768 2740 72777
rect 3056 72811 3108 72820
rect 3056 72777 3065 72811
rect 3065 72777 3099 72811
rect 3099 72777 3108 72811
rect 3056 72768 3108 72777
rect 3884 72811 3936 72820
rect 3884 72777 3893 72811
rect 3893 72777 3927 72811
rect 3927 72777 3936 72811
rect 3884 72768 3936 72777
rect 7012 72768 7064 72820
rect 8300 72768 8352 72820
rect 8576 72700 8628 72752
rect 10876 72700 10928 72752
rect 11336 72700 11388 72752
rect 4620 72632 4672 72684
rect 4712 72632 4764 72684
rect 5448 72632 5500 72684
rect 6092 72632 6144 72684
rect 10324 72675 10376 72684
rect 10324 72641 10333 72675
rect 10333 72641 10367 72675
rect 10367 72641 10376 72675
rect 10324 72632 10376 72641
rect 5264 72564 5316 72616
rect 6460 72564 6512 72616
rect 8024 72564 8076 72616
rect 10876 72607 10928 72616
rect 10876 72573 10885 72607
rect 10885 72573 10919 72607
rect 10919 72573 10928 72607
rect 10876 72564 10928 72573
rect 11612 72564 11664 72616
rect 11796 72607 11848 72616
rect 11796 72573 11805 72607
rect 11805 72573 11839 72607
rect 11839 72573 11848 72607
rect 11796 72564 11848 72573
rect 11980 72607 12032 72616
rect 11980 72573 11989 72607
rect 11989 72573 12023 72607
rect 12023 72573 12032 72607
rect 11980 72564 12032 72573
rect 12348 72564 12400 72616
rect 10048 72496 10100 72548
rect 3516 72428 3568 72480
rect 4068 72428 4120 72480
rect 5816 72471 5868 72480
rect 5816 72437 5825 72471
rect 5825 72437 5859 72471
rect 5859 72437 5868 72471
rect 5816 72428 5868 72437
rect 6184 72471 6236 72480
rect 6184 72437 6193 72471
rect 6193 72437 6227 72471
rect 6227 72437 6236 72471
rect 6184 72428 6236 72437
rect 9220 72471 9272 72480
rect 9220 72437 9229 72471
rect 9229 72437 9263 72471
rect 9263 72437 9272 72471
rect 9220 72428 9272 72437
rect 9680 72428 9732 72480
rect 10508 72428 10560 72480
rect 12532 72428 12584 72480
rect 7648 72326 7700 72378
rect 7712 72326 7764 72378
rect 7776 72326 7828 72378
rect 7840 72326 7892 72378
rect 14315 72326 14367 72378
rect 14379 72326 14431 72378
rect 14443 72326 14495 72378
rect 14507 72326 14559 72378
rect 4988 72267 5040 72276
rect 4988 72233 4997 72267
rect 4997 72233 5031 72267
rect 5031 72233 5040 72267
rect 4988 72224 5040 72233
rect 5540 72267 5592 72276
rect 5540 72233 5549 72267
rect 5549 72233 5583 72267
rect 5583 72233 5592 72267
rect 5540 72224 5592 72233
rect 6092 72224 6144 72276
rect 11980 72224 12032 72276
rect 2780 72088 2832 72140
rect 3240 72088 3292 72140
rect 3700 72088 3752 72140
rect 6552 72088 6604 72140
rect 6828 72088 6880 72140
rect 7104 72131 7156 72140
rect 7104 72097 7113 72131
rect 7113 72097 7147 72131
rect 7147 72097 7156 72131
rect 7104 72088 7156 72097
rect 9220 72088 9272 72140
rect 9312 72131 9364 72140
rect 9312 72097 9321 72131
rect 9321 72097 9355 72131
rect 9355 72097 9364 72131
rect 9680 72131 9732 72140
rect 9312 72088 9364 72097
rect 9680 72097 9689 72131
rect 9689 72097 9723 72131
rect 9723 72097 9732 72131
rect 9680 72088 9732 72097
rect 8116 72020 8168 72072
rect 8576 72063 8628 72072
rect 8576 72029 8585 72063
rect 8585 72029 8619 72063
rect 8619 72029 8628 72063
rect 8576 72020 8628 72029
rect 8852 72063 8904 72072
rect 8852 72029 8861 72063
rect 8861 72029 8895 72063
rect 8895 72029 8904 72063
rect 8852 72020 8904 72029
rect 5908 71952 5960 72004
rect 6736 71952 6788 72004
rect 7196 71952 7248 72004
rect 8944 71952 8996 72004
rect 8208 71884 8260 71936
rect 11336 71884 11388 71936
rect 4315 71782 4367 71834
rect 4379 71782 4431 71834
rect 4443 71782 4495 71834
rect 4507 71782 4559 71834
rect 10982 71782 11034 71834
rect 11046 71782 11098 71834
rect 11110 71782 11162 71834
rect 11174 71782 11226 71834
rect 17648 71782 17700 71834
rect 17712 71782 17764 71834
rect 17776 71782 17828 71834
rect 17840 71782 17892 71834
rect 3240 71723 3292 71732
rect 3240 71689 3249 71723
rect 3249 71689 3283 71723
rect 3283 71689 3292 71723
rect 3240 71680 3292 71689
rect 5264 71680 5316 71732
rect 6828 71723 6880 71732
rect 6828 71689 6837 71723
rect 6837 71689 6871 71723
rect 6871 71689 6880 71723
rect 6828 71680 6880 71689
rect 8668 71680 8720 71732
rect 9312 71680 9364 71732
rect 17500 71723 17552 71732
rect 17500 71689 17509 71723
rect 17509 71689 17543 71723
rect 17543 71689 17552 71723
rect 17500 71680 17552 71689
rect 5448 71544 5500 71596
rect 6092 71544 6144 71596
rect 6552 71544 6604 71596
rect 10600 71587 10652 71596
rect 5080 71519 5132 71528
rect 5080 71485 5089 71519
rect 5089 71485 5123 71519
rect 5123 71485 5132 71519
rect 5080 71476 5132 71485
rect 8208 71519 8260 71528
rect 3700 71383 3752 71392
rect 3700 71349 3709 71383
rect 3709 71349 3743 71383
rect 3743 71349 3752 71383
rect 3700 71340 3752 71349
rect 7472 71383 7524 71392
rect 7472 71349 7481 71383
rect 7481 71349 7515 71383
rect 7515 71349 7524 71383
rect 8208 71485 8217 71519
rect 8217 71485 8251 71519
rect 8251 71485 8260 71519
rect 8208 71476 8260 71485
rect 8392 71476 8444 71528
rect 10600 71553 10609 71587
rect 10609 71553 10643 71587
rect 10643 71553 10652 71587
rect 10600 71544 10652 71553
rect 8852 71476 8904 71528
rect 11336 71544 11388 71596
rect 11428 71519 11480 71528
rect 11428 71485 11437 71519
rect 11437 71485 11471 71519
rect 11471 71485 11480 71519
rect 11704 71519 11756 71528
rect 11428 71476 11480 71485
rect 11704 71485 11713 71519
rect 11713 71485 11747 71519
rect 11747 71485 11756 71519
rect 11704 71476 11756 71485
rect 11888 71519 11940 71528
rect 11888 71485 11897 71519
rect 11897 71485 11931 71519
rect 11931 71485 11940 71519
rect 11888 71476 11940 71485
rect 12808 71519 12860 71528
rect 12808 71485 12817 71519
rect 12817 71485 12851 71519
rect 12851 71485 12860 71519
rect 12808 71476 12860 71485
rect 16120 71519 16172 71528
rect 16120 71485 16129 71519
rect 16129 71485 16163 71519
rect 16163 71485 16172 71519
rect 16120 71476 16172 71485
rect 8760 71451 8812 71460
rect 8760 71417 8769 71451
rect 8769 71417 8803 71451
rect 8803 71417 8812 71451
rect 8760 71408 8812 71417
rect 11336 71408 11388 71460
rect 7472 71340 7524 71349
rect 9220 71340 9272 71392
rect 11704 71340 11756 71392
rect 16028 71383 16080 71392
rect 16028 71349 16037 71383
rect 16037 71349 16071 71383
rect 16071 71349 16080 71383
rect 16028 71340 16080 71349
rect 7648 71238 7700 71290
rect 7712 71238 7764 71290
rect 7776 71238 7828 71290
rect 7840 71238 7892 71290
rect 14315 71238 14367 71290
rect 14379 71238 14431 71290
rect 14443 71238 14495 71290
rect 14507 71238 14559 71290
rect 5448 71179 5500 71188
rect 5448 71145 5457 71179
rect 5457 71145 5491 71179
rect 5491 71145 5500 71179
rect 5448 71136 5500 71145
rect 8576 71136 8628 71188
rect 9588 71136 9640 71188
rect 11888 71136 11940 71188
rect 10784 71068 10836 71120
rect 11428 71068 11480 71120
rect 4528 71000 4580 71052
rect 4712 71043 4764 71052
rect 4712 71009 4721 71043
rect 4721 71009 4755 71043
rect 4755 71009 4764 71043
rect 4712 71000 4764 71009
rect 5080 71000 5132 71052
rect 6736 71000 6788 71052
rect 8116 71000 8168 71052
rect 8760 71000 8812 71052
rect 6828 70975 6880 70984
rect 6828 70941 6837 70975
rect 6837 70941 6871 70975
rect 6871 70941 6880 70975
rect 6828 70932 6880 70941
rect 9588 70975 9640 70984
rect 9588 70941 9597 70975
rect 9597 70941 9631 70975
rect 9631 70941 9640 70975
rect 9588 70932 9640 70941
rect 4160 70907 4212 70916
rect 4160 70873 4169 70907
rect 4169 70873 4203 70907
rect 4203 70873 4212 70907
rect 4160 70864 4212 70873
rect 8392 70796 8444 70848
rect 10140 70796 10192 70848
rect 10232 70839 10284 70848
rect 10232 70805 10241 70839
rect 10241 70805 10275 70839
rect 10275 70805 10284 70839
rect 10232 70796 10284 70805
rect 11980 70796 12032 70848
rect 16120 70839 16172 70848
rect 16120 70805 16129 70839
rect 16129 70805 16163 70839
rect 16163 70805 16172 70839
rect 16120 70796 16172 70805
rect 4315 70694 4367 70746
rect 4379 70694 4431 70746
rect 4443 70694 4495 70746
rect 4507 70694 4559 70746
rect 10982 70694 11034 70746
rect 11046 70694 11098 70746
rect 11110 70694 11162 70746
rect 11174 70694 11226 70746
rect 17648 70694 17700 70746
rect 17712 70694 17764 70746
rect 17776 70694 17828 70746
rect 17840 70694 17892 70746
rect 1492 70592 1544 70644
rect 2780 70592 2832 70644
rect 4712 70592 4764 70644
rect 5540 70592 5592 70644
rect 8576 70592 8628 70644
rect 10324 70592 10376 70644
rect 10784 70592 10836 70644
rect 11704 70592 11756 70644
rect 5724 70499 5776 70508
rect 5724 70465 5733 70499
rect 5733 70465 5767 70499
rect 5767 70465 5776 70499
rect 7840 70499 7892 70508
rect 5724 70456 5776 70465
rect 5908 70431 5960 70440
rect 5908 70397 5917 70431
rect 5917 70397 5951 70431
rect 5951 70397 5960 70431
rect 5908 70388 5960 70397
rect 7840 70465 7849 70499
rect 7849 70465 7883 70499
rect 7883 70465 7892 70499
rect 7840 70456 7892 70465
rect 8116 70456 8168 70508
rect 6828 70388 6880 70440
rect 8392 70388 8444 70440
rect 8576 70431 8628 70440
rect 8576 70397 8585 70431
rect 8585 70397 8619 70431
rect 8619 70397 8628 70431
rect 8576 70388 8628 70397
rect 9772 70388 9824 70440
rect 10232 70456 10284 70508
rect 10784 70499 10836 70508
rect 10140 70431 10192 70440
rect 10140 70397 10149 70431
rect 10149 70397 10183 70431
rect 10183 70397 10192 70431
rect 10140 70388 10192 70397
rect 10416 70388 10468 70440
rect 10784 70465 10793 70499
rect 10793 70465 10827 70499
rect 10827 70465 10836 70499
rect 10784 70456 10836 70465
rect 11704 70388 11756 70440
rect 11980 70431 12032 70440
rect 11980 70397 11989 70431
rect 11989 70397 12023 70431
rect 12023 70397 12032 70431
rect 11980 70388 12032 70397
rect 12072 70388 12124 70440
rect 1768 70252 1820 70304
rect 4068 70252 4120 70304
rect 4620 70295 4672 70304
rect 4620 70261 4629 70295
rect 4629 70261 4663 70295
rect 4663 70261 4672 70295
rect 4620 70252 4672 70261
rect 7472 70295 7524 70304
rect 7472 70261 7481 70295
rect 7481 70261 7515 70295
rect 7515 70261 7524 70295
rect 7472 70252 7524 70261
rect 8024 70252 8076 70304
rect 9588 70252 9640 70304
rect 10140 70252 10192 70304
rect 11796 70252 11848 70304
rect 7648 70150 7700 70202
rect 7712 70150 7764 70202
rect 7776 70150 7828 70202
rect 7840 70150 7892 70202
rect 14315 70150 14367 70202
rect 14379 70150 14431 70202
rect 14443 70150 14495 70202
rect 14507 70150 14559 70202
rect 6736 70048 6788 70100
rect 8760 70091 8812 70100
rect 8760 70057 8769 70091
rect 8769 70057 8803 70091
rect 8803 70057 8812 70091
rect 8760 70048 8812 70057
rect 1492 69955 1544 69964
rect 1492 69921 1501 69955
rect 1501 69921 1535 69955
rect 1535 69921 1544 69955
rect 1492 69912 1544 69921
rect 4804 69912 4856 69964
rect 7380 69912 7432 69964
rect 8208 69912 8260 69964
rect 9956 69980 10008 70032
rect 9680 69955 9732 69964
rect 9680 69921 9689 69955
rect 9689 69921 9723 69955
rect 9723 69921 9732 69955
rect 9680 69912 9732 69921
rect 1768 69887 1820 69896
rect 1768 69853 1777 69887
rect 1777 69853 1811 69887
rect 1811 69853 1820 69887
rect 1768 69844 1820 69853
rect 6552 69844 6604 69896
rect 9772 69887 9824 69896
rect 9772 69853 9781 69887
rect 9781 69853 9815 69887
rect 9815 69853 9824 69887
rect 9772 69844 9824 69853
rect 10140 69912 10192 69964
rect 10416 69912 10468 69964
rect 9864 69776 9916 69828
rect 11980 69776 12032 69828
rect 2504 69708 2556 69760
rect 4620 69708 4672 69760
rect 5264 69751 5316 69760
rect 5264 69717 5273 69751
rect 5273 69717 5307 69751
rect 5307 69717 5316 69751
rect 5264 69708 5316 69717
rect 5908 69708 5960 69760
rect 8392 69751 8444 69760
rect 8392 69717 8401 69751
rect 8401 69717 8435 69751
rect 8435 69717 8444 69751
rect 8392 69708 8444 69717
rect 10416 69708 10468 69760
rect 12072 69708 12124 69760
rect 4315 69606 4367 69658
rect 4379 69606 4431 69658
rect 4443 69606 4495 69658
rect 4507 69606 4559 69658
rect 10982 69606 11034 69658
rect 11046 69606 11098 69658
rect 11110 69606 11162 69658
rect 11174 69606 11226 69658
rect 17648 69606 17700 69658
rect 17712 69606 17764 69658
rect 17776 69606 17828 69658
rect 17840 69606 17892 69658
rect 5816 69504 5868 69556
rect 9496 69504 9548 69556
rect 4160 69479 4212 69488
rect 4160 69445 4169 69479
rect 4169 69445 4203 69479
rect 4203 69445 4212 69479
rect 4160 69436 4212 69445
rect 6736 69436 6788 69488
rect 2504 69368 2556 69420
rect 5816 69411 5868 69420
rect 5816 69377 5825 69411
rect 5825 69377 5859 69411
rect 5859 69377 5868 69411
rect 5816 69368 5868 69377
rect 12072 69436 12124 69488
rect 7472 69368 7524 69420
rect 11888 69368 11940 69420
rect 2596 69300 2648 69352
rect 4068 69343 4120 69352
rect 1768 69232 1820 69284
rect 2228 69164 2280 69216
rect 2596 69164 2648 69216
rect 3056 69207 3108 69216
rect 3056 69173 3065 69207
rect 3065 69173 3099 69207
rect 3099 69173 3108 69207
rect 3056 69164 3108 69173
rect 3608 69164 3660 69216
rect 3700 69164 3752 69216
rect 4068 69309 4077 69343
rect 4077 69309 4111 69343
rect 4111 69309 4120 69343
rect 4068 69300 4120 69309
rect 4620 69343 4672 69352
rect 4620 69309 4629 69343
rect 4629 69309 4663 69343
rect 4663 69309 4672 69343
rect 4620 69300 4672 69309
rect 6368 69343 6420 69352
rect 6368 69309 6377 69343
rect 6377 69309 6411 69343
rect 6411 69309 6420 69343
rect 6368 69300 6420 69309
rect 6644 69343 6696 69352
rect 6644 69309 6653 69343
rect 6653 69309 6687 69343
rect 6687 69309 6696 69343
rect 6644 69300 6696 69309
rect 7196 69300 7248 69352
rect 8208 69343 8260 69352
rect 8208 69309 8217 69343
rect 8217 69309 8251 69343
rect 8251 69309 8260 69343
rect 8208 69300 8260 69309
rect 9956 69343 10008 69352
rect 9956 69309 9965 69343
rect 9965 69309 9999 69343
rect 9999 69309 10008 69343
rect 9956 69300 10008 69309
rect 10140 69343 10192 69352
rect 10140 69309 10149 69343
rect 10149 69309 10183 69343
rect 10183 69309 10192 69343
rect 10140 69300 10192 69309
rect 9680 69232 9732 69284
rect 4804 69164 4856 69216
rect 7380 69164 7432 69216
rect 9496 69207 9548 69216
rect 9496 69173 9505 69207
rect 9505 69173 9539 69207
rect 9539 69173 9548 69207
rect 11980 69300 12032 69352
rect 11796 69232 11848 69284
rect 12348 69232 12400 69284
rect 9496 69164 9548 69173
rect 11060 69164 11112 69216
rect 7648 69062 7700 69114
rect 7712 69062 7764 69114
rect 7776 69062 7828 69114
rect 7840 69062 7892 69114
rect 14315 69062 14367 69114
rect 14379 69062 14431 69114
rect 14443 69062 14495 69114
rect 14507 69062 14559 69114
rect 5540 69003 5592 69012
rect 5540 68969 5549 69003
rect 5549 68969 5583 69003
rect 5583 68969 5592 69003
rect 5540 68960 5592 68969
rect 6000 68960 6052 69012
rect 6644 68960 6696 69012
rect 3516 68935 3568 68944
rect 3516 68901 3525 68935
rect 3525 68901 3559 68935
rect 3559 68901 3568 68935
rect 3516 68892 3568 68901
rect 9496 68892 9548 68944
rect 2228 68867 2280 68876
rect 2228 68833 2237 68867
rect 2237 68833 2271 68867
rect 2271 68833 2280 68867
rect 2228 68824 2280 68833
rect 2504 68867 2556 68876
rect 2504 68833 2513 68867
rect 2513 68833 2547 68867
rect 2547 68833 2556 68867
rect 2504 68824 2556 68833
rect 3884 68824 3936 68876
rect 5356 68867 5408 68876
rect 5356 68833 5365 68867
rect 5365 68833 5399 68867
rect 5399 68833 5408 68867
rect 5356 68824 5408 68833
rect 8024 68867 8076 68876
rect 8024 68833 8033 68867
rect 8033 68833 8067 68867
rect 8067 68833 8076 68867
rect 8024 68824 8076 68833
rect 8576 68824 8628 68876
rect 14096 68892 14148 68944
rect 1676 68799 1728 68808
rect 1676 68765 1685 68799
rect 1685 68765 1719 68799
rect 1719 68765 1728 68799
rect 1676 68756 1728 68765
rect 2780 68756 2832 68808
rect 4068 68799 4120 68808
rect 4068 68765 4077 68799
rect 4077 68765 4111 68799
rect 4111 68765 4120 68799
rect 4068 68756 4120 68765
rect 4988 68756 5040 68808
rect 7012 68756 7064 68808
rect 8300 68799 8352 68808
rect 5080 68688 5132 68740
rect 6368 68688 6420 68740
rect 6920 68688 6972 68740
rect 8300 68765 8309 68799
rect 8309 68765 8343 68799
rect 8343 68765 8352 68799
rect 8300 68756 8352 68765
rect 8024 68688 8076 68740
rect 10048 68799 10100 68808
rect 10048 68765 10057 68799
rect 10057 68765 10091 68799
rect 10091 68765 10100 68799
rect 10048 68756 10100 68765
rect 10508 68824 10560 68876
rect 12440 68867 12492 68876
rect 12440 68833 12449 68867
rect 12449 68833 12483 68867
rect 12483 68833 12492 68867
rect 12440 68824 12492 68833
rect 13912 68824 13964 68876
rect 15016 68756 15068 68808
rect 15936 68756 15988 68808
rect 16120 68756 16172 68808
rect 9956 68688 10008 68740
rect 10692 68688 10744 68740
rect 1768 68620 1820 68672
rect 2136 68620 2188 68672
rect 3608 68620 3660 68672
rect 6092 68620 6144 68672
rect 6552 68663 6604 68672
rect 6552 68629 6561 68663
rect 6561 68629 6595 68663
rect 6595 68629 6604 68663
rect 6552 68620 6604 68629
rect 7380 68620 7432 68672
rect 9220 68663 9272 68672
rect 9220 68629 9229 68663
rect 9229 68629 9263 68663
rect 9263 68629 9272 68663
rect 9220 68620 9272 68629
rect 9864 68620 9916 68672
rect 11428 68620 11480 68672
rect 11612 68663 11664 68672
rect 11612 68629 11621 68663
rect 11621 68629 11655 68663
rect 11655 68629 11664 68663
rect 11612 68620 11664 68629
rect 12072 68663 12124 68672
rect 12072 68629 12081 68663
rect 12081 68629 12115 68663
rect 12115 68629 12124 68663
rect 12072 68620 12124 68629
rect 12624 68663 12676 68672
rect 12624 68629 12633 68663
rect 12633 68629 12667 68663
rect 12667 68629 12676 68663
rect 12624 68620 12676 68629
rect 12808 68620 12860 68672
rect 13360 68663 13412 68672
rect 13360 68629 13369 68663
rect 13369 68629 13403 68663
rect 13403 68629 13412 68663
rect 13360 68620 13412 68629
rect 16120 68663 16172 68672
rect 16120 68629 16129 68663
rect 16129 68629 16163 68663
rect 16163 68629 16172 68663
rect 16120 68620 16172 68629
rect 4315 68518 4367 68570
rect 4379 68518 4431 68570
rect 4443 68518 4495 68570
rect 4507 68518 4559 68570
rect 10982 68518 11034 68570
rect 11046 68518 11098 68570
rect 11110 68518 11162 68570
rect 11174 68518 11226 68570
rect 17648 68518 17700 68570
rect 17712 68518 17764 68570
rect 17776 68518 17828 68570
rect 17840 68518 17892 68570
rect 6736 68459 6788 68468
rect 6736 68425 6745 68459
rect 6745 68425 6779 68459
rect 6779 68425 6788 68459
rect 6736 68416 6788 68425
rect 8576 68416 8628 68468
rect 17500 68459 17552 68468
rect 17500 68425 17509 68459
rect 17509 68425 17543 68459
rect 17543 68425 17552 68459
rect 17500 68416 17552 68425
rect 7932 68348 7984 68400
rect 9956 68348 10008 68400
rect 10324 68348 10376 68400
rect 10784 68348 10836 68400
rect 11244 68348 11296 68400
rect 11336 68348 11388 68400
rect 1492 68323 1544 68332
rect 1492 68289 1501 68323
rect 1501 68289 1535 68323
rect 1535 68289 1544 68323
rect 1492 68280 1544 68289
rect 1768 68323 1820 68332
rect 1768 68289 1777 68323
rect 1777 68289 1811 68323
rect 1811 68289 1820 68323
rect 1768 68280 1820 68289
rect 4988 68280 5040 68332
rect 10692 68280 10744 68332
rect 2780 68144 2832 68196
rect 5080 68212 5132 68264
rect 5632 68212 5684 68264
rect 7380 68212 7432 68264
rect 11612 68280 11664 68332
rect 5356 68144 5408 68196
rect 8484 68144 8536 68196
rect 8852 68144 8904 68196
rect 11152 68255 11204 68264
rect 11152 68221 11161 68255
rect 11161 68221 11195 68255
rect 11195 68221 11204 68255
rect 11152 68212 11204 68221
rect 11428 68212 11480 68264
rect 10140 68144 10192 68196
rect 10784 68144 10836 68196
rect 2872 68119 2924 68128
rect 2872 68085 2881 68119
rect 2881 68085 2915 68119
rect 2915 68085 2924 68119
rect 2872 68076 2924 68085
rect 3700 68076 3752 68128
rect 3884 68076 3936 68128
rect 8024 68119 8076 68128
rect 8024 68085 8033 68119
rect 8033 68085 8067 68119
rect 8067 68085 8076 68119
rect 8024 68076 8076 68085
rect 8392 68076 8444 68128
rect 9496 68119 9548 68128
rect 9496 68085 9505 68119
rect 9505 68085 9539 68119
rect 9539 68085 9548 68119
rect 9496 68076 9548 68085
rect 9772 68076 9824 68128
rect 11336 68076 11388 68128
rect 12624 68212 12676 68264
rect 12808 68255 12860 68264
rect 12808 68221 12817 68255
rect 12817 68221 12851 68255
rect 12851 68221 12860 68255
rect 12808 68212 12860 68221
rect 13176 68255 13228 68264
rect 13176 68221 13185 68255
rect 13185 68221 13219 68255
rect 13219 68221 13228 68255
rect 13176 68212 13228 68221
rect 13360 68255 13412 68264
rect 13360 68221 13369 68255
rect 13369 68221 13403 68255
rect 13403 68221 13412 68255
rect 13360 68212 13412 68221
rect 16120 68255 16172 68264
rect 16120 68221 16129 68255
rect 16129 68221 16163 68255
rect 16163 68221 16172 68255
rect 16120 68212 16172 68221
rect 16396 68255 16448 68264
rect 16396 68221 16405 68255
rect 16405 68221 16439 68255
rect 16439 68221 16448 68255
rect 16396 68212 16448 68221
rect 12440 68119 12492 68128
rect 12440 68085 12449 68119
rect 12449 68085 12483 68119
rect 12483 68085 12492 68119
rect 12440 68076 12492 68085
rect 13912 68119 13964 68128
rect 13912 68085 13921 68119
rect 13921 68085 13955 68119
rect 13955 68085 13964 68119
rect 13912 68076 13964 68085
rect 14096 68076 14148 68128
rect 15108 68076 15160 68128
rect 7648 67974 7700 68026
rect 7712 67974 7764 68026
rect 7776 67974 7828 68026
rect 7840 67974 7892 68026
rect 14315 67974 14367 68026
rect 14379 67974 14431 68026
rect 14443 67974 14495 68026
rect 14507 67974 14559 68026
rect 2228 67872 2280 67924
rect 3884 67872 3936 67924
rect 4068 67915 4120 67924
rect 4068 67881 4077 67915
rect 4077 67881 4111 67915
rect 4111 67881 4120 67915
rect 4068 67872 4120 67881
rect 4896 67915 4948 67924
rect 4896 67881 4905 67915
rect 4905 67881 4939 67915
rect 4939 67881 4948 67915
rect 4896 67872 4948 67881
rect 8300 67872 8352 67924
rect 8392 67872 8444 67924
rect 10416 67872 10468 67924
rect 1492 67804 1544 67856
rect 2504 67804 2556 67856
rect 2872 67736 2924 67788
rect 3332 67736 3384 67788
rect 3700 67736 3752 67788
rect 4068 67736 4120 67788
rect 1768 67711 1820 67720
rect 1768 67677 1777 67711
rect 1777 67677 1811 67711
rect 1811 67677 1820 67711
rect 1768 67668 1820 67677
rect 2320 67711 2372 67720
rect 2320 67677 2329 67711
rect 2329 67677 2363 67711
rect 2363 67677 2372 67711
rect 2320 67668 2372 67677
rect 2780 67711 2832 67720
rect 2780 67677 2789 67711
rect 2789 67677 2823 67711
rect 2823 67677 2832 67711
rect 2780 67668 2832 67677
rect 4896 67736 4948 67788
rect 8116 67804 8168 67856
rect 10140 67804 10192 67856
rect 10324 67804 10376 67856
rect 7472 67779 7524 67788
rect 7472 67745 7481 67779
rect 7481 67745 7515 67779
rect 7515 67745 7524 67779
rect 7472 67736 7524 67745
rect 8944 67736 8996 67788
rect 10692 67736 10744 67788
rect 11152 67804 11204 67856
rect 11612 67804 11664 67856
rect 11336 67779 11388 67788
rect 11336 67745 11345 67779
rect 11345 67745 11379 67779
rect 11379 67745 11388 67779
rect 11336 67736 11388 67745
rect 13176 67779 13228 67788
rect 3792 67643 3844 67652
rect 3792 67609 3801 67643
rect 3801 67609 3835 67643
rect 3835 67609 3844 67643
rect 3792 67600 3844 67609
rect 4712 67643 4764 67652
rect 4712 67609 4721 67643
rect 4721 67609 4755 67643
rect 4755 67609 4764 67643
rect 4712 67600 4764 67609
rect 5172 67532 5224 67584
rect 6184 67575 6236 67584
rect 6184 67541 6193 67575
rect 6193 67541 6227 67575
rect 6227 67541 6236 67575
rect 6184 67532 6236 67541
rect 8024 67532 8076 67584
rect 13176 67745 13185 67779
rect 13185 67745 13219 67779
rect 13219 67745 13228 67779
rect 13176 67736 13228 67745
rect 15292 67736 15344 67788
rect 13728 67668 13780 67720
rect 15936 67668 15988 67720
rect 17132 67711 17184 67720
rect 17132 67677 17141 67711
rect 17141 67677 17175 67711
rect 17175 67677 17184 67711
rect 17132 67668 17184 67677
rect 9864 67532 9916 67584
rect 10876 67532 10928 67584
rect 11336 67532 11388 67584
rect 13084 67532 13136 67584
rect 4315 67430 4367 67482
rect 4379 67430 4431 67482
rect 4443 67430 4495 67482
rect 4507 67430 4559 67482
rect 10982 67430 11034 67482
rect 11046 67430 11098 67482
rect 11110 67430 11162 67482
rect 11174 67430 11226 67482
rect 17648 67430 17700 67482
rect 17712 67430 17764 67482
rect 17776 67430 17828 67482
rect 17840 67430 17892 67482
rect 2872 67371 2924 67380
rect 2872 67337 2881 67371
rect 2881 67337 2915 67371
rect 2915 67337 2924 67371
rect 2872 67328 2924 67337
rect 4896 67371 4948 67380
rect 4896 67337 4905 67371
rect 4905 67337 4939 67371
rect 4939 67337 4948 67371
rect 4896 67328 4948 67337
rect 6736 67371 6788 67380
rect 6736 67337 6745 67371
rect 6745 67337 6779 67371
rect 6779 67337 6788 67371
rect 6736 67328 6788 67337
rect 6920 67328 6972 67380
rect 13176 67328 13228 67380
rect 3976 67192 4028 67244
rect 14372 67303 14424 67312
rect 14372 67269 14381 67303
rect 14381 67269 14415 67303
rect 14415 67269 14424 67303
rect 14372 67260 14424 67269
rect 10508 67235 10560 67244
rect 10508 67201 10517 67235
rect 10517 67201 10551 67235
rect 10551 67201 10560 67235
rect 10508 67192 10560 67201
rect 11980 67192 12032 67244
rect 1860 67167 1912 67176
rect 1860 67133 1869 67167
rect 1869 67133 1903 67167
rect 1903 67133 1912 67167
rect 1860 67124 1912 67133
rect 4252 67167 4304 67176
rect 4252 67133 4261 67167
rect 4261 67133 4295 67167
rect 4295 67133 4304 67167
rect 4252 67124 4304 67133
rect 5632 67124 5684 67176
rect 5908 67167 5960 67176
rect 5908 67133 5917 67167
rect 5917 67133 5951 67167
rect 5951 67133 5960 67167
rect 5908 67124 5960 67133
rect 6184 67167 6236 67176
rect 6184 67133 6193 67167
rect 6193 67133 6227 67167
rect 6227 67133 6236 67167
rect 6184 67124 6236 67133
rect 7196 67167 7248 67176
rect 7196 67133 7205 67167
rect 7205 67133 7239 67167
rect 7239 67133 7248 67167
rect 7196 67124 7248 67133
rect 2780 66988 2832 67040
rect 3332 66988 3384 67040
rect 6828 67056 6880 67108
rect 8024 67124 8076 67176
rect 9680 67167 9732 67176
rect 9680 67133 9689 67167
rect 9689 67133 9723 67167
rect 9723 67133 9732 67167
rect 9680 67124 9732 67133
rect 10416 67167 10468 67176
rect 5172 67031 5224 67040
rect 5172 66997 5181 67031
rect 5181 66997 5215 67031
rect 5215 66997 5224 67031
rect 5172 66988 5224 66997
rect 7472 66988 7524 67040
rect 8576 67031 8628 67040
rect 8576 66997 8585 67031
rect 8585 66997 8619 67031
rect 8619 66997 8628 67031
rect 8576 66988 8628 66997
rect 8944 66988 8996 67040
rect 9496 67031 9548 67040
rect 9496 66997 9505 67031
rect 9505 66997 9539 67031
rect 9539 66997 9548 67031
rect 10416 67133 10425 67167
rect 10425 67133 10459 67167
rect 10459 67133 10468 67167
rect 10416 67124 10468 67133
rect 12164 67167 12216 67176
rect 12164 67133 12173 67167
rect 12173 67133 12207 67167
rect 12207 67133 12216 67167
rect 12164 67124 12216 67133
rect 12256 67056 12308 67108
rect 12440 67056 12492 67108
rect 12992 67124 13044 67176
rect 15384 67124 15436 67176
rect 15936 67124 15988 67176
rect 16488 67124 16540 67176
rect 13268 67099 13320 67108
rect 13268 67065 13277 67099
rect 13277 67065 13311 67099
rect 13311 67065 13320 67099
rect 13268 67056 13320 67065
rect 9496 66988 9548 66997
rect 11336 66988 11388 67040
rect 11612 67031 11664 67040
rect 11612 66997 11621 67031
rect 11621 66997 11655 67031
rect 11655 66997 11664 67031
rect 11612 66988 11664 66997
rect 11980 67031 12032 67040
rect 11980 66997 11989 67031
rect 11989 66997 12023 67031
rect 12023 66997 12032 67031
rect 11980 66988 12032 66997
rect 13820 66988 13872 67040
rect 15292 66988 15344 67040
rect 17500 67031 17552 67040
rect 17500 66997 17509 67031
rect 17509 66997 17543 67031
rect 17543 66997 17552 67031
rect 17500 66988 17552 66997
rect 7648 66886 7700 66938
rect 7712 66886 7764 66938
rect 7776 66886 7828 66938
rect 7840 66886 7892 66938
rect 14315 66886 14367 66938
rect 14379 66886 14431 66938
rect 14443 66886 14495 66938
rect 14507 66886 14559 66938
rect 2320 66784 2372 66836
rect 2872 66784 2924 66836
rect 4252 66827 4304 66836
rect 4252 66793 4261 66827
rect 4261 66793 4295 66827
rect 4295 66793 4304 66827
rect 4252 66784 4304 66793
rect 8576 66784 8628 66836
rect 9680 66784 9732 66836
rect 15936 66784 15988 66836
rect 2136 66716 2188 66768
rect 11980 66716 12032 66768
rect 2596 66648 2648 66700
rect 3332 66648 3384 66700
rect 5264 66691 5316 66700
rect 5264 66657 5273 66691
rect 5273 66657 5307 66691
rect 5307 66657 5316 66691
rect 5264 66648 5316 66657
rect 5632 66648 5684 66700
rect 6552 66648 6604 66700
rect 6736 66648 6788 66700
rect 7104 66648 7156 66700
rect 7472 66691 7524 66700
rect 7472 66657 7481 66691
rect 7481 66657 7515 66691
rect 7515 66657 7524 66691
rect 7472 66648 7524 66657
rect 8208 66648 8260 66700
rect 9128 66648 9180 66700
rect 9588 66691 9640 66700
rect 9588 66657 9597 66691
rect 9597 66657 9631 66691
rect 9631 66657 9640 66691
rect 9588 66648 9640 66657
rect 9864 66691 9916 66700
rect 9864 66657 9873 66691
rect 9873 66657 9907 66691
rect 9907 66657 9916 66691
rect 9864 66648 9916 66657
rect 5908 66580 5960 66632
rect 9680 66623 9732 66632
rect 9680 66589 9689 66623
rect 9689 66589 9723 66623
rect 9723 66589 9732 66623
rect 9680 66580 9732 66589
rect 5080 66512 5132 66564
rect 6000 66512 6052 66564
rect 9220 66512 9272 66564
rect 12440 66691 12492 66700
rect 12440 66657 12449 66691
rect 12449 66657 12483 66691
rect 12483 66657 12492 66691
rect 12900 66691 12952 66700
rect 12440 66648 12492 66657
rect 12900 66657 12909 66691
rect 12909 66657 12943 66691
rect 12943 66657 12952 66691
rect 12900 66648 12952 66657
rect 14372 66648 14424 66700
rect 16120 66648 16172 66700
rect 12164 66580 12216 66632
rect 12532 66580 12584 66632
rect 12992 66580 13044 66632
rect 15200 66580 15252 66632
rect 16672 66623 16724 66632
rect 16672 66589 16681 66623
rect 16681 66589 16715 66623
rect 16715 66589 16724 66623
rect 16672 66580 16724 66589
rect 10416 66512 10468 66564
rect 1860 66444 1912 66496
rect 5172 66444 5224 66496
rect 6828 66444 6880 66496
rect 7288 66444 7340 66496
rect 8208 66444 8260 66496
rect 10692 66444 10744 66496
rect 12256 66487 12308 66496
rect 12256 66453 12265 66487
rect 12265 66453 12299 66487
rect 12299 66453 12308 66487
rect 12256 66444 12308 66453
rect 12532 66487 12584 66496
rect 12532 66453 12541 66487
rect 12541 66453 12575 66487
rect 12575 66453 12584 66487
rect 12532 66444 12584 66453
rect 4315 66342 4367 66394
rect 4379 66342 4431 66394
rect 4443 66342 4495 66394
rect 4507 66342 4559 66394
rect 10982 66342 11034 66394
rect 11046 66342 11098 66394
rect 11110 66342 11162 66394
rect 11174 66342 11226 66394
rect 17648 66342 17700 66394
rect 17712 66342 17764 66394
rect 17776 66342 17828 66394
rect 17840 66342 17892 66394
rect 2596 66240 2648 66292
rect 2872 66283 2924 66292
rect 2872 66249 2881 66283
rect 2881 66249 2915 66283
rect 2915 66249 2924 66283
rect 2872 66240 2924 66249
rect 5172 66240 5224 66292
rect 3424 66172 3476 66224
rect 7472 66240 7524 66292
rect 9496 66240 9548 66292
rect 10048 66240 10100 66292
rect 14004 66240 14056 66292
rect 14372 66283 14424 66292
rect 14372 66249 14381 66283
rect 14381 66249 14415 66283
rect 14415 66249 14424 66283
rect 14372 66240 14424 66249
rect 5632 66104 5684 66156
rect 9220 66172 9272 66224
rect 9864 66172 9916 66224
rect 2872 66036 2924 66088
rect 3608 66036 3660 66088
rect 5080 66079 5132 66088
rect 5080 66045 5089 66079
rect 5089 66045 5123 66079
rect 5123 66045 5132 66079
rect 5080 66036 5132 66045
rect 7288 66079 7340 66088
rect 7288 66045 7297 66079
rect 7297 66045 7331 66079
rect 7331 66045 7340 66079
rect 7288 66036 7340 66045
rect 8116 66079 8168 66088
rect 6828 65968 6880 66020
rect 8116 66045 8125 66079
rect 8125 66045 8159 66079
rect 8159 66045 8168 66079
rect 8116 66036 8168 66045
rect 8576 66079 8628 66088
rect 8576 66045 8585 66079
rect 8585 66045 8619 66079
rect 8619 66045 8628 66079
rect 8576 66036 8628 66045
rect 9588 66036 9640 66088
rect 10140 66172 10192 66224
rect 11060 66172 11112 66224
rect 11612 66172 11664 66224
rect 12440 66172 12492 66224
rect 13360 66104 13412 66156
rect 15476 66104 15528 66156
rect 8208 65968 8260 66020
rect 11980 66036 12032 66088
rect 12532 66036 12584 66088
rect 13268 66079 13320 66088
rect 13268 66045 13277 66079
rect 13277 66045 13311 66079
rect 13311 66045 13320 66079
rect 13268 66036 13320 66045
rect 15384 66036 15436 66088
rect 11796 65968 11848 66020
rect 12808 65968 12860 66020
rect 1860 65900 1912 65952
rect 2780 65900 2832 65952
rect 3332 65900 3384 65952
rect 4620 65900 4672 65952
rect 4896 65900 4948 65952
rect 7472 65900 7524 65952
rect 9128 65943 9180 65952
rect 9128 65909 9137 65943
rect 9137 65909 9171 65943
rect 9171 65909 9180 65943
rect 9128 65900 9180 65909
rect 9220 65900 9272 65952
rect 9680 65900 9732 65952
rect 9772 65900 9824 65952
rect 10048 65900 10100 65952
rect 10324 65943 10376 65952
rect 10324 65909 10333 65943
rect 10333 65909 10367 65943
rect 10367 65909 10376 65943
rect 10324 65900 10376 65909
rect 11244 65943 11296 65952
rect 11244 65909 11253 65943
rect 11253 65909 11287 65943
rect 11287 65909 11296 65943
rect 11244 65900 11296 65909
rect 11336 65900 11388 65952
rect 11612 65900 11664 65952
rect 12900 65900 12952 65952
rect 14740 65943 14792 65952
rect 14740 65909 14749 65943
rect 14749 65909 14783 65943
rect 14783 65909 14792 65943
rect 14740 65900 14792 65909
rect 15108 65900 15160 65952
rect 16580 65900 16632 65952
rect 7648 65798 7700 65850
rect 7712 65798 7764 65850
rect 7776 65798 7828 65850
rect 7840 65798 7892 65850
rect 14315 65798 14367 65850
rect 14379 65798 14431 65850
rect 14443 65798 14495 65850
rect 14507 65798 14559 65850
rect 2136 65696 2188 65748
rect 2320 65696 2372 65748
rect 8576 65696 8628 65748
rect 8760 65696 8812 65748
rect 10140 65696 10192 65748
rect 12532 65696 12584 65748
rect 13912 65696 13964 65748
rect 15384 65739 15436 65748
rect 15384 65705 15393 65739
rect 15393 65705 15427 65739
rect 15427 65705 15436 65739
rect 15384 65696 15436 65705
rect 16120 65739 16172 65748
rect 16120 65705 16129 65739
rect 16129 65705 16163 65739
rect 16163 65705 16172 65739
rect 16120 65696 16172 65705
rect 2504 65628 2556 65680
rect 2872 65628 2924 65680
rect 3332 65560 3384 65612
rect 9128 65628 9180 65680
rect 4804 65560 4856 65612
rect 7472 65603 7524 65612
rect 7472 65569 7481 65603
rect 7481 65569 7515 65603
rect 7515 65569 7524 65603
rect 7472 65560 7524 65569
rect 7932 65603 7984 65612
rect 7932 65569 7941 65603
rect 7941 65569 7975 65603
rect 7975 65569 7984 65603
rect 7932 65560 7984 65569
rect 5448 65492 5500 65544
rect 8116 65492 8168 65544
rect 3976 65424 4028 65476
rect 7472 65424 7524 65476
rect 8392 65560 8444 65612
rect 8760 65560 8812 65612
rect 10692 65560 10744 65612
rect 11336 65628 11388 65680
rect 13268 65628 13320 65680
rect 10600 65492 10652 65544
rect 12256 65560 12308 65612
rect 13176 65560 13228 65612
rect 14004 65560 14056 65612
rect 11520 65535 11572 65544
rect 11520 65501 11529 65535
rect 11529 65501 11563 65535
rect 11563 65501 11572 65535
rect 11520 65492 11572 65501
rect 11980 65492 12032 65544
rect 13636 65535 13688 65544
rect 13636 65501 13645 65535
rect 13645 65501 13679 65535
rect 13679 65501 13688 65535
rect 13636 65492 13688 65501
rect 10416 65424 10468 65476
rect 2228 65399 2280 65408
rect 2228 65365 2237 65399
rect 2237 65365 2271 65399
rect 2271 65365 2280 65399
rect 2228 65356 2280 65365
rect 3700 65399 3752 65408
rect 3700 65365 3709 65399
rect 3709 65365 3743 65399
rect 3743 65365 3752 65399
rect 3700 65356 3752 65365
rect 5080 65356 5132 65408
rect 5540 65399 5592 65408
rect 5540 65365 5549 65399
rect 5549 65365 5583 65399
rect 5583 65365 5592 65399
rect 5540 65356 5592 65365
rect 6092 65399 6144 65408
rect 6092 65365 6101 65399
rect 6101 65365 6135 65399
rect 6135 65365 6144 65399
rect 6092 65356 6144 65365
rect 9956 65356 10008 65408
rect 12256 65356 12308 65408
rect 4315 65254 4367 65306
rect 4379 65254 4431 65306
rect 4443 65254 4495 65306
rect 4507 65254 4559 65306
rect 10982 65254 11034 65306
rect 11046 65254 11098 65306
rect 11110 65254 11162 65306
rect 11174 65254 11226 65306
rect 17648 65254 17700 65306
rect 17712 65254 17764 65306
rect 17776 65254 17828 65306
rect 17840 65254 17892 65306
rect 3332 65152 3384 65204
rect 5264 65195 5316 65204
rect 5264 65161 5273 65195
rect 5273 65161 5307 65195
rect 5307 65161 5316 65195
rect 5264 65152 5316 65161
rect 4068 65084 4120 65136
rect 6092 65152 6144 65204
rect 6920 65152 6972 65204
rect 7932 65195 7984 65204
rect 7932 65161 7941 65195
rect 7941 65161 7975 65195
rect 7975 65161 7984 65195
rect 7932 65152 7984 65161
rect 9588 65152 9640 65204
rect 10600 65152 10652 65204
rect 13176 65195 13228 65204
rect 13176 65161 13185 65195
rect 13185 65161 13219 65195
rect 13219 65161 13228 65195
rect 13176 65152 13228 65161
rect 17500 65195 17552 65204
rect 17500 65161 17509 65195
rect 17509 65161 17543 65195
rect 17543 65161 17552 65195
rect 17500 65152 17552 65161
rect 2596 65016 2648 65068
rect 3700 65016 3752 65068
rect 1768 64948 1820 65000
rect 2228 64991 2280 65000
rect 2228 64957 2237 64991
rect 2237 64957 2271 64991
rect 2271 64957 2280 64991
rect 2228 64948 2280 64957
rect 5540 65016 5592 65068
rect 5816 65016 5868 65068
rect 2504 64880 2556 64932
rect 4712 64948 4764 65000
rect 8300 64948 8352 65000
rect 4896 64880 4948 64932
rect 8944 64948 8996 65000
rect 9956 64948 10008 65000
rect 10600 65059 10652 65068
rect 10600 65025 10609 65059
rect 10609 65025 10643 65059
rect 10643 65025 10652 65059
rect 10600 65016 10652 65025
rect 10692 64991 10744 65000
rect 10692 64957 10701 64991
rect 10701 64957 10735 64991
rect 10735 64957 10744 64991
rect 10692 64948 10744 64957
rect 8852 64880 8904 64932
rect 12348 64991 12400 65000
rect 12348 64957 12357 64991
rect 12357 64957 12391 64991
rect 12391 64957 12400 64991
rect 12348 64948 12400 64957
rect 14004 64948 14056 65000
rect 16120 64991 16172 65000
rect 16120 64957 16129 64991
rect 16129 64957 16163 64991
rect 16163 64957 16172 64991
rect 16120 64948 16172 64957
rect 16396 64991 16448 65000
rect 16396 64957 16405 64991
rect 16405 64957 16439 64991
rect 16439 64957 16448 64991
rect 16396 64948 16448 64957
rect 12716 64880 12768 64932
rect 12900 64880 12952 64932
rect 13636 64880 13688 64932
rect 15108 64880 15160 64932
rect 2872 64812 2924 64864
rect 7472 64812 7524 64864
rect 8484 64812 8536 64864
rect 8760 64855 8812 64864
rect 8760 64821 8769 64855
rect 8769 64821 8803 64855
rect 8803 64821 8812 64855
rect 8760 64812 8812 64821
rect 10140 64812 10192 64864
rect 7648 64710 7700 64762
rect 7712 64710 7764 64762
rect 7776 64710 7828 64762
rect 7840 64710 7892 64762
rect 14315 64710 14367 64762
rect 14379 64710 14431 64762
rect 14443 64710 14495 64762
rect 14507 64710 14559 64762
rect 3424 64608 3476 64660
rect 4068 64608 4120 64660
rect 6644 64651 6696 64660
rect 6644 64617 6653 64651
rect 6653 64617 6687 64651
rect 6687 64617 6696 64651
rect 6644 64608 6696 64617
rect 8392 64608 8444 64660
rect 9864 64608 9916 64660
rect 8484 64540 8536 64592
rect 2872 64472 2924 64524
rect 3884 64472 3936 64524
rect 3976 64472 4028 64524
rect 4620 64472 4672 64524
rect 7288 64472 7340 64524
rect 3056 64447 3108 64456
rect 3056 64413 3065 64447
rect 3065 64413 3099 64447
rect 3099 64413 3108 64447
rect 3056 64404 3108 64413
rect 6368 64404 6420 64456
rect 8300 64472 8352 64524
rect 8208 64404 8260 64456
rect 8576 64472 8628 64524
rect 9588 64472 9640 64524
rect 10140 64515 10192 64524
rect 10140 64481 10149 64515
rect 10149 64481 10183 64515
rect 10183 64481 10192 64515
rect 10140 64472 10192 64481
rect 10324 64515 10376 64524
rect 10324 64481 10333 64515
rect 10333 64481 10367 64515
rect 10367 64481 10376 64515
rect 10324 64472 10376 64481
rect 10784 64472 10836 64524
rect 13084 64472 13136 64524
rect 15108 64472 15160 64524
rect 16120 64472 16172 64524
rect 8668 64404 8720 64456
rect 11336 64404 11388 64456
rect 12992 64447 13044 64456
rect 12992 64413 13001 64447
rect 13001 64413 13035 64447
rect 13035 64413 13044 64447
rect 12992 64404 13044 64413
rect 14372 64447 14424 64456
rect 14372 64413 14381 64447
rect 14381 64413 14415 64447
rect 14415 64413 14424 64447
rect 14372 64404 14424 64413
rect 15660 64404 15712 64456
rect 16856 64447 16908 64456
rect 16856 64413 16865 64447
rect 16865 64413 16899 64447
rect 16899 64413 16908 64447
rect 16856 64404 16908 64413
rect 2688 64336 2740 64388
rect 7104 64336 7156 64388
rect 1768 64268 1820 64320
rect 2412 64268 2464 64320
rect 4896 64268 4948 64320
rect 5816 64311 5868 64320
rect 5816 64277 5825 64311
rect 5825 64277 5859 64311
rect 5859 64277 5868 64311
rect 5816 64268 5868 64277
rect 9312 64311 9364 64320
rect 9312 64277 9321 64311
rect 9321 64277 9355 64311
rect 9355 64277 9364 64311
rect 9312 64268 9364 64277
rect 9772 64311 9824 64320
rect 9772 64277 9781 64311
rect 9781 64277 9815 64311
rect 9815 64277 9824 64311
rect 9772 64268 9824 64277
rect 4315 64166 4367 64218
rect 4379 64166 4431 64218
rect 4443 64166 4495 64218
rect 4507 64166 4559 64218
rect 10982 64166 11034 64218
rect 11046 64166 11098 64218
rect 11110 64166 11162 64218
rect 11174 64166 11226 64218
rect 17648 64166 17700 64218
rect 17712 64166 17764 64218
rect 17776 64166 17828 64218
rect 17840 64166 17892 64218
rect 6368 64107 6420 64116
rect 6368 64073 6377 64107
rect 6377 64073 6411 64107
rect 6411 64073 6420 64107
rect 6368 64064 6420 64073
rect 10324 64064 10376 64116
rect 15108 64107 15160 64116
rect 15108 64073 15117 64107
rect 15117 64073 15151 64107
rect 15151 64073 15160 64107
rect 15108 64064 15160 64073
rect 2780 63996 2832 64048
rect 2688 63903 2740 63912
rect 2688 63869 2697 63903
rect 2697 63869 2731 63903
rect 2731 63869 2740 63903
rect 2688 63860 2740 63869
rect 4068 63996 4120 64048
rect 9312 63996 9364 64048
rect 10508 63996 10560 64048
rect 11336 63996 11388 64048
rect 4160 63928 4212 63980
rect 4712 63928 4764 63980
rect 6092 63928 6144 63980
rect 2136 63835 2188 63844
rect 2136 63801 2145 63835
rect 2145 63801 2179 63835
rect 2179 63801 2188 63835
rect 2136 63792 2188 63801
rect 2412 63792 2464 63844
rect 3608 63860 3660 63912
rect 5264 63903 5316 63912
rect 5264 63869 5273 63903
rect 5273 63869 5307 63903
rect 5307 63869 5316 63903
rect 5264 63860 5316 63869
rect 7104 63903 7156 63912
rect 3056 63792 3108 63844
rect 4068 63792 4120 63844
rect 4896 63792 4948 63844
rect 7104 63869 7113 63903
rect 7113 63869 7147 63903
rect 7147 63869 7156 63903
rect 7104 63860 7156 63869
rect 7932 63903 7984 63912
rect 7932 63869 7941 63903
rect 7941 63869 7975 63903
rect 7975 63869 7984 63903
rect 7932 63860 7984 63869
rect 8392 63928 8444 63980
rect 8208 63860 8260 63912
rect 8484 63903 8536 63912
rect 8484 63869 8493 63903
rect 8493 63869 8527 63903
rect 8527 63869 8536 63903
rect 8484 63860 8536 63869
rect 9772 63903 9824 63912
rect 9772 63869 9781 63903
rect 9781 63869 9815 63903
rect 9815 63869 9824 63903
rect 9772 63860 9824 63869
rect 10508 63903 10560 63912
rect 7196 63835 7248 63844
rect 7196 63801 7205 63835
rect 7205 63801 7239 63835
rect 7239 63801 7248 63835
rect 7196 63792 7248 63801
rect 1676 63767 1728 63776
rect 1676 63733 1685 63767
rect 1685 63733 1719 63767
rect 1719 63733 1728 63767
rect 1676 63724 1728 63733
rect 4620 63724 4672 63776
rect 5080 63767 5132 63776
rect 5080 63733 5089 63767
rect 5089 63733 5123 63767
rect 5123 63733 5132 63767
rect 5080 63724 5132 63733
rect 7472 63724 7524 63776
rect 9956 63792 10008 63844
rect 10508 63869 10517 63903
rect 10517 63869 10551 63903
rect 10551 63869 10560 63903
rect 10508 63860 10560 63869
rect 12072 63903 12124 63912
rect 12072 63869 12081 63903
rect 12081 63869 12115 63903
rect 12115 63869 12124 63903
rect 12072 63860 12124 63869
rect 15384 63928 15436 63980
rect 13084 63903 13136 63912
rect 13084 63869 13093 63903
rect 13093 63869 13127 63903
rect 13127 63869 13136 63903
rect 13084 63860 13136 63869
rect 14004 63903 14056 63912
rect 11060 63792 11112 63844
rect 8484 63724 8536 63776
rect 9404 63724 9456 63776
rect 9680 63724 9732 63776
rect 11152 63724 11204 63776
rect 12532 63792 12584 63844
rect 14004 63869 14013 63903
rect 14013 63869 14047 63903
rect 14047 63869 14056 63903
rect 14004 63860 14056 63869
rect 15568 63860 15620 63912
rect 16488 63860 16540 63912
rect 13268 63724 13320 63776
rect 15660 63724 15712 63776
rect 17500 63767 17552 63776
rect 17500 63733 17509 63767
rect 17509 63733 17543 63767
rect 17543 63733 17552 63767
rect 17500 63724 17552 63733
rect 7648 63622 7700 63674
rect 7712 63622 7764 63674
rect 7776 63622 7828 63674
rect 7840 63622 7892 63674
rect 14315 63622 14367 63674
rect 14379 63622 14431 63674
rect 14443 63622 14495 63674
rect 14507 63622 14559 63674
rect 5264 63520 5316 63572
rect 6092 63520 6144 63572
rect 6368 63520 6420 63572
rect 6644 63563 6696 63572
rect 6644 63529 6653 63563
rect 6653 63529 6687 63563
rect 6687 63529 6696 63563
rect 6644 63520 6696 63529
rect 8576 63520 8628 63572
rect 10140 63520 10192 63572
rect 10508 63520 10560 63572
rect 1768 63359 1820 63368
rect 1768 63325 1777 63359
rect 1777 63325 1811 63359
rect 1811 63325 1820 63359
rect 1768 63316 1820 63325
rect 2136 63316 2188 63368
rect 3884 63384 3936 63436
rect 3976 63316 4028 63368
rect 4528 63359 4580 63368
rect 4528 63325 4537 63359
rect 4537 63325 4571 63359
rect 4571 63325 4580 63359
rect 4528 63316 4580 63325
rect 8024 63384 8076 63436
rect 9864 63452 9916 63504
rect 11612 63520 11664 63572
rect 12072 63520 12124 63572
rect 15568 63563 15620 63572
rect 15568 63529 15577 63563
rect 15577 63529 15611 63563
rect 15611 63529 15620 63563
rect 15568 63520 15620 63529
rect 15752 63520 15804 63572
rect 9404 63427 9456 63436
rect 9404 63393 9413 63427
rect 9413 63393 9447 63427
rect 9447 63393 9456 63427
rect 9404 63384 9456 63393
rect 9588 63384 9640 63436
rect 9772 63427 9824 63436
rect 9772 63393 9781 63427
rect 9781 63393 9815 63427
rect 9815 63393 9824 63427
rect 9772 63384 9824 63393
rect 10692 63427 10744 63436
rect 7748 63316 7800 63368
rect 9036 63316 9088 63368
rect 10692 63393 10701 63427
rect 10701 63393 10735 63427
rect 10735 63393 10744 63427
rect 10692 63384 10744 63393
rect 12532 63384 12584 63436
rect 14740 63384 14792 63436
rect 15108 63384 15160 63436
rect 15568 63384 15620 63436
rect 10968 63316 11020 63368
rect 11428 63316 11480 63368
rect 2688 63248 2740 63300
rect 3424 63291 3476 63300
rect 3424 63257 3433 63291
rect 3433 63257 3467 63291
rect 3467 63257 3476 63291
rect 3424 63248 3476 63257
rect 9220 63291 9272 63300
rect 9220 63257 9229 63291
rect 9229 63257 9263 63291
rect 9263 63257 9272 63291
rect 9220 63248 9272 63257
rect 9680 63248 9732 63300
rect 10232 63248 10284 63300
rect 1676 63180 1728 63232
rect 2228 63180 2280 63232
rect 4068 63223 4120 63232
rect 4068 63189 4077 63223
rect 4077 63189 4111 63223
rect 4111 63189 4120 63223
rect 4068 63180 4120 63189
rect 8300 63223 8352 63232
rect 8300 63189 8309 63223
rect 8309 63189 8343 63223
rect 8343 63189 8352 63223
rect 8300 63180 8352 63189
rect 9588 63180 9640 63232
rect 10048 63180 10100 63232
rect 12992 63223 13044 63232
rect 12992 63189 13001 63223
rect 13001 63189 13035 63223
rect 13035 63189 13044 63223
rect 13360 63223 13412 63232
rect 12992 63180 13044 63189
rect 13360 63189 13369 63223
rect 13369 63189 13403 63223
rect 13403 63189 13412 63223
rect 13360 63180 13412 63189
rect 13728 63316 13780 63368
rect 14832 63180 14884 63232
rect 16212 63223 16264 63232
rect 16212 63189 16221 63223
rect 16221 63189 16255 63223
rect 16255 63189 16264 63223
rect 16212 63180 16264 63189
rect 4315 63078 4367 63130
rect 4379 63078 4431 63130
rect 4443 63078 4495 63130
rect 4507 63078 4559 63130
rect 10982 63078 11034 63130
rect 11046 63078 11098 63130
rect 11110 63078 11162 63130
rect 11174 63078 11226 63130
rect 17648 63078 17700 63130
rect 17712 63078 17764 63130
rect 17776 63078 17828 63130
rect 17840 63078 17892 63130
rect 2596 62976 2648 63028
rect 3976 62976 4028 63028
rect 4160 62976 4212 63028
rect 5448 62976 5500 63028
rect 9404 62976 9456 63028
rect 9956 63019 10008 63028
rect 9956 62985 9965 63019
rect 9965 62985 9999 63019
rect 9999 62985 10008 63019
rect 9956 62976 10008 62985
rect 9036 62908 9088 62960
rect 2228 62772 2280 62824
rect 2504 62815 2556 62824
rect 2504 62781 2513 62815
rect 2513 62781 2547 62815
rect 2547 62781 2556 62815
rect 2504 62772 2556 62781
rect 4804 62772 4856 62824
rect 5632 62772 5684 62824
rect 5816 62772 5868 62824
rect 6644 62815 6696 62824
rect 6644 62781 6653 62815
rect 6653 62781 6687 62815
rect 6687 62781 6696 62815
rect 6644 62772 6696 62781
rect 6828 62772 6880 62824
rect 7472 62772 7524 62824
rect 9404 62840 9456 62892
rect 1492 62747 1544 62756
rect 1492 62713 1501 62747
rect 1501 62713 1535 62747
rect 1535 62713 1544 62747
rect 1492 62704 1544 62713
rect 4068 62747 4120 62756
rect 4068 62713 4077 62747
rect 4077 62713 4111 62747
rect 4111 62713 4120 62747
rect 4068 62704 4120 62713
rect 4988 62704 5040 62756
rect 7748 62747 7800 62756
rect 7748 62713 7757 62747
rect 7757 62713 7791 62747
rect 7791 62713 7800 62747
rect 7748 62704 7800 62713
rect 8392 62704 8444 62756
rect 10692 62908 10744 62960
rect 12624 62976 12676 63028
rect 14740 63019 14792 63028
rect 14740 62985 14749 63019
rect 14749 62985 14783 63019
rect 14783 62985 14792 63019
rect 14740 62976 14792 62985
rect 15016 63019 15068 63028
rect 15016 62985 15025 63019
rect 15025 62985 15059 63019
rect 15059 62985 15068 63019
rect 15016 62976 15068 62985
rect 16948 63019 17000 63028
rect 16948 62985 16957 63019
rect 16957 62985 16991 63019
rect 16991 62985 17000 63019
rect 16948 62976 17000 62985
rect 10048 62815 10100 62824
rect 10048 62781 10057 62815
rect 10057 62781 10091 62815
rect 10091 62781 10100 62815
rect 10048 62772 10100 62781
rect 10232 62815 10284 62824
rect 10232 62781 10241 62815
rect 10241 62781 10275 62815
rect 10275 62781 10284 62815
rect 10232 62772 10284 62781
rect 10692 62815 10744 62824
rect 10692 62781 10701 62815
rect 10701 62781 10735 62815
rect 10735 62781 10744 62815
rect 10692 62772 10744 62781
rect 10968 62772 11020 62824
rect 4160 62636 4212 62688
rect 4712 62636 4764 62688
rect 4804 62636 4856 62688
rect 6552 62679 6604 62688
rect 6552 62645 6561 62679
rect 6561 62645 6595 62679
rect 6595 62645 6604 62679
rect 6552 62636 6604 62645
rect 7288 62679 7340 62688
rect 7288 62645 7297 62679
rect 7297 62645 7331 62679
rect 7331 62645 7340 62679
rect 7288 62636 7340 62645
rect 8760 62679 8812 62688
rect 8760 62645 8769 62679
rect 8769 62645 8803 62679
rect 8803 62645 8812 62679
rect 8760 62636 8812 62645
rect 12164 62636 12216 62688
rect 12532 62636 12584 62688
rect 13084 62772 13136 62824
rect 15016 62772 15068 62824
rect 15752 62772 15804 62824
rect 13360 62636 13412 62688
rect 13820 62636 13872 62688
rect 7648 62534 7700 62586
rect 7712 62534 7764 62586
rect 7776 62534 7828 62586
rect 7840 62534 7892 62586
rect 14315 62534 14367 62586
rect 14379 62534 14431 62586
rect 14443 62534 14495 62586
rect 14507 62534 14559 62586
rect 2412 62475 2464 62484
rect 2412 62441 2421 62475
rect 2421 62441 2455 62475
rect 2455 62441 2464 62475
rect 2412 62432 2464 62441
rect 3884 62432 3936 62484
rect 4804 62432 4856 62484
rect 1676 62296 1728 62348
rect 2872 62364 2924 62416
rect 9864 62432 9916 62484
rect 10232 62475 10284 62484
rect 10232 62441 10241 62475
rect 10241 62441 10275 62475
rect 10275 62441 10284 62475
rect 10232 62432 10284 62441
rect 12716 62432 12768 62484
rect 2136 62271 2188 62280
rect 2136 62237 2145 62271
rect 2145 62237 2179 62271
rect 2179 62237 2188 62271
rect 2136 62228 2188 62237
rect 3424 62228 3476 62280
rect 3976 62271 4028 62280
rect 3976 62237 3985 62271
rect 3985 62237 4019 62271
rect 4019 62237 4028 62271
rect 3976 62228 4028 62237
rect 2964 62160 3016 62212
rect 4068 62160 4120 62212
rect 8944 62296 8996 62348
rect 9864 62296 9916 62348
rect 11336 62339 11388 62348
rect 11336 62305 11345 62339
rect 11345 62305 11379 62339
rect 11379 62305 11388 62339
rect 11336 62296 11388 62305
rect 12440 62339 12492 62348
rect 12440 62305 12449 62339
rect 12449 62305 12483 62339
rect 12483 62305 12492 62339
rect 12440 62296 12492 62305
rect 13360 62296 13412 62348
rect 14280 62296 14332 62348
rect 11520 62271 11572 62280
rect 11520 62237 11529 62271
rect 11529 62237 11563 62271
rect 11563 62237 11572 62271
rect 11520 62228 11572 62237
rect 14004 62271 14056 62280
rect 14004 62237 14013 62271
rect 14013 62237 14047 62271
rect 14047 62237 14056 62271
rect 14004 62228 14056 62237
rect 15200 62271 15252 62280
rect 15200 62237 15209 62271
rect 15209 62237 15243 62271
rect 15243 62237 15252 62271
rect 15200 62228 15252 62237
rect 15568 62228 15620 62280
rect 4712 62160 4764 62212
rect 9772 62160 9824 62212
rect 10140 62160 10192 62212
rect 9496 62092 9548 62144
rect 10692 62135 10744 62144
rect 10692 62101 10701 62135
rect 10701 62101 10735 62135
rect 10735 62101 10744 62135
rect 10692 62092 10744 62101
rect 13728 62092 13780 62144
rect 15384 62092 15436 62144
rect 4315 61990 4367 62042
rect 4379 61990 4431 62042
rect 4443 61990 4495 62042
rect 4507 61990 4559 62042
rect 10982 61990 11034 62042
rect 11046 61990 11098 62042
rect 11110 61990 11162 62042
rect 11174 61990 11226 62042
rect 17648 61990 17700 62042
rect 17712 61990 17764 62042
rect 17776 61990 17828 62042
rect 17840 61990 17892 62042
rect 3976 61888 4028 61940
rect 6920 61888 6972 61940
rect 7104 61888 7156 61940
rect 8760 61888 8812 61940
rect 8944 61820 8996 61872
rect 2136 61752 2188 61804
rect 2504 61795 2556 61804
rect 1676 61684 1728 61736
rect 2504 61761 2513 61795
rect 2513 61761 2547 61795
rect 2547 61761 2556 61795
rect 2504 61752 2556 61761
rect 2688 61752 2740 61804
rect 3884 61752 3936 61804
rect 8484 61752 8536 61804
rect 9128 61752 9180 61804
rect 11336 61888 11388 61940
rect 11520 61888 11572 61940
rect 14740 61931 14792 61940
rect 14740 61897 14749 61931
rect 14749 61897 14783 61931
rect 14783 61897 14792 61931
rect 14740 61888 14792 61897
rect 13268 61820 13320 61872
rect 14280 61863 14332 61872
rect 14280 61829 14289 61863
rect 14289 61829 14323 61863
rect 14323 61829 14332 61863
rect 14280 61820 14332 61829
rect 14648 61820 14700 61872
rect 15016 61820 15068 61872
rect 1492 61659 1544 61668
rect 1492 61625 1501 61659
rect 1501 61625 1535 61659
rect 1535 61625 1544 61659
rect 1492 61616 1544 61625
rect 4712 61684 4764 61736
rect 13636 61752 13688 61804
rect 3056 61616 3108 61668
rect 10324 61684 10376 61736
rect 12716 61727 12768 61736
rect 10232 61616 10284 61668
rect 12716 61693 12725 61727
rect 12725 61693 12759 61727
rect 12759 61693 12768 61727
rect 12716 61684 12768 61693
rect 13268 61727 13320 61736
rect 13268 61693 13277 61727
rect 13277 61693 13311 61727
rect 13311 61693 13320 61727
rect 13268 61684 13320 61693
rect 14740 61684 14792 61736
rect 15568 61727 15620 61736
rect 12624 61616 12676 61668
rect 13728 61616 13780 61668
rect 3148 61591 3200 61600
rect 3148 61557 3157 61591
rect 3157 61557 3191 61591
rect 3191 61557 3200 61591
rect 3148 61548 3200 61557
rect 3424 61591 3476 61600
rect 3424 61557 3433 61591
rect 3433 61557 3467 61591
rect 3467 61557 3476 61591
rect 3424 61548 3476 61557
rect 5448 61591 5500 61600
rect 5448 61557 5457 61591
rect 5457 61557 5491 61591
rect 5491 61557 5500 61591
rect 5448 61548 5500 61557
rect 8484 61591 8536 61600
rect 8484 61557 8493 61591
rect 8493 61557 8527 61591
rect 8527 61557 8536 61591
rect 8484 61548 8536 61557
rect 10140 61548 10192 61600
rect 11520 61548 11572 61600
rect 11704 61548 11756 61600
rect 14004 61548 14056 61600
rect 14924 61548 14976 61600
rect 15568 61693 15577 61727
rect 15577 61693 15611 61727
rect 15611 61693 15620 61727
rect 15568 61684 15620 61693
rect 15936 61548 15988 61600
rect 16672 61591 16724 61600
rect 16672 61557 16681 61591
rect 16681 61557 16715 61591
rect 16715 61557 16724 61591
rect 16672 61548 16724 61557
rect 7648 61446 7700 61498
rect 7712 61446 7764 61498
rect 7776 61446 7828 61498
rect 7840 61446 7892 61498
rect 14315 61446 14367 61498
rect 14379 61446 14431 61498
rect 14443 61446 14495 61498
rect 14507 61446 14559 61498
rect 3056 61387 3108 61396
rect 3056 61353 3065 61387
rect 3065 61353 3099 61387
rect 3099 61353 3108 61387
rect 3056 61344 3108 61353
rect 3424 61344 3476 61396
rect 4804 61387 4856 61396
rect 4804 61353 4813 61387
rect 4813 61353 4847 61387
rect 4847 61353 4856 61387
rect 4804 61344 4856 61353
rect 9772 61387 9824 61396
rect 9772 61353 9781 61387
rect 9781 61353 9815 61387
rect 9815 61353 9824 61387
rect 9772 61344 9824 61353
rect 10232 61344 10284 61396
rect 4712 61276 4764 61328
rect 7380 61276 7432 61328
rect 7564 61276 7616 61328
rect 8024 61276 8076 61328
rect 1216 61208 1268 61260
rect 2688 61208 2740 61260
rect 3700 61208 3752 61260
rect 1768 61183 1820 61192
rect 1768 61149 1777 61183
rect 1777 61149 1811 61183
rect 1811 61149 1820 61183
rect 1768 61140 1820 61149
rect 3424 61072 3476 61124
rect 5448 61208 5500 61260
rect 8300 61251 8352 61260
rect 8300 61217 8309 61251
rect 8309 61217 8343 61251
rect 8343 61217 8352 61251
rect 8300 61208 8352 61217
rect 8760 61251 8812 61260
rect 8760 61217 8769 61251
rect 8769 61217 8803 61251
rect 8803 61217 8812 61251
rect 8760 61208 8812 61217
rect 9772 61208 9824 61260
rect 9864 61208 9916 61260
rect 11060 61251 11112 61260
rect 11060 61217 11069 61251
rect 11069 61217 11103 61251
rect 11103 61217 11112 61251
rect 11060 61208 11112 61217
rect 11428 61208 11480 61260
rect 13452 61276 13504 61328
rect 13176 61251 13228 61260
rect 13176 61217 13185 61251
rect 13185 61217 13219 61251
rect 13219 61217 13228 61251
rect 13176 61208 13228 61217
rect 13820 61208 13872 61260
rect 14648 61208 14700 61260
rect 7196 61140 7248 61192
rect 7380 61140 7432 61192
rect 9036 61140 9088 61192
rect 9496 61140 9548 61192
rect 10048 61140 10100 61192
rect 11336 61140 11388 61192
rect 13636 61140 13688 61192
rect 15016 61183 15068 61192
rect 15016 61149 15025 61183
rect 15025 61149 15059 61183
rect 15059 61149 15068 61183
rect 15016 61140 15068 61149
rect 4068 61004 4120 61056
rect 4620 61004 4672 61056
rect 8300 61047 8352 61056
rect 8300 61013 8309 61047
rect 8309 61013 8343 61047
rect 8343 61013 8352 61047
rect 8300 61004 8352 61013
rect 8668 61004 8720 61056
rect 10232 61004 10284 61056
rect 12348 61004 12400 61056
rect 16120 61047 16172 61056
rect 16120 61013 16129 61047
rect 16129 61013 16163 61047
rect 16163 61013 16172 61047
rect 16120 61004 16172 61013
rect 4315 60902 4367 60954
rect 4379 60902 4431 60954
rect 4443 60902 4495 60954
rect 4507 60902 4559 60954
rect 10982 60902 11034 60954
rect 11046 60902 11098 60954
rect 11110 60902 11162 60954
rect 11174 60902 11226 60954
rect 17648 60902 17700 60954
rect 17712 60902 17764 60954
rect 17776 60902 17828 60954
rect 17840 60902 17892 60954
rect 3424 60843 3476 60852
rect 3424 60809 3433 60843
rect 3433 60809 3467 60843
rect 3467 60809 3476 60843
rect 3424 60800 3476 60809
rect 3700 60800 3752 60852
rect 1952 60664 2004 60716
rect 5264 60800 5316 60852
rect 5540 60800 5592 60852
rect 8484 60800 8536 60852
rect 9864 60800 9916 60852
rect 10048 60800 10100 60852
rect 11428 60843 11480 60852
rect 2688 60639 2740 60648
rect 2688 60605 2697 60639
rect 2697 60605 2731 60639
rect 2731 60605 2740 60639
rect 2688 60596 2740 60605
rect 2872 60596 2924 60648
rect 3056 60596 3108 60648
rect 8944 60664 8996 60716
rect 9128 60664 9180 60716
rect 4620 60596 4672 60648
rect 8300 60639 8352 60648
rect 8300 60605 8309 60639
rect 8309 60605 8343 60639
rect 8343 60605 8352 60639
rect 8300 60596 8352 60605
rect 10416 60596 10468 60648
rect 10600 60639 10652 60648
rect 10600 60605 10609 60639
rect 10609 60605 10643 60639
rect 10643 60605 10652 60639
rect 10600 60596 10652 60605
rect 11428 60809 11437 60843
rect 11437 60809 11471 60843
rect 11471 60809 11480 60843
rect 11428 60800 11480 60809
rect 13176 60800 13228 60852
rect 11796 60732 11848 60784
rect 14648 60732 14700 60784
rect 11428 60664 11480 60716
rect 11980 60664 12032 60716
rect 12532 60707 12584 60716
rect 12532 60673 12541 60707
rect 12541 60673 12575 60707
rect 12575 60673 12584 60707
rect 12532 60664 12584 60673
rect 11796 60596 11848 60648
rect 1676 60503 1728 60512
rect 1676 60469 1685 60503
rect 1685 60469 1719 60503
rect 1719 60469 1728 60503
rect 1676 60460 1728 60469
rect 4344 60503 4396 60512
rect 4344 60469 4353 60503
rect 4353 60469 4387 60503
rect 4387 60469 4396 60503
rect 4344 60460 4396 60469
rect 8024 60460 8076 60512
rect 8392 60503 8444 60512
rect 8392 60469 8401 60503
rect 8401 60469 8435 60503
rect 8435 60469 8444 60503
rect 8392 60460 8444 60469
rect 9128 60460 9180 60512
rect 12440 60639 12492 60648
rect 12440 60605 12449 60639
rect 12449 60605 12483 60639
rect 12483 60605 12492 60639
rect 12716 60639 12768 60648
rect 12440 60596 12492 60605
rect 12716 60605 12725 60639
rect 12725 60605 12759 60639
rect 12759 60605 12768 60639
rect 12716 60596 12768 60605
rect 16120 60639 16172 60648
rect 16120 60605 16129 60639
rect 16129 60605 16163 60639
rect 16163 60605 16172 60639
rect 16120 60596 16172 60605
rect 16488 60596 16540 60648
rect 11980 60460 12032 60512
rect 13452 60503 13504 60512
rect 13452 60469 13461 60503
rect 13461 60469 13495 60503
rect 13495 60469 13504 60503
rect 13452 60460 13504 60469
rect 15016 60460 15068 60512
rect 17500 60503 17552 60512
rect 17500 60469 17509 60503
rect 17509 60469 17543 60503
rect 17543 60469 17552 60503
rect 17500 60460 17552 60469
rect 7648 60358 7700 60410
rect 7712 60358 7764 60410
rect 7776 60358 7828 60410
rect 7840 60358 7892 60410
rect 14315 60358 14367 60410
rect 14379 60358 14431 60410
rect 14443 60358 14495 60410
rect 14507 60358 14559 60410
rect 2688 60256 2740 60308
rect 4620 60299 4672 60308
rect 4620 60265 4629 60299
rect 4629 60265 4663 60299
rect 4663 60265 4672 60299
rect 4620 60256 4672 60265
rect 7380 60256 7432 60308
rect 8300 60256 8352 60308
rect 9772 60256 9824 60308
rect 10416 60256 10468 60308
rect 12716 60256 12768 60308
rect 2780 60120 2832 60172
rect 6460 60120 6512 60172
rect 8668 60120 8720 60172
rect 14740 60256 14792 60308
rect 16120 60299 16172 60308
rect 16120 60265 16129 60299
rect 16129 60265 16163 60299
rect 16163 60265 16172 60299
rect 16120 60256 16172 60265
rect 10876 60163 10928 60172
rect 10876 60129 10885 60163
rect 10885 60129 10919 60163
rect 10919 60129 10928 60163
rect 10876 60120 10928 60129
rect 12440 60120 12492 60172
rect 2872 60052 2924 60104
rect 3424 60052 3476 60104
rect 3700 60052 3752 60104
rect 9404 60095 9456 60104
rect 9404 60061 9413 60095
rect 9413 60061 9447 60095
rect 9447 60061 9456 60095
rect 9404 60052 9456 60061
rect 11704 60052 11756 60104
rect 6184 60027 6236 60036
rect 6184 59993 6193 60027
rect 6193 59993 6227 60027
rect 6227 59993 6236 60027
rect 6184 59984 6236 59993
rect 12716 59984 12768 60036
rect 13176 60163 13228 60172
rect 13176 60129 13185 60163
rect 13185 60129 13219 60163
rect 13219 60129 13228 60163
rect 13176 60120 13228 60129
rect 12992 60095 13044 60104
rect 12992 60061 13001 60095
rect 13001 60061 13035 60095
rect 13035 60061 13044 60095
rect 12992 60052 13044 60061
rect 14004 59984 14056 60036
rect 1768 59916 1820 59968
rect 1952 59916 2004 59968
rect 2688 59916 2740 59968
rect 8300 59959 8352 59968
rect 8300 59925 8309 59959
rect 8309 59925 8343 59959
rect 8343 59925 8352 59959
rect 8300 59916 8352 59925
rect 8576 59916 8628 59968
rect 10600 59959 10652 59968
rect 10600 59925 10609 59959
rect 10609 59925 10643 59959
rect 10643 59925 10652 59959
rect 10600 59916 10652 59925
rect 11520 59916 11572 59968
rect 14832 59916 14884 59968
rect 4315 59814 4367 59866
rect 4379 59814 4431 59866
rect 4443 59814 4495 59866
rect 4507 59814 4559 59866
rect 10982 59814 11034 59866
rect 11046 59814 11098 59866
rect 11110 59814 11162 59866
rect 11174 59814 11226 59866
rect 17648 59814 17700 59866
rect 17712 59814 17764 59866
rect 17776 59814 17828 59866
rect 17840 59814 17892 59866
rect 3700 59755 3752 59764
rect 3700 59721 3709 59755
rect 3709 59721 3743 59755
rect 3743 59721 3752 59755
rect 3700 59712 3752 59721
rect 4804 59712 4856 59764
rect 5632 59755 5684 59764
rect 5632 59721 5641 59755
rect 5641 59721 5675 59755
rect 5675 59721 5684 59755
rect 5632 59712 5684 59721
rect 6276 59755 6328 59764
rect 6276 59721 6285 59755
rect 6285 59721 6319 59755
rect 6319 59721 6328 59755
rect 6276 59712 6328 59721
rect 6736 59712 6788 59764
rect 1492 59644 1544 59696
rect 6184 59644 6236 59696
rect 9036 59712 9088 59764
rect 2688 59508 2740 59560
rect 6460 59576 6512 59628
rect 6920 59576 6972 59628
rect 2872 59372 2924 59424
rect 3424 59372 3476 59424
rect 5816 59508 5868 59560
rect 6000 59508 6052 59560
rect 7288 59551 7340 59560
rect 7288 59517 7297 59551
rect 7297 59517 7331 59551
rect 7331 59517 7340 59551
rect 7288 59508 7340 59517
rect 10600 59712 10652 59764
rect 10784 59619 10836 59628
rect 7196 59440 7248 59492
rect 10416 59508 10468 59560
rect 10784 59585 10793 59619
rect 10793 59585 10827 59619
rect 10827 59585 10836 59619
rect 10784 59576 10836 59585
rect 10692 59551 10744 59560
rect 10692 59517 10701 59551
rect 10701 59517 10735 59551
rect 10735 59517 10744 59551
rect 10692 59508 10744 59517
rect 8484 59440 8536 59492
rect 8944 59440 8996 59492
rect 9772 59440 9824 59492
rect 8668 59415 8720 59424
rect 8668 59381 8677 59415
rect 8677 59381 8711 59415
rect 8711 59381 8720 59415
rect 8668 59372 8720 59381
rect 10692 59372 10744 59424
rect 13176 59712 13228 59764
rect 13452 59755 13504 59764
rect 13452 59721 13461 59755
rect 13461 59721 13495 59755
rect 13495 59721 13504 59755
rect 13452 59712 13504 59721
rect 14004 59755 14056 59764
rect 14004 59721 14013 59755
rect 14013 59721 14047 59755
rect 14047 59721 14056 59755
rect 14004 59712 14056 59721
rect 14096 59712 14148 59764
rect 13544 59644 13596 59696
rect 12532 59551 12584 59560
rect 12532 59517 12541 59551
rect 12541 59517 12575 59551
rect 12575 59517 12584 59551
rect 12532 59508 12584 59517
rect 12716 59551 12768 59560
rect 12716 59517 12725 59551
rect 12725 59517 12759 59551
rect 12759 59517 12768 59551
rect 12716 59508 12768 59517
rect 12992 59551 13044 59560
rect 12992 59517 13001 59551
rect 13001 59517 13035 59551
rect 13035 59517 13044 59551
rect 12992 59508 13044 59517
rect 13544 59551 13596 59560
rect 13544 59517 13553 59551
rect 13553 59517 13587 59551
rect 13587 59517 13596 59551
rect 13544 59508 13596 59517
rect 15936 59508 15988 59560
rect 16396 59551 16448 59560
rect 16396 59517 16405 59551
rect 16405 59517 16439 59551
rect 16439 59517 16448 59551
rect 16396 59508 16448 59517
rect 12348 59440 12400 59492
rect 13268 59372 13320 59424
rect 13452 59372 13504 59424
rect 7648 59270 7700 59322
rect 7712 59270 7764 59322
rect 7776 59270 7828 59322
rect 7840 59270 7892 59322
rect 14315 59270 14367 59322
rect 14379 59270 14431 59322
rect 14443 59270 14495 59322
rect 14507 59270 14559 59322
rect 1584 59143 1636 59152
rect 1584 59109 1593 59143
rect 1593 59109 1627 59143
rect 1627 59109 1636 59143
rect 1584 59100 1636 59109
rect 1768 59100 1820 59152
rect 1492 59075 1544 59084
rect 1492 59041 1501 59075
rect 1501 59041 1535 59075
rect 1535 59041 1544 59075
rect 1492 59032 1544 59041
rect 2872 59168 2924 59220
rect 4804 59168 4856 59220
rect 10600 59168 10652 59220
rect 10876 59211 10928 59220
rect 10876 59177 10885 59211
rect 10885 59177 10919 59211
rect 10919 59177 10928 59211
rect 10876 59168 10928 59177
rect 11612 59168 11664 59220
rect 12348 59168 12400 59220
rect 5448 59100 5500 59152
rect 1676 58964 1728 59016
rect 2228 58964 2280 59016
rect 4620 59032 4672 59084
rect 4988 59032 5040 59084
rect 5724 59075 5776 59084
rect 5724 59041 5733 59075
rect 5733 59041 5767 59075
rect 5767 59041 5776 59075
rect 5724 59032 5776 59041
rect 6828 59032 6880 59084
rect 7380 59032 7432 59084
rect 8392 59100 8444 59152
rect 12716 59100 12768 59152
rect 13268 59100 13320 59152
rect 8484 59075 8536 59084
rect 8484 59041 8493 59075
rect 8493 59041 8527 59075
rect 8527 59041 8536 59075
rect 8484 59032 8536 59041
rect 8668 59007 8720 59016
rect 8668 58973 8677 59007
rect 8677 58973 8711 59007
rect 8711 58973 8720 59007
rect 8668 58964 8720 58973
rect 9128 59032 9180 59084
rect 9772 59075 9824 59084
rect 9772 59041 9781 59075
rect 9781 59041 9815 59075
rect 9815 59041 9824 59075
rect 9772 59032 9824 59041
rect 11612 59032 11664 59084
rect 12164 59032 12216 59084
rect 9496 58964 9548 59016
rect 4068 58896 4120 58948
rect 6000 58896 6052 58948
rect 12440 58896 12492 58948
rect 13820 59168 13872 59220
rect 13912 58964 13964 59016
rect 14832 59007 14884 59016
rect 14832 58973 14841 59007
rect 14841 58973 14875 59007
rect 14875 58973 14884 59007
rect 14832 58964 14884 58973
rect 6644 58871 6696 58880
rect 6644 58837 6653 58871
rect 6653 58837 6687 58871
rect 6687 58837 6696 58871
rect 6644 58828 6696 58837
rect 7196 58828 7248 58880
rect 8300 58871 8352 58880
rect 8300 58837 8309 58871
rect 8309 58837 8343 58871
rect 8343 58837 8352 58871
rect 8300 58828 8352 58837
rect 12808 58871 12860 58880
rect 12808 58837 12817 58871
rect 12817 58837 12851 58871
rect 12851 58837 12860 58871
rect 12808 58828 12860 58837
rect 14648 58828 14700 58880
rect 15936 58828 15988 58880
rect 4315 58726 4367 58778
rect 4379 58726 4431 58778
rect 4443 58726 4495 58778
rect 4507 58726 4559 58778
rect 10982 58726 11034 58778
rect 11046 58726 11098 58778
rect 11110 58726 11162 58778
rect 11174 58726 11226 58778
rect 17648 58726 17700 58778
rect 17712 58726 17764 58778
rect 17776 58726 17828 58778
rect 17840 58726 17892 58778
rect 2780 58624 2832 58676
rect 4620 58667 4672 58676
rect 4620 58633 4629 58667
rect 4629 58633 4663 58667
rect 4663 58633 4672 58667
rect 4620 58624 4672 58633
rect 4988 58667 5040 58676
rect 4988 58633 4997 58667
rect 4997 58633 5031 58667
rect 5031 58633 5040 58667
rect 4988 58624 5040 58633
rect 8024 58624 8076 58676
rect 14648 58667 14700 58676
rect 14648 58633 14657 58667
rect 14657 58633 14691 58667
rect 14691 58633 14700 58667
rect 14648 58624 14700 58633
rect 4068 58556 4120 58608
rect 1216 58488 1268 58540
rect 1768 58531 1820 58540
rect 1768 58497 1777 58531
rect 1777 58497 1811 58531
rect 1811 58497 1820 58531
rect 1768 58488 1820 58497
rect 4620 58420 4672 58472
rect 6828 58488 6880 58540
rect 9680 58556 9732 58608
rect 10416 58599 10468 58608
rect 10416 58565 10425 58599
rect 10425 58565 10459 58599
rect 10459 58565 10468 58599
rect 10416 58556 10468 58565
rect 11244 58556 11296 58608
rect 11428 58556 11480 58608
rect 12164 58488 12216 58540
rect 6000 58463 6052 58472
rect 6000 58429 6009 58463
rect 6009 58429 6043 58463
rect 6043 58429 6052 58463
rect 6000 58420 6052 58429
rect 6368 58463 6420 58472
rect 6368 58429 6377 58463
rect 6377 58429 6411 58463
rect 6411 58429 6420 58463
rect 6368 58420 6420 58429
rect 1768 58284 1820 58336
rect 3056 58284 3108 58336
rect 3424 58284 3476 58336
rect 5080 58284 5132 58336
rect 8300 58420 8352 58472
rect 8576 58463 8628 58472
rect 8576 58429 8585 58463
rect 8585 58429 8619 58463
rect 8619 58429 8628 58463
rect 8576 58420 8628 58429
rect 9680 58463 9732 58472
rect 9680 58429 9689 58463
rect 9689 58429 9723 58463
rect 9723 58429 9732 58463
rect 9680 58420 9732 58429
rect 6920 58352 6972 58404
rect 10600 58420 10652 58472
rect 12440 58463 12492 58472
rect 12440 58429 12449 58463
rect 12449 58429 12483 58463
rect 12483 58429 12492 58463
rect 12440 58420 12492 58429
rect 12808 58420 12860 58472
rect 13636 58420 13688 58472
rect 8024 58284 8076 58336
rect 8208 58284 8260 58336
rect 9128 58327 9180 58336
rect 9128 58293 9137 58327
rect 9137 58293 9171 58327
rect 9171 58293 9180 58327
rect 9128 58284 9180 58293
rect 9496 58327 9548 58336
rect 9496 58293 9505 58327
rect 9505 58293 9539 58327
rect 9539 58293 9548 58327
rect 9496 58284 9548 58293
rect 11428 58284 11480 58336
rect 11612 58284 11664 58336
rect 12072 58327 12124 58336
rect 12072 58293 12081 58327
rect 12081 58293 12115 58327
rect 12115 58293 12124 58327
rect 12072 58284 12124 58293
rect 12256 58327 12308 58336
rect 12256 58293 12265 58327
rect 12265 58293 12299 58327
rect 12299 58293 12308 58327
rect 12256 58284 12308 58293
rect 14096 58327 14148 58336
rect 14096 58293 14105 58327
rect 14105 58293 14139 58327
rect 14139 58293 14148 58327
rect 14096 58284 14148 58293
rect 7648 58182 7700 58234
rect 7712 58182 7764 58234
rect 7776 58182 7828 58234
rect 7840 58182 7892 58234
rect 14315 58182 14367 58234
rect 14379 58182 14431 58234
rect 14443 58182 14495 58234
rect 14507 58182 14559 58234
rect 1308 58080 1360 58132
rect 1400 58012 1452 58064
rect 6276 58080 6328 58132
rect 6460 58123 6512 58132
rect 6460 58089 6469 58123
rect 6469 58089 6503 58123
rect 6503 58089 6512 58123
rect 6460 58080 6512 58089
rect 6736 58080 6788 58132
rect 11152 58123 11204 58132
rect 11152 58089 11161 58123
rect 11161 58089 11195 58123
rect 11195 58089 11204 58123
rect 11152 58080 11204 58089
rect 12256 58080 12308 58132
rect 15936 58123 15988 58132
rect 15936 58089 15945 58123
rect 15945 58089 15979 58123
rect 15979 58089 15988 58123
rect 15936 58080 15988 58089
rect 1492 57919 1544 57928
rect 1492 57885 1501 57919
rect 1501 57885 1535 57919
rect 1535 57885 1544 57919
rect 1492 57876 1544 57885
rect 2228 57876 2280 57928
rect 1400 57808 1452 57860
rect 1952 57808 2004 57860
rect 3700 57876 3752 57928
rect 4804 57987 4856 57996
rect 4804 57953 4813 57987
rect 4813 57953 4847 57987
rect 4847 57953 4856 57987
rect 4804 57944 4856 57953
rect 5724 58012 5776 58064
rect 7932 58012 7984 58064
rect 8576 58012 8628 58064
rect 6460 57944 6512 57996
rect 7656 57944 7708 57996
rect 7840 57987 7892 57996
rect 7840 57953 7849 57987
rect 7849 57953 7883 57987
rect 7883 57953 7892 57987
rect 7840 57944 7892 57953
rect 9772 57944 9824 57996
rect 12532 57987 12584 57996
rect 4620 57876 4672 57928
rect 3516 57808 3568 57860
rect 6184 57876 6236 57928
rect 8392 57876 8444 57928
rect 9312 57876 9364 57928
rect 6736 57808 6788 57860
rect 10692 57876 10744 57928
rect 10876 57876 10928 57928
rect 12532 57953 12541 57987
rect 12541 57953 12575 57987
rect 12575 57953 12584 57987
rect 12532 57944 12584 57953
rect 12808 57987 12860 57996
rect 12808 57953 12817 57987
rect 12817 57953 12851 57987
rect 12851 57953 12860 57987
rect 12808 57944 12860 57953
rect 13176 57987 13228 57996
rect 13176 57953 13185 57987
rect 13185 57953 13219 57987
rect 13219 57953 13228 57987
rect 13176 57944 13228 57953
rect 11704 57919 11756 57928
rect 11704 57885 11713 57919
rect 11713 57885 11747 57919
rect 11747 57885 11756 57919
rect 11704 57876 11756 57885
rect 12256 57876 12308 57928
rect 13544 57919 13596 57928
rect 13544 57885 13553 57919
rect 13553 57885 13587 57919
rect 13587 57885 13596 57919
rect 13544 57876 13596 57885
rect 13820 57876 13872 57928
rect 11244 57808 11296 57860
rect 11612 57808 11664 57860
rect 3056 57740 3108 57792
rect 6276 57783 6328 57792
rect 6276 57749 6285 57783
rect 6285 57749 6319 57783
rect 6319 57749 6328 57783
rect 6276 57740 6328 57749
rect 7840 57740 7892 57792
rect 8576 57783 8628 57792
rect 8576 57749 8585 57783
rect 8585 57749 8619 57783
rect 8619 57749 8628 57783
rect 8576 57740 8628 57749
rect 9036 57740 9088 57792
rect 9680 57740 9732 57792
rect 10692 57740 10744 57792
rect 13912 57740 13964 57792
rect 15568 57740 15620 57792
rect 4315 57638 4367 57690
rect 4379 57638 4431 57690
rect 4443 57638 4495 57690
rect 4507 57638 4559 57690
rect 10982 57638 11034 57690
rect 11046 57638 11098 57690
rect 11110 57638 11162 57690
rect 11174 57638 11226 57690
rect 17648 57638 17700 57690
rect 17712 57638 17764 57690
rect 17776 57638 17828 57690
rect 17840 57638 17892 57690
rect 5448 57536 5500 57588
rect 9312 57536 9364 57588
rect 9588 57536 9640 57588
rect 10324 57536 10376 57588
rect 12808 57536 12860 57588
rect 6368 57468 6420 57520
rect 7564 57468 7616 57520
rect 2044 57400 2096 57452
rect 3700 57400 3752 57452
rect 3056 57332 3108 57384
rect 6736 57400 6788 57452
rect 9864 57400 9916 57452
rect 10876 57400 10928 57452
rect 6828 57332 6880 57384
rect 7288 57332 7340 57384
rect 2228 57196 2280 57248
rect 6644 57264 6696 57316
rect 10324 57332 10376 57384
rect 10968 57332 11020 57384
rect 14648 57468 14700 57520
rect 11796 57443 11848 57452
rect 11796 57409 11805 57443
rect 11805 57409 11839 57443
rect 11839 57409 11848 57443
rect 11796 57400 11848 57409
rect 12256 57400 12308 57452
rect 7656 57264 7708 57316
rect 9772 57264 9824 57316
rect 3700 57196 3752 57248
rect 4620 57196 4672 57248
rect 5448 57196 5500 57248
rect 5724 57196 5776 57248
rect 7380 57196 7432 57248
rect 8392 57239 8444 57248
rect 8392 57205 8401 57239
rect 8401 57205 8435 57239
rect 8435 57205 8444 57239
rect 8392 57196 8444 57205
rect 9864 57196 9916 57248
rect 12532 57332 12584 57384
rect 15936 57375 15988 57384
rect 12716 57264 12768 57316
rect 13176 57264 13228 57316
rect 15936 57341 15945 57375
rect 15945 57341 15979 57375
rect 15979 57341 15988 57375
rect 15936 57332 15988 57341
rect 16212 57375 16264 57384
rect 16212 57341 16221 57375
rect 16221 57341 16255 57375
rect 16255 57341 16264 57375
rect 16212 57332 16264 57341
rect 12256 57196 12308 57248
rect 12808 57196 12860 57248
rect 13452 57239 13504 57248
rect 13452 57205 13461 57239
rect 13461 57205 13495 57239
rect 13495 57205 13504 57239
rect 13452 57196 13504 57205
rect 17316 57239 17368 57248
rect 17316 57205 17325 57239
rect 17325 57205 17359 57239
rect 17359 57205 17368 57239
rect 17316 57196 17368 57205
rect 7648 57094 7700 57146
rect 7712 57094 7764 57146
rect 7776 57094 7828 57146
rect 7840 57094 7892 57146
rect 14315 57094 14367 57146
rect 14379 57094 14431 57146
rect 14443 57094 14495 57146
rect 14507 57094 14559 57146
rect 4804 56992 4856 57044
rect 6184 57035 6236 57044
rect 6184 57001 6193 57035
rect 6193 57001 6227 57035
rect 6227 57001 6236 57035
rect 6184 56992 6236 57001
rect 9680 56992 9732 57044
rect 12072 56992 12124 57044
rect 12532 56992 12584 57044
rect 3056 56924 3108 56976
rect 3424 56924 3476 56976
rect 6828 56924 6880 56976
rect 1676 56856 1728 56908
rect 3516 56856 3568 56908
rect 4804 56856 4856 56908
rect 6184 56856 6236 56908
rect 8576 56924 8628 56976
rect 9312 56924 9364 56976
rect 12440 56967 12492 56976
rect 12440 56933 12449 56967
rect 12449 56933 12483 56967
rect 12483 56933 12492 56967
rect 12440 56924 12492 56933
rect 8852 56856 8904 56908
rect 9496 56856 9548 56908
rect 9680 56856 9732 56908
rect 10600 56856 10652 56908
rect 11704 56899 11756 56908
rect 1768 56788 1820 56840
rect 6276 56788 6328 56840
rect 7840 56788 7892 56840
rect 8208 56788 8260 56840
rect 10416 56788 10468 56840
rect 11704 56865 11713 56899
rect 11713 56865 11747 56899
rect 11747 56865 11756 56899
rect 11704 56856 11756 56865
rect 12624 56856 12676 56908
rect 12992 56899 13044 56908
rect 12992 56865 13001 56899
rect 13001 56865 13035 56899
rect 13035 56865 13044 56899
rect 12992 56856 13044 56865
rect 7472 56720 7524 56772
rect 15660 56788 15712 56840
rect 2688 56652 2740 56704
rect 3516 56652 3568 56704
rect 5724 56652 5776 56704
rect 6736 56652 6788 56704
rect 8576 56652 8628 56704
rect 12256 56652 12308 56704
rect 12808 56652 12860 56704
rect 14188 56652 14240 56704
rect 16672 56695 16724 56704
rect 16672 56661 16681 56695
rect 16681 56661 16715 56695
rect 16715 56661 16724 56695
rect 16672 56652 16724 56661
rect 4315 56550 4367 56602
rect 4379 56550 4431 56602
rect 4443 56550 4495 56602
rect 4507 56550 4559 56602
rect 10982 56550 11034 56602
rect 11046 56550 11098 56602
rect 11110 56550 11162 56602
rect 11174 56550 11226 56602
rect 17648 56550 17700 56602
rect 17712 56550 17764 56602
rect 17776 56550 17828 56602
rect 17840 56550 17892 56602
rect 1492 56448 1544 56500
rect 4804 56448 4856 56500
rect 4988 56448 5040 56500
rect 5632 56491 5684 56500
rect 3516 56380 3568 56432
rect 4068 56380 4120 56432
rect 2688 56312 2740 56364
rect 3700 56312 3752 56364
rect 4988 56312 5040 56364
rect 2872 56287 2924 56296
rect 2872 56253 2881 56287
rect 2881 56253 2915 56287
rect 2915 56253 2924 56287
rect 2872 56244 2924 56253
rect 4344 56287 4396 56296
rect 4344 56253 4353 56287
rect 4353 56253 4387 56287
rect 4387 56253 4396 56287
rect 4344 56244 4396 56253
rect 4068 56108 4120 56160
rect 4804 56108 4856 56160
rect 5632 56457 5641 56491
rect 5641 56457 5675 56491
rect 5675 56457 5684 56491
rect 5632 56448 5684 56457
rect 7104 56448 7156 56500
rect 7288 56448 7340 56500
rect 7840 56448 7892 56500
rect 7012 56380 7064 56432
rect 6368 56244 6420 56296
rect 6736 56244 6788 56296
rect 7012 56287 7064 56296
rect 7012 56253 7021 56287
rect 7021 56253 7055 56287
rect 7055 56253 7064 56287
rect 7012 56244 7064 56253
rect 8300 56244 8352 56296
rect 8668 56448 8720 56500
rect 11888 56491 11940 56500
rect 11888 56457 11897 56491
rect 11897 56457 11931 56491
rect 11931 56457 11940 56491
rect 11888 56448 11940 56457
rect 10416 56380 10468 56432
rect 12072 56380 12124 56432
rect 9864 56244 9916 56296
rect 7472 56176 7524 56228
rect 10416 56176 10468 56228
rect 11152 56287 11204 56296
rect 11152 56253 11161 56287
rect 11161 56253 11195 56287
rect 11195 56253 11204 56287
rect 12532 56287 12584 56296
rect 11152 56244 11204 56253
rect 12532 56253 12541 56287
rect 12541 56253 12575 56287
rect 12575 56253 12584 56287
rect 12532 56244 12584 56253
rect 11888 56176 11940 56228
rect 13728 56176 13780 56228
rect 6184 56108 6236 56160
rect 6736 56108 6788 56160
rect 8944 56108 8996 56160
rect 9312 56151 9364 56160
rect 9312 56117 9321 56151
rect 9321 56117 9355 56151
rect 9355 56117 9364 56151
rect 9312 56108 9364 56117
rect 12532 56151 12584 56160
rect 12532 56117 12541 56151
rect 12541 56117 12575 56151
rect 12575 56117 12584 56151
rect 12532 56108 12584 56117
rect 12992 56108 13044 56160
rect 14188 56151 14240 56160
rect 14188 56117 14197 56151
rect 14197 56117 14231 56151
rect 14231 56117 14240 56151
rect 16396 56287 16448 56296
rect 16396 56253 16405 56287
rect 16405 56253 16439 56287
rect 16439 56253 16448 56287
rect 16396 56244 16448 56253
rect 14188 56108 14240 56117
rect 15660 56108 15712 56160
rect 17500 56151 17552 56160
rect 17500 56117 17509 56151
rect 17509 56117 17543 56151
rect 17543 56117 17552 56151
rect 17500 56108 17552 56117
rect 7648 56006 7700 56058
rect 7712 56006 7764 56058
rect 7776 56006 7828 56058
rect 7840 56006 7892 56058
rect 14315 56006 14367 56058
rect 14379 56006 14431 56058
rect 14443 56006 14495 56058
rect 14507 56006 14559 56058
rect 1676 55947 1728 55956
rect 1676 55913 1685 55947
rect 1685 55913 1719 55947
rect 1719 55913 1728 55947
rect 1676 55904 1728 55913
rect 2688 55904 2740 55956
rect 6276 55904 6328 55956
rect 6460 55947 6512 55956
rect 6460 55913 6469 55947
rect 6469 55913 6503 55947
rect 6503 55913 6512 55947
rect 6460 55904 6512 55913
rect 8300 55947 8352 55956
rect 8300 55913 8309 55947
rect 8309 55913 8343 55947
rect 8343 55913 8352 55947
rect 8300 55904 8352 55913
rect 8852 55947 8904 55956
rect 8852 55913 8861 55947
rect 8861 55913 8895 55947
rect 8895 55913 8904 55947
rect 8852 55904 8904 55913
rect 9496 55904 9548 55956
rect 1768 55836 1820 55888
rect 2412 55768 2464 55820
rect 2688 55768 2740 55820
rect 4896 55836 4948 55888
rect 6920 55836 6972 55888
rect 9680 55904 9732 55956
rect 10968 55904 11020 55956
rect 11152 55904 11204 55956
rect 12164 55904 12216 55956
rect 17316 55904 17368 55956
rect 4988 55811 5040 55820
rect 4988 55777 4997 55811
rect 4997 55777 5031 55811
rect 5031 55777 5040 55811
rect 4988 55768 5040 55777
rect 5172 55811 5224 55820
rect 5172 55777 5181 55811
rect 5181 55777 5215 55811
rect 5215 55777 5224 55811
rect 5172 55768 5224 55777
rect 4344 55632 4396 55684
rect 6184 55632 6236 55684
rect 7012 55768 7064 55820
rect 7472 55768 7524 55820
rect 6920 55743 6972 55752
rect 6920 55709 6929 55743
rect 6929 55709 6963 55743
rect 6963 55709 6972 55743
rect 6920 55700 6972 55709
rect 7288 55700 7340 55752
rect 9680 55768 9732 55820
rect 8852 55632 8904 55684
rect 9864 55768 9916 55820
rect 10324 55768 10376 55820
rect 12532 55836 12584 55888
rect 12716 55836 12768 55888
rect 13084 55836 13136 55888
rect 13728 55836 13780 55888
rect 12808 55768 12860 55820
rect 10508 55700 10560 55752
rect 10600 55743 10652 55752
rect 10600 55709 10609 55743
rect 10609 55709 10643 55743
rect 10643 55709 10652 55743
rect 10600 55700 10652 55709
rect 12072 55700 12124 55752
rect 12164 55700 12216 55752
rect 13084 55700 13136 55752
rect 14188 55768 14240 55820
rect 15384 55768 15436 55820
rect 17408 55768 17460 55820
rect 13912 55743 13964 55752
rect 13912 55709 13921 55743
rect 13921 55709 13955 55743
rect 13955 55709 13964 55743
rect 13912 55700 13964 55709
rect 15476 55700 15528 55752
rect 16304 55700 16356 55752
rect 17132 55743 17184 55752
rect 17132 55709 17141 55743
rect 17141 55709 17175 55743
rect 17175 55709 17184 55743
rect 17132 55700 17184 55709
rect 10876 55632 10928 55684
rect 4712 55564 4764 55616
rect 5724 55607 5776 55616
rect 5724 55573 5733 55607
rect 5733 55573 5767 55607
rect 5767 55573 5776 55607
rect 5724 55564 5776 55573
rect 6276 55564 6328 55616
rect 11888 55607 11940 55616
rect 11888 55573 11897 55607
rect 11897 55573 11931 55607
rect 11931 55573 11940 55607
rect 11888 55564 11940 55573
rect 12072 55564 12124 55616
rect 15292 55564 15344 55616
rect 4315 55462 4367 55514
rect 4379 55462 4431 55514
rect 4443 55462 4495 55514
rect 4507 55462 4559 55514
rect 10982 55462 11034 55514
rect 11046 55462 11098 55514
rect 11110 55462 11162 55514
rect 11174 55462 11226 55514
rect 17648 55462 17700 55514
rect 17712 55462 17764 55514
rect 17776 55462 17828 55514
rect 17840 55462 17892 55514
rect 1768 55360 1820 55412
rect 3148 55360 3200 55412
rect 3424 55403 3476 55412
rect 3424 55369 3433 55403
rect 3433 55369 3467 55403
rect 3467 55369 3476 55403
rect 3424 55360 3476 55369
rect 3516 55360 3568 55412
rect 3148 55156 3200 55208
rect 6092 55360 6144 55412
rect 8852 55360 8904 55412
rect 10324 55360 10376 55412
rect 10508 55403 10560 55412
rect 10508 55369 10517 55403
rect 10517 55369 10551 55403
rect 10551 55369 10560 55403
rect 10508 55360 10560 55369
rect 11520 55360 11572 55412
rect 12164 55360 12216 55412
rect 13912 55360 13964 55412
rect 5540 55292 5592 55344
rect 5172 55224 5224 55276
rect 5724 55224 5776 55276
rect 6092 55156 6144 55208
rect 6276 55199 6328 55208
rect 6276 55165 6285 55199
rect 6285 55165 6319 55199
rect 6319 55165 6328 55199
rect 6276 55156 6328 55165
rect 7012 55224 7064 55276
rect 9496 55292 9548 55344
rect 14188 55292 14240 55344
rect 8300 55224 8352 55276
rect 8668 55224 8720 55276
rect 8852 55224 8904 55276
rect 9312 55224 9364 55276
rect 11520 55267 11572 55276
rect 4712 55088 4764 55140
rect 5540 55088 5592 55140
rect 5724 55088 5776 55140
rect 7380 55131 7432 55140
rect 7380 55097 7389 55131
rect 7389 55097 7423 55131
rect 7423 55097 7432 55131
rect 7380 55088 7432 55097
rect 8392 55199 8444 55208
rect 8392 55165 8401 55199
rect 8401 55165 8435 55199
rect 8435 55165 8444 55199
rect 8392 55156 8444 55165
rect 11520 55233 11529 55267
rect 11529 55233 11563 55267
rect 11563 55233 11572 55267
rect 11520 55224 11572 55233
rect 9956 55156 10008 55208
rect 10876 55156 10928 55208
rect 12072 55224 12124 55276
rect 13820 55224 13872 55276
rect 16304 55360 16356 55412
rect 17132 55360 17184 55412
rect 2228 55020 2280 55072
rect 4436 55063 4488 55072
rect 4436 55029 4445 55063
rect 4445 55029 4479 55063
rect 4479 55029 4488 55063
rect 4436 55020 4488 55029
rect 4804 55020 4856 55072
rect 7288 55063 7340 55072
rect 7288 55029 7297 55063
rect 7297 55029 7331 55063
rect 7331 55029 7340 55063
rect 11980 55156 12032 55208
rect 14372 55199 14424 55208
rect 7288 55020 7340 55029
rect 9588 55020 9640 55072
rect 11428 55020 11480 55072
rect 11612 55020 11664 55072
rect 11888 55020 11940 55072
rect 13268 55088 13320 55140
rect 14372 55165 14381 55199
rect 14381 55165 14415 55199
rect 14415 55165 14424 55199
rect 14372 55156 14424 55165
rect 15384 55156 15436 55208
rect 17408 55224 17460 55276
rect 18144 55156 18196 55208
rect 12808 55063 12860 55072
rect 12808 55029 12817 55063
rect 12817 55029 12851 55063
rect 12851 55029 12860 55063
rect 12808 55020 12860 55029
rect 14740 55063 14792 55072
rect 14740 55029 14749 55063
rect 14749 55029 14783 55063
rect 14783 55029 14792 55063
rect 14740 55020 14792 55029
rect 16764 55020 16816 55072
rect 7648 54918 7700 54970
rect 7712 54918 7764 54970
rect 7776 54918 7828 54970
rect 7840 54918 7892 54970
rect 14315 54918 14367 54970
rect 14379 54918 14431 54970
rect 14443 54918 14495 54970
rect 14507 54918 14559 54970
rect 4896 54816 4948 54868
rect 11796 54859 11848 54868
rect 11796 54825 11805 54859
rect 11805 54825 11839 54859
rect 11839 54825 11848 54859
rect 11796 54816 11848 54825
rect 12716 54816 12768 54868
rect 12900 54816 12952 54868
rect 13820 54816 13872 54868
rect 9772 54748 9824 54800
rect 2412 54723 2464 54732
rect 2412 54689 2421 54723
rect 2421 54689 2455 54723
rect 2455 54689 2464 54723
rect 2412 54680 2464 54689
rect 2872 54723 2924 54732
rect 2872 54689 2881 54723
rect 2881 54689 2915 54723
rect 2915 54689 2924 54723
rect 2872 54680 2924 54689
rect 5540 54723 5592 54732
rect 5540 54689 5549 54723
rect 5549 54689 5583 54723
rect 5583 54689 5592 54723
rect 5540 54680 5592 54689
rect 8208 54680 8260 54732
rect 8392 54680 8444 54732
rect 8852 54723 8904 54732
rect 8852 54689 8861 54723
rect 8861 54689 8895 54723
rect 8895 54689 8904 54723
rect 8852 54680 8904 54689
rect 9036 54680 9088 54732
rect 10784 54680 10836 54732
rect 13084 54680 13136 54732
rect 7288 54655 7340 54664
rect 7288 54621 7297 54655
rect 7297 54621 7331 54655
rect 7331 54621 7340 54655
rect 7288 54612 7340 54621
rect 9496 54655 9548 54664
rect 9496 54621 9505 54655
rect 9505 54621 9539 54655
rect 9539 54621 9548 54655
rect 9496 54612 9548 54621
rect 10600 54612 10652 54664
rect 11428 54655 11480 54664
rect 11428 54621 11437 54655
rect 11437 54621 11471 54655
rect 11471 54621 11480 54655
rect 11428 54612 11480 54621
rect 16856 54723 16908 54732
rect 13728 54612 13780 54664
rect 16120 54655 16172 54664
rect 16120 54621 16129 54655
rect 16129 54621 16163 54655
rect 16163 54621 16172 54655
rect 16120 54612 16172 54621
rect 16856 54689 16865 54723
rect 16865 54689 16899 54723
rect 16899 54689 16908 54723
rect 16856 54680 16908 54689
rect 17132 54612 17184 54664
rect 1492 54544 1544 54596
rect 5816 54544 5868 54596
rect 6920 54544 6972 54596
rect 12900 54544 12952 54596
rect 13268 54544 13320 54596
rect 16396 54544 16448 54596
rect 16948 54587 17000 54596
rect 16948 54553 16957 54587
rect 16957 54553 16991 54587
rect 16991 54553 17000 54587
rect 16948 54544 17000 54553
rect 1768 54476 1820 54528
rect 4068 54476 4120 54528
rect 5724 54476 5776 54528
rect 6368 54476 6420 54528
rect 6736 54476 6788 54528
rect 8300 54519 8352 54528
rect 8300 54485 8309 54519
rect 8309 54485 8343 54519
rect 8343 54485 8352 54519
rect 8300 54476 8352 54485
rect 8576 54476 8628 54528
rect 9036 54476 9088 54528
rect 9496 54476 9548 54528
rect 9772 54476 9824 54528
rect 10876 54476 10928 54528
rect 12624 54519 12676 54528
rect 12624 54485 12633 54519
rect 12633 54485 12667 54519
rect 12667 54485 12676 54519
rect 12624 54476 12676 54485
rect 13452 54476 13504 54528
rect 15936 54476 15988 54528
rect 4315 54374 4367 54426
rect 4379 54374 4431 54426
rect 4443 54374 4495 54426
rect 4507 54374 4559 54426
rect 10982 54374 11034 54426
rect 11046 54374 11098 54426
rect 11110 54374 11162 54426
rect 11174 54374 11226 54426
rect 17648 54374 17700 54426
rect 17712 54374 17764 54426
rect 17776 54374 17828 54426
rect 17840 54374 17892 54426
rect 2872 54315 2924 54324
rect 2872 54281 2881 54315
rect 2881 54281 2915 54315
rect 2915 54281 2924 54315
rect 2872 54272 2924 54281
rect 5540 54272 5592 54324
rect 6184 54272 6236 54324
rect 9220 54272 9272 54324
rect 6736 54204 6788 54256
rect 1584 54179 1636 54188
rect 1584 54145 1593 54179
rect 1593 54145 1627 54179
rect 1627 54145 1636 54179
rect 1584 54136 1636 54145
rect 1676 54136 1728 54188
rect 2228 54136 2280 54188
rect 6920 54136 6972 54188
rect 1492 54111 1544 54120
rect 1492 54077 1501 54111
rect 1501 54077 1535 54111
rect 1535 54077 1544 54111
rect 1492 54068 1544 54077
rect 1768 54068 1820 54120
rect 3516 54068 3568 54120
rect 4712 54068 4764 54120
rect 6184 54068 6236 54120
rect 6460 54068 6512 54120
rect 7840 54068 7892 54120
rect 8300 54136 8352 54188
rect 10784 54272 10836 54324
rect 11980 54272 12032 54324
rect 12532 54272 12584 54324
rect 16856 54272 16908 54324
rect 9772 54204 9824 54256
rect 10140 54204 10192 54256
rect 10324 54204 10376 54256
rect 12532 54179 12584 54188
rect 12532 54145 12541 54179
rect 12541 54145 12575 54179
rect 12575 54145 12584 54179
rect 12532 54136 12584 54145
rect 15844 54179 15896 54188
rect 15844 54145 15853 54179
rect 15853 54145 15887 54179
rect 15887 54145 15896 54179
rect 15844 54136 15896 54145
rect 4528 54000 4580 54052
rect 8392 54068 8444 54120
rect 9496 54068 9548 54120
rect 9680 54068 9732 54120
rect 10140 54068 10192 54120
rect 11704 54068 11756 54120
rect 11888 54068 11940 54120
rect 12164 54068 12216 54120
rect 12348 54068 12400 54120
rect 12624 54111 12676 54120
rect 12624 54077 12633 54111
rect 12633 54077 12667 54111
rect 12667 54077 12676 54111
rect 12624 54068 12676 54077
rect 12900 54111 12952 54120
rect 12900 54077 12909 54111
rect 12909 54077 12943 54111
rect 12943 54077 12952 54111
rect 12900 54068 12952 54077
rect 14096 54111 14148 54120
rect 14096 54077 14105 54111
rect 14105 54077 14139 54111
rect 14139 54077 14148 54111
rect 14096 54068 14148 54077
rect 15292 54111 15344 54120
rect 15292 54077 15301 54111
rect 15301 54077 15335 54111
rect 15335 54077 15344 54111
rect 15292 54068 15344 54077
rect 15936 54111 15988 54120
rect 15936 54077 15945 54111
rect 15945 54077 15979 54111
rect 15979 54077 15988 54111
rect 15936 54068 15988 54077
rect 16396 54068 16448 54120
rect 16672 54111 16724 54120
rect 16672 54077 16681 54111
rect 16681 54077 16715 54111
rect 16715 54077 16724 54111
rect 16672 54068 16724 54077
rect 8300 54000 8352 54052
rect 4252 53932 4304 53984
rect 6184 53975 6236 53984
rect 6184 53941 6193 53975
rect 6193 53941 6227 53975
rect 6227 53941 6236 53975
rect 6184 53932 6236 53941
rect 8576 53975 8628 53984
rect 8576 53941 8585 53975
rect 8585 53941 8619 53975
rect 8619 53941 8628 53975
rect 8576 53932 8628 53941
rect 10600 53932 10652 53984
rect 11152 53975 11204 53984
rect 11152 53941 11161 53975
rect 11161 53941 11195 53975
rect 11195 53941 11204 53975
rect 11152 53932 11204 53941
rect 12440 53932 12492 53984
rect 13728 53932 13780 53984
rect 14004 53932 14056 53984
rect 15108 53975 15160 53984
rect 15108 53941 15117 53975
rect 15117 53941 15151 53975
rect 15151 53941 15160 53975
rect 15108 53932 15160 53941
rect 16120 53932 16172 53984
rect 17132 53932 17184 53984
rect 7648 53830 7700 53882
rect 7712 53830 7764 53882
rect 7776 53830 7828 53882
rect 7840 53830 7892 53882
rect 14315 53830 14367 53882
rect 14379 53830 14431 53882
rect 14443 53830 14495 53882
rect 14507 53830 14559 53882
rect 1676 53771 1728 53780
rect 1676 53737 1685 53771
rect 1685 53737 1719 53771
rect 1719 53737 1728 53771
rect 1676 53728 1728 53737
rect 6460 53728 6512 53780
rect 2228 53660 2280 53712
rect 2872 53660 2924 53712
rect 3056 53592 3108 53644
rect 4252 53660 4304 53712
rect 4528 53660 4580 53712
rect 5172 53660 5224 53712
rect 5540 53660 5592 53712
rect 8668 53728 8720 53780
rect 9680 53728 9732 53780
rect 11152 53728 11204 53780
rect 11428 53728 11480 53780
rect 12256 53728 12308 53780
rect 12532 53728 12584 53780
rect 14188 53728 14240 53780
rect 4896 53635 4948 53644
rect 3608 53524 3660 53576
rect 4896 53601 4905 53635
rect 4905 53601 4939 53635
rect 4939 53601 4948 53635
rect 4896 53592 4948 53601
rect 5816 53592 5868 53644
rect 6184 53592 6236 53644
rect 9588 53660 9640 53712
rect 10876 53660 10928 53712
rect 8668 53635 8720 53644
rect 2412 53388 2464 53440
rect 2780 53431 2832 53440
rect 2780 53397 2789 53431
rect 2789 53397 2823 53431
rect 2823 53397 2832 53431
rect 2780 53388 2832 53397
rect 3148 53388 3200 53440
rect 5540 53524 5592 53576
rect 6920 53524 6972 53576
rect 8668 53601 8677 53635
rect 8677 53601 8711 53635
rect 8711 53601 8720 53635
rect 8668 53592 8720 53601
rect 8852 53635 8904 53644
rect 8852 53601 8861 53635
rect 8861 53601 8895 53635
rect 8895 53601 8904 53635
rect 8852 53592 8904 53601
rect 9496 53635 9548 53644
rect 9496 53601 9505 53635
rect 9505 53601 9539 53635
rect 9539 53601 9548 53635
rect 9496 53592 9548 53601
rect 10600 53635 10652 53644
rect 10600 53601 10609 53635
rect 10609 53601 10643 53635
rect 10643 53601 10652 53635
rect 10600 53592 10652 53601
rect 10784 53635 10836 53644
rect 10784 53601 10793 53635
rect 10793 53601 10827 53635
rect 10827 53601 10836 53635
rect 10784 53592 10836 53601
rect 11612 53592 11664 53644
rect 12808 53635 12860 53644
rect 8116 53524 8168 53576
rect 10140 53567 10192 53576
rect 10140 53533 10149 53567
rect 10149 53533 10183 53567
rect 10183 53533 10192 53567
rect 10140 53524 10192 53533
rect 11888 53524 11940 53576
rect 12072 53524 12124 53576
rect 12808 53601 12817 53635
rect 12817 53601 12851 53635
rect 12851 53601 12860 53635
rect 12808 53592 12860 53601
rect 12900 53567 12952 53576
rect 12900 53533 12909 53567
rect 12909 53533 12943 53567
rect 12943 53533 12952 53567
rect 12900 53524 12952 53533
rect 4344 53499 4396 53508
rect 4344 53465 4353 53499
rect 4353 53465 4387 53499
rect 4387 53465 4396 53499
rect 4344 53456 4396 53465
rect 7472 53456 7524 53508
rect 4988 53431 5040 53440
rect 4988 53397 4997 53431
rect 4997 53397 5031 53431
rect 5031 53397 5040 53431
rect 4988 53388 5040 53397
rect 6092 53431 6144 53440
rect 6092 53397 6101 53431
rect 6101 53397 6135 53431
rect 6135 53397 6144 53431
rect 6092 53388 6144 53397
rect 6644 53431 6696 53440
rect 6644 53397 6653 53431
rect 6653 53397 6687 53431
rect 6687 53397 6696 53431
rect 6644 53388 6696 53397
rect 7380 53388 7432 53440
rect 9220 53456 9272 53508
rect 9588 53456 9640 53508
rect 12440 53456 12492 53508
rect 12808 53456 12860 53508
rect 8392 53388 8444 53440
rect 10140 53388 10192 53440
rect 10324 53388 10376 53440
rect 12900 53388 12952 53440
rect 13084 53592 13136 53644
rect 14648 53592 14700 53644
rect 15292 53635 15344 53644
rect 15292 53601 15301 53635
rect 15301 53601 15335 53635
rect 15335 53601 15344 53635
rect 15292 53592 15344 53601
rect 15936 53635 15988 53644
rect 15936 53601 15945 53635
rect 15945 53601 15979 53635
rect 15979 53601 15988 53635
rect 15936 53592 15988 53601
rect 16212 53635 16264 53644
rect 16212 53601 16221 53635
rect 16221 53601 16255 53635
rect 16255 53601 16264 53635
rect 16212 53592 16264 53601
rect 16672 53524 16724 53576
rect 14096 53456 14148 53508
rect 15108 53499 15160 53508
rect 15108 53465 15117 53499
rect 15117 53465 15151 53499
rect 15151 53465 15160 53499
rect 15108 53456 15160 53465
rect 14648 53388 14700 53440
rect 16580 53388 16632 53440
rect 17040 53431 17092 53440
rect 17040 53397 17049 53431
rect 17049 53397 17083 53431
rect 17083 53397 17092 53431
rect 17040 53388 17092 53397
rect 4315 53286 4367 53338
rect 4379 53286 4431 53338
rect 4443 53286 4495 53338
rect 4507 53286 4559 53338
rect 10982 53286 11034 53338
rect 11046 53286 11098 53338
rect 11110 53286 11162 53338
rect 11174 53286 11226 53338
rect 17648 53286 17700 53338
rect 17712 53286 17764 53338
rect 17776 53286 17828 53338
rect 17840 53286 17892 53338
rect 2412 53184 2464 53236
rect 4896 53184 4948 53236
rect 8116 53184 8168 53236
rect 8668 53184 8720 53236
rect 8852 53227 8904 53236
rect 8852 53193 8861 53227
rect 8861 53193 8895 53227
rect 8895 53193 8904 53227
rect 8852 53184 8904 53193
rect 9496 53184 9548 53236
rect 10600 53184 10652 53236
rect 6920 53159 6972 53168
rect 6920 53125 6929 53159
rect 6929 53125 6963 53159
rect 6963 53125 6972 53159
rect 6920 53116 6972 53125
rect 7380 53116 7432 53168
rect 11428 53184 11480 53236
rect 11244 53116 11296 53168
rect 1676 53048 1728 53100
rect 6644 53048 6696 53100
rect 7472 53048 7524 53100
rect 10232 53091 10284 53100
rect 10232 53057 10241 53091
rect 10241 53057 10275 53091
rect 10275 53057 10284 53091
rect 10232 53048 10284 53057
rect 11796 53116 11848 53168
rect 17040 53184 17092 53236
rect 14648 53116 14700 53168
rect 13176 53091 13228 53100
rect 2412 52980 2464 53032
rect 4068 52980 4120 53032
rect 4528 53023 4580 53032
rect 4528 52989 4537 53023
rect 4537 52989 4571 53023
rect 4571 52989 4580 53023
rect 4528 52980 4580 52989
rect 3148 52844 3200 52896
rect 3516 52887 3568 52896
rect 3516 52853 3525 52887
rect 3525 52853 3559 52887
rect 3559 52853 3568 52887
rect 3516 52844 3568 52853
rect 4068 52844 4120 52896
rect 5540 52844 5592 52896
rect 5632 52844 5684 52896
rect 7012 52980 7064 53032
rect 7104 52980 7156 53032
rect 6644 52912 6696 52964
rect 6828 52912 6880 52964
rect 9220 52912 9272 52964
rect 11612 52980 11664 53032
rect 11796 52980 11848 53032
rect 13176 53057 13185 53091
rect 13185 53057 13219 53091
rect 13219 53057 13228 53091
rect 13176 53048 13228 53057
rect 6368 52844 6420 52896
rect 6552 52844 6604 52896
rect 7380 52844 7432 52896
rect 8208 52844 8260 52896
rect 10600 52844 10652 52896
rect 11336 52912 11388 52964
rect 11520 52912 11572 52964
rect 12072 52844 12124 52896
rect 12532 52844 12584 52896
rect 13176 52912 13228 52964
rect 14188 53048 14240 53100
rect 14740 53048 14792 53100
rect 15292 53048 15344 53100
rect 14556 52980 14608 53032
rect 15568 53023 15620 53032
rect 15568 52989 15577 53023
rect 15577 52989 15611 53023
rect 15611 52989 15620 53023
rect 15568 52980 15620 52989
rect 15936 53023 15988 53032
rect 15936 52989 15945 53023
rect 15945 52989 15979 53023
rect 15979 52989 15988 53023
rect 15936 52980 15988 52989
rect 16672 53023 16724 53032
rect 15016 52912 15068 52964
rect 16672 52989 16681 53023
rect 16681 52989 16715 53023
rect 16715 52989 16724 53023
rect 16672 52980 16724 52989
rect 17960 53023 18012 53032
rect 17960 52989 17969 53023
rect 17969 52989 18003 53023
rect 18003 52989 18012 53023
rect 17960 52980 18012 52989
rect 13084 52844 13136 52896
rect 14188 52887 14240 52896
rect 14188 52853 14197 52887
rect 14197 52853 14231 52887
rect 14231 52853 14240 52887
rect 14188 52844 14240 52853
rect 15936 52844 15988 52896
rect 17960 52844 18012 52896
rect 7648 52742 7700 52794
rect 7712 52742 7764 52794
rect 7776 52742 7828 52794
rect 7840 52742 7892 52794
rect 14315 52742 14367 52794
rect 14379 52742 14431 52794
rect 14443 52742 14495 52794
rect 14507 52742 14559 52794
rect 3056 52640 3108 52692
rect 1676 52615 1728 52624
rect 1676 52581 1685 52615
rect 1685 52581 1719 52615
rect 1719 52581 1728 52615
rect 1676 52572 1728 52581
rect 3148 52547 3200 52556
rect 3148 52513 3157 52547
rect 3157 52513 3191 52547
rect 3191 52513 3200 52547
rect 3148 52504 3200 52513
rect 3056 52436 3108 52488
rect 3516 52640 3568 52692
rect 4712 52683 4764 52692
rect 4712 52649 4721 52683
rect 4721 52649 4755 52683
rect 4755 52649 4764 52683
rect 4712 52640 4764 52649
rect 5172 52683 5224 52692
rect 5172 52649 5181 52683
rect 5181 52649 5215 52683
rect 5215 52649 5224 52683
rect 5172 52640 5224 52649
rect 5540 52640 5592 52692
rect 6368 52640 6420 52692
rect 7472 52640 7524 52692
rect 9220 52640 9272 52692
rect 10784 52640 10836 52692
rect 12164 52640 12216 52692
rect 16212 52683 16264 52692
rect 4528 52572 4580 52624
rect 8208 52572 8260 52624
rect 11244 52572 11296 52624
rect 11704 52572 11756 52624
rect 3516 52436 3568 52488
rect 7104 52436 7156 52488
rect 7472 52479 7524 52488
rect 7472 52445 7481 52479
rect 7481 52445 7515 52479
rect 7515 52445 7524 52479
rect 7472 52436 7524 52445
rect 8208 52436 8260 52488
rect 8392 52504 8444 52556
rect 8852 52504 8904 52556
rect 9956 52504 10008 52556
rect 10784 52547 10836 52556
rect 10784 52513 10793 52547
rect 10793 52513 10827 52547
rect 10827 52513 10836 52547
rect 10784 52504 10836 52513
rect 10876 52504 10928 52556
rect 11428 52504 11480 52556
rect 13268 52572 13320 52624
rect 13912 52572 13964 52624
rect 13452 52504 13504 52556
rect 14648 52547 14700 52556
rect 14648 52513 14657 52547
rect 14657 52513 14691 52547
rect 14691 52513 14700 52547
rect 14648 52504 14700 52513
rect 15016 52547 15068 52556
rect 15016 52513 15025 52547
rect 15025 52513 15059 52547
rect 15059 52513 15068 52547
rect 15016 52504 15068 52513
rect 15108 52504 15160 52556
rect 10140 52479 10192 52488
rect 10140 52445 10149 52479
rect 10149 52445 10183 52479
rect 10183 52445 10192 52479
rect 10140 52436 10192 52445
rect 8392 52368 8444 52420
rect 8760 52368 8812 52420
rect 10508 52368 10560 52420
rect 2412 52300 2464 52352
rect 6092 52343 6144 52352
rect 6092 52309 6101 52343
rect 6101 52309 6135 52343
rect 6135 52309 6144 52343
rect 6092 52300 6144 52309
rect 9956 52300 10008 52352
rect 11888 52436 11940 52488
rect 12256 52436 12308 52488
rect 12900 52436 12952 52488
rect 15476 52436 15528 52488
rect 11796 52368 11848 52420
rect 13268 52368 13320 52420
rect 13452 52368 13504 52420
rect 14096 52368 14148 52420
rect 16212 52649 16221 52683
rect 16221 52649 16255 52683
rect 16255 52649 16264 52683
rect 16212 52640 16264 52649
rect 16856 52504 16908 52556
rect 17132 52411 17184 52420
rect 17132 52377 17141 52411
rect 17141 52377 17175 52411
rect 17175 52377 17184 52411
rect 17132 52368 17184 52377
rect 12256 52300 12308 52352
rect 14280 52300 14332 52352
rect 14740 52300 14792 52352
rect 15936 52300 15988 52352
rect 4315 52198 4367 52250
rect 4379 52198 4431 52250
rect 4443 52198 4495 52250
rect 4507 52198 4559 52250
rect 10982 52198 11034 52250
rect 11046 52198 11098 52250
rect 11110 52198 11162 52250
rect 11174 52198 11226 52250
rect 17648 52198 17700 52250
rect 17712 52198 17764 52250
rect 17776 52198 17828 52250
rect 17840 52198 17892 52250
rect 4160 51960 4212 52012
rect 4988 51960 5040 52012
rect 6552 52096 6604 52148
rect 8392 52139 8444 52148
rect 8392 52105 8401 52139
rect 8401 52105 8435 52139
rect 8435 52105 8444 52139
rect 8392 52096 8444 52105
rect 8852 52096 8904 52148
rect 9036 52096 9088 52148
rect 10876 52096 10928 52148
rect 11336 52096 11388 52148
rect 13912 52096 13964 52148
rect 14004 52096 14056 52148
rect 15108 52096 15160 52148
rect 16856 52096 16908 52148
rect 17960 52139 18012 52148
rect 17960 52105 17969 52139
rect 17969 52105 18003 52139
rect 18003 52105 18012 52139
rect 17960 52096 18012 52105
rect 5540 51960 5592 52012
rect 6184 52028 6236 52080
rect 6828 52028 6880 52080
rect 7012 52071 7064 52080
rect 7012 52037 7021 52071
rect 7021 52037 7055 52071
rect 7055 52037 7064 52071
rect 7012 52028 7064 52037
rect 8760 52028 8812 52080
rect 11244 52028 11296 52080
rect 11612 52028 11664 52080
rect 13820 52028 13872 52080
rect 4528 51892 4580 51944
rect 6092 51935 6144 51944
rect 6092 51901 6101 51935
rect 6101 51901 6135 51935
rect 6135 51901 6144 51935
rect 6092 51892 6144 51901
rect 6552 51935 6604 51944
rect 6552 51901 6561 51935
rect 6561 51901 6595 51935
rect 6595 51901 6604 51935
rect 6552 51892 6604 51901
rect 4160 51824 4212 51876
rect 5080 51824 5132 51876
rect 6828 51824 6880 51876
rect 2780 51799 2832 51808
rect 2780 51765 2789 51799
rect 2789 51765 2823 51799
rect 2823 51765 2832 51799
rect 2780 51756 2832 51765
rect 4712 51756 4764 51808
rect 4804 51756 4856 51808
rect 5264 51756 5316 51808
rect 6460 51756 6512 51808
rect 9588 51892 9640 51944
rect 9956 51892 10008 51944
rect 10232 51892 10284 51944
rect 10876 51892 10928 51944
rect 11428 51935 11480 51944
rect 11428 51901 11437 51935
rect 11437 51901 11471 51935
rect 11471 51901 11480 51935
rect 11428 51892 11480 51901
rect 12256 51960 12308 52012
rect 12900 52003 12952 52012
rect 12900 51969 12909 52003
rect 12909 51969 12943 52003
rect 12943 51969 12952 52003
rect 16304 52028 16356 52080
rect 16672 52028 16724 52080
rect 12900 51960 12952 51969
rect 10600 51867 10652 51876
rect 10600 51833 10609 51867
rect 10609 51833 10643 51867
rect 10643 51833 10652 51867
rect 10600 51824 10652 51833
rect 10968 51824 11020 51876
rect 13176 51892 13228 51944
rect 13912 51935 13964 51944
rect 13912 51901 13921 51935
rect 13921 51901 13955 51935
rect 13955 51901 13964 51935
rect 13912 51892 13964 51901
rect 14648 51960 14700 52012
rect 14280 51892 14332 51944
rect 15384 51892 15436 51944
rect 15568 51892 15620 51944
rect 15936 51960 15988 52012
rect 16212 51935 16264 51944
rect 16212 51901 16221 51935
rect 16221 51901 16255 51935
rect 16255 51901 16264 51935
rect 16212 51892 16264 51901
rect 16764 51935 16816 51944
rect 8208 51756 8260 51808
rect 8392 51756 8444 51808
rect 10784 51756 10836 51808
rect 11428 51756 11480 51808
rect 11612 51756 11664 51808
rect 13728 51824 13780 51876
rect 16764 51901 16773 51935
rect 16773 51901 16807 51935
rect 16807 51901 16816 51935
rect 16764 51892 16816 51901
rect 17408 51824 17460 51876
rect 7648 51654 7700 51706
rect 7712 51654 7764 51706
rect 7776 51654 7828 51706
rect 7840 51654 7892 51706
rect 14315 51654 14367 51706
rect 14379 51654 14431 51706
rect 14443 51654 14495 51706
rect 14507 51654 14559 51706
rect 1584 51552 1636 51604
rect 3148 51595 3200 51604
rect 3148 51561 3157 51595
rect 3157 51561 3191 51595
rect 3191 51561 3200 51595
rect 3148 51552 3200 51561
rect 6184 51595 6236 51604
rect 6184 51561 6193 51595
rect 6193 51561 6227 51595
rect 6227 51561 6236 51595
rect 6184 51552 6236 51561
rect 8944 51552 8996 51604
rect 9956 51552 10008 51604
rect 10324 51552 10376 51604
rect 10968 51552 11020 51604
rect 7012 51484 7064 51536
rect 7564 51484 7616 51536
rect 8116 51484 8168 51536
rect 8668 51484 8720 51536
rect 9036 51484 9088 51536
rect 3148 51416 3200 51468
rect 3792 51416 3844 51468
rect 5172 51459 5224 51468
rect 5172 51425 5181 51459
rect 5181 51425 5215 51459
rect 5215 51425 5224 51459
rect 5172 51416 5224 51425
rect 4068 51348 4120 51400
rect 3056 51280 3108 51332
rect 3792 51280 3844 51332
rect 3516 51212 3568 51264
rect 4528 51280 4580 51332
rect 5080 51280 5132 51332
rect 5448 51416 5500 51468
rect 6092 51416 6144 51468
rect 7748 51416 7800 51468
rect 7932 51459 7984 51468
rect 7932 51425 7941 51459
rect 7941 51425 7975 51459
rect 7975 51425 7984 51459
rect 7932 51416 7984 51425
rect 9220 51459 9272 51468
rect 6828 51348 6880 51400
rect 7012 51348 7064 51400
rect 8116 51348 8168 51400
rect 9220 51425 9229 51459
rect 9229 51425 9263 51459
rect 9263 51425 9272 51459
rect 9220 51416 9272 51425
rect 9588 51484 9640 51536
rect 9772 51484 9824 51536
rect 10508 51484 10560 51536
rect 10324 51416 10376 51468
rect 10968 51459 11020 51468
rect 10968 51425 10977 51459
rect 10977 51425 11011 51459
rect 11011 51425 11020 51459
rect 10968 51416 11020 51425
rect 5448 51280 5500 51332
rect 7472 51280 7524 51332
rect 5540 51212 5592 51264
rect 6368 51212 6420 51264
rect 7748 51212 7800 51264
rect 8760 51212 8812 51264
rect 10140 51348 10192 51400
rect 9772 51280 9824 51332
rect 11336 51552 11388 51604
rect 12164 51527 12216 51536
rect 11336 51416 11388 51468
rect 12164 51493 12173 51527
rect 12173 51493 12207 51527
rect 12207 51493 12216 51527
rect 12164 51484 12216 51493
rect 12440 51484 12492 51536
rect 13912 51552 13964 51604
rect 15016 51552 15068 51604
rect 17132 51595 17184 51604
rect 17132 51561 17141 51595
rect 17141 51561 17175 51595
rect 17175 51561 17184 51595
rect 17132 51552 17184 51561
rect 17500 51595 17552 51604
rect 17500 51561 17509 51595
rect 17509 51561 17543 51595
rect 17543 51561 17552 51595
rect 17500 51552 17552 51561
rect 12900 51484 12952 51536
rect 11612 51348 11664 51400
rect 12256 51416 12308 51468
rect 12532 51416 12584 51468
rect 17040 51484 17092 51536
rect 15568 51459 15620 51468
rect 15568 51425 15577 51459
rect 15577 51425 15611 51459
rect 15611 51425 15620 51459
rect 15568 51416 15620 51425
rect 16028 51459 16080 51468
rect 16028 51425 16037 51459
rect 16037 51425 16071 51459
rect 16071 51425 16080 51459
rect 16028 51416 16080 51425
rect 16212 51459 16264 51468
rect 16212 51425 16221 51459
rect 16221 51425 16255 51459
rect 16255 51425 16264 51459
rect 16212 51416 16264 51425
rect 16396 51416 16448 51468
rect 16764 51459 16816 51468
rect 16764 51425 16773 51459
rect 16773 51425 16807 51459
rect 16807 51425 16816 51459
rect 16764 51416 16816 51425
rect 17316 51416 17368 51468
rect 12900 51391 12952 51400
rect 12900 51357 12909 51391
rect 12909 51357 12943 51391
rect 12943 51357 12952 51391
rect 12900 51348 12952 51357
rect 13176 51391 13228 51400
rect 13176 51357 13185 51391
rect 13185 51357 13219 51391
rect 13219 51357 13228 51391
rect 13176 51348 13228 51357
rect 15384 51348 15436 51400
rect 12072 51212 12124 51264
rect 12624 51212 12676 51264
rect 13268 51212 13320 51264
rect 15384 51212 15436 51264
rect 4315 51110 4367 51162
rect 4379 51110 4431 51162
rect 4443 51110 4495 51162
rect 4507 51110 4559 51162
rect 10982 51110 11034 51162
rect 11046 51110 11098 51162
rect 11110 51110 11162 51162
rect 11174 51110 11226 51162
rect 17648 51110 17700 51162
rect 17712 51110 17764 51162
rect 17776 51110 17828 51162
rect 17840 51110 17892 51162
rect 3240 51008 3292 51060
rect 4068 51008 4120 51060
rect 4528 50940 4580 50992
rect 5172 51008 5224 51060
rect 5724 51008 5776 51060
rect 6092 51008 6144 51060
rect 7564 51008 7616 51060
rect 7840 51008 7892 51060
rect 5540 50940 5592 50992
rect 7472 50940 7524 50992
rect 7932 50940 7984 50992
rect 8208 51008 8260 51060
rect 9220 51008 9272 51060
rect 9680 51008 9732 51060
rect 9772 51008 9824 51060
rect 10324 51008 10376 51060
rect 11980 51008 12032 51060
rect 12440 51051 12492 51060
rect 12440 51017 12449 51051
rect 12449 51017 12483 51051
rect 12483 51017 12492 51051
rect 12440 51008 12492 51017
rect 12808 51008 12860 51060
rect 13176 51051 13228 51060
rect 13176 51017 13185 51051
rect 13185 51017 13219 51051
rect 13219 51017 13228 51051
rect 13176 51008 13228 51017
rect 13452 51008 13504 51060
rect 13728 51008 13780 51060
rect 15292 51008 15344 51060
rect 1584 50804 1636 50856
rect 1768 50847 1820 50856
rect 1768 50813 1777 50847
rect 1777 50813 1811 50847
rect 1811 50813 1820 50847
rect 1768 50804 1820 50813
rect 2228 50804 2280 50856
rect 5172 50804 5224 50856
rect 5816 50872 5868 50924
rect 7196 50872 7248 50924
rect 5632 50804 5684 50856
rect 6460 50804 6512 50856
rect 7012 50804 7064 50856
rect 7472 50804 7524 50856
rect 7748 50847 7800 50856
rect 7748 50813 7757 50847
rect 7757 50813 7791 50847
rect 7791 50813 7800 50847
rect 7748 50804 7800 50813
rect 8576 50872 8628 50924
rect 11612 50872 11664 50924
rect 8760 50847 8812 50856
rect 2412 50668 2464 50720
rect 4252 50711 4304 50720
rect 4252 50677 4261 50711
rect 4261 50677 4295 50711
rect 4295 50677 4304 50711
rect 4252 50668 4304 50677
rect 6736 50736 6788 50788
rect 5632 50711 5684 50720
rect 5632 50677 5641 50711
rect 5641 50677 5675 50711
rect 5675 50677 5684 50711
rect 5632 50668 5684 50677
rect 7380 50736 7432 50788
rect 8208 50736 8260 50788
rect 8760 50813 8769 50847
rect 8769 50813 8803 50847
rect 8803 50813 8812 50847
rect 8760 50804 8812 50813
rect 7012 50711 7064 50720
rect 7012 50677 7021 50711
rect 7021 50677 7055 50711
rect 7055 50677 7064 50711
rect 7012 50668 7064 50677
rect 7288 50711 7340 50720
rect 7288 50677 7297 50711
rect 7297 50677 7331 50711
rect 7331 50677 7340 50711
rect 7288 50668 7340 50677
rect 8484 50668 8536 50720
rect 8944 50711 8996 50720
rect 8944 50677 8953 50711
rect 8953 50677 8987 50711
rect 8987 50677 8996 50711
rect 8944 50668 8996 50677
rect 9772 50668 9824 50720
rect 10324 50804 10376 50856
rect 10508 50847 10560 50856
rect 10508 50813 10517 50847
rect 10517 50813 10551 50847
rect 10551 50813 10560 50847
rect 10508 50804 10560 50813
rect 11244 50847 11296 50856
rect 10692 50736 10744 50788
rect 11244 50813 11253 50847
rect 11253 50813 11287 50847
rect 11287 50813 11296 50847
rect 11244 50804 11296 50813
rect 17040 50940 17092 50992
rect 13176 50872 13228 50924
rect 15016 50872 15068 50924
rect 15108 50872 15160 50924
rect 15752 50872 15804 50924
rect 17316 50872 17368 50924
rect 13728 50804 13780 50856
rect 13912 50847 13964 50856
rect 13912 50813 13921 50847
rect 13921 50813 13955 50847
rect 13955 50813 13964 50847
rect 13912 50804 13964 50813
rect 16580 50804 16632 50856
rect 17132 50847 17184 50856
rect 13268 50736 13320 50788
rect 10324 50711 10376 50720
rect 10324 50677 10333 50711
rect 10333 50677 10367 50711
rect 10367 50677 10376 50711
rect 10324 50668 10376 50677
rect 12808 50668 12860 50720
rect 12900 50668 12952 50720
rect 14832 50668 14884 50720
rect 15292 50668 15344 50720
rect 15476 50711 15528 50720
rect 15476 50677 15485 50711
rect 15485 50677 15519 50711
rect 15519 50677 15528 50711
rect 15476 50668 15528 50677
rect 16580 50711 16632 50720
rect 16580 50677 16589 50711
rect 16589 50677 16623 50711
rect 16623 50677 16632 50711
rect 17132 50813 17141 50847
rect 17141 50813 17175 50847
rect 17175 50813 17184 50847
rect 17132 50804 17184 50813
rect 17500 50847 17552 50856
rect 17500 50813 17509 50847
rect 17509 50813 17543 50847
rect 17543 50813 17552 50847
rect 17500 50804 17552 50813
rect 18052 50711 18104 50720
rect 16580 50668 16632 50677
rect 18052 50677 18061 50711
rect 18061 50677 18095 50711
rect 18095 50677 18104 50711
rect 18052 50668 18104 50677
rect 7648 50566 7700 50618
rect 7712 50566 7764 50618
rect 7776 50566 7828 50618
rect 7840 50566 7892 50618
rect 14315 50566 14367 50618
rect 14379 50566 14431 50618
rect 14443 50566 14495 50618
rect 14507 50566 14559 50618
rect 4896 50464 4948 50516
rect 5172 50464 5224 50516
rect 5540 50507 5592 50516
rect 5540 50473 5549 50507
rect 5549 50473 5583 50507
rect 5583 50473 5592 50507
rect 5540 50464 5592 50473
rect 7380 50464 7432 50516
rect 8208 50464 8260 50516
rect 8300 50464 8352 50516
rect 3700 50396 3752 50448
rect 6828 50396 6880 50448
rect 7196 50396 7248 50448
rect 9404 50464 9456 50516
rect 10784 50507 10836 50516
rect 10784 50473 10793 50507
rect 10793 50473 10827 50507
rect 10827 50473 10836 50507
rect 10784 50464 10836 50473
rect 11244 50464 11296 50516
rect 4068 50371 4120 50380
rect 4068 50337 4077 50371
rect 4077 50337 4111 50371
rect 4111 50337 4120 50371
rect 4068 50328 4120 50337
rect 4160 50371 4212 50380
rect 4160 50337 4169 50371
rect 4169 50337 4203 50371
rect 4203 50337 4212 50371
rect 4160 50328 4212 50337
rect 3240 50303 3292 50312
rect 3240 50269 3249 50303
rect 3249 50269 3283 50303
rect 3283 50269 3292 50303
rect 3240 50260 3292 50269
rect 3516 50260 3568 50312
rect 3700 50260 3752 50312
rect 4252 50260 4304 50312
rect 6368 50260 6420 50312
rect 7196 50260 7248 50312
rect 10140 50396 10192 50448
rect 7472 50192 7524 50244
rect 8300 50192 8352 50244
rect 9220 50371 9272 50380
rect 9220 50337 9229 50371
rect 9229 50337 9263 50371
rect 9263 50337 9272 50371
rect 9220 50328 9272 50337
rect 9404 50371 9456 50380
rect 9404 50337 9413 50371
rect 9413 50337 9447 50371
rect 9447 50337 9456 50371
rect 9404 50328 9456 50337
rect 10968 50328 11020 50380
rect 11520 50328 11572 50380
rect 8944 50260 8996 50312
rect 13176 50464 13228 50516
rect 16028 50464 16080 50516
rect 17132 50464 17184 50516
rect 14832 50396 14884 50448
rect 16212 50396 16264 50448
rect 13176 50328 13228 50380
rect 13360 50371 13412 50380
rect 13360 50337 13369 50371
rect 13369 50337 13403 50371
rect 13403 50337 13412 50371
rect 13360 50328 13412 50337
rect 15568 50371 15620 50380
rect 15568 50337 15577 50371
rect 15577 50337 15611 50371
rect 15611 50337 15620 50371
rect 15568 50328 15620 50337
rect 15752 50328 15804 50380
rect 12440 50260 12492 50312
rect 12808 50260 12860 50312
rect 15844 50303 15896 50312
rect 11888 50192 11940 50244
rect 12256 50192 12308 50244
rect 15844 50269 15853 50303
rect 15853 50269 15887 50303
rect 15887 50269 15896 50303
rect 15844 50260 15896 50269
rect 16212 50260 16264 50312
rect 17132 50328 17184 50380
rect 17316 50328 17368 50380
rect 18052 50192 18104 50244
rect 1768 50124 1820 50176
rect 7748 50124 7800 50176
rect 8944 50124 8996 50176
rect 10784 50124 10836 50176
rect 14004 50124 14056 50176
rect 4315 50022 4367 50074
rect 4379 50022 4431 50074
rect 4443 50022 4495 50074
rect 4507 50022 4559 50074
rect 10982 50022 11034 50074
rect 11046 50022 11098 50074
rect 11110 50022 11162 50074
rect 11174 50022 11226 50074
rect 17648 50022 17700 50074
rect 17712 50022 17764 50074
rect 17776 50022 17828 50074
rect 17840 50022 17892 50074
rect 2228 49963 2280 49972
rect 2228 49929 2237 49963
rect 2237 49929 2271 49963
rect 2271 49929 2280 49963
rect 2228 49920 2280 49929
rect 4160 49920 4212 49972
rect 5816 49920 5868 49972
rect 6460 49920 6512 49972
rect 7932 49920 7984 49972
rect 9220 49963 9272 49972
rect 9220 49929 9229 49963
rect 9229 49929 9263 49963
rect 9263 49929 9272 49963
rect 9220 49920 9272 49929
rect 9588 49920 9640 49972
rect 10140 49920 10192 49972
rect 11888 49963 11940 49972
rect 5172 49852 5224 49904
rect 6092 49895 6144 49904
rect 6092 49861 6101 49895
rect 6101 49861 6135 49895
rect 6135 49861 6144 49895
rect 6092 49852 6144 49861
rect 7012 49852 7064 49904
rect 2504 49759 2556 49768
rect 2504 49725 2513 49759
rect 2513 49725 2547 49759
rect 2547 49725 2556 49759
rect 2504 49716 2556 49725
rect 3240 49784 3292 49836
rect 4988 49759 5040 49768
rect 4988 49725 4997 49759
rect 4997 49725 5031 49759
rect 5031 49725 5040 49759
rect 4988 49716 5040 49725
rect 5172 49759 5224 49768
rect 5172 49725 5181 49759
rect 5181 49725 5215 49759
rect 5215 49725 5224 49759
rect 5172 49716 5224 49725
rect 5816 49716 5868 49768
rect 6368 49716 6420 49768
rect 6092 49648 6144 49700
rect 6276 49648 6328 49700
rect 6828 49648 6880 49700
rect 7012 49716 7064 49768
rect 7472 49716 7524 49768
rect 7748 49759 7800 49768
rect 7748 49725 7757 49759
rect 7757 49725 7791 49759
rect 7791 49725 7800 49759
rect 7748 49716 7800 49725
rect 7840 49759 7892 49768
rect 7840 49725 7849 49759
rect 7849 49725 7883 49759
rect 7883 49725 7892 49759
rect 8116 49784 8168 49836
rect 8484 49852 8536 49904
rect 8576 49852 8628 49904
rect 8852 49852 8904 49904
rect 10140 49827 10192 49836
rect 10140 49793 10149 49827
rect 10149 49793 10183 49827
rect 10183 49793 10192 49827
rect 10140 49784 10192 49793
rect 7840 49716 7892 49725
rect 8208 49759 8260 49768
rect 8208 49725 8217 49759
rect 8217 49725 8251 49759
rect 8251 49725 8260 49759
rect 8208 49716 8260 49725
rect 8484 49759 8536 49768
rect 2320 49580 2372 49632
rect 2872 49580 2924 49632
rect 8484 49725 8493 49759
rect 8493 49725 8527 49759
rect 8527 49725 8536 49759
rect 8484 49716 8536 49725
rect 9404 49716 9456 49768
rect 9680 49759 9732 49768
rect 9680 49725 9689 49759
rect 9689 49725 9723 49759
rect 9723 49725 9732 49759
rect 9680 49716 9732 49725
rect 10324 49759 10376 49768
rect 8760 49648 8812 49700
rect 10324 49725 10333 49759
rect 10333 49725 10367 49759
rect 10367 49725 10376 49759
rect 10324 49716 10376 49725
rect 8852 49580 8904 49632
rect 9680 49580 9732 49632
rect 11888 49929 11897 49963
rect 11897 49929 11931 49963
rect 11931 49929 11940 49963
rect 11888 49920 11940 49929
rect 12440 49963 12492 49972
rect 12440 49929 12449 49963
rect 12449 49929 12483 49963
rect 12483 49929 12492 49963
rect 12440 49920 12492 49929
rect 13360 49920 13412 49972
rect 13912 49920 13964 49972
rect 14832 49920 14884 49972
rect 16028 49920 16080 49972
rect 16396 49920 16448 49972
rect 11060 49784 11112 49836
rect 11980 49852 12032 49904
rect 10600 49759 10652 49768
rect 10600 49725 10609 49759
rect 10609 49725 10643 49759
rect 10643 49725 10652 49759
rect 10600 49716 10652 49725
rect 10784 49716 10836 49768
rect 11520 49759 11572 49768
rect 11520 49725 11529 49759
rect 11529 49725 11563 49759
rect 11563 49725 11572 49759
rect 11520 49716 11572 49725
rect 12072 49759 12124 49768
rect 12072 49725 12081 49759
rect 12081 49725 12115 49759
rect 12115 49725 12124 49759
rect 12072 49716 12124 49725
rect 16212 49895 16264 49904
rect 16212 49861 16221 49895
rect 16221 49861 16255 49895
rect 16255 49861 16264 49895
rect 16212 49852 16264 49861
rect 12440 49784 12492 49836
rect 12808 49784 12860 49836
rect 12900 49784 12952 49836
rect 13176 49784 13228 49836
rect 14096 49784 14148 49836
rect 15384 49784 15436 49836
rect 15108 49716 15160 49768
rect 16304 49716 16356 49768
rect 16672 49852 16724 49904
rect 14832 49648 14884 49700
rect 16212 49648 16264 49700
rect 17224 49759 17276 49768
rect 10508 49580 10560 49632
rect 13636 49580 13688 49632
rect 15016 49623 15068 49632
rect 15016 49589 15025 49623
rect 15025 49589 15059 49623
rect 15059 49589 15068 49623
rect 15016 49580 15068 49589
rect 17224 49725 17233 49759
rect 17233 49725 17267 49759
rect 17267 49725 17276 49759
rect 17224 49716 17276 49725
rect 17500 49759 17552 49768
rect 17500 49725 17509 49759
rect 17509 49725 17543 49759
rect 17543 49725 17552 49759
rect 17500 49716 17552 49725
rect 16764 49580 16816 49632
rect 7648 49478 7700 49530
rect 7712 49478 7764 49530
rect 7776 49478 7828 49530
rect 7840 49478 7892 49530
rect 14315 49478 14367 49530
rect 14379 49478 14431 49530
rect 14443 49478 14495 49530
rect 14507 49478 14559 49530
rect 2504 49419 2556 49428
rect 2504 49385 2513 49419
rect 2513 49385 2547 49419
rect 2547 49385 2556 49419
rect 2504 49376 2556 49385
rect 6276 49419 6328 49428
rect 6276 49385 6285 49419
rect 6285 49385 6319 49419
rect 6319 49385 6328 49419
rect 6276 49376 6328 49385
rect 6828 49376 6880 49428
rect 8760 49419 8812 49428
rect 8760 49385 8769 49419
rect 8769 49385 8803 49419
rect 8803 49385 8812 49419
rect 8760 49376 8812 49385
rect 9956 49376 10008 49428
rect 10140 49376 10192 49428
rect 11060 49376 11112 49428
rect 12072 49419 12124 49428
rect 12072 49385 12081 49419
rect 12081 49385 12115 49419
rect 12115 49385 12124 49419
rect 14096 49419 14148 49428
rect 12072 49376 12124 49385
rect 3516 49240 3568 49292
rect 4068 49240 4120 49292
rect 6920 49240 6972 49292
rect 7012 49240 7064 49292
rect 9588 49308 9640 49360
rect 10600 49308 10652 49360
rect 10692 49308 10744 49360
rect 14096 49385 14105 49419
rect 14105 49385 14139 49419
rect 14139 49385 14148 49419
rect 14096 49376 14148 49385
rect 15568 49376 15620 49428
rect 17500 49419 17552 49428
rect 17500 49385 17509 49419
rect 17509 49385 17543 49419
rect 17543 49385 17552 49419
rect 17500 49376 17552 49385
rect 13728 49308 13780 49360
rect 14740 49351 14792 49360
rect 14740 49317 14749 49351
rect 14749 49317 14783 49351
rect 14783 49317 14792 49351
rect 14740 49308 14792 49317
rect 8116 49240 8168 49292
rect 8852 49283 8904 49292
rect 8852 49249 8861 49283
rect 8861 49249 8895 49283
rect 8895 49249 8904 49283
rect 8852 49240 8904 49249
rect 10048 49240 10100 49292
rect 11980 49240 12032 49292
rect 12256 49240 12308 49292
rect 12716 49283 12768 49292
rect 12716 49249 12725 49283
rect 12725 49249 12759 49283
rect 12759 49249 12768 49283
rect 12716 49240 12768 49249
rect 14096 49240 14148 49292
rect 2412 49172 2464 49224
rect 7564 49215 7616 49224
rect 7564 49181 7573 49215
rect 7573 49181 7607 49215
rect 7607 49181 7616 49215
rect 7564 49172 7616 49181
rect 7932 49215 7984 49224
rect 7932 49181 7941 49215
rect 7941 49181 7975 49215
rect 7975 49181 7984 49215
rect 7932 49172 7984 49181
rect 9680 49172 9732 49224
rect 11428 49172 11480 49224
rect 12532 49172 12584 49224
rect 12808 49172 12860 49224
rect 14280 49172 14332 49224
rect 15016 49308 15068 49360
rect 15292 49351 15344 49360
rect 15292 49317 15301 49351
rect 15301 49317 15335 49351
rect 15335 49317 15344 49351
rect 15292 49308 15344 49317
rect 15384 49308 15436 49360
rect 15752 49308 15804 49360
rect 16672 49308 16724 49360
rect 16764 49240 16816 49292
rect 17500 49240 17552 49292
rect 15016 49172 15068 49224
rect 16672 49215 16724 49224
rect 16672 49181 16681 49215
rect 16681 49181 16715 49215
rect 16715 49181 16724 49215
rect 16672 49172 16724 49181
rect 5540 49147 5592 49156
rect 5540 49113 5549 49147
rect 5549 49113 5583 49147
rect 5583 49113 5592 49147
rect 5540 49104 5592 49113
rect 10692 49104 10744 49156
rect 10968 49104 11020 49156
rect 1584 49079 1636 49088
rect 1584 49045 1593 49079
rect 1593 49045 1627 49079
rect 1627 49045 1636 49079
rect 1584 49036 1636 49045
rect 5172 49079 5224 49088
rect 5172 49045 5181 49079
rect 5181 49045 5215 49079
rect 5215 49045 5224 49079
rect 5172 49036 5224 49045
rect 8300 49036 8352 49088
rect 10324 49036 10376 49088
rect 11612 49079 11664 49088
rect 11612 49045 11621 49079
rect 11621 49045 11655 49079
rect 11655 49045 11664 49079
rect 11612 49036 11664 49045
rect 12900 49079 12952 49088
rect 12900 49045 12909 49079
rect 12909 49045 12943 49079
rect 12943 49045 12952 49079
rect 12900 49036 12952 49045
rect 13636 49079 13688 49088
rect 13636 49045 13645 49079
rect 13645 49045 13679 49079
rect 13679 49045 13688 49079
rect 13636 49036 13688 49045
rect 13912 49036 13964 49088
rect 14556 49079 14608 49088
rect 14556 49045 14565 49079
rect 14565 49045 14599 49079
rect 14599 49045 14608 49079
rect 14556 49036 14608 49045
rect 4315 48934 4367 48986
rect 4379 48934 4431 48986
rect 4443 48934 4495 48986
rect 4507 48934 4559 48986
rect 10982 48934 11034 48986
rect 11046 48934 11098 48986
rect 11110 48934 11162 48986
rect 11174 48934 11226 48986
rect 17648 48934 17700 48986
rect 17712 48934 17764 48986
rect 17776 48934 17828 48986
rect 17840 48934 17892 48986
rect 3240 48832 3292 48884
rect 3516 48875 3568 48884
rect 3516 48841 3525 48875
rect 3525 48841 3559 48875
rect 3559 48841 3568 48875
rect 3516 48832 3568 48841
rect 5080 48832 5132 48884
rect 7288 48832 7340 48884
rect 10508 48832 10560 48884
rect 10600 48832 10652 48884
rect 6000 48764 6052 48816
rect 6276 48764 6328 48816
rect 1676 48696 1728 48748
rect 3700 48696 3752 48748
rect 5080 48696 5132 48748
rect 5172 48696 5224 48748
rect 6920 48696 6972 48748
rect 7564 48764 7616 48816
rect 11060 48764 11112 48816
rect 10600 48739 10652 48748
rect 10600 48705 10609 48739
rect 10609 48705 10643 48739
rect 10643 48705 10652 48739
rect 10600 48696 10652 48705
rect 1584 48628 1636 48680
rect 2044 48628 2096 48680
rect 4896 48671 4948 48680
rect 4896 48637 4905 48671
rect 4905 48637 4939 48671
rect 4939 48637 4948 48671
rect 4896 48628 4948 48637
rect 5356 48671 5408 48680
rect 5356 48637 5365 48671
rect 5365 48637 5399 48671
rect 5399 48637 5408 48671
rect 5356 48628 5408 48637
rect 6828 48628 6880 48680
rect 7288 48628 7340 48680
rect 7748 48671 7800 48680
rect 7748 48637 7757 48671
rect 7757 48637 7791 48671
rect 7791 48637 7800 48671
rect 7748 48628 7800 48637
rect 7932 48628 7984 48680
rect 9588 48628 9640 48680
rect 9864 48671 9916 48680
rect 9864 48637 9873 48671
rect 9873 48637 9907 48671
rect 9907 48637 9916 48671
rect 9864 48628 9916 48637
rect 10140 48671 10192 48680
rect 10140 48637 10149 48671
rect 10149 48637 10183 48671
rect 10183 48637 10192 48671
rect 10140 48628 10192 48637
rect 10324 48628 10376 48680
rect 10968 48628 11020 48680
rect 11244 48671 11296 48680
rect 11244 48637 11253 48671
rect 11253 48637 11287 48671
rect 11287 48637 11296 48671
rect 11244 48628 11296 48637
rect 11428 48832 11480 48884
rect 12072 48832 12124 48884
rect 12440 48832 12492 48884
rect 12900 48832 12952 48884
rect 14740 48832 14792 48884
rect 14832 48832 14884 48884
rect 15568 48832 15620 48884
rect 12440 48696 12492 48748
rect 13360 48696 13412 48748
rect 14832 48696 14884 48748
rect 16672 48696 16724 48748
rect 17316 48739 17368 48748
rect 17316 48705 17325 48739
rect 17325 48705 17359 48739
rect 17359 48705 17368 48739
rect 17316 48696 17368 48705
rect 17500 48696 17552 48748
rect 12256 48628 12308 48680
rect 15292 48671 15344 48680
rect 15292 48637 15301 48671
rect 15301 48637 15335 48671
rect 15335 48637 15344 48671
rect 15292 48628 15344 48637
rect 16304 48628 16356 48680
rect 11980 48560 12032 48612
rect 14556 48560 14608 48612
rect 16672 48560 16724 48612
rect 17500 48560 17552 48612
rect 2412 48492 2464 48544
rect 6920 48492 6972 48544
rect 8852 48492 8904 48544
rect 9588 48492 9640 48544
rect 13544 48492 13596 48544
rect 14096 48492 14148 48544
rect 14740 48492 14792 48544
rect 16580 48535 16632 48544
rect 16580 48501 16589 48535
rect 16589 48501 16623 48535
rect 16623 48501 16632 48535
rect 16580 48492 16632 48501
rect 7648 48390 7700 48442
rect 7712 48390 7764 48442
rect 7776 48390 7828 48442
rect 7840 48390 7892 48442
rect 14315 48390 14367 48442
rect 14379 48390 14431 48442
rect 14443 48390 14495 48442
rect 14507 48390 14559 48442
rect 3424 48288 3476 48340
rect 3700 48288 3752 48340
rect 7380 48288 7432 48340
rect 8116 48288 8168 48340
rect 8392 48288 8444 48340
rect 8852 48288 8904 48340
rect 10140 48288 10192 48340
rect 10324 48288 10376 48340
rect 10692 48288 10744 48340
rect 7012 48220 7064 48272
rect 7196 48263 7248 48272
rect 7196 48229 7205 48263
rect 7205 48229 7239 48263
rect 7239 48229 7248 48263
rect 7196 48220 7248 48229
rect 9404 48220 9456 48272
rect 9588 48220 9640 48272
rect 11244 48288 11296 48340
rect 12716 48331 12768 48340
rect 12716 48297 12725 48331
rect 12725 48297 12759 48331
rect 12759 48297 12768 48331
rect 12716 48288 12768 48297
rect 14096 48288 14148 48340
rect 5172 48152 5224 48204
rect 5816 48195 5868 48204
rect 5816 48161 5825 48195
rect 5825 48161 5859 48195
rect 5859 48161 5868 48195
rect 5816 48152 5868 48161
rect 7380 48195 7432 48204
rect 7380 48161 7389 48195
rect 7389 48161 7423 48195
rect 7423 48161 7432 48195
rect 7380 48152 7432 48161
rect 8392 48152 8444 48204
rect 9128 48152 9180 48204
rect 5356 48084 5408 48136
rect 6092 48084 6144 48136
rect 6920 48084 6972 48136
rect 7196 48084 7248 48136
rect 8208 48084 8260 48136
rect 7472 48059 7524 48068
rect 7472 48025 7481 48059
rect 7481 48025 7515 48059
rect 7515 48025 7524 48059
rect 7472 48016 7524 48025
rect 11796 48220 11848 48272
rect 12624 48220 12676 48272
rect 17316 48288 17368 48340
rect 16304 48220 16356 48272
rect 16488 48220 16540 48272
rect 17592 48220 17644 48272
rect 10416 48195 10468 48204
rect 10416 48161 10425 48195
rect 10425 48161 10459 48195
rect 10459 48161 10468 48195
rect 10416 48152 10468 48161
rect 10508 48195 10560 48204
rect 10508 48161 10517 48195
rect 10517 48161 10551 48195
rect 10551 48161 10560 48195
rect 10508 48152 10560 48161
rect 10692 48152 10744 48204
rect 15936 48195 15988 48204
rect 15936 48161 15945 48195
rect 15945 48161 15979 48195
rect 15979 48161 15988 48195
rect 15936 48152 15988 48161
rect 17316 48152 17368 48204
rect 10140 48084 10192 48136
rect 11060 48084 11112 48136
rect 12900 48084 12952 48136
rect 13268 48127 13320 48136
rect 13268 48093 13277 48127
rect 13277 48093 13311 48127
rect 13311 48093 13320 48127
rect 13268 48084 13320 48093
rect 15476 48084 15528 48136
rect 15752 48084 15804 48136
rect 10600 48016 10652 48068
rect 1584 47991 1636 48000
rect 1584 47957 1593 47991
rect 1593 47957 1627 47991
rect 1627 47957 1636 47991
rect 1584 47948 1636 47957
rect 4896 47991 4948 48000
rect 4896 47957 4905 47991
rect 4905 47957 4939 47991
rect 4939 47957 4948 47991
rect 4896 47948 4948 47957
rect 5356 47948 5408 48000
rect 6920 47948 6972 48000
rect 7564 47948 7616 48000
rect 8024 47948 8076 48000
rect 8300 47948 8352 48000
rect 8760 47948 8812 48000
rect 10048 47948 10100 48000
rect 10784 47991 10836 48000
rect 10784 47957 10793 47991
rect 10793 47957 10827 47991
rect 10827 47957 10836 47991
rect 10784 47948 10836 47957
rect 13912 47948 13964 48000
rect 15476 47948 15528 48000
rect 4315 47846 4367 47898
rect 4379 47846 4431 47898
rect 4443 47846 4495 47898
rect 4507 47846 4559 47898
rect 10982 47846 11034 47898
rect 11046 47846 11098 47898
rect 11110 47846 11162 47898
rect 11174 47846 11226 47898
rect 17648 47846 17700 47898
rect 17712 47846 17764 47898
rect 17776 47846 17828 47898
rect 17840 47846 17892 47898
rect 2964 47744 3016 47796
rect 5172 47744 5224 47796
rect 1676 47608 1728 47660
rect 2044 47540 2096 47592
rect 5816 47676 5868 47728
rect 6644 47744 6696 47796
rect 8484 47787 8536 47796
rect 8484 47753 8493 47787
rect 8493 47753 8527 47787
rect 8527 47753 8536 47787
rect 8484 47744 8536 47753
rect 9128 47787 9180 47796
rect 9128 47753 9137 47787
rect 9137 47753 9171 47787
rect 9171 47753 9180 47787
rect 9128 47744 9180 47753
rect 6092 47540 6144 47592
rect 6920 47583 6972 47592
rect 6920 47549 6929 47583
rect 6929 47549 6963 47583
rect 6963 47549 6972 47583
rect 6920 47540 6972 47549
rect 8300 47583 8352 47592
rect 8300 47549 8309 47583
rect 8309 47549 8343 47583
rect 8343 47549 8352 47583
rect 8300 47540 8352 47549
rect 10416 47744 10468 47796
rect 13268 47744 13320 47796
rect 16304 47744 16356 47796
rect 16396 47608 16448 47660
rect 17960 47608 18012 47660
rect 9128 47472 9180 47524
rect 10600 47540 10652 47592
rect 11796 47583 11848 47592
rect 11796 47549 11805 47583
rect 11805 47549 11839 47583
rect 11839 47549 11848 47583
rect 11796 47540 11848 47549
rect 11888 47540 11940 47592
rect 12256 47540 12308 47592
rect 11520 47515 11572 47524
rect 11520 47481 11529 47515
rect 11529 47481 11563 47515
rect 11563 47481 11572 47515
rect 12716 47515 12768 47524
rect 11520 47472 11572 47481
rect 12716 47481 12725 47515
rect 12725 47481 12759 47515
rect 12759 47481 12768 47515
rect 12716 47472 12768 47481
rect 15844 47583 15896 47592
rect 15844 47549 15853 47583
rect 15853 47549 15887 47583
rect 15887 47549 15896 47583
rect 15844 47540 15896 47549
rect 15568 47472 15620 47524
rect 16488 47472 16540 47524
rect 4712 47404 4764 47456
rect 4896 47404 4948 47456
rect 5172 47404 5224 47456
rect 5816 47404 5868 47456
rect 7196 47404 7248 47456
rect 7380 47404 7432 47456
rect 8208 47404 8260 47456
rect 9680 47404 9732 47456
rect 10508 47404 10560 47456
rect 12900 47404 12952 47456
rect 15476 47447 15528 47456
rect 15476 47413 15485 47447
rect 15485 47413 15519 47447
rect 15519 47413 15528 47447
rect 15476 47404 15528 47413
rect 15844 47404 15896 47456
rect 16120 47404 16172 47456
rect 7648 47302 7700 47354
rect 7712 47302 7764 47354
rect 7776 47302 7828 47354
rect 7840 47302 7892 47354
rect 14315 47302 14367 47354
rect 14379 47302 14431 47354
rect 14443 47302 14495 47354
rect 14507 47302 14559 47354
rect 6644 47200 6696 47252
rect 3516 47107 3568 47116
rect 3516 47073 3525 47107
rect 3525 47073 3559 47107
rect 3559 47073 3568 47107
rect 3516 47064 3568 47073
rect 3608 47064 3660 47116
rect 1676 47039 1728 47048
rect 1676 47005 1685 47039
rect 1685 47005 1719 47039
rect 1719 47005 1728 47039
rect 1676 46996 1728 47005
rect 2412 46996 2464 47048
rect 3240 46996 3292 47048
rect 5632 47107 5684 47116
rect 5632 47073 5641 47107
rect 5641 47073 5675 47107
rect 5675 47073 5684 47107
rect 5632 47064 5684 47073
rect 3976 47039 4028 47048
rect 3976 47005 3985 47039
rect 3985 47005 4019 47039
rect 4019 47005 4028 47039
rect 3976 46996 4028 47005
rect 4068 46996 4120 47048
rect 8392 47200 8444 47252
rect 12808 47243 12860 47252
rect 9036 47132 9088 47184
rect 12808 47209 12817 47243
rect 12817 47209 12851 47243
rect 12851 47209 12860 47243
rect 12808 47200 12860 47209
rect 14096 47200 14148 47252
rect 15936 47200 15988 47252
rect 15568 47132 15620 47184
rect 2044 46971 2096 46980
rect 2044 46937 2053 46971
rect 2053 46937 2087 46971
rect 2087 46937 2096 46971
rect 2044 46928 2096 46937
rect 2504 46928 2556 46980
rect 5540 46928 5592 46980
rect 6644 46928 6696 46980
rect 8576 47107 8628 47116
rect 8300 47039 8352 47048
rect 8300 47005 8309 47039
rect 8309 47005 8343 47039
rect 8343 47005 8352 47039
rect 8300 46996 8352 47005
rect 8576 47073 8585 47107
rect 8585 47073 8619 47107
rect 8619 47073 8628 47107
rect 8576 47064 8628 47073
rect 8760 47107 8812 47116
rect 8760 47073 8769 47107
rect 8769 47073 8803 47107
rect 8803 47073 8812 47107
rect 8760 47064 8812 47073
rect 9220 47064 9272 47116
rect 10600 47064 10652 47116
rect 10968 47107 11020 47116
rect 10968 47073 10977 47107
rect 10977 47073 11011 47107
rect 11011 47073 11020 47107
rect 10968 47064 11020 47073
rect 16856 47064 16908 47116
rect 17132 47064 17184 47116
rect 9864 46996 9916 47048
rect 12900 46996 12952 47048
rect 13268 47039 13320 47048
rect 13268 47005 13277 47039
rect 13277 47005 13311 47039
rect 13311 47005 13320 47039
rect 13268 46996 13320 47005
rect 7748 46928 7800 46980
rect 8392 46928 8444 46980
rect 10692 46928 10744 46980
rect 11520 46928 11572 46980
rect 12256 46928 12308 46980
rect 14740 46928 14792 46980
rect 15476 46928 15528 46980
rect 16856 46928 16908 46980
rect 8300 46860 8352 46912
rect 9864 46860 9916 46912
rect 10140 46860 10192 46912
rect 4315 46758 4367 46810
rect 4379 46758 4431 46810
rect 4443 46758 4495 46810
rect 4507 46758 4559 46810
rect 10982 46758 11034 46810
rect 11046 46758 11098 46810
rect 11110 46758 11162 46810
rect 11174 46758 11226 46810
rect 17648 46758 17700 46810
rect 17712 46758 17764 46810
rect 17776 46758 17828 46810
rect 17840 46758 17892 46810
rect 3608 46656 3660 46708
rect 4068 46656 4120 46708
rect 5632 46699 5684 46708
rect 5632 46665 5641 46699
rect 5641 46665 5675 46699
rect 5675 46665 5684 46699
rect 5632 46656 5684 46665
rect 7748 46699 7800 46708
rect 7748 46665 7757 46699
rect 7757 46665 7791 46699
rect 7791 46665 7800 46699
rect 7748 46656 7800 46665
rect 9220 46656 9272 46708
rect 9680 46656 9732 46708
rect 9772 46656 9824 46708
rect 10140 46656 10192 46708
rect 10600 46699 10652 46708
rect 10600 46665 10609 46699
rect 10609 46665 10643 46699
rect 10643 46665 10652 46699
rect 10600 46656 10652 46665
rect 11428 46656 11480 46708
rect 13176 46656 13228 46708
rect 17316 46656 17368 46708
rect 3240 46588 3292 46640
rect 5540 46588 5592 46640
rect 10968 46588 11020 46640
rect 1676 46520 1728 46572
rect 4528 46520 4580 46572
rect 4712 46520 4764 46572
rect 5172 46520 5224 46572
rect 12900 46520 12952 46572
rect 13176 46520 13228 46572
rect 5632 46495 5684 46504
rect 1492 46384 1544 46436
rect 3516 46316 3568 46368
rect 4068 46316 4120 46368
rect 5632 46461 5641 46495
rect 5641 46461 5675 46495
rect 5675 46461 5684 46495
rect 5632 46452 5684 46461
rect 4712 46384 4764 46436
rect 5264 46384 5316 46436
rect 6092 46452 6144 46504
rect 6920 46495 6972 46504
rect 6920 46461 6929 46495
rect 6929 46461 6963 46495
rect 6963 46461 6972 46495
rect 6920 46452 6972 46461
rect 9956 46452 10008 46504
rect 11428 46495 11480 46504
rect 11428 46461 11437 46495
rect 11437 46461 11471 46495
rect 11471 46461 11480 46495
rect 11428 46452 11480 46461
rect 12808 46452 12860 46504
rect 13268 46452 13320 46504
rect 17040 46495 17092 46504
rect 8760 46384 8812 46436
rect 17040 46461 17049 46495
rect 17049 46461 17083 46495
rect 17083 46461 17092 46495
rect 17040 46452 17092 46461
rect 18144 46384 18196 46436
rect 5172 46316 5224 46368
rect 5816 46316 5868 46368
rect 8576 46316 8628 46368
rect 9404 46316 9456 46368
rect 12256 46316 12308 46368
rect 13912 46316 13964 46368
rect 16212 46359 16264 46368
rect 16212 46325 16221 46359
rect 16221 46325 16255 46359
rect 16255 46325 16264 46359
rect 16212 46316 16264 46325
rect 17132 46316 17184 46368
rect 7648 46214 7700 46266
rect 7712 46214 7764 46266
rect 7776 46214 7828 46266
rect 7840 46214 7892 46266
rect 14315 46214 14367 46266
rect 14379 46214 14431 46266
rect 14443 46214 14495 46266
rect 14507 46214 14559 46266
rect 1676 46112 1728 46164
rect 2320 46112 2372 46164
rect 4068 46112 4120 46164
rect 5632 46112 5684 46164
rect 6736 46112 6788 46164
rect 7012 46155 7064 46164
rect 7012 46121 7021 46155
rect 7021 46121 7055 46155
rect 7055 46121 7064 46155
rect 7012 46112 7064 46121
rect 9128 46112 9180 46164
rect 9312 46112 9364 46164
rect 9956 46112 10008 46164
rect 10784 46112 10836 46164
rect 11612 46112 11664 46164
rect 12256 46155 12308 46164
rect 12256 46121 12265 46155
rect 12265 46121 12299 46155
rect 12299 46121 12308 46155
rect 12256 46112 12308 46121
rect 12716 46112 12768 46164
rect 13084 46112 13136 46164
rect 13636 46112 13688 46164
rect 16580 46112 16632 46164
rect 17132 46112 17184 46164
rect 17316 46112 17368 46164
rect 2504 45976 2556 46028
rect 3516 45908 3568 45960
rect 4068 45951 4120 45960
rect 4068 45917 4077 45951
rect 4077 45917 4111 45951
rect 4111 45917 4120 45951
rect 4068 45908 4120 45917
rect 6552 45908 6604 45960
rect 8484 46044 8536 46096
rect 10692 46087 10744 46096
rect 10692 46053 10701 46087
rect 10701 46053 10735 46087
rect 10735 46053 10744 46087
rect 10692 46044 10744 46053
rect 10876 46044 10928 46096
rect 7288 45976 7340 46028
rect 8024 46019 8076 46028
rect 8024 45985 8033 46019
rect 8033 45985 8067 46019
rect 8067 45985 8076 46019
rect 8024 45976 8076 45985
rect 8116 45976 8168 46028
rect 9680 45976 9732 46028
rect 10416 45976 10468 46028
rect 12716 46019 12768 46028
rect 12716 45985 12725 46019
rect 12725 45985 12759 46019
rect 12759 45985 12768 46019
rect 12716 45976 12768 45985
rect 13176 46044 13228 46096
rect 8392 45908 8444 45960
rect 8852 45908 8904 45960
rect 9036 45908 9088 45960
rect 9864 45908 9916 45960
rect 12900 45908 12952 45960
rect 12992 45908 13044 45960
rect 13176 45951 13228 45960
rect 13176 45917 13185 45951
rect 13185 45917 13219 45951
rect 13219 45917 13228 45951
rect 13176 45908 13228 45917
rect 12348 45840 12400 45892
rect 1492 45772 1544 45824
rect 5632 45772 5684 45824
rect 6644 45772 6696 45824
rect 6920 45772 6972 45824
rect 7288 45815 7340 45824
rect 7288 45781 7297 45815
rect 7297 45781 7331 45815
rect 7331 45781 7340 45815
rect 7288 45772 7340 45781
rect 9680 45772 9732 45824
rect 9864 45815 9916 45824
rect 9864 45781 9873 45815
rect 9873 45781 9907 45815
rect 9907 45781 9916 45815
rect 9864 45772 9916 45781
rect 10232 45772 10284 45824
rect 11428 45815 11480 45824
rect 11428 45781 11437 45815
rect 11437 45781 11471 45815
rect 11471 45781 11480 45815
rect 11428 45772 11480 45781
rect 12440 45772 12492 45824
rect 14556 46044 14608 46096
rect 15108 46044 15160 46096
rect 14648 46019 14700 46028
rect 14648 45985 14657 46019
rect 14657 45985 14691 46019
rect 14691 45985 14700 46019
rect 14648 45976 14700 45985
rect 16580 45976 16632 46028
rect 15476 45908 15528 45960
rect 15936 45908 15988 45960
rect 18420 45908 18472 45960
rect 4315 45670 4367 45722
rect 4379 45670 4431 45722
rect 4443 45670 4495 45722
rect 4507 45670 4559 45722
rect 10982 45670 11034 45722
rect 11046 45670 11098 45722
rect 11110 45670 11162 45722
rect 11174 45670 11226 45722
rect 17648 45670 17700 45722
rect 17712 45670 17764 45722
rect 17776 45670 17828 45722
rect 17840 45670 17892 45722
rect 3516 45568 3568 45620
rect 5632 45568 5684 45620
rect 6184 45568 6236 45620
rect 8024 45568 8076 45620
rect 8392 45568 8444 45620
rect 10784 45568 10836 45620
rect 9864 45500 9916 45552
rect 2228 45432 2280 45484
rect 3424 45432 3476 45484
rect 9404 45432 9456 45484
rect 1584 45364 1636 45416
rect 5632 45407 5684 45416
rect 5632 45373 5641 45407
rect 5641 45373 5675 45407
rect 5675 45373 5684 45407
rect 5632 45364 5684 45373
rect 6092 45364 6144 45416
rect 6644 45364 6696 45416
rect 9772 45364 9824 45416
rect 10232 45364 10284 45416
rect 10416 45500 10468 45552
rect 10692 45500 10744 45552
rect 12256 45568 12308 45620
rect 12532 45568 12584 45620
rect 12900 45611 12952 45620
rect 12900 45577 12909 45611
rect 12909 45577 12943 45611
rect 12943 45577 12952 45611
rect 12900 45568 12952 45577
rect 15292 45568 15344 45620
rect 15660 45568 15712 45620
rect 12808 45500 12860 45552
rect 15752 45500 15804 45552
rect 13544 45432 13596 45484
rect 16580 45432 16632 45484
rect 11428 45407 11480 45416
rect 11428 45373 11437 45407
rect 11437 45373 11471 45407
rect 11471 45373 11480 45407
rect 11428 45364 11480 45373
rect 11612 45364 11664 45416
rect 11888 45364 11940 45416
rect 12808 45364 12860 45416
rect 12992 45296 13044 45348
rect 14648 45407 14700 45416
rect 14648 45373 14657 45407
rect 14657 45373 14691 45407
rect 14691 45373 14700 45407
rect 14648 45364 14700 45373
rect 15476 45407 15528 45416
rect 15476 45373 15485 45407
rect 15485 45373 15519 45407
rect 15519 45373 15528 45407
rect 15476 45364 15528 45373
rect 17592 45407 17644 45416
rect 17592 45373 17601 45407
rect 17601 45373 17635 45407
rect 17635 45373 17644 45407
rect 17592 45364 17644 45373
rect 15568 45296 15620 45348
rect 2964 45228 3016 45280
rect 4068 45228 4120 45280
rect 5816 45228 5868 45280
rect 8024 45228 8076 45280
rect 12532 45228 12584 45280
rect 14004 45271 14056 45280
rect 14004 45237 14013 45271
rect 14013 45237 14047 45271
rect 14047 45237 14056 45271
rect 14004 45228 14056 45237
rect 14832 45228 14884 45280
rect 15384 45228 15436 45280
rect 16856 45296 16908 45348
rect 17316 45296 17368 45348
rect 18236 45228 18288 45280
rect 7648 45126 7700 45178
rect 7712 45126 7764 45178
rect 7776 45126 7828 45178
rect 7840 45126 7892 45178
rect 14315 45126 14367 45178
rect 14379 45126 14431 45178
rect 14443 45126 14495 45178
rect 14507 45126 14559 45178
rect 2320 45024 2372 45076
rect 4252 45067 4304 45076
rect 4252 45033 4261 45067
rect 4261 45033 4295 45067
rect 4295 45033 4304 45067
rect 4252 45024 4304 45033
rect 8116 45067 8168 45076
rect 8116 45033 8125 45067
rect 8125 45033 8159 45067
rect 8159 45033 8168 45067
rect 8116 45024 8168 45033
rect 9680 45024 9732 45076
rect 9864 45024 9916 45076
rect 11428 45024 11480 45076
rect 12072 45024 12124 45076
rect 12716 45067 12768 45076
rect 12716 45033 12725 45067
rect 12725 45033 12759 45067
rect 12759 45033 12768 45067
rect 12716 45024 12768 45033
rect 12992 45067 13044 45076
rect 12992 45033 13001 45067
rect 13001 45033 13035 45067
rect 13035 45033 13044 45067
rect 12992 45024 13044 45033
rect 15568 45067 15620 45076
rect 15568 45033 15577 45067
rect 15577 45033 15611 45067
rect 15611 45033 15620 45067
rect 15568 45024 15620 45033
rect 16212 45024 16264 45076
rect 17592 45024 17644 45076
rect 18328 45024 18380 45076
rect 1952 44956 2004 45008
rect 2228 44956 2280 45008
rect 7104 44956 7156 45008
rect 8668 44956 8720 45008
rect 1308 44888 1360 44940
rect 2412 44888 2464 44940
rect 3976 44888 4028 44940
rect 4068 44820 4120 44872
rect 6184 44888 6236 44940
rect 5264 44820 5316 44872
rect 6920 44820 6972 44872
rect 7288 44820 7340 44872
rect 6092 44752 6144 44804
rect 7104 44752 7156 44804
rect 8300 44888 8352 44940
rect 12900 44956 12952 45008
rect 14832 44956 14884 45008
rect 15936 44956 15988 45008
rect 9772 44888 9824 44940
rect 10876 44931 10928 44940
rect 9588 44820 9640 44872
rect 10876 44897 10885 44931
rect 10885 44897 10919 44931
rect 10919 44897 10928 44931
rect 10876 44888 10928 44897
rect 11612 44888 11664 44940
rect 12164 44888 12216 44940
rect 13544 44888 13596 44940
rect 15752 44931 15804 44940
rect 15752 44897 15761 44931
rect 15761 44897 15795 44931
rect 15795 44897 15804 44931
rect 15752 44888 15804 44897
rect 16672 44931 16724 44940
rect 16672 44897 16681 44931
rect 16681 44897 16715 44931
rect 16715 44897 16724 44931
rect 16672 44888 16724 44897
rect 12440 44820 12492 44872
rect 12532 44820 12584 44872
rect 12900 44820 12952 44872
rect 9220 44752 9272 44804
rect 10968 44752 11020 44804
rect 11520 44752 11572 44804
rect 1584 44727 1636 44736
rect 1584 44693 1593 44727
rect 1593 44693 1627 44727
rect 1627 44693 1636 44727
rect 1584 44684 1636 44693
rect 6276 44684 6328 44736
rect 11796 44727 11848 44736
rect 11796 44693 11805 44727
rect 11805 44693 11839 44727
rect 11839 44693 11848 44727
rect 11796 44684 11848 44693
rect 14556 44727 14608 44736
rect 14556 44693 14565 44727
rect 14565 44693 14599 44727
rect 14599 44693 14608 44727
rect 14556 44684 14608 44693
rect 15844 44684 15896 44736
rect 4315 44582 4367 44634
rect 4379 44582 4431 44634
rect 4443 44582 4495 44634
rect 4507 44582 4559 44634
rect 10982 44582 11034 44634
rect 11046 44582 11098 44634
rect 11110 44582 11162 44634
rect 11174 44582 11226 44634
rect 17648 44582 17700 44634
rect 17712 44582 17764 44634
rect 17776 44582 17828 44634
rect 17840 44582 17892 44634
rect 1676 44523 1728 44532
rect 1676 44489 1685 44523
rect 1685 44489 1719 44523
rect 1719 44489 1728 44523
rect 1676 44480 1728 44489
rect 2320 44480 2372 44532
rect 3976 44480 4028 44532
rect 7196 44523 7248 44532
rect 7196 44489 7205 44523
rect 7205 44489 7239 44523
rect 7239 44489 7248 44523
rect 7196 44480 7248 44489
rect 8116 44480 8168 44532
rect 9036 44480 9088 44532
rect 4068 44412 4120 44464
rect 4252 44412 4304 44464
rect 6000 44412 6052 44464
rect 7380 44455 7432 44464
rect 7380 44421 7389 44455
rect 7389 44421 7423 44455
rect 7423 44421 7432 44455
rect 7380 44412 7432 44421
rect 9220 44412 9272 44464
rect 3976 44276 4028 44328
rect 5264 44276 5316 44328
rect 5632 44276 5684 44328
rect 6276 44319 6328 44328
rect 6276 44285 6285 44319
rect 6285 44285 6319 44319
rect 6319 44285 6328 44319
rect 6276 44276 6328 44285
rect 8024 44344 8076 44396
rect 8300 44344 8352 44396
rect 8116 44319 8168 44328
rect 6000 44208 6052 44260
rect 6552 44208 6604 44260
rect 7012 44208 7064 44260
rect 8116 44285 8125 44319
rect 8125 44285 8159 44319
rect 8159 44285 8168 44319
rect 8116 44276 8168 44285
rect 11612 44480 11664 44532
rect 13544 44480 13596 44532
rect 11520 44455 11572 44464
rect 11520 44421 11529 44455
rect 11529 44421 11563 44455
rect 11563 44421 11572 44455
rect 11520 44412 11572 44421
rect 12440 44412 12492 44464
rect 14096 44412 14148 44464
rect 9680 44344 9732 44396
rect 10232 44319 10284 44328
rect 10232 44285 10241 44319
rect 10241 44285 10275 44319
rect 10275 44285 10284 44319
rect 10232 44276 10284 44285
rect 8024 44208 8076 44260
rect 9772 44208 9824 44260
rect 9864 44208 9916 44260
rect 10876 44276 10928 44328
rect 12716 44387 12768 44396
rect 12716 44353 12725 44387
rect 12725 44353 12759 44387
rect 12759 44353 12768 44387
rect 12716 44344 12768 44353
rect 12348 44276 12400 44328
rect 12532 44276 12584 44328
rect 13728 44276 13780 44328
rect 12716 44208 12768 44260
rect 13360 44208 13412 44260
rect 13820 44208 13872 44260
rect 14096 44276 14148 44328
rect 14924 44480 14976 44532
rect 14924 44344 14976 44396
rect 16948 44480 17000 44532
rect 16672 44412 16724 44464
rect 15752 44276 15804 44328
rect 15384 44208 15436 44260
rect 16396 44208 16448 44260
rect 17316 44276 17368 44328
rect 17592 44319 17644 44328
rect 17592 44285 17601 44319
rect 17601 44285 17635 44319
rect 17635 44285 17644 44319
rect 17592 44276 17644 44285
rect 14740 44140 14792 44192
rect 15660 44140 15712 44192
rect 16580 44140 16632 44192
rect 7648 44038 7700 44090
rect 7712 44038 7764 44090
rect 7776 44038 7828 44090
rect 7840 44038 7892 44090
rect 14315 44038 14367 44090
rect 14379 44038 14431 44090
rect 14443 44038 14495 44090
rect 14507 44038 14559 44090
rect 7104 43936 7156 43988
rect 8300 43979 8352 43988
rect 8300 43945 8309 43979
rect 8309 43945 8343 43979
rect 8343 43945 8352 43979
rect 8300 43936 8352 43945
rect 3240 43868 3292 43920
rect 4160 43911 4212 43920
rect 4160 43877 4169 43911
rect 4169 43877 4203 43911
rect 4203 43877 4212 43911
rect 4160 43868 4212 43877
rect 4988 43868 5040 43920
rect 3976 43800 4028 43852
rect 6920 43843 6972 43852
rect 6920 43809 6929 43843
rect 6929 43809 6963 43843
rect 6963 43809 6972 43843
rect 6920 43800 6972 43809
rect 7104 43800 7156 43852
rect 7472 43800 7524 43852
rect 8300 43800 8352 43852
rect 10324 43936 10376 43988
rect 11888 43936 11940 43988
rect 12440 43936 12492 43988
rect 12716 43936 12768 43988
rect 13268 43936 13320 43988
rect 15568 43979 15620 43988
rect 15568 43945 15577 43979
rect 15577 43945 15611 43979
rect 15611 43945 15620 43979
rect 15568 43936 15620 43945
rect 14188 43868 14240 43920
rect 14372 43868 14424 43920
rect 17592 43868 17644 43920
rect 9680 43800 9732 43852
rect 10324 43843 10376 43852
rect 10324 43809 10333 43843
rect 10333 43809 10367 43843
rect 10367 43809 10376 43843
rect 10324 43800 10376 43809
rect 11520 43800 11572 43852
rect 13084 43800 13136 43852
rect 13544 43800 13596 43852
rect 14280 43800 14332 43852
rect 15752 43843 15804 43852
rect 15752 43809 15761 43843
rect 15761 43809 15795 43843
rect 15795 43809 15804 43843
rect 15752 43800 15804 43809
rect 16028 43843 16080 43852
rect 16028 43809 16037 43843
rect 16037 43809 16071 43843
rect 16071 43809 16080 43843
rect 16028 43800 16080 43809
rect 16396 43843 16448 43852
rect 16396 43809 16405 43843
rect 16405 43809 16439 43843
rect 16439 43809 16448 43843
rect 16396 43800 16448 43809
rect 16948 43843 17000 43852
rect 16948 43809 16957 43843
rect 16957 43809 16991 43843
rect 16991 43809 17000 43843
rect 16948 43800 17000 43809
rect 1676 43732 1728 43784
rect 1952 43732 2004 43784
rect 4068 43775 4120 43784
rect 4068 43741 4077 43775
rect 4077 43741 4111 43775
rect 4111 43741 4120 43775
rect 4068 43732 4120 43741
rect 4988 43775 5040 43784
rect 4988 43741 4997 43775
rect 4997 43741 5031 43775
rect 5031 43741 5040 43775
rect 4988 43732 5040 43741
rect 9864 43732 9916 43784
rect 10416 43775 10468 43784
rect 10416 43741 10425 43775
rect 10425 43741 10459 43775
rect 10459 43741 10468 43775
rect 10416 43732 10468 43741
rect 12532 43732 12584 43784
rect 12900 43732 12952 43784
rect 16120 43775 16172 43784
rect 16120 43741 16129 43775
rect 16129 43741 16163 43775
rect 16163 43741 16172 43775
rect 16120 43732 16172 43741
rect 6644 43664 6696 43716
rect 6920 43664 6972 43716
rect 3516 43639 3568 43648
rect 3516 43605 3525 43639
rect 3525 43605 3559 43639
rect 3559 43605 3568 43639
rect 3516 43596 3568 43605
rect 6460 43596 6512 43648
rect 6828 43596 6880 43648
rect 8668 43596 8720 43648
rect 12716 43596 12768 43648
rect 14832 43596 14884 43648
rect 15016 43596 15068 43648
rect 15936 43596 15988 43648
rect 4315 43494 4367 43546
rect 4379 43494 4431 43546
rect 4443 43494 4495 43546
rect 4507 43494 4559 43546
rect 10982 43494 11034 43546
rect 11046 43494 11098 43546
rect 11110 43494 11162 43546
rect 11174 43494 11226 43546
rect 17648 43494 17700 43546
rect 17712 43494 17764 43546
rect 17776 43494 17828 43546
rect 17840 43494 17892 43546
rect 3700 43392 3752 43444
rect 3976 43392 4028 43444
rect 4068 43392 4120 43444
rect 7012 43392 7064 43444
rect 7472 43392 7524 43444
rect 8300 43435 8352 43444
rect 8300 43401 8309 43435
rect 8309 43401 8343 43435
rect 8343 43401 8352 43435
rect 8300 43392 8352 43401
rect 8484 43392 8536 43444
rect 4896 43324 4948 43376
rect 5540 43324 5592 43376
rect 1676 43256 1728 43308
rect 3608 43256 3660 43308
rect 1584 43188 1636 43240
rect 3700 43188 3752 43240
rect 4896 43188 4948 43240
rect 6184 43324 6236 43376
rect 7288 43324 7340 43376
rect 6276 43299 6328 43308
rect 6276 43265 6285 43299
rect 6285 43265 6319 43299
rect 6319 43265 6328 43299
rect 6276 43256 6328 43265
rect 9864 43299 9916 43308
rect 9864 43265 9873 43299
rect 9873 43265 9907 43299
rect 9907 43265 9916 43299
rect 9864 43256 9916 43265
rect 5816 43052 5868 43104
rect 6092 43188 6144 43240
rect 6644 43188 6696 43240
rect 7196 43188 7248 43240
rect 8576 43231 8628 43240
rect 8576 43197 8585 43231
rect 8585 43197 8619 43231
rect 8619 43197 8628 43231
rect 8576 43188 8628 43197
rect 10324 43188 10376 43240
rect 10784 43392 10836 43444
rect 11520 43435 11572 43444
rect 11520 43401 11529 43435
rect 11529 43401 11563 43435
rect 11563 43401 11572 43435
rect 11520 43392 11572 43401
rect 12624 43392 12676 43444
rect 13544 43435 13596 43444
rect 13544 43401 13553 43435
rect 13553 43401 13587 43435
rect 13587 43401 13596 43435
rect 13544 43392 13596 43401
rect 13820 43392 13872 43444
rect 16028 43392 16080 43444
rect 14280 43324 14332 43376
rect 13728 43256 13780 43308
rect 14188 43256 14240 43308
rect 16948 43256 17000 43308
rect 10784 43120 10836 43172
rect 13820 43188 13872 43240
rect 15936 43188 15988 43240
rect 16672 43231 16724 43240
rect 16672 43197 16681 43231
rect 16681 43197 16715 43231
rect 16715 43197 16724 43231
rect 16672 43188 16724 43197
rect 18420 43256 18472 43308
rect 12072 43052 12124 43104
rect 12624 43120 12676 43172
rect 14372 43120 14424 43172
rect 14832 43120 14884 43172
rect 13084 43052 13136 43104
rect 13544 43052 13596 43104
rect 14924 43052 14976 43104
rect 15384 43052 15436 43104
rect 17316 43052 17368 43104
rect 18052 43052 18104 43104
rect 7648 42950 7700 43002
rect 7712 42950 7764 43002
rect 7776 42950 7828 43002
rect 7840 42950 7892 43002
rect 14315 42950 14367 43002
rect 14379 42950 14431 43002
rect 14443 42950 14495 43002
rect 14507 42950 14559 43002
rect 1676 42848 1728 42900
rect 3792 42848 3844 42900
rect 4068 42848 4120 42900
rect 4988 42891 5040 42900
rect 4988 42857 4997 42891
rect 4997 42857 5031 42891
rect 5031 42857 5040 42891
rect 4988 42848 5040 42857
rect 6184 42848 6236 42900
rect 8392 42848 8444 42900
rect 8576 42848 8628 42900
rect 10232 42848 10284 42900
rect 12440 42848 12492 42900
rect 12716 42848 12768 42900
rect 15108 42848 15160 42900
rect 16672 42891 16724 42900
rect 7196 42780 7248 42832
rect 7932 42780 7984 42832
rect 8116 42780 8168 42832
rect 3516 42712 3568 42764
rect 4896 42712 4948 42764
rect 8392 42755 8444 42764
rect 1952 42687 2004 42696
rect 1952 42653 1961 42687
rect 1961 42653 1995 42687
rect 1995 42653 2004 42687
rect 1952 42644 2004 42653
rect 3424 42687 3476 42696
rect 3424 42653 3433 42687
rect 3433 42653 3467 42687
rect 3467 42653 3476 42687
rect 3424 42644 3476 42653
rect 8392 42721 8401 42755
rect 8401 42721 8435 42755
rect 8435 42721 8444 42755
rect 8392 42712 8444 42721
rect 8484 42712 8536 42764
rect 9588 42712 9640 42764
rect 8300 42644 8352 42696
rect 9772 42644 9824 42696
rect 6092 42576 6144 42628
rect 8668 42576 8720 42628
rect 10784 42780 10836 42832
rect 11520 42823 11572 42832
rect 11520 42789 11529 42823
rect 11529 42789 11563 42823
rect 11563 42789 11572 42823
rect 11520 42780 11572 42789
rect 13268 42780 13320 42832
rect 10232 42755 10284 42764
rect 10232 42721 10241 42755
rect 10241 42721 10275 42755
rect 10275 42721 10284 42755
rect 10232 42712 10284 42721
rect 10692 42712 10744 42764
rect 13544 42755 13596 42764
rect 13544 42721 13553 42755
rect 13553 42721 13587 42755
rect 13587 42721 13596 42755
rect 13544 42712 13596 42721
rect 13820 42755 13872 42764
rect 13820 42721 13829 42755
rect 13829 42721 13863 42755
rect 13863 42721 13872 42755
rect 13820 42712 13872 42721
rect 15568 42780 15620 42832
rect 13084 42644 13136 42696
rect 14188 42644 14240 42696
rect 10508 42619 10560 42628
rect 1492 42508 1544 42560
rect 7012 42551 7064 42560
rect 7012 42517 7021 42551
rect 7021 42517 7055 42551
rect 7055 42517 7064 42551
rect 7012 42508 7064 42517
rect 7748 42551 7800 42560
rect 7748 42517 7757 42551
rect 7757 42517 7791 42551
rect 7791 42517 7800 42551
rect 7748 42508 7800 42517
rect 8116 42508 8168 42560
rect 10508 42585 10517 42619
rect 10517 42585 10551 42619
rect 10551 42585 10560 42619
rect 10508 42576 10560 42585
rect 10784 42619 10836 42628
rect 10784 42585 10793 42619
rect 10793 42585 10827 42619
rect 10827 42585 10836 42619
rect 10784 42576 10836 42585
rect 14924 42576 14976 42628
rect 15936 42755 15988 42764
rect 15936 42721 15945 42755
rect 15945 42721 15979 42755
rect 15979 42721 15988 42755
rect 15936 42712 15988 42721
rect 16672 42857 16681 42891
rect 16681 42857 16715 42891
rect 16715 42857 16724 42891
rect 16672 42848 16724 42857
rect 15292 42644 15344 42696
rect 15568 42576 15620 42628
rect 16672 42576 16724 42628
rect 9404 42508 9456 42560
rect 9772 42508 9824 42560
rect 10692 42551 10744 42560
rect 10692 42517 10701 42551
rect 10701 42517 10735 42551
rect 10735 42517 10744 42551
rect 10692 42508 10744 42517
rect 13176 42508 13228 42560
rect 14832 42508 14884 42560
rect 15936 42508 15988 42560
rect 16028 42508 16080 42560
rect 16396 42508 16448 42560
rect 4315 42406 4367 42458
rect 4379 42406 4431 42458
rect 4443 42406 4495 42458
rect 4507 42406 4559 42458
rect 10982 42406 11034 42458
rect 11046 42406 11098 42458
rect 11110 42406 11162 42458
rect 11174 42406 11226 42458
rect 17648 42406 17700 42458
rect 17712 42406 17764 42458
rect 17776 42406 17828 42458
rect 17840 42406 17892 42458
rect 2872 42347 2924 42356
rect 2872 42313 2881 42347
rect 2881 42313 2915 42347
rect 2915 42313 2924 42347
rect 2872 42304 2924 42313
rect 3516 42347 3568 42356
rect 3516 42313 3525 42347
rect 3525 42313 3559 42347
rect 3559 42313 3568 42347
rect 3516 42304 3568 42313
rect 4160 42304 4212 42356
rect 1676 42168 1728 42220
rect 6000 42304 6052 42356
rect 8392 42304 8444 42356
rect 8944 42304 8996 42356
rect 9404 42304 9456 42356
rect 4896 42236 4948 42288
rect 7564 42279 7616 42288
rect 7564 42245 7573 42279
rect 7573 42245 7607 42279
rect 7607 42245 7616 42279
rect 7564 42236 7616 42245
rect 7748 42211 7800 42220
rect 1584 42100 1636 42152
rect 5172 42143 5224 42152
rect 5172 42109 5181 42143
rect 5181 42109 5215 42143
rect 5215 42109 5224 42143
rect 5172 42100 5224 42109
rect 7748 42177 7757 42211
rect 7757 42177 7791 42211
rect 7791 42177 7800 42211
rect 7748 42168 7800 42177
rect 9588 42304 9640 42356
rect 10232 42347 10284 42356
rect 10232 42313 10241 42347
rect 10241 42313 10275 42347
rect 10275 42313 10284 42347
rect 10232 42304 10284 42313
rect 10692 42304 10744 42356
rect 11428 42304 11480 42356
rect 13084 42347 13136 42356
rect 13084 42313 13093 42347
rect 13093 42313 13127 42347
rect 13127 42313 13136 42347
rect 13084 42304 13136 42313
rect 14004 42304 14056 42356
rect 14188 42304 14240 42356
rect 14832 42304 14884 42356
rect 15292 42304 15344 42356
rect 15568 42347 15620 42356
rect 15568 42313 15577 42347
rect 15577 42313 15611 42347
rect 15611 42313 15620 42347
rect 15568 42304 15620 42313
rect 6000 42100 6052 42152
rect 6276 42100 6328 42152
rect 7472 42032 7524 42084
rect 7932 42032 7984 42084
rect 8944 42100 8996 42152
rect 9864 42168 9916 42220
rect 10232 42100 10284 42152
rect 13544 42236 13596 42288
rect 15936 42236 15988 42288
rect 17776 42236 17828 42288
rect 18328 42236 18380 42288
rect 12164 42168 12216 42220
rect 12992 42168 13044 42220
rect 13268 42168 13320 42220
rect 10692 42143 10744 42152
rect 10692 42109 10701 42143
rect 10701 42109 10735 42143
rect 10735 42109 10744 42143
rect 10692 42100 10744 42109
rect 4252 41964 4304 42016
rect 5264 41964 5316 42016
rect 9036 42032 9088 42084
rect 11612 42100 11664 42152
rect 11980 42100 12032 42152
rect 13544 42100 13596 42152
rect 13820 42100 13872 42152
rect 15844 42143 15896 42152
rect 15844 42109 15853 42143
rect 15853 42109 15887 42143
rect 15887 42109 15896 42143
rect 15844 42100 15896 42109
rect 16396 42100 16448 42152
rect 17316 42168 17368 42220
rect 17960 42168 18012 42220
rect 15108 42032 15160 42084
rect 15752 42032 15804 42084
rect 16948 42100 17000 42152
rect 9496 41964 9548 42016
rect 12532 42007 12584 42016
rect 12532 41973 12541 42007
rect 12541 41973 12575 42007
rect 12575 41973 12584 42007
rect 12532 41964 12584 41973
rect 7648 41862 7700 41914
rect 7712 41862 7764 41914
rect 7776 41862 7828 41914
rect 7840 41862 7892 41914
rect 14315 41862 14367 41914
rect 14379 41862 14431 41914
rect 14443 41862 14495 41914
rect 14507 41862 14559 41914
rect 1676 41760 1728 41812
rect 3424 41803 3476 41812
rect 3424 41769 3433 41803
rect 3433 41769 3467 41803
rect 3467 41769 3476 41803
rect 3424 41760 3476 41769
rect 5172 41760 5224 41812
rect 4160 41692 4212 41744
rect 4988 41692 5040 41744
rect 6184 41760 6236 41812
rect 7196 41760 7248 41812
rect 8300 41803 8352 41812
rect 8300 41769 8309 41803
rect 8309 41769 8343 41803
rect 8343 41769 8352 41803
rect 8300 41760 8352 41769
rect 8484 41760 8536 41812
rect 10324 41803 10376 41812
rect 10324 41769 10333 41803
rect 10333 41769 10367 41803
rect 10367 41769 10376 41803
rect 10324 41760 10376 41769
rect 10784 41760 10836 41812
rect 13820 41760 13872 41812
rect 5724 41692 5776 41744
rect 7012 41692 7064 41744
rect 5264 41624 5316 41676
rect 6000 41624 6052 41676
rect 7104 41624 7156 41676
rect 8116 41624 8168 41676
rect 9220 41624 9272 41676
rect 9496 41667 9548 41676
rect 9496 41633 9505 41667
rect 9505 41633 9539 41667
rect 9539 41633 9548 41667
rect 9496 41624 9548 41633
rect 9680 41624 9732 41676
rect 14740 41692 14792 41744
rect 11520 41667 11572 41676
rect 11520 41633 11529 41667
rect 11529 41633 11563 41667
rect 11563 41633 11572 41667
rect 11520 41624 11572 41633
rect 11980 41624 12032 41676
rect 12992 41667 13044 41676
rect 12992 41633 13001 41667
rect 13001 41633 13035 41667
rect 13035 41633 13044 41667
rect 12992 41624 13044 41633
rect 13728 41624 13780 41676
rect 15568 41760 15620 41812
rect 15844 41760 15896 41812
rect 16948 41803 17000 41812
rect 16948 41769 16957 41803
rect 16957 41769 16991 41803
rect 16991 41769 17000 41803
rect 16948 41760 17000 41769
rect 15752 41692 15804 41744
rect 15384 41624 15436 41676
rect 15936 41667 15988 41676
rect 15936 41633 15945 41667
rect 15945 41633 15979 41667
rect 15979 41633 15988 41667
rect 15936 41624 15988 41633
rect 16396 41624 16448 41676
rect 16764 41624 16816 41676
rect 6184 41556 6236 41608
rect 8944 41556 8996 41608
rect 9036 41556 9088 41608
rect 12164 41556 12216 41608
rect 12532 41599 12584 41608
rect 12532 41565 12541 41599
rect 12541 41565 12575 41599
rect 12575 41565 12584 41599
rect 12532 41556 12584 41565
rect 13176 41556 13228 41608
rect 15752 41599 15804 41608
rect 15752 41565 15761 41599
rect 15761 41565 15795 41599
rect 15795 41565 15804 41599
rect 15752 41556 15804 41565
rect 5632 41488 5684 41540
rect 6000 41488 6052 41540
rect 15936 41488 15988 41540
rect 17500 41488 17552 41540
rect 18328 41488 18380 41540
rect 1584 41463 1636 41472
rect 1584 41429 1593 41463
rect 1593 41429 1627 41463
rect 1627 41429 1636 41463
rect 1584 41420 1636 41429
rect 6828 41420 6880 41472
rect 8484 41420 8536 41472
rect 12716 41420 12768 41472
rect 13544 41420 13596 41472
rect 14004 41463 14056 41472
rect 14004 41429 14013 41463
rect 14013 41429 14047 41463
rect 14047 41429 14056 41463
rect 14004 41420 14056 41429
rect 4315 41318 4367 41370
rect 4379 41318 4431 41370
rect 4443 41318 4495 41370
rect 4507 41318 4559 41370
rect 10982 41318 11034 41370
rect 11046 41318 11098 41370
rect 11110 41318 11162 41370
rect 11174 41318 11226 41370
rect 17648 41318 17700 41370
rect 17712 41318 17764 41370
rect 17776 41318 17828 41370
rect 17840 41318 17892 41370
rect 1768 41216 1820 41268
rect 2504 41216 2556 41268
rect 3240 41216 3292 41268
rect 6184 41259 6236 41268
rect 1676 41080 1728 41132
rect 6184 41225 6193 41259
rect 6193 41225 6227 41259
rect 6227 41225 6236 41259
rect 6184 41216 6236 41225
rect 7012 41216 7064 41268
rect 9220 41216 9272 41268
rect 5540 41191 5592 41200
rect 5540 41157 5549 41191
rect 5549 41157 5583 41191
rect 5583 41157 5592 41191
rect 5540 41148 5592 41157
rect 1584 41012 1636 41064
rect 4620 41012 4672 41064
rect 5080 41055 5132 41064
rect 5080 41021 5089 41055
rect 5089 41021 5123 41055
rect 5123 41021 5132 41055
rect 5080 41012 5132 41021
rect 5632 41055 5684 41064
rect 5632 41021 5641 41055
rect 5641 41021 5675 41055
rect 5675 41021 5684 41055
rect 5632 41012 5684 41021
rect 6184 41012 6236 41064
rect 6828 41148 6880 41200
rect 7472 41191 7524 41200
rect 7472 41157 7481 41191
rect 7481 41157 7515 41191
rect 7515 41157 7524 41191
rect 7472 41148 7524 41157
rect 8576 41148 8628 41200
rect 8944 41148 8996 41200
rect 9220 41080 9272 41132
rect 6920 41012 6972 41064
rect 8300 41012 8352 41064
rect 8760 41012 8812 41064
rect 8944 41012 8996 41064
rect 9680 41148 9732 41200
rect 10232 41080 10284 41132
rect 7012 40876 7064 40928
rect 8116 40919 8168 40928
rect 8116 40885 8125 40919
rect 8125 40885 8159 40919
rect 8159 40885 8168 40919
rect 8116 40876 8168 40885
rect 8576 40876 8628 40928
rect 10324 41012 10376 41064
rect 11428 41080 11480 41132
rect 11888 41216 11940 41268
rect 12256 41216 12308 41268
rect 15384 41216 15436 41268
rect 16396 41216 16448 41268
rect 16948 41216 17000 41268
rect 17960 41259 18012 41268
rect 17960 41225 17969 41259
rect 17969 41225 18003 41259
rect 18003 41225 18012 41259
rect 17960 41216 18012 41225
rect 11612 41080 11664 41132
rect 14004 41148 14056 41200
rect 15660 41148 15712 41200
rect 16856 41148 16908 41200
rect 17408 41148 17460 41200
rect 18328 41148 18380 41200
rect 11980 41080 12032 41132
rect 12624 41123 12676 41132
rect 12624 41089 12633 41123
rect 12633 41089 12667 41123
rect 12667 41089 12676 41123
rect 12624 41080 12676 41089
rect 13820 41123 13872 41132
rect 13820 41089 13829 41123
rect 13829 41089 13863 41123
rect 13863 41089 13872 41123
rect 13820 41080 13872 41089
rect 14556 41080 14608 41132
rect 15476 41080 15528 41132
rect 12164 41055 12216 41064
rect 9864 40944 9916 40996
rect 10876 40944 10928 40996
rect 12164 41021 12173 41055
rect 12173 41021 12207 41055
rect 12207 41021 12216 41055
rect 12164 41012 12216 41021
rect 11980 40944 12032 40996
rect 12716 41012 12768 41064
rect 12992 41055 13044 41064
rect 12992 41021 13001 41055
rect 13001 41021 13035 41055
rect 13035 41021 13044 41055
rect 12992 41012 13044 41021
rect 12624 40944 12676 40996
rect 14740 41012 14792 41064
rect 15936 41012 15988 41064
rect 16396 41080 16448 41132
rect 16304 40944 16356 40996
rect 10324 40876 10376 40928
rect 14832 40876 14884 40928
rect 15016 40919 15068 40928
rect 15016 40885 15025 40919
rect 15025 40885 15059 40919
rect 15059 40885 15068 40919
rect 15016 40876 15068 40885
rect 15476 40919 15528 40928
rect 15476 40885 15485 40919
rect 15485 40885 15519 40919
rect 15519 40885 15528 40919
rect 15476 40876 15528 40885
rect 15660 40876 15712 40928
rect 16672 41012 16724 41064
rect 17592 41012 17644 41064
rect 17316 40876 17368 40928
rect 7648 40774 7700 40826
rect 7712 40774 7764 40826
rect 7776 40774 7828 40826
rect 7840 40774 7892 40826
rect 14315 40774 14367 40826
rect 14379 40774 14431 40826
rect 14443 40774 14495 40826
rect 14507 40774 14559 40826
rect 4988 40672 5040 40724
rect 6184 40672 6236 40724
rect 6920 40672 6972 40724
rect 7472 40672 7524 40724
rect 9128 40672 9180 40724
rect 5264 40604 5316 40656
rect 8116 40604 8168 40656
rect 4252 40536 4304 40588
rect 7472 40536 7524 40588
rect 9036 40579 9088 40588
rect 5264 40468 5316 40520
rect 5632 40400 5684 40452
rect 6920 40400 6972 40452
rect 9036 40545 9045 40579
rect 9045 40545 9079 40579
rect 9079 40545 9088 40579
rect 9036 40536 9088 40545
rect 11704 40672 11756 40724
rect 16764 40715 16816 40724
rect 16764 40681 16773 40715
rect 16773 40681 16807 40715
rect 16807 40681 16816 40715
rect 16764 40672 16816 40681
rect 17592 40672 17644 40724
rect 8852 40511 8904 40520
rect 8852 40477 8861 40511
rect 8861 40477 8895 40511
rect 8895 40477 8904 40511
rect 8852 40468 8904 40477
rect 9588 40536 9640 40588
rect 10324 40536 10376 40588
rect 10784 40579 10836 40588
rect 10784 40545 10793 40579
rect 10793 40545 10827 40579
rect 10827 40545 10836 40579
rect 10784 40536 10836 40545
rect 10876 40579 10928 40588
rect 10876 40545 10885 40579
rect 10885 40545 10919 40579
rect 10919 40545 10928 40579
rect 10876 40536 10928 40545
rect 12164 40536 12216 40588
rect 12440 40536 12492 40588
rect 13084 40579 13136 40588
rect 13084 40545 13093 40579
rect 13093 40545 13127 40579
rect 13127 40545 13136 40579
rect 13084 40536 13136 40545
rect 13820 40536 13872 40588
rect 15200 40604 15252 40656
rect 13636 40468 13688 40520
rect 9036 40400 9088 40452
rect 9220 40400 9272 40452
rect 13820 40400 13872 40452
rect 14648 40536 14700 40588
rect 14924 40536 14976 40588
rect 15844 40579 15896 40588
rect 15844 40545 15853 40579
rect 15853 40545 15887 40579
rect 15887 40545 15896 40579
rect 15844 40536 15896 40545
rect 18144 40536 18196 40588
rect 14648 40400 14700 40452
rect 15476 40400 15528 40452
rect 16856 40400 16908 40452
rect 1584 40375 1636 40384
rect 1584 40341 1593 40375
rect 1593 40341 1627 40375
rect 1627 40341 1636 40375
rect 1584 40332 1636 40341
rect 1676 40332 1728 40384
rect 8300 40332 8352 40384
rect 9864 40332 9916 40384
rect 12624 40332 12676 40384
rect 16304 40332 16356 40384
rect 17316 40375 17368 40384
rect 17316 40341 17325 40375
rect 17325 40341 17359 40375
rect 17359 40341 17368 40375
rect 17316 40332 17368 40341
rect 4315 40230 4367 40282
rect 4379 40230 4431 40282
rect 4443 40230 4495 40282
rect 4507 40230 4559 40282
rect 10982 40230 11034 40282
rect 11046 40230 11098 40282
rect 11110 40230 11162 40282
rect 11174 40230 11226 40282
rect 17648 40230 17700 40282
rect 17712 40230 17764 40282
rect 17776 40230 17828 40282
rect 17840 40230 17892 40282
rect 3700 40128 3752 40180
rect 11980 40171 12032 40180
rect 11980 40137 11989 40171
rect 11989 40137 12023 40171
rect 12023 40137 12032 40171
rect 11980 40128 12032 40137
rect 12164 40128 12216 40180
rect 12348 40128 12400 40180
rect 4896 40060 4948 40112
rect 7472 40060 7524 40112
rect 9036 40060 9088 40112
rect 6920 39992 6972 40044
rect 10048 40060 10100 40112
rect 10232 40060 10284 40112
rect 10968 40060 11020 40112
rect 14924 40128 14976 40180
rect 15200 40128 15252 40180
rect 15936 40128 15988 40180
rect 17224 40171 17276 40180
rect 17224 40137 17233 40171
rect 17233 40137 17267 40171
rect 17267 40137 17276 40171
rect 17224 40128 17276 40137
rect 18144 40128 18196 40180
rect 4620 39924 4672 39976
rect 4436 39856 4488 39908
rect 6000 39924 6052 39976
rect 7196 39967 7248 39976
rect 4896 39856 4948 39908
rect 4344 39831 4396 39840
rect 4344 39797 4353 39831
rect 4353 39797 4387 39831
rect 4387 39797 4396 39831
rect 4344 39788 4396 39797
rect 5724 39831 5776 39840
rect 5724 39797 5733 39831
rect 5733 39797 5767 39831
rect 5767 39797 5776 39831
rect 5724 39788 5776 39797
rect 6184 39856 6236 39908
rect 7196 39933 7205 39967
rect 7205 39933 7239 39967
rect 7239 39933 7248 39967
rect 7196 39924 7248 39933
rect 11428 39992 11480 40044
rect 6920 39856 6972 39908
rect 9588 39856 9640 39908
rect 6644 39788 6696 39840
rect 8576 39788 8628 39840
rect 9220 39788 9272 39840
rect 10048 39788 10100 39840
rect 10876 39831 10928 39840
rect 10876 39797 10885 39831
rect 10885 39797 10919 39831
rect 10919 39797 10928 39831
rect 10876 39788 10928 39797
rect 11244 39831 11296 39840
rect 11244 39797 11253 39831
rect 11253 39797 11287 39831
rect 11287 39797 11296 39831
rect 11244 39788 11296 39797
rect 11704 39967 11756 39976
rect 11704 39933 11713 39967
rect 11713 39933 11747 39967
rect 11747 39933 11756 39967
rect 11704 39924 11756 39933
rect 11888 39967 11940 39976
rect 11888 39933 11897 39967
rect 11897 39933 11931 39967
rect 11931 39933 11940 39967
rect 11888 39924 11940 39933
rect 12532 39967 12584 39976
rect 12532 39933 12541 39967
rect 12541 39933 12575 39967
rect 12575 39933 12584 39967
rect 12532 39924 12584 39933
rect 13544 39924 13596 39976
rect 16304 39967 16356 39976
rect 16304 39933 16313 39967
rect 16313 39933 16347 39967
rect 16347 39933 16356 39967
rect 16304 39924 16356 39933
rect 16764 39967 16816 39976
rect 15200 39856 15252 39908
rect 15844 39899 15896 39908
rect 15844 39865 15853 39899
rect 15853 39865 15887 39899
rect 15887 39865 15896 39899
rect 16764 39933 16773 39967
rect 16773 39933 16807 39967
rect 16807 39933 16816 39967
rect 16764 39924 16816 39933
rect 16856 39924 16908 39976
rect 15844 39856 15896 39865
rect 12164 39788 12216 39840
rect 13084 39788 13136 39840
rect 13268 39788 13320 39840
rect 17132 39788 17184 39840
rect 18420 39788 18472 39840
rect 7648 39686 7700 39738
rect 7712 39686 7764 39738
rect 7776 39686 7828 39738
rect 7840 39686 7892 39738
rect 14315 39686 14367 39738
rect 14379 39686 14431 39738
rect 14443 39686 14495 39738
rect 14507 39686 14559 39738
rect 2136 39584 2188 39636
rect 2320 39584 2372 39636
rect 4436 39584 4488 39636
rect 4620 39627 4672 39636
rect 4620 39593 4629 39627
rect 4629 39593 4663 39627
rect 4663 39593 4672 39627
rect 4620 39584 4672 39593
rect 5264 39584 5316 39636
rect 7196 39584 7248 39636
rect 9588 39584 9640 39636
rect 11888 39627 11940 39636
rect 2964 39516 3016 39568
rect 3332 39516 3384 39568
rect 3240 39491 3292 39500
rect 3240 39457 3249 39491
rect 3249 39457 3283 39491
rect 3283 39457 3292 39491
rect 3608 39516 3660 39568
rect 8116 39516 8168 39568
rect 9404 39516 9456 39568
rect 11888 39593 11897 39627
rect 11897 39593 11931 39627
rect 11931 39593 11940 39627
rect 11888 39584 11940 39593
rect 12348 39584 12400 39636
rect 14648 39584 14700 39636
rect 17316 39627 17368 39636
rect 17316 39593 17325 39627
rect 17325 39593 17359 39627
rect 17359 39593 17368 39627
rect 17316 39584 17368 39593
rect 3700 39491 3752 39500
rect 3240 39448 3292 39457
rect 3700 39457 3709 39491
rect 3709 39457 3743 39491
rect 3743 39457 3752 39491
rect 3700 39448 3752 39457
rect 4620 39491 4672 39500
rect 4620 39457 4629 39491
rect 4629 39457 4663 39491
rect 4663 39457 4672 39491
rect 4620 39448 4672 39457
rect 5356 39448 5408 39500
rect 7656 39491 7708 39500
rect 3332 39423 3384 39432
rect 3332 39389 3341 39423
rect 3341 39389 3375 39423
rect 3375 39389 3384 39423
rect 3332 39380 3384 39389
rect 7656 39457 7665 39491
rect 7665 39457 7699 39491
rect 7699 39457 7708 39491
rect 7656 39448 7708 39457
rect 10876 39491 10928 39500
rect 7564 39380 7616 39432
rect 6644 39287 6696 39296
rect 6644 39253 6653 39287
rect 6653 39253 6687 39287
rect 6687 39253 6696 39287
rect 6644 39244 6696 39253
rect 10876 39457 10885 39491
rect 10885 39457 10919 39491
rect 10919 39457 10928 39491
rect 10876 39448 10928 39457
rect 11244 39448 11296 39500
rect 12440 39516 12492 39568
rect 14188 39559 14240 39568
rect 14188 39525 14197 39559
rect 14197 39525 14231 39559
rect 14231 39525 14240 39559
rect 14188 39516 14240 39525
rect 14372 39516 14424 39568
rect 15292 39516 15344 39568
rect 11980 39448 12032 39500
rect 13176 39448 13228 39500
rect 13452 39448 13504 39500
rect 15660 39448 15712 39500
rect 15936 39491 15988 39500
rect 15936 39457 15945 39491
rect 15945 39457 15979 39491
rect 15979 39457 15988 39491
rect 15936 39448 15988 39457
rect 16304 39491 16356 39500
rect 16304 39457 16313 39491
rect 16313 39457 16347 39491
rect 16347 39457 16356 39491
rect 16304 39448 16356 39457
rect 16856 39491 16908 39500
rect 16856 39457 16865 39491
rect 16865 39457 16899 39491
rect 16899 39457 16908 39491
rect 16856 39448 16908 39457
rect 11612 39380 11664 39432
rect 12716 39380 12768 39432
rect 12900 39380 12952 39432
rect 15292 39380 15344 39432
rect 16764 39380 16816 39432
rect 11244 39312 11296 39364
rect 9496 39244 9548 39296
rect 13452 39244 13504 39296
rect 15200 39244 15252 39296
rect 15476 39244 15528 39296
rect 4315 39142 4367 39194
rect 4379 39142 4431 39194
rect 4443 39142 4495 39194
rect 4507 39142 4559 39194
rect 10982 39142 11034 39194
rect 11046 39142 11098 39194
rect 11110 39142 11162 39194
rect 11174 39142 11226 39194
rect 17648 39142 17700 39194
rect 17712 39142 17764 39194
rect 17776 39142 17828 39194
rect 17840 39142 17892 39194
rect 2688 39083 2740 39092
rect 2688 39049 2697 39083
rect 2697 39049 2731 39083
rect 2731 39049 2740 39083
rect 2688 39040 2740 39049
rect 3240 39040 3292 39092
rect 3332 39040 3384 39092
rect 3792 39083 3844 39092
rect 3792 39049 3801 39083
rect 3801 39049 3835 39083
rect 3835 39049 3844 39083
rect 3792 39040 3844 39049
rect 5356 39040 5408 39092
rect 5724 39040 5776 39092
rect 6920 39083 6972 39092
rect 6920 39049 6929 39083
rect 6929 39049 6963 39083
rect 6963 39049 6972 39083
rect 6920 39040 6972 39049
rect 8392 39083 8444 39092
rect 5632 38972 5684 39024
rect 4712 38904 4764 38956
rect 3332 38836 3384 38888
rect 3792 38836 3844 38888
rect 5080 38879 5132 38888
rect 5080 38845 5089 38879
rect 5089 38845 5123 38879
rect 5123 38845 5132 38879
rect 5080 38836 5132 38845
rect 6184 38836 6236 38888
rect 7472 38879 7524 38888
rect 7472 38845 7481 38879
rect 7481 38845 7515 38879
rect 7515 38845 7524 38879
rect 7472 38836 7524 38845
rect 8392 39049 8401 39083
rect 8401 39049 8435 39083
rect 8435 39049 8444 39083
rect 8392 39040 8444 39049
rect 10324 39040 10376 39092
rect 10232 38972 10284 39024
rect 10600 38947 10652 38956
rect 10600 38913 10609 38947
rect 10609 38913 10643 38947
rect 10643 38913 10652 38947
rect 10600 38904 10652 38913
rect 8484 38879 8536 38888
rect 8484 38845 8493 38879
rect 8493 38845 8527 38879
rect 8527 38845 8536 38879
rect 8484 38836 8536 38845
rect 8852 38879 8904 38888
rect 8852 38845 8861 38879
rect 8861 38845 8895 38879
rect 8895 38845 8904 38879
rect 8852 38836 8904 38845
rect 9588 38836 9640 38888
rect 9956 38836 10008 38888
rect 10232 38836 10284 38888
rect 10416 38879 10468 38888
rect 10416 38845 10425 38879
rect 10425 38845 10459 38879
rect 10459 38845 10468 38879
rect 10416 38836 10468 38845
rect 3700 38768 3752 38820
rect 6736 38768 6788 38820
rect 7656 38768 7708 38820
rect 8116 38768 8168 38820
rect 10600 38768 10652 38820
rect 12532 39040 12584 39092
rect 12716 39040 12768 39092
rect 13636 39083 13688 39092
rect 13636 39049 13645 39083
rect 13645 39049 13679 39083
rect 13679 39049 13688 39083
rect 13636 39040 13688 39049
rect 14372 39083 14424 39092
rect 14372 39049 14381 39083
rect 14381 39049 14415 39083
rect 14415 39049 14424 39083
rect 14372 39040 14424 39049
rect 15384 39040 15436 39092
rect 16488 39040 16540 39092
rect 18236 39083 18288 39092
rect 18236 39049 18245 39083
rect 18245 39049 18279 39083
rect 18279 39049 18288 39083
rect 18236 39040 18288 39049
rect 12348 38972 12400 39024
rect 10968 38904 11020 38956
rect 12992 38947 13044 38956
rect 12992 38913 13001 38947
rect 13001 38913 13035 38947
rect 13035 38913 13044 38947
rect 12992 38904 13044 38913
rect 11060 38879 11112 38888
rect 11060 38845 11069 38879
rect 11069 38845 11103 38879
rect 11103 38845 11112 38879
rect 11060 38836 11112 38845
rect 11980 38879 12032 38888
rect 11980 38845 11989 38879
rect 11989 38845 12023 38879
rect 12023 38845 12032 38879
rect 11980 38836 12032 38845
rect 12164 38879 12216 38888
rect 12164 38845 12173 38879
rect 12173 38845 12207 38879
rect 12207 38845 12216 38879
rect 12164 38836 12216 38845
rect 13636 38904 13688 38956
rect 16212 39015 16264 39024
rect 16212 38981 16221 39015
rect 16221 38981 16255 39015
rect 16255 38981 16264 39015
rect 16212 38972 16264 38981
rect 13544 38836 13596 38888
rect 13728 38768 13780 38820
rect 8852 38700 8904 38752
rect 12440 38700 12492 38752
rect 13452 38700 13504 38752
rect 15292 38836 15344 38888
rect 16304 38879 16356 38888
rect 16304 38845 16313 38879
rect 16313 38845 16347 38879
rect 16347 38845 16356 38879
rect 16304 38836 16356 38845
rect 16488 38879 16540 38888
rect 16488 38845 16497 38879
rect 16497 38845 16531 38879
rect 16531 38845 16540 38879
rect 16488 38836 16540 38845
rect 15936 38768 15988 38820
rect 16764 38768 16816 38820
rect 16948 38836 17000 38888
rect 18052 38768 18104 38820
rect 7648 38598 7700 38650
rect 7712 38598 7764 38650
rect 7776 38598 7828 38650
rect 7840 38598 7892 38650
rect 14315 38598 14367 38650
rect 14379 38598 14431 38650
rect 14443 38598 14495 38650
rect 14507 38598 14559 38650
rect 4620 38496 4672 38548
rect 5540 38496 5592 38548
rect 3976 38428 4028 38480
rect 1584 38360 1636 38412
rect 3516 38360 3568 38412
rect 5356 38360 5408 38412
rect 1676 38292 1728 38344
rect 3976 38335 4028 38344
rect 3976 38301 3985 38335
rect 3985 38301 4019 38335
rect 4019 38301 4028 38335
rect 3976 38292 4028 38301
rect 6828 38496 6880 38548
rect 8116 38496 8168 38548
rect 9312 38496 9364 38548
rect 10508 38496 10560 38548
rect 10784 38496 10836 38548
rect 10876 38496 10928 38548
rect 12440 38496 12492 38548
rect 12808 38496 12860 38548
rect 13728 38496 13780 38548
rect 8484 38428 8536 38480
rect 6828 38403 6880 38412
rect 6828 38369 6837 38403
rect 6837 38369 6871 38403
rect 6871 38369 6880 38403
rect 6828 38360 6880 38369
rect 10968 38428 11020 38480
rect 12348 38428 12400 38480
rect 8392 38292 8444 38344
rect 8944 38360 8996 38412
rect 8576 38224 8628 38276
rect 9772 38360 9824 38412
rect 10784 38403 10836 38412
rect 10784 38369 10793 38403
rect 10793 38369 10827 38403
rect 10827 38369 10836 38403
rect 10784 38360 10836 38369
rect 10876 38360 10928 38412
rect 10416 38292 10468 38344
rect 13636 38360 13688 38412
rect 13728 38292 13780 38344
rect 14740 38403 14792 38412
rect 14740 38369 14749 38403
rect 14749 38369 14783 38403
rect 14783 38369 14792 38403
rect 14740 38360 14792 38369
rect 15292 38496 15344 38548
rect 15844 38496 15896 38548
rect 16856 38496 16908 38548
rect 17316 38496 17368 38548
rect 15568 38403 15620 38412
rect 15568 38369 15577 38403
rect 15577 38369 15611 38403
rect 15611 38369 15620 38403
rect 15568 38360 15620 38369
rect 16856 38403 16908 38412
rect 16856 38369 16865 38403
rect 16865 38369 16899 38403
rect 16899 38369 16908 38403
rect 16856 38360 16908 38369
rect 16304 38292 16356 38344
rect 9772 38224 9824 38276
rect 11244 38224 11296 38276
rect 12808 38224 12860 38276
rect 13544 38224 13596 38276
rect 15660 38224 15712 38276
rect 5080 38156 5132 38208
rect 6184 38199 6236 38208
rect 6184 38165 6193 38199
rect 6193 38165 6227 38199
rect 6227 38165 6236 38199
rect 6184 38156 6236 38165
rect 9220 38199 9272 38208
rect 9220 38165 9229 38199
rect 9229 38165 9263 38199
rect 9263 38165 9272 38199
rect 9220 38156 9272 38165
rect 9956 38156 10008 38208
rect 10416 38156 10468 38208
rect 14648 38199 14700 38208
rect 14648 38165 14657 38199
rect 14657 38165 14691 38199
rect 14691 38165 14700 38199
rect 14648 38156 14700 38165
rect 4315 38054 4367 38106
rect 4379 38054 4431 38106
rect 4443 38054 4495 38106
rect 4507 38054 4559 38106
rect 10982 38054 11034 38106
rect 11046 38054 11098 38106
rect 11110 38054 11162 38106
rect 11174 38054 11226 38106
rect 17648 38054 17700 38106
rect 17712 38054 17764 38106
rect 17776 38054 17828 38106
rect 17840 38054 17892 38106
rect 1676 37952 1728 38004
rect 3240 37952 3292 38004
rect 3516 37995 3568 38004
rect 3516 37961 3525 37995
rect 3525 37961 3559 37995
rect 3559 37961 3568 37995
rect 3516 37952 3568 37961
rect 9312 37952 9364 38004
rect 13636 37952 13688 38004
rect 15016 37952 15068 38004
rect 7380 37927 7432 37936
rect 7380 37893 7389 37927
rect 7389 37893 7423 37927
rect 7423 37893 7432 37927
rect 7380 37884 7432 37893
rect 7472 37884 7524 37936
rect 8116 37884 8168 37936
rect 10416 37884 10468 37936
rect 5540 37816 5592 37868
rect 6000 37816 6052 37868
rect 1860 37748 1912 37800
rect 3608 37748 3660 37800
rect 3976 37748 4028 37800
rect 1768 37612 1820 37664
rect 3792 37655 3844 37664
rect 3792 37621 3801 37655
rect 3801 37621 3835 37655
rect 3835 37621 3844 37655
rect 6736 37791 6788 37800
rect 6736 37757 6745 37791
rect 6745 37757 6779 37791
rect 6779 37757 6788 37791
rect 6736 37748 6788 37757
rect 6920 37791 6972 37800
rect 6920 37757 6929 37791
rect 6929 37757 6963 37791
rect 6963 37757 6972 37791
rect 6920 37748 6972 37757
rect 7472 37791 7524 37800
rect 7472 37757 7481 37791
rect 7481 37757 7515 37791
rect 7515 37757 7524 37791
rect 7472 37748 7524 37757
rect 10140 37816 10192 37868
rect 9128 37748 9180 37800
rect 6000 37680 6052 37732
rect 6828 37680 6880 37732
rect 9864 37723 9916 37732
rect 9864 37689 9873 37723
rect 9873 37689 9907 37723
rect 9907 37689 9916 37723
rect 9864 37680 9916 37689
rect 11428 37816 11480 37868
rect 11888 37816 11940 37868
rect 12624 37859 12676 37868
rect 11980 37791 12032 37800
rect 11980 37757 11989 37791
rect 11989 37757 12023 37791
rect 12023 37757 12032 37791
rect 11980 37748 12032 37757
rect 12072 37748 12124 37800
rect 12624 37825 12633 37859
rect 12633 37825 12667 37859
rect 12667 37825 12676 37859
rect 12624 37816 12676 37825
rect 10968 37680 11020 37732
rect 12440 37680 12492 37732
rect 14924 37748 14976 37800
rect 15568 37952 15620 38004
rect 16488 37952 16540 38004
rect 16856 37952 16908 38004
rect 17960 37952 18012 38004
rect 16856 37859 16908 37868
rect 16856 37825 16865 37859
rect 16865 37825 16899 37859
rect 16899 37825 16908 37859
rect 16856 37816 16908 37825
rect 15568 37748 15620 37800
rect 15936 37748 15988 37800
rect 14740 37680 14792 37732
rect 15660 37680 15712 37732
rect 16304 37680 16356 37732
rect 16488 37748 16540 37800
rect 17316 37791 17368 37800
rect 17316 37757 17325 37791
rect 17325 37757 17359 37791
rect 17359 37757 17368 37791
rect 17316 37748 17368 37757
rect 3792 37612 3844 37621
rect 7012 37612 7064 37664
rect 7472 37612 7524 37664
rect 8392 37612 8444 37664
rect 8484 37612 8536 37664
rect 9312 37612 9364 37664
rect 10416 37612 10468 37664
rect 10784 37655 10836 37664
rect 10784 37621 10793 37655
rect 10793 37621 10827 37655
rect 10827 37621 10836 37655
rect 10784 37612 10836 37621
rect 10876 37612 10928 37664
rect 11888 37655 11940 37664
rect 11888 37621 11897 37655
rect 11897 37621 11931 37655
rect 11931 37621 11940 37655
rect 11888 37612 11940 37621
rect 13728 37612 13780 37664
rect 14096 37612 14148 37664
rect 15936 37612 15988 37664
rect 7648 37510 7700 37562
rect 7712 37510 7764 37562
rect 7776 37510 7828 37562
rect 7840 37510 7892 37562
rect 14315 37510 14367 37562
rect 14379 37510 14431 37562
rect 14443 37510 14495 37562
rect 14507 37510 14559 37562
rect 5080 37408 5132 37460
rect 6920 37408 6972 37460
rect 9312 37408 9364 37460
rect 11244 37408 11296 37460
rect 12348 37408 12400 37460
rect 6736 37340 6788 37392
rect 9036 37340 9088 37392
rect 1492 37272 1544 37324
rect 1860 37272 1912 37324
rect 3700 37272 3752 37324
rect 6184 37272 6236 37324
rect 6828 37315 6880 37324
rect 3608 37247 3660 37256
rect 1768 37068 1820 37120
rect 3240 37068 3292 37120
rect 3608 37213 3617 37247
rect 3617 37213 3651 37247
rect 3651 37213 3660 37247
rect 3608 37204 3660 37213
rect 3976 37204 4028 37256
rect 6828 37281 6837 37315
rect 6837 37281 6871 37315
rect 6871 37281 6880 37315
rect 6828 37272 6880 37281
rect 6920 37272 6972 37324
rect 7196 37272 7248 37324
rect 8576 37272 8628 37324
rect 8760 37315 8812 37324
rect 8760 37281 8769 37315
rect 8769 37281 8803 37315
rect 8803 37281 8812 37315
rect 8760 37272 8812 37281
rect 9128 37315 9180 37324
rect 9128 37281 9137 37315
rect 9137 37281 9171 37315
rect 9171 37281 9180 37315
rect 9128 37272 9180 37281
rect 9312 37315 9364 37324
rect 9312 37281 9321 37315
rect 9321 37281 9355 37315
rect 9355 37281 9364 37315
rect 9312 37272 9364 37281
rect 9588 37272 9640 37324
rect 11980 37340 12032 37392
rect 12440 37340 12492 37392
rect 14924 37408 14976 37460
rect 7380 37204 7432 37256
rect 8300 37204 8352 37256
rect 11336 37272 11388 37324
rect 12072 37315 12124 37324
rect 12072 37281 12081 37315
rect 12081 37281 12115 37315
rect 12115 37281 12124 37315
rect 12072 37272 12124 37281
rect 13084 37272 13136 37324
rect 14096 37272 14148 37324
rect 14556 37272 14608 37324
rect 15384 37408 15436 37460
rect 17408 37451 17460 37460
rect 17408 37417 17417 37451
rect 17417 37417 17451 37451
rect 17451 37417 17460 37451
rect 17408 37408 17460 37417
rect 12164 37204 12216 37256
rect 14648 37204 14700 37256
rect 15108 37247 15160 37256
rect 15108 37213 15117 37247
rect 15117 37213 15151 37247
rect 15151 37213 15160 37247
rect 15108 37204 15160 37213
rect 15936 37340 15988 37392
rect 15568 37315 15620 37324
rect 15568 37281 15577 37315
rect 15577 37281 15611 37315
rect 15611 37281 15620 37315
rect 15568 37272 15620 37281
rect 15660 37272 15712 37324
rect 15936 37204 15988 37256
rect 16120 37247 16172 37256
rect 16120 37213 16129 37247
rect 16129 37213 16163 37247
rect 16163 37213 16172 37247
rect 16120 37204 16172 37213
rect 6276 37136 6328 37188
rect 10968 37136 11020 37188
rect 5632 37111 5684 37120
rect 5632 37077 5641 37111
rect 5641 37077 5675 37111
rect 5675 37077 5684 37111
rect 5632 37068 5684 37077
rect 8116 37068 8168 37120
rect 8484 37068 8536 37120
rect 10784 37068 10836 37120
rect 14188 37068 14240 37120
rect 15108 37068 15160 37120
rect 17132 37247 17184 37256
rect 17132 37213 17141 37247
rect 17141 37213 17175 37247
rect 17175 37213 17184 37247
rect 17132 37204 17184 37213
rect 17408 37136 17460 37188
rect 18052 37068 18104 37120
rect 4315 36966 4367 37018
rect 4379 36966 4431 37018
rect 4443 36966 4495 37018
rect 4507 36966 4559 37018
rect 10982 36966 11034 37018
rect 11046 36966 11098 37018
rect 11110 36966 11162 37018
rect 11174 36966 11226 37018
rect 17648 36966 17700 37018
rect 17712 36966 17764 37018
rect 17776 36966 17828 37018
rect 17840 36966 17892 37018
rect 4896 36864 4948 36916
rect 3976 36796 4028 36848
rect 6276 36864 6328 36916
rect 8300 36864 8352 36916
rect 9312 36864 9364 36916
rect 10232 36907 10284 36916
rect 10232 36873 10241 36907
rect 10241 36873 10275 36907
rect 10275 36873 10284 36907
rect 10232 36864 10284 36873
rect 10508 36864 10560 36916
rect 10876 36907 10928 36916
rect 10876 36873 10885 36907
rect 10885 36873 10919 36907
rect 10919 36873 10928 36907
rect 10876 36864 10928 36873
rect 12348 36864 12400 36916
rect 12808 36907 12860 36916
rect 12808 36873 12817 36907
rect 12817 36873 12851 36907
rect 12851 36873 12860 36907
rect 12808 36864 12860 36873
rect 13636 36864 13688 36916
rect 14556 36864 14608 36916
rect 15200 36864 15252 36916
rect 18052 36907 18104 36916
rect 18052 36873 18061 36907
rect 18061 36873 18095 36907
rect 18095 36873 18104 36907
rect 18052 36864 18104 36873
rect 5264 36660 5316 36712
rect 5632 36796 5684 36848
rect 5908 36796 5960 36848
rect 6184 36796 6236 36848
rect 9128 36796 9180 36848
rect 10140 36796 10192 36848
rect 12900 36796 12952 36848
rect 10232 36728 10284 36780
rect 15292 36796 15344 36848
rect 16488 36796 16540 36848
rect 16764 36796 16816 36848
rect 17408 36796 17460 36848
rect 14004 36728 14056 36780
rect 16396 36728 16448 36780
rect 6276 36703 6328 36712
rect 6276 36669 6285 36703
rect 6285 36669 6319 36703
rect 6319 36669 6328 36703
rect 6276 36660 6328 36669
rect 7472 36660 7524 36712
rect 7932 36660 7984 36712
rect 8116 36703 8168 36712
rect 8116 36669 8125 36703
rect 8125 36669 8159 36703
rect 8159 36669 8168 36703
rect 8116 36660 8168 36669
rect 9956 36660 10008 36712
rect 10140 36660 10192 36712
rect 10508 36660 10560 36712
rect 12440 36660 12492 36712
rect 11520 36592 11572 36644
rect 11980 36592 12032 36644
rect 12256 36592 12308 36644
rect 14096 36660 14148 36712
rect 15844 36660 15896 36712
rect 16580 36635 16632 36644
rect 16580 36601 16589 36635
rect 16589 36601 16623 36635
rect 16623 36601 16632 36635
rect 17408 36660 17460 36712
rect 16580 36592 16632 36601
rect 17684 36592 17736 36644
rect 17868 36592 17920 36644
rect 1768 36524 1820 36576
rect 3240 36567 3292 36576
rect 3240 36533 3249 36567
rect 3249 36533 3283 36567
rect 3283 36533 3292 36567
rect 3240 36524 3292 36533
rect 4896 36524 4948 36576
rect 5540 36524 5592 36576
rect 5816 36524 5868 36576
rect 6276 36524 6328 36576
rect 6828 36524 6880 36576
rect 7012 36567 7064 36576
rect 7012 36533 7021 36567
rect 7021 36533 7055 36567
rect 7055 36533 7064 36567
rect 7012 36524 7064 36533
rect 11336 36524 11388 36576
rect 14924 36524 14976 36576
rect 16120 36567 16172 36576
rect 16120 36533 16129 36567
rect 16129 36533 16163 36567
rect 16163 36533 16172 36567
rect 16120 36524 16172 36533
rect 7648 36422 7700 36474
rect 7712 36422 7764 36474
rect 7776 36422 7828 36474
rect 7840 36422 7892 36474
rect 14315 36422 14367 36474
rect 14379 36422 14431 36474
rect 14443 36422 14495 36474
rect 14507 36422 14559 36474
rect 5264 36320 5316 36372
rect 6736 36320 6788 36372
rect 8760 36320 8812 36372
rect 9312 36363 9364 36372
rect 9312 36329 9321 36363
rect 9321 36329 9355 36363
rect 9355 36329 9364 36363
rect 9312 36320 9364 36329
rect 10508 36320 10560 36372
rect 10876 36320 10928 36372
rect 12164 36363 12216 36372
rect 12164 36329 12173 36363
rect 12173 36329 12207 36363
rect 12207 36329 12216 36363
rect 12164 36320 12216 36329
rect 12716 36363 12768 36372
rect 12716 36329 12725 36363
rect 12725 36329 12759 36363
rect 12759 36329 12768 36363
rect 12716 36320 12768 36329
rect 13452 36363 13504 36372
rect 13452 36329 13461 36363
rect 13461 36329 13495 36363
rect 13495 36329 13504 36363
rect 13452 36320 13504 36329
rect 14096 36363 14148 36372
rect 14096 36329 14105 36363
rect 14105 36329 14139 36363
rect 14139 36329 14148 36363
rect 14096 36320 14148 36329
rect 14648 36320 14700 36372
rect 15200 36320 15252 36372
rect 16396 36363 16448 36372
rect 16396 36329 16405 36363
rect 16405 36329 16439 36363
rect 16439 36329 16448 36363
rect 16396 36320 16448 36329
rect 16580 36320 16632 36372
rect 17408 36363 17460 36372
rect 17408 36329 17417 36363
rect 17417 36329 17451 36363
rect 17451 36329 17460 36363
rect 17408 36320 17460 36329
rect 4896 36295 4948 36304
rect 4896 36261 4905 36295
rect 4905 36261 4939 36295
rect 4939 36261 4948 36295
rect 4896 36252 4948 36261
rect 8116 36252 8168 36304
rect 11796 36252 11848 36304
rect 12808 36252 12860 36304
rect 14556 36252 14608 36304
rect 5356 36227 5408 36236
rect 5356 36193 5365 36227
rect 5365 36193 5399 36227
rect 5399 36193 5408 36227
rect 5356 36184 5408 36193
rect 7196 36227 7248 36236
rect 7196 36193 7205 36227
rect 7205 36193 7239 36227
rect 7239 36193 7248 36227
rect 7196 36184 7248 36193
rect 7288 36184 7340 36236
rect 9220 36227 9272 36236
rect 9220 36193 9229 36227
rect 9229 36193 9263 36227
rect 9263 36193 9272 36227
rect 9220 36184 9272 36193
rect 11336 36227 11388 36236
rect 11336 36193 11345 36227
rect 11345 36193 11379 36227
rect 11379 36193 11388 36227
rect 11336 36184 11388 36193
rect 13084 36227 13136 36236
rect 13084 36193 13093 36227
rect 13093 36193 13127 36227
rect 13127 36193 13136 36227
rect 13084 36184 13136 36193
rect 14740 36227 14792 36236
rect 14740 36193 14749 36227
rect 14749 36193 14783 36227
rect 14783 36193 14792 36227
rect 14740 36184 14792 36193
rect 14924 36227 14976 36236
rect 14924 36193 14933 36227
rect 14933 36193 14967 36227
rect 14967 36193 14976 36227
rect 14924 36184 14976 36193
rect 16488 36252 16540 36304
rect 8300 36116 8352 36168
rect 14280 36116 14332 36168
rect 17960 36184 18012 36236
rect 16396 36116 16448 36168
rect 1860 35980 1912 36032
rect 2044 35980 2096 36032
rect 2320 35980 2372 36032
rect 5908 35980 5960 36032
rect 6460 35980 6512 36032
rect 16580 35980 16632 36032
rect 4315 35878 4367 35930
rect 4379 35878 4431 35930
rect 4443 35878 4495 35930
rect 4507 35878 4559 35930
rect 10982 35878 11034 35930
rect 11046 35878 11098 35930
rect 11110 35878 11162 35930
rect 11174 35878 11226 35930
rect 17648 35878 17700 35930
rect 17712 35878 17764 35930
rect 17776 35878 17828 35930
rect 17840 35878 17892 35930
rect 3884 35776 3936 35828
rect 5356 35776 5408 35828
rect 6368 35819 6420 35828
rect 6368 35785 6377 35819
rect 6377 35785 6411 35819
rect 6411 35785 6420 35819
rect 6368 35776 6420 35785
rect 7288 35776 7340 35828
rect 8484 35776 8536 35828
rect 9220 35776 9272 35828
rect 9588 35776 9640 35828
rect 11336 35776 11388 35828
rect 12532 35819 12584 35828
rect 12532 35785 12541 35819
rect 12541 35785 12575 35819
rect 12575 35785 12584 35819
rect 12532 35776 12584 35785
rect 13084 35819 13136 35828
rect 13084 35785 13093 35819
rect 13093 35785 13127 35819
rect 13127 35785 13136 35819
rect 13084 35776 13136 35785
rect 14280 35776 14332 35828
rect 14924 35776 14976 35828
rect 15660 35776 15712 35828
rect 15844 35819 15896 35828
rect 15844 35785 15853 35819
rect 15853 35785 15887 35819
rect 15887 35785 15896 35819
rect 15844 35776 15896 35785
rect 16488 35776 16540 35828
rect 18144 35819 18196 35828
rect 18144 35785 18153 35819
rect 18153 35785 18187 35819
rect 18187 35785 18196 35819
rect 18144 35776 18196 35785
rect 8300 35708 8352 35760
rect 9404 35708 9456 35760
rect 1860 35640 1912 35692
rect 2504 35640 2556 35692
rect 1584 35572 1636 35624
rect 6828 35572 6880 35624
rect 9956 35615 10008 35624
rect 9956 35581 9965 35615
rect 9965 35581 9999 35615
rect 9999 35581 10008 35615
rect 9956 35572 10008 35581
rect 12164 35708 12216 35760
rect 13544 35708 13596 35760
rect 15292 35708 15344 35760
rect 17500 35751 17552 35760
rect 17500 35717 17509 35751
rect 17509 35717 17543 35751
rect 17543 35717 17552 35751
rect 17500 35708 17552 35717
rect 12348 35640 12400 35692
rect 11428 35572 11480 35624
rect 11796 35572 11848 35624
rect 11980 35615 12032 35624
rect 11980 35581 11989 35615
rect 11989 35581 12023 35615
rect 12023 35581 12032 35615
rect 11980 35572 12032 35581
rect 14188 35615 14240 35624
rect 14188 35581 14197 35615
rect 14197 35581 14231 35615
rect 14231 35581 14240 35615
rect 14188 35572 14240 35581
rect 15844 35572 15896 35624
rect 16580 35572 16632 35624
rect 14556 35504 14608 35556
rect 14924 35504 14976 35556
rect 15936 35504 15988 35556
rect 5724 35436 5776 35488
rect 6000 35436 6052 35488
rect 7196 35479 7248 35488
rect 7196 35445 7205 35479
rect 7205 35445 7239 35479
rect 7239 35445 7248 35479
rect 7196 35436 7248 35445
rect 13268 35436 13320 35488
rect 13544 35436 13596 35488
rect 13728 35479 13780 35488
rect 13728 35445 13737 35479
rect 13737 35445 13771 35479
rect 13771 35445 13780 35479
rect 13728 35436 13780 35445
rect 14740 35436 14792 35488
rect 7648 35334 7700 35386
rect 7712 35334 7764 35386
rect 7776 35334 7828 35386
rect 7840 35334 7892 35386
rect 14315 35334 14367 35386
rect 14379 35334 14431 35386
rect 14443 35334 14495 35386
rect 14507 35334 14559 35386
rect 6184 35232 6236 35284
rect 14188 35275 14240 35284
rect 14188 35241 14197 35275
rect 14197 35241 14231 35275
rect 14231 35241 14240 35275
rect 14188 35232 14240 35241
rect 14924 35232 14976 35284
rect 17408 35275 17460 35284
rect 17408 35241 17417 35275
rect 17417 35241 17451 35275
rect 17451 35241 17460 35275
rect 17408 35232 17460 35241
rect 2320 35164 2372 35216
rect 6000 35096 6052 35148
rect 6920 35096 6972 35148
rect 9680 35164 9732 35216
rect 13084 35164 13136 35216
rect 2504 35028 2556 35080
rect 3976 35071 4028 35080
rect 3976 35037 3985 35071
rect 3985 35037 4019 35071
rect 4019 35037 4028 35071
rect 3976 35028 4028 35037
rect 7288 35028 7340 35080
rect 4620 34960 4672 35012
rect 8484 35096 8536 35148
rect 9956 35096 10008 35148
rect 13636 35096 13688 35148
rect 14740 35139 14792 35148
rect 14740 35105 14749 35139
rect 14749 35105 14783 35139
rect 14783 35105 14792 35139
rect 14740 35096 14792 35105
rect 16212 35139 16264 35148
rect 16212 35105 16221 35139
rect 16221 35105 16255 35139
rect 16255 35105 16264 35139
rect 16212 35096 16264 35105
rect 16488 35096 16540 35148
rect 1584 34935 1636 34944
rect 1584 34901 1593 34935
rect 1593 34901 1627 34935
rect 1627 34901 1636 34935
rect 1584 34892 1636 34901
rect 5080 34892 5132 34944
rect 6736 34892 6788 34944
rect 9772 34892 9824 34944
rect 16304 35028 16356 35080
rect 17132 35071 17184 35080
rect 17132 35037 17141 35071
rect 17141 35037 17175 35071
rect 17175 35037 17184 35071
rect 17132 35028 17184 35037
rect 14648 34960 14700 35012
rect 16396 34960 16448 35012
rect 15936 34892 15988 34944
rect 4315 34790 4367 34842
rect 4379 34790 4431 34842
rect 4443 34790 4495 34842
rect 4507 34790 4559 34842
rect 10982 34790 11034 34842
rect 11046 34790 11098 34842
rect 11110 34790 11162 34842
rect 11174 34790 11226 34842
rect 17648 34790 17700 34842
rect 17712 34790 17764 34842
rect 17776 34790 17828 34842
rect 17840 34790 17892 34842
rect 6000 34688 6052 34740
rect 7932 34688 7984 34740
rect 14740 34731 14792 34740
rect 14740 34697 14749 34731
rect 14749 34697 14783 34731
rect 14783 34697 14792 34731
rect 14740 34688 14792 34697
rect 15568 34731 15620 34740
rect 15568 34697 15577 34731
rect 15577 34697 15611 34731
rect 15611 34697 15620 34731
rect 15568 34688 15620 34697
rect 16212 34731 16264 34740
rect 16212 34697 16221 34731
rect 16221 34697 16255 34731
rect 16255 34697 16264 34731
rect 16212 34688 16264 34697
rect 16304 34688 16356 34740
rect 2320 34663 2372 34672
rect 2320 34629 2329 34663
rect 2329 34629 2363 34663
rect 2363 34629 2372 34663
rect 2320 34620 2372 34629
rect 15292 34620 15344 34672
rect 4620 34552 4672 34604
rect 1492 34484 1544 34536
rect 2504 34484 2556 34536
rect 4988 34552 5040 34604
rect 5448 34595 5500 34604
rect 5080 34484 5132 34536
rect 5448 34561 5457 34595
rect 5457 34561 5491 34595
rect 5491 34561 5500 34595
rect 5448 34552 5500 34561
rect 6184 34552 6236 34604
rect 5816 34484 5868 34536
rect 6368 34484 6420 34536
rect 6736 34527 6788 34536
rect 6736 34493 6745 34527
rect 6745 34493 6779 34527
rect 6779 34493 6788 34527
rect 6736 34484 6788 34493
rect 14648 34552 14700 34604
rect 14924 34552 14976 34604
rect 7932 34527 7984 34536
rect 7932 34493 7941 34527
rect 7941 34493 7975 34527
rect 7975 34493 7984 34527
rect 7932 34484 7984 34493
rect 8484 34527 8536 34536
rect 8484 34493 8493 34527
rect 8493 34493 8527 34527
rect 8527 34493 8536 34527
rect 8484 34484 8536 34493
rect 8944 34484 8996 34536
rect 9772 34484 9824 34536
rect 13636 34484 13688 34536
rect 14740 34484 14792 34536
rect 17500 34663 17552 34672
rect 16856 34595 16908 34604
rect 16856 34561 16865 34595
rect 16865 34561 16899 34595
rect 16899 34561 16908 34595
rect 16856 34552 16908 34561
rect 17500 34629 17509 34663
rect 17509 34629 17543 34663
rect 17543 34629 17552 34663
rect 17500 34620 17552 34629
rect 17408 34484 17460 34536
rect 6828 34416 6880 34468
rect 8300 34416 8352 34468
rect 8576 34416 8628 34468
rect 7472 34348 7524 34400
rect 7648 34246 7700 34298
rect 7712 34246 7764 34298
rect 7776 34246 7828 34298
rect 7840 34246 7892 34298
rect 14315 34246 14367 34298
rect 14379 34246 14431 34298
rect 14443 34246 14495 34298
rect 14507 34246 14559 34298
rect 6920 34144 6972 34196
rect 14832 34144 14884 34196
rect 15660 34144 15712 34196
rect 16856 34144 16908 34196
rect 6368 34119 6420 34128
rect 6368 34085 6377 34119
rect 6377 34085 6411 34119
rect 6411 34085 6420 34119
rect 6368 34076 6420 34085
rect 16304 34076 16356 34128
rect 3516 34051 3568 34060
rect 3516 34017 3525 34051
rect 3525 34017 3559 34051
rect 3559 34017 3568 34051
rect 3516 34008 3568 34017
rect 6828 34051 6880 34060
rect 6828 34017 6837 34051
rect 6837 34017 6871 34051
rect 6871 34017 6880 34051
rect 6828 34008 6880 34017
rect 7288 34008 7340 34060
rect 7472 34008 7524 34060
rect 9588 34051 9640 34060
rect 9588 34017 9597 34051
rect 9597 34017 9631 34051
rect 9631 34017 9640 34051
rect 9588 34008 9640 34017
rect 9680 34051 9732 34060
rect 9680 34017 9689 34051
rect 9689 34017 9723 34051
rect 9723 34017 9732 34051
rect 10048 34051 10100 34060
rect 9680 34008 9732 34017
rect 10048 34017 10057 34051
rect 10057 34017 10091 34051
rect 10091 34017 10100 34051
rect 10048 34008 10100 34017
rect 10232 34008 10284 34060
rect 14188 34051 14240 34060
rect 14188 34017 14197 34051
rect 14197 34017 14231 34051
rect 14231 34017 14240 34051
rect 14188 34008 14240 34017
rect 14832 34051 14884 34060
rect 14832 34017 14841 34051
rect 14841 34017 14875 34051
rect 14875 34017 14884 34051
rect 14832 34008 14884 34017
rect 15844 34008 15896 34060
rect 16488 34051 16540 34060
rect 16488 34017 16497 34051
rect 16497 34017 16531 34051
rect 16531 34017 16540 34051
rect 16488 34008 16540 34017
rect 3240 33983 3292 33992
rect 3240 33949 3249 33983
rect 3249 33949 3283 33983
rect 3283 33949 3292 33983
rect 3240 33940 3292 33949
rect 4896 33983 4948 33992
rect 4896 33949 4905 33983
rect 4905 33949 4939 33983
rect 4939 33949 4948 33983
rect 4896 33940 4948 33949
rect 9128 33940 9180 33992
rect 14924 33983 14976 33992
rect 6736 33872 6788 33924
rect 9680 33872 9732 33924
rect 14924 33949 14933 33983
rect 14933 33949 14967 33983
rect 14967 33949 14976 33983
rect 14924 33940 14976 33949
rect 16212 33983 16264 33992
rect 16212 33949 16221 33983
rect 16221 33949 16255 33983
rect 16255 33949 16264 33983
rect 16212 33940 16264 33949
rect 17132 33983 17184 33992
rect 17132 33949 17141 33983
rect 17141 33949 17175 33983
rect 17175 33949 17184 33983
rect 17132 33940 17184 33949
rect 4315 33702 4367 33754
rect 4379 33702 4431 33754
rect 4443 33702 4495 33754
rect 4507 33702 4559 33754
rect 10982 33702 11034 33754
rect 11046 33702 11098 33754
rect 11110 33702 11162 33754
rect 11174 33702 11226 33754
rect 17648 33702 17700 33754
rect 17712 33702 17764 33754
rect 17776 33702 17828 33754
rect 17840 33702 17892 33754
rect 2596 33600 2648 33652
rect 3516 33600 3568 33652
rect 5632 33600 5684 33652
rect 6000 33600 6052 33652
rect 6828 33600 6880 33652
rect 8300 33643 8352 33652
rect 8300 33609 8309 33643
rect 8309 33609 8343 33643
rect 8343 33609 8352 33643
rect 8300 33600 8352 33609
rect 8760 33600 8812 33652
rect 9128 33600 9180 33652
rect 10048 33600 10100 33652
rect 1676 33532 1728 33584
rect 5632 33464 5684 33516
rect 2780 33396 2832 33448
rect 3976 33396 4028 33448
rect 2688 33328 2740 33380
rect 3240 33328 3292 33380
rect 1768 33260 1820 33312
rect 3792 33303 3844 33312
rect 3792 33269 3801 33303
rect 3801 33269 3835 33303
rect 3835 33269 3844 33303
rect 6552 33439 6604 33448
rect 6552 33405 6561 33439
rect 6561 33405 6595 33439
rect 6595 33405 6604 33439
rect 6552 33396 6604 33405
rect 10508 33600 10560 33652
rect 14832 33643 14884 33652
rect 14832 33609 14841 33643
rect 14841 33609 14875 33643
rect 14875 33609 14884 33643
rect 14832 33600 14884 33609
rect 15568 33643 15620 33652
rect 15568 33609 15577 33643
rect 15577 33609 15611 33643
rect 15611 33609 15620 33643
rect 15568 33600 15620 33609
rect 15844 33643 15896 33652
rect 15844 33609 15853 33643
rect 15853 33609 15887 33643
rect 15887 33609 15896 33643
rect 15844 33600 15896 33609
rect 17500 33575 17552 33584
rect 17500 33541 17509 33575
rect 17509 33541 17543 33575
rect 17543 33541 17552 33575
rect 17500 33532 17552 33541
rect 5724 33371 5776 33380
rect 5724 33337 5733 33371
rect 5733 33337 5767 33371
rect 5767 33337 5776 33371
rect 5724 33328 5776 33337
rect 5816 33328 5868 33380
rect 3792 33260 3844 33269
rect 6920 33260 6972 33312
rect 15568 33396 15620 33448
rect 17040 33439 17092 33448
rect 9588 33328 9640 33380
rect 9956 33260 10008 33312
rect 14096 33303 14148 33312
rect 14096 33269 14105 33303
rect 14105 33269 14139 33303
rect 14139 33269 14148 33303
rect 14096 33260 14148 33269
rect 14188 33260 14240 33312
rect 14832 33260 14884 33312
rect 15936 33260 15988 33312
rect 16212 33303 16264 33312
rect 16212 33269 16221 33303
rect 16221 33269 16255 33303
rect 16255 33269 16264 33303
rect 16212 33260 16264 33269
rect 16580 33303 16632 33312
rect 16580 33269 16589 33303
rect 16589 33269 16623 33303
rect 16623 33269 16632 33303
rect 17040 33405 17049 33439
rect 17049 33405 17083 33439
rect 17083 33405 17092 33439
rect 17040 33396 17092 33405
rect 18052 33303 18104 33312
rect 16580 33260 16632 33269
rect 18052 33269 18061 33303
rect 18061 33269 18095 33303
rect 18095 33269 18104 33303
rect 18052 33260 18104 33269
rect 7648 33158 7700 33210
rect 7712 33158 7764 33210
rect 7776 33158 7828 33210
rect 7840 33158 7892 33210
rect 14315 33158 14367 33210
rect 14379 33158 14431 33210
rect 14443 33158 14495 33210
rect 14507 33158 14559 33210
rect 2964 33099 3016 33108
rect 2964 33065 2973 33099
rect 2973 33065 3007 33099
rect 3007 33065 3016 33099
rect 2964 33056 3016 33065
rect 6552 33056 6604 33108
rect 4712 32963 4764 32972
rect 4712 32929 4721 32963
rect 4721 32929 4755 32963
rect 4755 32929 4764 32963
rect 4712 32920 4764 32929
rect 5816 32988 5868 33040
rect 1400 32895 1452 32904
rect 1400 32861 1409 32895
rect 1409 32861 1443 32895
rect 1443 32861 1452 32895
rect 1400 32852 1452 32861
rect 1860 32852 1912 32904
rect 4160 32852 4212 32904
rect 6368 32920 6420 32972
rect 6828 33056 6880 33108
rect 7288 33056 7340 33108
rect 7472 33099 7524 33108
rect 7472 33065 7481 33099
rect 7481 33065 7515 33099
rect 7515 33065 7524 33099
rect 7472 33056 7524 33065
rect 15200 33056 15252 33108
rect 15844 33099 15896 33108
rect 15844 33065 15853 33099
rect 15853 33065 15887 33099
rect 15887 33065 15896 33099
rect 15844 33056 15896 33065
rect 9128 32988 9180 33040
rect 9864 32988 9916 33040
rect 9588 32963 9640 32972
rect 9588 32929 9597 32963
rect 9597 32929 9631 32963
rect 9631 32929 9640 32963
rect 9588 32920 9640 32929
rect 10324 32988 10376 33040
rect 14096 32988 14148 33040
rect 5356 32852 5408 32904
rect 5632 32852 5684 32904
rect 9864 32895 9916 32904
rect 9864 32861 9873 32895
rect 9873 32861 9907 32895
rect 9907 32861 9916 32895
rect 9864 32852 9916 32861
rect 9312 32784 9364 32836
rect 10232 32920 10284 32972
rect 13636 32920 13688 32972
rect 14188 32920 14240 32972
rect 14648 32963 14700 32972
rect 14648 32929 14657 32963
rect 14657 32929 14691 32963
rect 14691 32929 14700 32963
rect 14648 32920 14700 32929
rect 14924 32988 14976 33040
rect 17132 33031 17184 33040
rect 15752 32920 15804 32972
rect 17132 32997 17141 33031
rect 17141 32997 17175 33031
rect 17175 32997 17184 33031
rect 17132 32988 17184 32997
rect 17408 33031 17460 33040
rect 17408 32997 17417 33031
rect 17417 32997 17451 33031
rect 17451 32997 17460 33031
rect 17408 32988 17460 32997
rect 16304 32852 16356 32904
rect 18420 32852 18472 32904
rect 13912 32784 13964 32836
rect 14188 32784 14240 32836
rect 15936 32784 15988 32836
rect 3516 32716 3568 32768
rect 9128 32759 9180 32768
rect 9128 32725 9137 32759
rect 9137 32725 9171 32759
rect 9171 32725 9180 32759
rect 9128 32716 9180 32725
rect 9772 32716 9824 32768
rect 9956 32716 10008 32768
rect 10232 32716 10284 32768
rect 11336 32716 11388 32768
rect 4315 32614 4367 32666
rect 4379 32614 4431 32666
rect 4443 32614 4495 32666
rect 4507 32614 4559 32666
rect 10982 32614 11034 32666
rect 11046 32614 11098 32666
rect 11110 32614 11162 32666
rect 11174 32614 11226 32666
rect 17648 32614 17700 32666
rect 17712 32614 17764 32666
rect 17776 32614 17828 32666
rect 17840 32614 17892 32666
rect 2872 32555 2924 32564
rect 2872 32521 2881 32555
rect 2881 32521 2915 32555
rect 2915 32521 2924 32555
rect 2872 32512 2924 32521
rect 3516 32555 3568 32564
rect 3516 32521 3525 32555
rect 3525 32521 3559 32555
rect 3559 32521 3568 32555
rect 3516 32512 3568 32521
rect 5080 32555 5132 32564
rect 5080 32521 5089 32555
rect 5089 32521 5123 32555
rect 5123 32521 5132 32555
rect 5080 32512 5132 32521
rect 8024 32555 8076 32564
rect 8024 32521 8033 32555
rect 8033 32521 8067 32555
rect 8067 32521 8076 32555
rect 8024 32512 8076 32521
rect 8300 32512 8352 32564
rect 8576 32512 8628 32564
rect 10324 32512 10376 32564
rect 14648 32512 14700 32564
rect 15752 32512 15804 32564
rect 18420 32555 18472 32564
rect 18420 32521 18429 32555
rect 18429 32521 18463 32555
rect 18463 32521 18472 32555
rect 18420 32512 18472 32521
rect 8484 32444 8536 32496
rect 8852 32444 8904 32496
rect 9312 32487 9364 32496
rect 9312 32453 9321 32487
rect 9321 32453 9355 32487
rect 9355 32453 9364 32487
rect 9312 32444 9364 32453
rect 1768 32419 1820 32428
rect 1768 32385 1777 32419
rect 1777 32385 1811 32419
rect 1811 32385 1820 32419
rect 1768 32376 1820 32385
rect 5632 32376 5684 32428
rect 11060 32419 11112 32428
rect 1400 32308 1452 32360
rect 2688 32308 2740 32360
rect 4988 32351 5040 32360
rect 4988 32317 4997 32351
rect 4997 32317 5031 32351
rect 5031 32317 5040 32351
rect 4988 32308 5040 32317
rect 5356 32351 5408 32360
rect 5356 32317 5365 32351
rect 5365 32317 5399 32351
rect 5399 32317 5408 32351
rect 5356 32308 5408 32317
rect 5816 32351 5868 32360
rect 5816 32317 5825 32351
rect 5825 32317 5859 32351
rect 5859 32317 5868 32351
rect 5816 32308 5868 32317
rect 6368 32351 6420 32360
rect 6368 32317 6377 32351
rect 6377 32317 6411 32351
rect 6411 32317 6420 32351
rect 6368 32308 6420 32317
rect 8024 32308 8076 32360
rect 9128 32308 9180 32360
rect 9312 32308 9364 32360
rect 10232 32308 10284 32360
rect 11060 32385 11069 32419
rect 11069 32385 11103 32419
rect 11103 32385 11112 32419
rect 11060 32376 11112 32385
rect 11888 32376 11940 32428
rect 10324 32240 10376 32292
rect 11704 32308 11756 32360
rect 15200 32308 15252 32360
rect 15384 32308 15436 32360
rect 2688 32172 2740 32224
rect 3516 32172 3568 32224
rect 11336 32172 11388 32224
rect 13268 32240 13320 32292
rect 14096 32240 14148 32292
rect 15292 32283 15344 32292
rect 15292 32249 15301 32283
rect 15301 32249 15335 32283
rect 15335 32249 15344 32283
rect 15292 32240 15344 32249
rect 12900 32172 12952 32224
rect 13636 32215 13688 32224
rect 13636 32181 13645 32215
rect 13645 32181 13679 32215
rect 13679 32181 13688 32215
rect 13636 32172 13688 32181
rect 15568 32215 15620 32224
rect 15568 32181 15577 32215
rect 15577 32181 15611 32215
rect 15611 32181 15620 32215
rect 15568 32172 15620 32181
rect 16580 32215 16632 32224
rect 16580 32181 16589 32215
rect 16589 32181 16623 32215
rect 16623 32181 16632 32215
rect 17408 32308 17460 32360
rect 18052 32351 18104 32360
rect 16856 32240 16908 32292
rect 18052 32317 18061 32351
rect 18061 32317 18095 32351
rect 18095 32317 18104 32351
rect 18052 32308 18104 32317
rect 17776 32283 17828 32292
rect 17776 32249 17785 32283
rect 17785 32249 17819 32283
rect 17819 32249 17828 32283
rect 17776 32240 17828 32249
rect 16580 32172 16632 32181
rect 17408 32172 17460 32224
rect 17960 32172 18012 32224
rect 7648 32070 7700 32122
rect 7712 32070 7764 32122
rect 7776 32070 7828 32122
rect 7840 32070 7892 32122
rect 14315 32070 14367 32122
rect 14379 32070 14431 32122
rect 14443 32070 14495 32122
rect 14507 32070 14559 32122
rect 3332 31968 3384 32020
rect 3516 31968 3568 32020
rect 5356 32011 5408 32020
rect 5356 31977 5365 32011
rect 5365 31977 5399 32011
rect 5399 31977 5408 32011
rect 5356 31968 5408 31977
rect 6644 31968 6696 32020
rect 7288 31968 7340 32020
rect 9588 31968 9640 32020
rect 9864 32011 9916 32020
rect 9864 31977 9873 32011
rect 9873 31977 9907 32011
rect 9907 31977 9916 32011
rect 9864 31968 9916 31977
rect 12624 32011 12676 32020
rect 12624 31977 12633 32011
rect 12633 31977 12667 32011
rect 12667 31977 12676 32011
rect 12624 31968 12676 31977
rect 15476 31968 15528 32020
rect 15752 31968 15804 32020
rect 3148 31943 3200 31952
rect 3148 31909 3157 31943
rect 3157 31909 3191 31943
rect 3191 31909 3200 31943
rect 3148 31900 3200 31909
rect 6368 31900 6420 31952
rect 15844 31900 15896 31952
rect 17500 31900 17552 31952
rect 1584 31832 1636 31884
rect 4988 31832 5040 31884
rect 5816 31875 5868 31884
rect 5816 31841 5825 31875
rect 5825 31841 5859 31875
rect 5859 31841 5868 31875
rect 5816 31832 5868 31841
rect 6000 31832 6052 31884
rect 8024 31832 8076 31884
rect 1492 31807 1544 31816
rect 1492 31773 1501 31807
rect 1501 31773 1535 31807
rect 1535 31773 1544 31807
rect 1492 31764 1544 31773
rect 7472 31764 7524 31816
rect 8760 31832 8812 31884
rect 10600 31832 10652 31884
rect 11060 31875 11112 31884
rect 11060 31841 11069 31875
rect 11069 31841 11103 31875
rect 11103 31841 11112 31875
rect 11060 31832 11112 31841
rect 11520 31832 11572 31884
rect 12440 31875 12492 31884
rect 12440 31841 12449 31875
rect 12449 31841 12483 31875
rect 12483 31841 12492 31875
rect 12440 31832 12492 31841
rect 13728 31832 13780 31884
rect 14556 31875 14608 31884
rect 14556 31841 14565 31875
rect 14565 31841 14599 31875
rect 14599 31841 14608 31875
rect 14556 31832 14608 31841
rect 14648 31875 14700 31884
rect 14648 31841 14657 31875
rect 14657 31841 14691 31875
rect 14691 31841 14700 31875
rect 14832 31875 14884 31884
rect 14648 31832 14700 31841
rect 14832 31841 14841 31875
rect 14841 31841 14875 31875
rect 14875 31841 14884 31875
rect 14832 31832 14884 31841
rect 16304 31875 16356 31884
rect 16304 31841 16313 31875
rect 16313 31841 16347 31875
rect 16347 31841 16356 31875
rect 16304 31832 16356 31841
rect 8852 31764 8904 31816
rect 3332 31696 3384 31748
rect 4068 31696 4120 31748
rect 9864 31696 9916 31748
rect 10692 31696 10744 31748
rect 15936 31764 15988 31816
rect 17316 31764 17368 31816
rect 10876 31628 10928 31680
rect 11336 31628 11388 31680
rect 4315 31526 4367 31578
rect 4379 31526 4431 31578
rect 4443 31526 4495 31578
rect 4507 31526 4559 31578
rect 10982 31526 11034 31578
rect 11046 31526 11098 31578
rect 11110 31526 11162 31578
rect 11174 31526 11226 31578
rect 17648 31526 17700 31578
rect 17712 31526 17764 31578
rect 17776 31526 17828 31578
rect 17840 31526 17892 31578
rect 1860 31424 1912 31476
rect 6000 31424 6052 31476
rect 6552 31424 6604 31476
rect 7472 31467 7524 31476
rect 7472 31433 7481 31467
rect 7481 31433 7515 31467
rect 7515 31433 7524 31467
rect 7472 31424 7524 31433
rect 8760 31424 8812 31476
rect 14648 31424 14700 31476
rect 15936 31424 15988 31476
rect 1492 31356 1544 31408
rect 8024 31356 8076 31408
rect 14832 31356 14884 31408
rect 2136 31220 2188 31272
rect 2320 31220 2372 31272
rect 6276 31263 6328 31272
rect 1584 31195 1636 31204
rect 1584 31161 1593 31195
rect 1593 31161 1627 31195
rect 1627 31161 1636 31195
rect 1584 31152 1636 31161
rect 6000 31084 6052 31136
rect 6276 31229 6285 31263
rect 6285 31229 6319 31263
rect 6319 31229 6328 31263
rect 6276 31220 6328 31229
rect 7932 31220 7984 31272
rect 9496 31263 9548 31272
rect 7472 31152 7524 31204
rect 9496 31229 9505 31263
rect 9505 31229 9539 31263
rect 9539 31229 9548 31263
rect 9496 31220 9548 31229
rect 9864 31263 9916 31272
rect 9864 31229 9873 31263
rect 9873 31229 9907 31263
rect 9907 31229 9916 31263
rect 9864 31220 9916 31229
rect 9956 31220 10008 31272
rect 10784 31288 10836 31340
rect 15292 31288 15344 31340
rect 15844 31331 15896 31340
rect 15844 31297 15853 31331
rect 15853 31297 15887 31331
rect 15887 31297 15896 31331
rect 15844 31288 15896 31297
rect 11336 31220 11388 31272
rect 9956 31127 10008 31136
rect 9956 31093 9965 31127
rect 9965 31093 9999 31127
rect 9999 31093 10008 31127
rect 9956 31084 10008 31093
rect 11060 31084 11112 31136
rect 12440 31152 12492 31204
rect 15384 31220 15436 31272
rect 16120 31220 16172 31272
rect 16580 31220 16632 31272
rect 17316 31220 17368 31272
rect 17500 31263 17552 31272
rect 17500 31229 17509 31263
rect 17509 31229 17543 31263
rect 17543 31229 17552 31263
rect 17500 31220 17552 31229
rect 12072 31127 12124 31136
rect 12072 31093 12081 31127
rect 12081 31093 12115 31127
rect 12115 31093 12124 31127
rect 12072 31084 12124 31093
rect 14648 31127 14700 31136
rect 14648 31093 14657 31127
rect 14657 31093 14691 31127
rect 14691 31093 14700 31127
rect 14648 31084 14700 31093
rect 15844 31152 15896 31204
rect 17776 31195 17828 31204
rect 17776 31161 17785 31195
rect 17785 31161 17819 31195
rect 17819 31161 17828 31195
rect 17776 31152 17828 31161
rect 16120 31127 16172 31136
rect 16120 31093 16129 31127
rect 16129 31093 16163 31127
rect 16163 31093 16172 31127
rect 16120 31084 16172 31093
rect 7648 30982 7700 31034
rect 7712 30982 7764 31034
rect 7776 30982 7828 31034
rect 7840 30982 7892 31034
rect 14315 30982 14367 31034
rect 14379 30982 14431 31034
rect 14443 30982 14495 31034
rect 14507 30982 14559 31034
rect 3424 30812 3476 30864
rect 1768 30744 1820 30796
rect 6552 30880 6604 30932
rect 8024 30923 8076 30932
rect 8024 30889 8033 30923
rect 8033 30889 8067 30923
rect 8067 30889 8076 30923
rect 8024 30880 8076 30889
rect 9864 30923 9916 30932
rect 9864 30889 9873 30923
rect 9873 30889 9907 30923
rect 9907 30889 9916 30923
rect 9864 30880 9916 30889
rect 10600 30923 10652 30932
rect 10600 30889 10609 30923
rect 10609 30889 10643 30923
rect 10643 30889 10652 30923
rect 10600 30880 10652 30889
rect 15568 30880 15620 30932
rect 16304 30923 16356 30932
rect 16304 30889 16313 30923
rect 16313 30889 16347 30923
rect 16347 30889 16356 30923
rect 16304 30880 16356 30889
rect 16948 30880 17000 30932
rect 6184 30812 6236 30864
rect 10692 30812 10744 30864
rect 11336 30812 11388 30864
rect 5632 30787 5684 30796
rect 5632 30753 5641 30787
rect 5641 30753 5675 30787
rect 5675 30753 5684 30787
rect 5632 30744 5684 30753
rect 15752 30812 15804 30864
rect 16856 30855 16908 30864
rect 16856 30821 16865 30855
rect 16865 30821 16899 30855
rect 16899 30821 16908 30855
rect 16856 30812 16908 30821
rect 2136 30676 2188 30728
rect 2688 30676 2740 30728
rect 4988 30719 5040 30728
rect 4988 30685 4997 30719
rect 4997 30685 5031 30719
rect 5031 30685 5040 30719
rect 4988 30676 5040 30685
rect 15476 30676 15528 30728
rect 15936 30676 15988 30728
rect 11336 30608 11388 30660
rect 11612 30608 11664 30660
rect 15384 30651 15436 30660
rect 15384 30617 15393 30651
rect 15393 30617 15427 30651
rect 15427 30617 15436 30651
rect 15384 30608 15436 30617
rect 16488 30608 16540 30660
rect 16856 30608 16908 30660
rect 7656 30583 7708 30592
rect 7656 30549 7665 30583
rect 7665 30549 7699 30583
rect 7699 30549 7708 30583
rect 7656 30540 7708 30549
rect 12716 30583 12768 30592
rect 12716 30549 12725 30583
rect 12725 30549 12759 30583
rect 12759 30549 12768 30583
rect 12716 30540 12768 30549
rect 15200 30540 15252 30592
rect 16580 30540 16632 30592
rect 4315 30438 4367 30490
rect 4379 30438 4431 30490
rect 4443 30438 4495 30490
rect 4507 30438 4559 30490
rect 10982 30438 11034 30490
rect 11046 30438 11098 30490
rect 11110 30438 11162 30490
rect 11174 30438 11226 30490
rect 17648 30438 17700 30490
rect 17712 30438 17764 30490
rect 17776 30438 17828 30490
rect 17840 30438 17892 30490
rect 4988 30336 5040 30388
rect 6920 30268 6972 30320
rect 12900 30311 12952 30320
rect 12900 30277 12909 30311
rect 12909 30277 12943 30311
rect 12943 30277 12952 30311
rect 12900 30268 12952 30277
rect 15476 30336 15528 30388
rect 16304 30336 16356 30388
rect 15108 30311 15160 30320
rect 15108 30277 15117 30311
rect 15117 30277 15151 30311
rect 15151 30277 15160 30311
rect 15108 30268 15160 30277
rect 15844 30311 15896 30320
rect 15844 30277 15853 30311
rect 15853 30277 15887 30311
rect 15887 30277 15896 30311
rect 15844 30268 15896 30277
rect 15936 30268 15988 30320
rect 4436 30200 4488 30252
rect 5632 30200 5684 30252
rect 8944 30200 8996 30252
rect 17868 30200 17920 30252
rect 4896 30132 4948 30184
rect 5356 30132 5408 30184
rect 5448 30175 5500 30184
rect 5448 30141 5457 30175
rect 5457 30141 5491 30175
rect 5491 30141 5500 30175
rect 5448 30132 5500 30141
rect 5724 30132 5776 30184
rect 5908 30132 5960 30184
rect 6920 30132 6972 30184
rect 7196 30132 7248 30184
rect 8392 30175 8444 30184
rect 1676 30039 1728 30048
rect 1676 30005 1685 30039
rect 1685 30005 1719 30039
rect 1719 30005 1728 30039
rect 1676 29996 1728 30005
rect 2136 30039 2188 30048
rect 2136 30005 2145 30039
rect 2145 30005 2179 30039
rect 2179 30005 2188 30039
rect 2136 29996 2188 30005
rect 6552 29996 6604 30048
rect 8392 30141 8401 30175
rect 8401 30141 8435 30175
rect 8435 30141 8444 30175
rect 8392 30132 8444 30141
rect 8760 30132 8812 30184
rect 9128 30132 9180 30184
rect 10508 30132 10560 30184
rect 12716 30132 12768 30184
rect 13176 30132 13228 30184
rect 8300 29996 8352 30048
rect 12072 30039 12124 30048
rect 12072 30005 12081 30039
rect 12081 30005 12115 30039
rect 12115 30005 12124 30039
rect 12072 29996 12124 30005
rect 12532 30039 12584 30048
rect 12532 30005 12541 30039
rect 12541 30005 12575 30039
rect 12575 30005 12584 30039
rect 15200 30132 15252 30184
rect 16120 30175 16172 30184
rect 16120 30141 16129 30175
rect 16129 30141 16163 30175
rect 16163 30141 16172 30175
rect 16120 30132 16172 30141
rect 16580 30132 16632 30184
rect 16948 30132 17000 30184
rect 17500 30175 17552 30184
rect 17500 30141 17509 30175
rect 17509 30141 17543 30175
rect 17543 30141 17552 30175
rect 17500 30132 17552 30141
rect 12532 29996 12584 30005
rect 7648 29894 7700 29946
rect 7712 29894 7764 29946
rect 7776 29894 7828 29946
rect 7840 29894 7892 29946
rect 14315 29894 14367 29946
rect 14379 29894 14431 29946
rect 14443 29894 14495 29946
rect 14507 29894 14559 29946
rect 2044 29792 2096 29844
rect 4528 29835 4580 29844
rect 4528 29801 4537 29835
rect 4537 29801 4571 29835
rect 4571 29801 4580 29835
rect 4528 29792 4580 29801
rect 5724 29792 5776 29844
rect 13268 29792 13320 29844
rect 15292 29835 15344 29844
rect 15292 29801 15301 29835
rect 15301 29801 15335 29835
rect 15335 29801 15344 29835
rect 15292 29792 15344 29801
rect 16028 29792 16080 29844
rect 17132 29835 17184 29844
rect 17132 29801 17141 29835
rect 17141 29801 17175 29835
rect 17175 29801 17184 29835
rect 17132 29792 17184 29801
rect 3700 29767 3752 29776
rect 3700 29733 3709 29767
rect 3709 29733 3743 29767
rect 3743 29733 3752 29767
rect 3700 29724 3752 29733
rect 4436 29767 4488 29776
rect 4436 29733 4445 29767
rect 4445 29733 4479 29767
rect 4479 29733 4488 29767
rect 4436 29724 4488 29733
rect 5632 29724 5684 29776
rect 5908 29767 5960 29776
rect 5908 29733 5917 29767
rect 5917 29733 5951 29767
rect 5951 29733 5960 29767
rect 5908 29724 5960 29733
rect 1492 29656 1544 29708
rect 2136 29656 2188 29708
rect 4712 29699 4764 29708
rect 4712 29665 4721 29699
rect 4721 29665 4755 29699
rect 4755 29665 4764 29699
rect 4712 29656 4764 29665
rect 6828 29699 6880 29708
rect 6828 29665 6837 29699
rect 6837 29665 6871 29699
rect 6871 29665 6880 29699
rect 6828 29656 6880 29665
rect 8300 29699 8352 29708
rect 8300 29665 8309 29699
rect 8309 29665 8343 29699
rect 8343 29665 8352 29699
rect 8300 29656 8352 29665
rect 9128 29699 9180 29708
rect 9128 29665 9137 29699
rect 9137 29665 9171 29699
rect 9171 29665 9180 29699
rect 9128 29656 9180 29665
rect 9496 29656 9548 29708
rect 10140 29656 10192 29708
rect 10232 29656 10284 29708
rect 10968 29656 11020 29708
rect 8392 29588 8444 29640
rect 12624 29588 12676 29640
rect 12440 29520 12492 29572
rect 14372 29699 14424 29708
rect 14372 29665 14381 29699
rect 14381 29665 14415 29699
rect 14415 29665 14424 29699
rect 14372 29656 14424 29665
rect 16304 29656 16356 29708
rect 13176 29631 13228 29640
rect 13176 29597 13185 29631
rect 13185 29597 13219 29631
rect 13219 29597 13228 29631
rect 13176 29588 13228 29597
rect 15936 29588 15988 29640
rect 9404 29495 9456 29504
rect 9404 29461 9413 29495
rect 9413 29461 9447 29495
rect 9447 29461 9456 29495
rect 10692 29495 10744 29504
rect 9404 29452 9456 29461
rect 10692 29461 10701 29495
rect 10701 29461 10735 29495
rect 10735 29461 10744 29495
rect 10692 29452 10744 29461
rect 12256 29495 12308 29504
rect 12256 29461 12265 29495
rect 12265 29461 12299 29495
rect 12299 29461 12308 29495
rect 12256 29452 12308 29461
rect 13636 29452 13688 29504
rect 16212 29495 16264 29504
rect 16212 29461 16221 29495
rect 16221 29461 16255 29495
rect 16255 29461 16264 29495
rect 16212 29452 16264 29461
rect 16580 29452 16632 29504
rect 17500 29495 17552 29504
rect 17500 29461 17509 29495
rect 17509 29461 17543 29495
rect 17543 29461 17552 29495
rect 17500 29452 17552 29461
rect 4315 29350 4367 29402
rect 4379 29350 4431 29402
rect 4443 29350 4495 29402
rect 4507 29350 4559 29402
rect 10982 29350 11034 29402
rect 11046 29350 11098 29402
rect 11110 29350 11162 29402
rect 11174 29350 11226 29402
rect 17648 29350 17700 29402
rect 17712 29350 17764 29402
rect 17776 29350 17828 29402
rect 17840 29350 17892 29402
rect 7196 29248 7248 29300
rect 9496 29291 9548 29300
rect 1492 29155 1544 29164
rect 1492 29121 1501 29155
rect 1501 29121 1535 29155
rect 1535 29121 1544 29155
rect 1492 29112 1544 29121
rect 2596 29112 2648 29164
rect 5724 29112 5776 29164
rect 6184 29112 6236 29164
rect 6828 29155 6880 29164
rect 6828 29121 6837 29155
rect 6837 29121 6871 29155
rect 6871 29121 6880 29155
rect 6828 29112 6880 29121
rect 9496 29257 9505 29291
rect 9505 29257 9539 29291
rect 9539 29257 9548 29291
rect 9496 29248 9548 29257
rect 10232 29248 10284 29300
rect 10876 29248 10928 29300
rect 14372 29291 14424 29300
rect 14372 29257 14381 29291
rect 14381 29257 14415 29291
rect 14415 29257 14424 29291
rect 14372 29248 14424 29257
rect 15936 29248 15988 29300
rect 2044 29044 2096 29096
rect 3148 29019 3200 29028
rect 3148 28985 3157 29019
rect 3157 28985 3191 29019
rect 3191 28985 3200 29019
rect 3148 28976 3200 28985
rect 4896 28976 4948 29028
rect 5632 29019 5684 29028
rect 5632 28985 5641 29019
rect 5641 28985 5675 29019
rect 5675 28985 5684 29019
rect 5632 28976 5684 28985
rect 6368 29044 6420 29096
rect 12256 29112 12308 29164
rect 14648 29112 14700 29164
rect 8392 29044 8444 29096
rect 3424 28951 3476 28960
rect 3424 28917 3433 28951
rect 3433 28917 3467 28951
rect 3467 28917 3476 28951
rect 3424 28908 3476 28917
rect 5908 28976 5960 29028
rect 6552 28976 6604 29028
rect 9496 29044 9548 29096
rect 10140 29044 10192 29096
rect 12624 29087 12676 29096
rect 12624 29053 12633 29087
rect 12633 29053 12667 29087
rect 12667 29053 12676 29087
rect 12624 29044 12676 29053
rect 13636 29087 13688 29096
rect 11796 29019 11848 29028
rect 8024 28908 8076 28960
rect 8116 28908 8168 28960
rect 11796 28985 11805 29019
rect 11805 28985 11839 29019
rect 11839 28985 11848 29019
rect 13636 29053 13645 29087
rect 13645 29053 13679 29087
rect 13679 29053 13688 29087
rect 13636 29044 13688 29053
rect 15384 29087 15436 29096
rect 15384 29053 15393 29087
rect 15393 29053 15427 29087
rect 15427 29053 15436 29087
rect 15384 29044 15436 29053
rect 17132 29087 17184 29096
rect 15844 29019 15896 29028
rect 11796 28976 11848 28985
rect 15844 28985 15853 29019
rect 15853 28985 15887 29019
rect 15887 28985 15896 29019
rect 15844 28976 15896 28985
rect 12072 28908 12124 28960
rect 12624 28908 12676 28960
rect 16580 28951 16632 28960
rect 16580 28917 16589 28951
rect 16589 28917 16623 28951
rect 16623 28917 16632 28951
rect 17132 29053 17141 29087
rect 17141 29053 17175 29087
rect 17175 29053 17184 29087
rect 17132 29044 17184 29053
rect 17500 29087 17552 29096
rect 17500 29053 17509 29087
rect 17509 29053 17543 29087
rect 17543 29053 17552 29087
rect 17500 29044 17552 29053
rect 17776 29087 17828 29096
rect 17776 29053 17785 29087
rect 17785 29053 17819 29087
rect 17819 29053 17828 29087
rect 17776 29044 17828 29053
rect 16580 28908 16632 28917
rect 7648 28806 7700 28858
rect 7712 28806 7764 28858
rect 7776 28806 7828 28858
rect 7840 28806 7892 28858
rect 14315 28806 14367 28858
rect 14379 28806 14431 28858
rect 14443 28806 14495 28858
rect 14507 28806 14559 28858
rect 2136 28704 2188 28756
rect 2596 28747 2648 28756
rect 2596 28713 2605 28747
rect 2605 28713 2639 28747
rect 2639 28713 2648 28747
rect 3424 28747 3476 28756
rect 2596 28704 2648 28713
rect 3424 28713 3433 28747
rect 3433 28713 3467 28747
rect 3467 28713 3476 28747
rect 3424 28704 3476 28713
rect 6736 28704 6788 28756
rect 7104 28747 7156 28756
rect 7104 28713 7113 28747
rect 7113 28713 7147 28747
rect 7147 28713 7156 28747
rect 7104 28704 7156 28713
rect 8116 28704 8168 28756
rect 10416 28704 10468 28756
rect 12348 28704 12400 28756
rect 12716 28747 12768 28756
rect 12716 28713 12725 28747
rect 12725 28713 12759 28747
rect 12759 28713 12768 28747
rect 12716 28704 12768 28713
rect 13084 28704 13136 28756
rect 13912 28747 13964 28756
rect 13912 28713 13921 28747
rect 13921 28713 13955 28747
rect 13955 28713 13964 28747
rect 13912 28704 13964 28713
rect 14740 28704 14792 28756
rect 16028 28704 16080 28756
rect 1676 28636 1728 28688
rect 1584 28611 1636 28620
rect 1584 28577 1593 28611
rect 1593 28577 1627 28611
rect 1627 28577 1636 28611
rect 1584 28568 1636 28577
rect 3608 28611 3660 28620
rect 3608 28577 3617 28611
rect 3617 28577 3651 28611
rect 3651 28577 3660 28611
rect 3608 28568 3660 28577
rect 1952 28543 2004 28552
rect 1952 28509 1961 28543
rect 1961 28509 1995 28543
rect 1995 28509 2004 28543
rect 1952 28500 2004 28509
rect 4712 28568 4764 28620
rect 5264 28611 5316 28620
rect 5264 28577 5273 28611
rect 5273 28577 5307 28611
rect 5307 28577 5316 28611
rect 5264 28568 5316 28577
rect 5816 28568 5868 28620
rect 7012 28568 7064 28620
rect 8024 28611 8076 28620
rect 8024 28577 8033 28611
rect 8033 28577 8067 28611
rect 8067 28577 8076 28611
rect 8024 28568 8076 28577
rect 8668 28568 8720 28620
rect 8852 28611 8904 28620
rect 8852 28577 8861 28611
rect 8861 28577 8895 28611
rect 8895 28577 8904 28611
rect 8852 28568 8904 28577
rect 10140 28611 10192 28620
rect 10140 28577 10149 28611
rect 10149 28577 10183 28611
rect 10183 28577 10192 28611
rect 12624 28636 12676 28688
rect 13176 28636 13228 28688
rect 15108 28679 15160 28688
rect 15108 28645 15117 28679
rect 15117 28645 15151 28679
rect 15151 28645 15160 28679
rect 15108 28636 15160 28645
rect 16304 28636 16356 28688
rect 10140 28568 10192 28577
rect 12440 28611 12492 28620
rect 12440 28577 12449 28611
rect 12449 28577 12483 28611
rect 12483 28577 12492 28611
rect 12440 28568 12492 28577
rect 12072 28500 12124 28552
rect 14648 28611 14700 28620
rect 14648 28577 14657 28611
rect 14657 28577 14691 28611
rect 14691 28577 14700 28611
rect 14648 28568 14700 28577
rect 16304 28500 16356 28552
rect 16580 28704 16632 28756
rect 16672 28636 16724 28688
rect 17224 28636 17276 28688
rect 16580 28568 16632 28620
rect 17500 28568 17552 28620
rect 5724 28432 5776 28484
rect 8300 28432 8352 28484
rect 12532 28432 12584 28484
rect 12072 28364 12124 28416
rect 17408 28407 17460 28416
rect 17408 28373 17417 28407
rect 17417 28373 17451 28407
rect 17451 28373 17460 28407
rect 17408 28364 17460 28373
rect 4315 28262 4367 28314
rect 4379 28262 4431 28314
rect 4443 28262 4495 28314
rect 4507 28262 4559 28314
rect 10982 28262 11034 28314
rect 11046 28262 11098 28314
rect 11110 28262 11162 28314
rect 11174 28262 11226 28314
rect 17648 28262 17700 28314
rect 17712 28262 17764 28314
rect 17776 28262 17828 28314
rect 17840 28262 17892 28314
rect 1584 28160 1636 28212
rect 2596 28160 2648 28212
rect 3608 28160 3660 28212
rect 8024 28160 8076 28212
rect 8668 28160 8720 28212
rect 8852 28160 8904 28212
rect 9404 28203 9456 28212
rect 9404 28169 9413 28203
rect 9413 28169 9447 28203
rect 9447 28169 9456 28203
rect 9404 28160 9456 28169
rect 15936 28160 15988 28212
rect 1676 28067 1728 28076
rect 1676 28033 1685 28067
rect 1685 28033 1719 28067
rect 1719 28033 1728 28067
rect 1676 28024 1728 28033
rect 6736 28024 6788 28076
rect 8392 28092 8444 28144
rect 12348 28024 12400 28076
rect 4712 27999 4764 28008
rect 4712 27965 4721 27999
rect 4721 27965 4755 27999
rect 4755 27965 4764 27999
rect 4712 27956 4764 27965
rect 5908 27956 5960 28008
rect 6092 27956 6144 28008
rect 9036 27956 9088 28008
rect 11888 27999 11940 28008
rect 11888 27965 11897 27999
rect 11897 27965 11931 27999
rect 11931 27965 11940 27999
rect 11888 27956 11940 27965
rect 12440 27956 12492 28008
rect 12900 27999 12952 28008
rect 12900 27965 12909 27999
rect 12909 27965 12943 27999
rect 12943 27965 12952 27999
rect 12900 27956 12952 27965
rect 13360 28024 13412 28076
rect 13268 27956 13320 28008
rect 17776 28067 17828 28076
rect 17776 28033 17785 28067
rect 17785 28033 17819 28067
rect 17819 28033 17828 28067
rect 17776 28024 17828 28033
rect 13912 27999 13964 28008
rect 7472 27888 7524 27940
rect 13912 27965 13921 27999
rect 13921 27965 13955 27999
rect 13955 27965 13964 27999
rect 13912 27956 13964 27965
rect 15384 27999 15436 28008
rect 15384 27965 15393 27999
rect 15393 27965 15427 27999
rect 15427 27965 15436 27999
rect 15384 27956 15436 27965
rect 15844 27931 15896 27940
rect 15844 27897 15853 27931
rect 15853 27897 15887 27931
rect 15887 27897 15896 27931
rect 15844 27888 15896 27897
rect 16304 27888 16356 27940
rect 17316 27956 17368 28008
rect 17408 27956 17460 28008
rect 4344 27863 4396 27872
rect 4344 27829 4353 27863
rect 4353 27829 4387 27863
rect 4387 27829 4396 27863
rect 4344 27820 4396 27829
rect 5264 27863 5316 27872
rect 5264 27829 5273 27863
rect 5273 27829 5307 27863
rect 5307 27829 5316 27863
rect 5264 27820 5316 27829
rect 5632 27820 5684 27872
rect 9220 27820 9272 27872
rect 10140 27863 10192 27872
rect 10140 27829 10149 27863
rect 10149 27829 10183 27863
rect 10183 27829 10192 27863
rect 10140 27820 10192 27829
rect 12624 27820 12676 27872
rect 12992 27820 13044 27872
rect 13820 27820 13872 27872
rect 14648 27820 14700 27872
rect 7648 27718 7700 27770
rect 7712 27718 7764 27770
rect 7776 27718 7828 27770
rect 7840 27718 7892 27770
rect 14315 27718 14367 27770
rect 14379 27718 14431 27770
rect 14443 27718 14495 27770
rect 14507 27718 14559 27770
rect 5908 27616 5960 27668
rect 7012 27659 7064 27668
rect 7012 27625 7021 27659
rect 7021 27625 7055 27659
rect 7055 27625 7064 27659
rect 7012 27616 7064 27625
rect 4160 27548 4212 27600
rect 4344 27548 4396 27600
rect 5172 27548 5224 27600
rect 7104 27548 7156 27600
rect 2044 27480 2096 27532
rect 3516 27480 3568 27532
rect 4712 27523 4764 27532
rect 4712 27489 4721 27523
rect 4721 27489 4755 27523
rect 4755 27489 4764 27523
rect 4712 27480 4764 27489
rect 7932 27548 7984 27600
rect 8024 27523 8076 27532
rect 1676 27455 1728 27464
rect 1676 27421 1685 27455
rect 1685 27421 1719 27455
rect 1719 27421 1728 27455
rect 1676 27412 1728 27421
rect 2596 27412 2648 27464
rect 2780 27412 2832 27464
rect 8024 27489 8033 27523
rect 8033 27489 8067 27523
rect 8067 27489 8076 27523
rect 8300 27616 8352 27668
rect 8392 27659 8444 27668
rect 8392 27625 8401 27659
rect 8401 27625 8435 27659
rect 8435 27625 8444 27659
rect 8392 27616 8444 27625
rect 9036 27616 9088 27668
rect 11336 27616 11388 27668
rect 12900 27616 12952 27668
rect 15384 27659 15436 27668
rect 15384 27625 15393 27659
rect 15393 27625 15427 27659
rect 15427 27625 15436 27659
rect 15384 27616 15436 27625
rect 16304 27616 16356 27668
rect 16856 27616 16908 27668
rect 13268 27591 13320 27600
rect 13268 27557 13277 27591
rect 13277 27557 13311 27591
rect 13311 27557 13320 27591
rect 13268 27548 13320 27557
rect 16212 27548 16264 27600
rect 10324 27523 10376 27532
rect 8024 27480 8076 27489
rect 10324 27489 10333 27523
rect 10333 27489 10367 27523
rect 10367 27489 10376 27523
rect 10324 27480 10376 27489
rect 11336 27523 11388 27532
rect 11336 27489 11345 27523
rect 11345 27489 11379 27523
rect 11379 27489 11388 27523
rect 11336 27480 11388 27489
rect 12716 27523 12768 27532
rect 12716 27489 12725 27523
rect 12725 27489 12759 27523
rect 12759 27489 12768 27523
rect 12716 27480 12768 27489
rect 13820 27480 13872 27532
rect 14188 27480 14240 27532
rect 15016 27480 15068 27532
rect 17132 27548 17184 27600
rect 17592 27548 17644 27600
rect 14648 27455 14700 27464
rect 14648 27421 14657 27455
rect 14657 27421 14691 27455
rect 14691 27421 14700 27455
rect 14648 27412 14700 27421
rect 17408 27480 17460 27532
rect 17316 27412 17368 27464
rect 12716 27344 12768 27396
rect 16028 27344 16080 27396
rect 16488 27344 16540 27396
rect 16580 27344 16632 27396
rect 3424 27276 3476 27328
rect 6092 27319 6144 27328
rect 6092 27285 6101 27319
rect 6101 27285 6135 27319
rect 6135 27285 6144 27319
rect 6092 27276 6144 27285
rect 7380 27319 7432 27328
rect 7380 27285 7389 27319
rect 7389 27285 7423 27319
rect 7423 27285 7432 27319
rect 7380 27276 7432 27285
rect 8300 27276 8352 27328
rect 8760 27276 8812 27328
rect 10508 27319 10560 27328
rect 10508 27285 10517 27319
rect 10517 27285 10551 27319
rect 10551 27285 10560 27319
rect 10508 27276 10560 27285
rect 11888 27319 11940 27328
rect 11888 27285 11897 27319
rect 11897 27285 11931 27319
rect 11931 27285 11940 27319
rect 11888 27276 11940 27285
rect 13360 27276 13412 27328
rect 13912 27319 13964 27328
rect 13912 27285 13921 27319
rect 13921 27285 13955 27319
rect 13955 27285 13964 27319
rect 13912 27276 13964 27285
rect 4315 27174 4367 27226
rect 4379 27174 4431 27226
rect 4443 27174 4495 27226
rect 4507 27174 4559 27226
rect 10982 27174 11034 27226
rect 11046 27174 11098 27226
rect 11110 27174 11162 27226
rect 11174 27174 11226 27226
rect 17648 27174 17700 27226
rect 17712 27174 17764 27226
rect 17776 27174 17828 27226
rect 17840 27174 17892 27226
rect 2044 27072 2096 27124
rect 3516 27115 3568 27124
rect 3516 27081 3525 27115
rect 3525 27081 3559 27115
rect 3559 27081 3568 27115
rect 3516 27072 3568 27081
rect 4712 27072 4764 27124
rect 8024 27072 8076 27124
rect 10324 27072 10376 27124
rect 12716 27115 12768 27124
rect 12716 27081 12725 27115
rect 12725 27081 12759 27115
rect 12759 27081 12768 27115
rect 12716 27072 12768 27081
rect 13544 27115 13596 27124
rect 13544 27081 13553 27115
rect 13553 27081 13587 27115
rect 13587 27081 13596 27115
rect 13544 27072 13596 27081
rect 14188 27072 14240 27124
rect 17132 27072 17184 27124
rect 3332 27004 3384 27056
rect 6092 27004 6144 27056
rect 7932 27004 7984 27056
rect 11796 27004 11848 27056
rect 16488 27004 16540 27056
rect 17500 27047 17552 27056
rect 17500 27013 17509 27047
rect 17509 27013 17543 27047
rect 17543 27013 17552 27047
rect 17500 27004 17552 27013
rect 2780 26979 2832 26988
rect 2780 26945 2789 26979
rect 2789 26945 2823 26979
rect 2823 26945 2832 26979
rect 2780 26936 2832 26945
rect 2872 26868 2924 26920
rect 8668 26936 8720 26988
rect 3608 26868 3660 26920
rect 4160 26868 4212 26920
rect 4988 26868 5040 26920
rect 7472 26911 7524 26920
rect 7472 26877 7481 26911
rect 7481 26877 7515 26911
rect 7515 26877 7524 26911
rect 7472 26868 7524 26877
rect 13268 26936 13320 26988
rect 16856 26979 16908 26988
rect 16856 26945 16865 26979
rect 16865 26945 16899 26979
rect 16899 26945 16908 26979
rect 16856 26936 16908 26945
rect 5724 26800 5776 26852
rect 7104 26800 7156 26852
rect 11152 26868 11204 26920
rect 13912 26911 13964 26920
rect 13912 26877 13921 26911
rect 13921 26877 13955 26911
rect 13955 26877 13964 26911
rect 13912 26868 13964 26877
rect 14188 26911 14240 26920
rect 14188 26877 14197 26911
rect 14197 26877 14231 26911
rect 14231 26877 14240 26911
rect 14188 26868 14240 26877
rect 17040 26911 17092 26920
rect 11888 26843 11940 26852
rect 11888 26809 11897 26843
rect 11897 26809 11931 26843
rect 11931 26809 11940 26843
rect 11888 26800 11940 26809
rect 15016 26800 15068 26852
rect 17040 26877 17049 26911
rect 17049 26877 17083 26911
rect 17083 26877 17092 26911
rect 17040 26868 17092 26877
rect 17408 26868 17460 26920
rect 10876 26775 10928 26784
rect 10876 26741 10885 26775
rect 10885 26741 10919 26775
rect 10919 26741 10928 26775
rect 10876 26732 10928 26741
rect 11796 26732 11848 26784
rect 13268 26732 13320 26784
rect 13820 26732 13872 26784
rect 16028 26732 16080 26784
rect 17316 26732 17368 26784
rect 7648 26630 7700 26682
rect 7712 26630 7764 26682
rect 7776 26630 7828 26682
rect 7840 26630 7892 26682
rect 14315 26630 14367 26682
rect 14379 26630 14431 26682
rect 14443 26630 14495 26682
rect 14507 26630 14559 26682
rect 3608 26503 3660 26512
rect 1584 26435 1636 26444
rect 1584 26401 1593 26435
rect 1593 26401 1627 26435
rect 1627 26401 1636 26435
rect 1584 26392 1636 26401
rect 1676 26392 1728 26444
rect 2320 26392 2372 26444
rect 3608 26469 3617 26503
rect 3617 26469 3651 26503
rect 3651 26469 3660 26503
rect 3608 26460 3660 26469
rect 2044 26324 2096 26376
rect 3516 26392 3568 26444
rect 4620 26528 4672 26580
rect 5632 26528 5684 26580
rect 6460 26528 6512 26580
rect 7472 26528 7524 26580
rect 8484 26571 8536 26580
rect 8484 26537 8493 26571
rect 8493 26537 8527 26571
rect 8527 26537 8536 26571
rect 8484 26528 8536 26537
rect 8668 26571 8720 26580
rect 8668 26537 8677 26571
rect 8677 26537 8711 26571
rect 8711 26537 8720 26571
rect 8668 26528 8720 26537
rect 11520 26571 11572 26580
rect 11520 26537 11529 26571
rect 11529 26537 11563 26571
rect 11563 26537 11572 26571
rect 11520 26528 11572 26537
rect 16212 26528 16264 26580
rect 5172 26503 5224 26512
rect 5172 26469 5181 26503
rect 5181 26469 5215 26503
rect 5215 26469 5224 26503
rect 5172 26460 5224 26469
rect 7656 26460 7708 26512
rect 8392 26460 8444 26512
rect 16580 26460 16632 26512
rect 3240 26367 3292 26376
rect 3240 26333 3249 26367
rect 3249 26333 3283 26367
rect 3283 26333 3292 26367
rect 3240 26324 3292 26333
rect 7104 26392 7156 26444
rect 8116 26392 8168 26444
rect 8760 26435 8812 26444
rect 8760 26401 8769 26435
rect 8769 26401 8803 26435
rect 8803 26401 8812 26435
rect 8760 26392 8812 26401
rect 9312 26435 9364 26444
rect 9312 26401 9321 26435
rect 9321 26401 9355 26435
rect 9355 26401 9364 26435
rect 9312 26392 9364 26401
rect 11428 26392 11480 26444
rect 13360 26435 13412 26444
rect 13360 26401 13369 26435
rect 13369 26401 13403 26435
rect 13403 26401 13412 26435
rect 13360 26392 13412 26401
rect 14096 26435 14148 26444
rect 8668 26324 8720 26376
rect 12716 26324 12768 26376
rect 12992 26324 13044 26376
rect 14096 26401 14105 26435
rect 14105 26401 14139 26435
rect 14139 26401 14148 26435
rect 14096 26392 14148 26401
rect 16856 26528 16908 26580
rect 14188 26324 14240 26376
rect 15108 26324 15160 26376
rect 11152 26299 11204 26308
rect 4160 26188 4212 26240
rect 11152 26265 11161 26299
rect 11161 26265 11195 26299
rect 11195 26265 11204 26299
rect 11152 26256 11204 26265
rect 11888 26299 11940 26308
rect 11888 26265 11897 26299
rect 11897 26265 11931 26299
rect 11931 26265 11940 26299
rect 11888 26256 11940 26265
rect 13728 26256 13780 26308
rect 8576 26188 8628 26240
rect 10140 26188 10192 26240
rect 10692 26188 10744 26240
rect 15752 26188 15804 26240
rect 17316 26324 17368 26376
rect 4315 26086 4367 26138
rect 4379 26086 4431 26138
rect 4443 26086 4495 26138
rect 4507 26086 4559 26138
rect 10982 26086 11034 26138
rect 11046 26086 11098 26138
rect 11110 26086 11162 26138
rect 11174 26086 11226 26138
rect 17648 26086 17700 26138
rect 17712 26086 17764 26138
rect 17776 26086 17828 26138
rect 17840 26086 17892 26138
rect 1676 26027 1728 26036
rect 1676 25993 1685 26027
rect 1685 25993 1719 26027
rect 1719 25993 1728 26027
rect 1676 25984 1728 25993
rect 2044 26027 2096 26036
rect 2044 25993 2053 26027
rect 2053 25993 2087 26027
rect 2087 25993 2096 26027
rect 2044 25984 2096 25993
rect 2872 25984 2924 26036
rect 3332 25984 3384 26036
rect 3516 25984 3568 26036
rect 4160 26027 4212 26036
rect 4160 25993 4169 26027
rect 4169 25993 4203 26027
rect 4203 25993 4212 26027
rect 4160 25984 4212 25993
rect 7104 26027 7156 26036
rect 7104 25993 7113 26027
rect 7113 25993 7147 26027
rect 7147 25993 7156 26027
rect 7104 25984 7156 25993
rect 7656 26027 7708 26036
rect 7656 25993 7665 26027
rect 7665 25993 7699 26027
rect 7699 25993 7708 26027
rect 7656 25984 7708 25993
rect 9312 25984 9364 26036
rect 12808 26027 12860 26036
rect 12808 25993 12817 26027
rect 12817 25993 12851 26027
rect 12851 25993 12860 26027
rect 12808 25984 12860 25993
rect 15476 25984 15528 26036
rect 15752 25984 15804 26036
rect 16028 25984 16080 26036
rect 16856 25984 16908 26036
rect 4712 25916 4764 25968
rect 8760 25916 8812 25968
rect 17500 25959 17552 25968
rect 17500 25925 17509 25959
rect 17509 25925 17543 25959
rect 17543 25925 17552 25959
rect 17500 25916 17552 25925
rect 6460 25891 6512 25900
rect 3700 25780 3752 25832
rect 6460 25857 6469 25891
rect 6469 25857 6503 25891
rect 6503 25857 6512 25891
rect 6460 25848 6512 25857
rect 9864 25891 9916 25900
rect 9864 25857 9873 25891
rect 9873 25857 9907 25891
rect 9907 25857 9916 25891
rect 9864 25848 9916 25857
rect 16856 25891 16908 25900
rect 16856 25857 16865 25891
rect 16865 25857 16899 25891
rect 16899 25857 16908 25891
rect 16856 25848 16908 25857
rect 5908 25780 5960 25832
rect 6368 25823 6420 25832
rect 6368 25789 6377 25823
rect 6377 25789 6411 25823
rect 6411 25789 6420 25823
rect 6368 25780 6420 25789
rect 7656 25780 7708 25832
rect 8484 25780 8536 25832
rect 8576 25823 8628 25832
rect 8576 25789 8585 25823
rect 8585 25789 8619 25823
rect 8619 25789 8628 25823
rect 8576 25780 8628 25789
rect 9772 25823 9824 25832
rect 9772 25789 9781 25823
rect 9781 25789 9815 25823
rect 9815 25789 9824 25823
rect 9772 25780 9824 25789
rect 10140 25823 10192 25832
rect 10140 25789 10149 25823
rect 10149 25789 10183 25823
rect 10183 25789 10192 25823
rect 10140 25780 10192 25789
rect 10416 25780 10468 25832
rect 12072 25780 12124 25832
rect 12992 25823 13044 25832
rect 12992 25789 13001 25823
rect 13001 25789 13035 25823
rect 13035 25789 13044 25823
rect 12992 25780 13044 25789
rect 13360 25823 13412 25832
rect 13360 25789 13369 25823
rect 13369 25789 13403 25823
rect 13403 25789 13412 25823
rect 13360 25780 13412 25789
rect 10876 25712 10928 25764
rect 12532 25712 12584 25764
rect 13820 25780 13872 25832
rect 15660 25823 15712 25832
rect 15660 25789 15669 25823
rect 15669 25789 15703 25823
rect 15703 25789 15712 25823
rect 15660 25780 15712 25789
rect 17040 25823 17092 25832
rect 17040 25789 17049 25823
rect 17049 25789 17083 25823
rect 17083 25789 17092 25823
rect 17040 25780 17092 25789
rect 17408 25780 17460 25832
rect 14096 25712 14148 25764
rect 11428 25687 11480 25696
rect 11428 25653 11437 25687
rect 11437 25653 11471 25687
rect 11471 25653 11480 25687
rect 11428 25644 11480 25653
rect 12164 25687 12216 25696
rect 12164 25653 12173 25687
rect 12173 25653 12207 25687
rect 12207 25653 12216 25687
rect 12164 25644 12216 25653
rect 12716 25644 12768 25696
rect 17316 25644 17368 25696
rect 7648 25542 7700 25594
rect 7712 25542 7764 25594
rect 7776 25542 7828 25594
rect 7840 25542 7892 25594
rect 14315 25542 14367 25594
rect 14379 25542 14431 25594
rect 14443 25542 14495 25594
rect 14507 25542 14559 25594
rect 6552 25440 6604 25492
rect 8668 25483 8720 25492
rect 8668 25449 8677 25483
rect 8677 25449 8711 25483
rect 8711 25449 8720 25483
rect 8668 25440 8720 25449
rect 8760 25440 8812 25492
rect 9496 25483 9548 25492
rect 9496 25449 9505 25483
rect 9505 25449 9539 25483
rect 9539 25449 9548 25483
rect 9496 25440 9548 25449
rect 10416 25440 10468 25492
rect 12072 25440 12124 25492
rect 13636 25483 13688 25492
rect 13636 25449 13645 25483
rect 13645 25449 13679 25483
rect 13679 25449 13688 25483
rect 13636 25440 13688 25449
rect 15292 25440 15344 25492
rect 7104 25372 7156 25424
rect 3884 25304 3936 25356
rect 4620 25347 4672 25356
rect 4620 25313 4629 25347
rect 4629 25313 4663 25347
rect 4663 25313 4672 25347
rect 4620 25304 4672 25313
rect 5908 25304 5960 25356
rect 7380 25304 7432 25356
rect 7472 25347 7524 25356
rect 7472 25313 7481 25347
rect 7481 25313 7515 25347
rect 7515 25313 7524 25347
rect 10048 25372 10100 25424
rect 7472 25304 7524 25313
rect 9036 25304 9088 25356
rect 9404 25304 9456 25356
rect 12624 25372 12676 25424
rect 12716 25347 12768 25356
rect 12716 25313 12725 25347
rect 12725 25313 12759 25347
rect 12759 25313 12768 25347
rect 12716 25304 12768 25313
rect 12900 25347 12952 25356
rect 12900 25313 12909 25347
rect 12909 25313 12943 25347
rect 12943 25313 12952 25347
rect 12900 25304 12952 25313
rect 13268 25347 13320 25356
rect 13268 25313 13277 25347
rect 13277 25313 13311 25347
rect 13311 25313 13320 25347
rect 13268 25304 13320 25313
rect 15200 25347 15252 25356
rect 15200 25313 15209 25347
rect 15209 25313 15243 25347
rect 15243 25313 15252 25347
rect 15200 25304 15252 25313
rect 15568 25347 15620 25356
rect 15568 25313 15577 25347
rect 15577 25313 15611 25347
rect 15611 25313 15620 25347
rect 15568 25304 15620 25313
rect 15752 25304 15804 25356
rect 6644 25236 6696 25288
rect 9864 25236 9916 25288
rect 13360 25236 13412 25288
rect 17040 25236 17092 25288
rect 3792 25168 3844 25220
rect 6368 25168 6420 25220
rect 10416 25211 10468 25220
rect 10416 25177 10425 25211
rect 10425 25177 10459 25211
rect 10459 25177 10468 25211
rect 10416 25168 10468 25177
rect 1400 25100 1452 25152
rect 3700 25143 3752 25152
rect 3700 25109 3709 25143
rect 3709 25109 3743 25143
rect 3743 25109 3752 25143
rect 3700 25100 3752 25109
rect 4620 25143 4672 25152
rect 4620 25109 4629 25143
rect 4629 25109 4663 25143
rect 4663 25109 4672 25143
rect 4620 25100 4672 25109
rect 13544 25143 13596 25152
rect 13544 25109 13553 25143
rect 13553 25109 13587 25143
rect 13587 25109 13596 25143
rect 13544 25100 13596 25109
rect 16764 25100 16816 25152
rect 17408 25143 17460 25152
rect 17408 25109 17417 25143
rect 17417 25109 17451 25143
rect 17451 25109 17460 25143
rect 17408 25100 17460 25109
rect 4315 24998 4367 25050
rect 4379 24998 4431 25050
rect 4443 24998 4495 25050
rect 4507 24998 4559 25050
rect 10982 24998 11034 25050
rect 11046 24998 11098 25050
rect 11110 24998 11162 25050
rect 11174 24998 11226 25050
rect 17648 24998 17700 25050
rect 17712 24998 17764 25050
rect 17776 24998 17828 25050
rect 17840 24998 17892 25050
rect 3700 24896 3752 24948
rect 9036 24939 9088 24948
rect 9036 24905 9045 24939
rect 9045 24905 9079 24939
rect 9079 24905 9088 24939
rect 9036 24896 9088 24905
rect 15108 24939 15160 24948
rect 15108 24905 15117 24939
rect 15117 24905 15151 24939
rect 15151 24905 15160 24939
rect 15108 24896 15160 24905
rect 15568 24896 15620 24948
rect 3884 24871 3936 24880
rect 3884 24837 3893 24871
rect 3893 24837 3927 24871
rect 3927 24837 3936 24871
rect 3884 24828 3936 24837
rect 1860 24760 1912 24812
rect 1400 24735 1452 24744
rect 1400 24701 1409 24735
rect 1409 24701 1443 24735
rect 1443 24701 1452 24735
rect 1400 24692 1452 24701
rect 3884 24692 3936 24744
rect 7380 24828 7432 24880
rect 8024 24803 8076 24812
rect 8024 24769 8033 24803
rect 8033 24769 8067 24803
rect 8067 24769 8076 24803
rect 8024 24760 8076 24769
rect 4620 24692 4672 24744
rect 6644 24692 6696 24744
rect 7196 24692 7248 24744
rect 7380 24692 7432 24744
rect 8300 24828 8352 24880
rect 9864 24828 9916 24880
rect 12992 24828 13044 24880
rect 3516 24624 3568 24676
rect 7012 24624 7064 24676
rect 8300 24692 8352 24744
rect 8852 24692 8904 24744
rect 10232 24735 10284 24744
rect 10232 24701 10241 24735
rect 10241 24701 10275 24735
rect 10275 24701 10284 24735
rect 10232 24692 10284 24701
rect 13912 24760 13964 24812
rect 15200 24828 15252 24880
rect 17500 24871 17552 24880
rect 17500 24837 17509 24871
rect 17509 24837 17543 24871
rect 17543 24837 17552 24871
rect 17500 24828 17552 24837
rect 10784 24692 10836 24744
rect 14188 24735 14240 24744
rect 12624 24624 12676 24676
rect 13268 24624 13320 24676
rect 14188 24701 14197 24735
rect 14197 24701 14231 24735
rect 14231 24701 14240 24735
rect 14188 24692 14240 24701
rect 14832 24692 14884 24744
rect 14004 24624 14056 24676
rect 15752 24760 15804 24812
rect 16580 24803 16632 24812
rect 16580 24769 16589 24803
rect 16589 24769 16623 24803
rect 16623 24769 16632 24803
rect 16580 24760 16632 24769
rect 15660 24735 15712 24744
rect 15660 24701 15669 24735
rect 15669 24701 15703 24735
rect 15703 24701 15712 24735
rect 15660 24692 15712 24701
rect 17040 24735 17092 24744
rect 17040 24701 17049 24735
rect 17049 24701 17083 24735
rect 17083 24701 17092 24735
rect 17040 24692 17092 24701
rect 17408 24692 17460 24744
rect 5908 24556 5960 24608
rect 6368 24556 6420 24608
rect 11520 24556 11572 24608
rect 12716 24556 12768 24608
rect 12992 24556 13044 24608
rect 13820 24556 13872 24608
rect 16212 24624 16264 24676
rect 7648 24454 7700 24506
rect 7712 24454 7764 24506
rect 7776 24454 7828 24506
rect 7840 24454 7892 24506
rect 14315 24454 14367 24506
rect 14379 24454 14431 24506
rect 14443 24454 14495 24506
rect 14507 24454 14559 24506
rect 1860 24352 1912 24404
rect 4988 24395 5040 24404
rect 4988 24361 4997 24395
rect 4997 24361 5031 24395
rect 5031 24361 5040 24395
rect 4988 24352 5040 24361
rect 5540 24352 5592 24404
rect 6552 24352 6604 24404
rect 7104 24395 7156 24404
rect 7104 24361 7113 24395
rect 7113 24361 7147 24395
rect 7147 24361 7156 24395
rect 7104 24352 7156 24361
rect 7380 24352 7432 24404
rect 8300 24395 8352 24404
rect 8300 24361 8309 24395
rect 8309 24361 8343 24395
rect 8343 24361 8352 24395
rect 8300 24352 8352 24361
rect 10048 24352 10100 24404
rect 14004 24352 14056 24404
rect 14188 24395 14240 24404
rect 14188 24361 14197 24395
rect 14197 24361 14231 24395
rect 14231 24361 14240 24395
rect 14188 24352 14240 24361
rect 16672 24395 16724 24404
rect 16672 24361 16681 24395
rect 16681 24361 16715 24395
rect 16715 24361 16724 24395
rect 16672 24352 16724 24361
rect 16856 24352 16908 24404
rect 2780 24259 2832 24268
rect 2780 24225 2789 24259
rect 2789 24225 2823 24259
rect 2823 24225 2832 24259
rect 6644 24284 6696 24336
rect 10232 24284 10284 24336
rect 13452 24327 13504 24336
rect 13452 24293 13461 24327
rect 13461 24293 13495 24327
rect 13495 24293 13504 24327
rect 13452 24284 13504 24293
rect 17224 24284 17276 24336
rect 2780 24216 2832 24225
rect 1860 24148 1912 24200
rect 5356 24080 5408 24132
rect 4068 24055 4120 24064
rect 4068 24021 4077 24055
rect 4077 24021 4111 24055
rect 4111 24021 4120 24055
rect 4068 24012 4120 24021
rect 5080 24012 5132 24064
rect 5908 24216 5960 24268
rect 7012 24259 7064 24268
rect 7012 24225 7021 24259
rect 7021 24225 7055 24259
rect 7055 24225 7064 24259
rect 7012 24216 7064 24225
rect 8944 24216 8996 24268
rect 10048 24259 10100 24268
rect 10048 24225 10057 24259
rect 10057 24225 10091 24259
rect 10091 24225 10100 24259
rect 10048 24216 10100 24225
rect 10876 24216 10928 24268
rect 11336 24216 11388 24268
rect 12900 24259 12952 24268
rect 12900 24225 12909 24259
rect 12909 24225 12943 24259
rect 12943 24225 12952 24259
rect 12900 24216 12952 24225
rect 13176 24216 13228 24268
rect 14556 24216 14608 24268
rect 17040 24259 17092 24268
rect 17040 24225 17049 24259
rect 17049 24225 17083 24259
rect 17083 24225 17092 24259
rect 17040 24216 17092 24225
rect 9036 24148 9088 24200
rect 12808 24148 12860 24200
rect 15108 24148 15160 24200
rect 8024 24080 8076 24132
rect 8668 24123 8720 24132
rect 8668 24089 8677 24123
rect 8677 24089 8711 24123
rect 8711 24089 8720 24123
rect 8668 24080 8720 24089
rect 9864 24080 9916 24132
rect 6644 24055 6696 24064
rect 6644 24021 6653 24055
rect 6653 24021 6687 24055
rect 6687 24021 6696 24055
rect 6644 24012 6696 24021
rect 4315 23910 4367 23962
rect 4379 23910 4431 23962
rect 4443 23910 4495 23962
rect 4507 23910 4559 23962
rect 10982 23910 11034 23962
rect 11046 23910 11098 23962
rect 11110 23910 11162 23962
rect 11174 23910 11226 23962
rect 17648 23910 17700 23962
rect 17712 23910 17764 23962
rect 17776 23910 17828 23962
rect 17840 23910 17892 23962
rect 11336 23851 11388 23860
rect 11336 23817 11345 23851
rect 11345 23817 11379 23851
rect 11379 23817 11388 23851
rect 11336 23808 11388 23817
rect 11980 23808 12032 23860
rect 14556 23808 14608 23860
rect 10876 23740 10928 23792
rect 15936 23740 15988 23792
rect 16948 23740 17000 23792
rect 1768 23715 1820 23724
rect 1768 23681 1777 23715
rect 1777 23681 1811 23715
rect 1811 23681 1820 23715
rect 1768 23672 1820 23681
rect 6000 23672 6052 23724
rect 7012 23672 7064 23724
rect 8484 23672 8536 23724
rect 10048 23672 10100 23724
rect 16764 23715 16816 23724
rect 16764 23681 16773 23715
rect 16773 23681 16807 23715
rect 16807 23681 16816 23715
rect 16764 23672 16816 23681
rect 17408 23672 17460 23724
rect 1860 23604 1912 23656
rect 5448 23604 5500 23656
rect 6552 23647 6604 23656
rect 6552 23613 6561 23647
rect 6561 23613 6595 23647
rect 6595 23613 6604 23647
rect 6552 23604 6604 23613
rect 7104 23647 7156 23656
rect 7104 23613 7113 23647
rect 7113 23613 7147 23647
rect 7147 23613 7156 23647
rect 7104 23604 7156 23613
rect 7288 23647 7340 23656
rect 7288 23613 7297 23647
rect 7297 23613 7331 23647
rect 7331 23613 7340 23647
rect 7288 23604 7340 23613
rect 7380 23604 7432 23656
rect 8024 23647 8076 23656
rect 8024 23613 8033 23647
rect 8033 23613 8067 23647
rect 8067 23613 8076 23647
rect 8024 23604 8076 23613
rect 3148 23579 3200 23588
rect 3148 23545 3157 23579
rect 3157 23545 3191 23579
rect 3191 23545 3200 23579
rect 3148 23536 3200 23545
rect 5172 23579 5224 23588
rect 5172 23545 5181 23579
rect 5181 23545 5215 23579
rect 5215 23545 5224 23579
rect 5172 23536 5224 23545
rect 12072 23647 12124 23656
rect 10140 23536 10192 23588
rect 12072 23613 12081 23647
rect 12081 23613 12115 23647
rect 12115 23613 12124 23647
rect 12072 23604 12124 23613
rect 12900 23647 12952 23656
rect 12900 23613 12909 23647
rect 12909 23613 12943 23647
rect 12943 23613 12952 23647
rect 12900 23604 12952 23613
rect 13636 23647 13688 23656
rect 13636 23613 13645 23647
rect 13645 23613 13679 23647
rect 13679 23613 13688 23647
rect 13636 23604 13688 23613
rect 14096 23604 14148 23656
rect 12624 23536 12676 23588
rect 15108 23604 15160 23656
rect 15844 23604 15896 23656
rect 17132 23604 17184 23656
rect 16764 23536 16816 23588
rect 16856 23536 16908 23588
rect 5080 23511 5132 23520
rect 5080 23477 5089 23511
rect 5089 23477 5123 23511
rect 5123 23477 5132 23511
rect 5080 23468 5132 23477
rect 9036 23511 9088 23520
rect 9036 23477 9045 23511
rect 9045 23477 9079 23511
rect 9079 23477 9088 23511
rect 9036 23468 9088 23477
rect 15936 23511 15988 23520
rect 15936 23477 15945 23511
rect 15945 23477 15979 23511
rect 15979 23477 15988 23511
rect 15936 23468 15988 23477
rect 16212 23468 16264 23520
rect 17040 23468 17092 23520
rect 17316 23468 17368 23520
rect 7648 23366 7700 23418
rect 7712 23366 7764 23418
rect 7776 23366 7828 23418
rect 7840 23366 7892 23418
rect 14315 23366 14367 23418
rect 14379 23366 14431 23418
rect 14443 23366 14495 23418
rect 14507 23366 14559 23418
rect 1768 23264 1820 23316
rect 2688 23264 2740 23316
rect 1860 22992 1912 23044
rect 3884 23264 3936 23316
rect 3792 23128 3844 23180
rect 7380 23264 7432 23316
rect 8484 23307 8536 23316
rect 8484 23273 8493 23307
rect 8493 23273 8527 23307
rect 8527 23273 8536 23307
rect 8484 23264 8536 23273
rect 8944 23264 8996 23316
rect 11060 23307 11112 23316
rect 11060 23273 11069 23307
rect 11069 23273 11103 23307
rect 11103 23273 11112 23307
rect 11060 23264 11112 23273
rect 13636 23307 13688 23316
rect 13636 23273 13645 23307
rect 13645 23273 13679 23307
rect 13679 23273 13688 23307
rect 13636 23264 13688 23273
rect 5264 23196 5316 23248
rect 12348 23196 12400 23248
rect 14924 23196 14976 23248
rect 15016 23196 15068 23248
rect 4712 23128 4764 23180
rect 5356 23128 5408 23180
rect 6552 23128 6604 23180
rect 7288 23128 7340 23180
rect 7564 23128 7616 23180
rect 4160 23060 4212 23112
rect 5908 23060 5960 23112
rect 7380 23060 7432 23112
rect 9956 23128 10008 23180
rect 10416 23128 10468 23180
rect 10600 23171 10652 23180
rect 10600 23137 10609 23171
rect 10609 23137 10643 23171
rect 10643 23137 10652 23171
rect 10600 23128 10652 23137
rect 11888 23128 11940 23180
rect 12440 23171 12492 23180
rect 12440 23137 12449 23171
rect 12449 23137 12483 23171
rect 12483 23137 12492 23171
rect 12900 23171 12952 23180
rect 12440 23128 12492 23137
rect 12900 23137 12909 23171
rect 12909 23137 12943 23171
rect 12943 23137 12952 23171
rect 12900 23128 12952 23137
rect 13912 23128 13964 23180
rect 14556 23171 14608 23180
rect 14556 23137 14565 23171
rect 14565 23137 14599 23171
rect 14599 23137 14608 23171
rect 14556 23128 14608 23137
rect 16580 23171 16632 23180
rect 11428 23060 11480 23112
rect 13268 23103 13320 23112
rect 13268 23069 13277 23103
rect 13277 23069 13311 23103
rect 13311 23069 13320 23103
rect 16580 23137 16589 23171
rect 16589 23137 16623 23171
rect 16623 23137 16632 23171
rect 16580 23128 16632 23137
rect 17040 23171 17092 23180
rect 17040 23137 17049 23171
rect 17049 23137 17083 23171
rect 17083 23137 17092 23171
rect 17040 23128 17092 23137
rect 13268 23060 13320 23069
rect 16120 23060 16172 23112
rect 15476 22992 15528 23044
rect 5356 22967 5408 22976
rect 5356 22933 5365 22967
rect 5365 22933 5399 22967
rect 5399 22933 5408 22967
rect 5356 22924 5408 22933
rect 9496 22967 9548 22976
rect 9496 22933 9505 22967
rect 9505 22933 9539 22967
rect 9539 22933 9548 22967
rect 9496 22924 9548 22933
rect 12716 22924 12768 22976
rect 16028 22967 16080 22976
rect 16028 22933 16037 22967
rect 16037 22933 16071 22967
rect 16071 22933 16080 22967
rect 16028 22924 16080 22933
rect 17040 22924 17092 22976
rect 17408 22967 17460 22976
rect 17408 22933 17417 22967
rect 17417 22933 17451 22967
rect 17451 22933 17460 22967
rect 17408 22924 17460 22933
rect 4315 22822 4367 22874
rect 4379 22822 4431 22874
rect 4443 22822 4495 22874
rect 4507 22822 4559 22874
rect 10982 22822 11034 22874
rect 11046 22822 11098 22874
rect 11110 22822 11162 22874
rect 11174 22822 11226 22874
rect 17648 22822 17700 22874
rect 17712 22822 17764 22874
rect 17776 22822 17828 22874
rect 17840 22822 17892 22874
rect 4068 22720 4120 22772
rect 6552 22763 6604 22772
rect 6552 22729 6561 22763
rect 6561 22729 6595 22763
rect 6595 22729 6604 22763
rect 6552 22720 6604 22729
rect 6736 22720 6788 22772
rect 8116 22720 8168 22772
rect 10416 22720 10468 22772
rect 10600 22720 10652 22772
rect 11428 22763 11480 22772
rect 11428 22729 11437 22763
rect 11437 22729 11471 22763
rect 11471 22729 11480 22763
rect 11428 22720 11480 22729
rect 9956 22652 10008 22704
rect 10968 22652 11020 22704
rect 5356 22584 5408 22636
rect 9496 22584 9548 22636
rect 13084 22720 13136 22772
rect 4988 22559 5040 22568
rect 4988 22525 4997 22559
rect 4997 22525 5031 22559
rect 5031 22525 5040 22559
rect 4988 22516 5040 22525
rect 5172 22559 5224 22568
rect 5172 22525 5181 22559
rect 5181 22525 5215 22559
rect 5215 22525 5224 22559
rect 5172 22516 5224 22525
rect 8116 22559 8168 22568
rect 8116 22525 8125 22559
rect 8125 22525 8159 22559
rect 8159 22525 8168 22559
rect 8116 22516 8168 22525
rect 8300 22516 8352 22568
rect 3792 22423 3844 22432
rect 3792 22389 3801 22423
rect 3801 22389 3835 22423
rect 3835 22389 3844 22423
rect 3792 22380 3844 22389
rect 4804 22423 4856 22432
rect 4804 22389 4813 22423
rect 4813 22389 4847 22423
rect 4847 22389 4856 22423
rect 4804 22380 4856 22389
rect 7104 22423 7156 22432
rect 7104 22389 7113 22423
rect 7113 22389 7147 22423
rect 7147 22389 7156 22423
rect 7564 22448 7616 22500
rect 8484 22448 8536 22500
rect 10508 22559 10560 22568
rect 10508 22525 10517 22559
rect 10517 22525 10551 22559
rect 10551 22525 10560 22559
rect 13636 22695 13688 22704
rect 13636 22661 13645 22695
rect 13645 22661 13679 22695
rect 13679 22661 13688 22695
rect 13636 22652 13688 22661
rect 12900 22584 12952 22636
rect 14832 22720 14884 22772
rect 16120 22720 16172 22772
rect 14924 22652 14976 22704
rect 17500 22695 17552 22704
rect 10508 22516 10560 22525
rect 13084 22516 13136 22568
rect 13360 22516 13412 22568
rect 13452 22516 13504 22568
rect 14556 22584 14608 22636
rect 17500 22661 17509 22695
rect 17509 22661 17543 22695
rect 17543 22661 17552 22695
rect 17500 22652 17552 22661
rect 15200 22584 15252 22636
rect 16764 22584 16816 22636
rect 16672 22559 16724 22568
rect 16672 22525 16681 22559
rect 16681 22525 16715 22559
rect 16715 22525 16724 22559
rect 16672 22516 16724 22525
rect 9864 22448 9916 22500
rect 16856 22448 16908 22500
rect 7104 22380 7156 22389
rect 7380 22380 7432 22432
rect 9772 22423 9824 22432
rect 9772 22389 9781 22423
rect 9781 22389 9815 22423
rect 9815 22389 9824 22423
rect 9772 22380 9824 22389
rect 11336 22380 11388 22432
rect 12440 22380 12492 22432
rect 7648 22278 7700 22330
rect 7712 22278 7764 22330
rect 7776 22278 7828 22330
rect 7840 22278 7892 22330
rect 14315 22278 14367 22330
rect 14379 22278 14431 22330
rect 14443 22278 14495 22330
rect 14507 22278 14559 22330
rect 3792 22176 3844 22228
rect 3884 22108 3936 22160
rect 1860 22083 1912 22092
rect 1860 22049 1869 22083
rect 1869 22049 1903 22083
rect 1903 22049 1912 22083
rect 1860 22040 1912 22049
rect 2136 22083 2188 22092
rect 2136 22049 2145 22083
rect 2145 22049 2179 22083
rect 2179 22049 2188 22083
rect 2136 22040 2188 22049
rect 4712 22176 4764 22228
rect 4988 22176 5040 22228
rect 6184 22176 6236 22228
rect 6460 22219 6512 22228
rect 6460 22185 6469 22219
rect 6469 22185 6503 22219
rect 6503 22185 6512 22219
rect 6460 22176 6512 22185
rect 8484 22219 8536 22228
rect 8484 22185 8493 22219
rect 8493 22185 8527 22219
rect 8527 22185 8536 22219
rect 8484 22176 8536 22185
rect 14648 22176 14700 22228
rect 6736 22108 6788 22160
rect 9680 22151 9732 22160
rect 9680 22117 9689 22151
rect 9689 22117 9723 22151
rect 9723 22117 9732 22151
rect 9680 22108 9732 22117
rect 5080 21904 5132 21956
rect 5724 22083 5776 22092
rect 5724 22049 5733 22083
rect 5733 22049 5767 22083
rect 5767 22049 5776 22083
rect 5724 22040 5776 22049
rect 7012 22083 7064 22092
rect 7012 22049 7021 22083
rect 7021 22049 7055 22083
rect 7055 22049 7064 22083
rect 7012 22040 7064 22049
rect 7104 22040 7156 22092
rect 9864 22040 9916 22092
rect 10048 22040 10100 22092
rect 10968 22040 11020 22092
rect 12716 22040 12768 22092
rect 15016 22083 15068 22092
rect 6368 21972 6420 22024
rect 8116 22015 8168 22024
rect 8116 21981 8125 22015
rect 8125 21981 8159 22015
rect 8159 21981 8168 22015
rect 8116 21972 8168 21981
rect 8576 21972 8628 22024
rect 10232 22015 10284 22024
rect 10232 21981 10241 22015
rect 10241 21981 10275 22015
rect 10275 21981 10284 22015
rect 10232 21972 10284 21981
rect 10692 22015 10744 22024
rect 10692 21981 10701 22015
rect 10701 21981 10735 22015
rect 10735 21981 10744 22015
rect 10692 21972 10744 21981
rect 11520 21972 11572 22024
rect 15016 22049 15025 22083
rect 15025 22049 15059 22083
rect 15059 22049 15068 22083
rect 15016 22040 15068 22049
rect 15660 22108 15712 22160
rect 16212 22040 16264 22092
rect 16672 22040 16724 22092
rect 16856 22083 16908 22092
rect 16856 22049 16865 22083
rect 16865 22049 16899 22083
rect 16899 22049 16908 22083
rect 16856 22040 16908 22049
rect 14924 21972 14976 22024
rect 15660 21972 15712 22024
rect 16764 21972 16816 22024
rect 13636 21904 13688 21956
rect 15384 21904 15436 21956
rect 16488 21904 16540 21956
rect 3424 21879 3476 21888
rect 3424 21845 3433 21879
rect 3433 21845 3467 21879
rect 3467 21845 3476 21879
rect 3424 21836 3476 21845
rect 7380 21879 7432 21888
rect 7380 21845 7389 21879
rect 7389 21845 7423 21879
rect 7423 21845 7432 21879
rect 7380 21836 7432 21845
rect 13452 21879 13504 21888
rect 13452 21845 13461 21879
rect 13461 21845 13495 21879
rect 13495 21845 13504 21879
rect 13452 21836 13504 21845
rect 13912 21879 13964 21888
rect 13912 21845 13921 21879
rect 13921 21845 13955 21879
rect 13955 21845 13964 21879
rect 13912 21836 13964 21845
rect 15568 21836 15620 21888
rect 16580 21836 16632 21888
rect 4315 21734 4367 21786
rect 4379 21734 4431 21786
rect 4443 21734 4495 21786
rect 4507 21734 4559 21786
rect 10982 21734 11034 21786
rect 11046 21734 11098 21786
rect 11110 21734 11162 21786
rect 11174 21734 11226 21786
rect 17648 21734 17700 21786
rect 17712 21734 17764 21786
rect 17776 21734 17828 21786
rect 17840 21734 17892 21786
rect 2136 21632 2188 21684
rect 7380 21632 7432 21684
rect 8300 21632 8352 21684
rect 10048 21632 10100 21684
rect 10232 21675 10284 21684
rect 10232 21641 10241 21675
rect 10241 21641 10275 21675
rect 10275 21641 10284 21675
rect 10232 21632 10284 21641
rect 1860 21564 1912 21616
rect 10692 21564 10744 21616
rect 5540 21496 5592 21548
rect 6644 21539 6696 21548
rect 6644 21505 6653 21539
rect 6653 21505 6687 21539
rect 6687 21505 6696 21539
rect 6644 21496 6696 21505
rect 6368 21428 6420 21480
rect 7288 21471 7340 21480
rect 7288 21437 7297 21471
rect 7297 21437 7331 21471
rect 7331 21437 7340 21471
rect 7288 21428 7340 21437
rect 8208 21471 8260 21480
rect 8208 21437 8217 21471
rect 8217 21437 8251 21471
rect 8251 21437 8260 21471
rect 8208 21428 8260 21437
rect 12348 21632 12400 21684
rect 12532 21675 12584 21684
rect 12532 21641 12541 21675
rect 12541 21641 12575 21675
rect 12575 21641 12584 21675
rect 12532 21632 12584 21641
rect 15016 21632 15068 21684
rect 15660 21675 15712 21684
rect 15660 21641 15669 21675
rect 15669 21641 15703 21675
rect 15703 21641 15712 21675
rect 15660 21632 15712 21641
rect 14188 21564 14240 21616
rect 15292 21564 15344 21616
rect 17040 21564 17092 21616
rect 14372 21539 14424 21548
rect 14372 21505 14381 21539
rect 14381 21505 14415 21539
rect 14415 21505 14424 21539
rect 14372 21496 14424 21505
rect 14648 21539 14700 21548
rect 14648 21505 14657 21539
rect 14657 21505 14691 21539
rect 14691 21505 14700 21539
rect 14648 21496 14700 21505
rect 15016 21496 15068 21548
rect 17224 21496 17276 21548
rect 5724 21360 5776 21412
rect 6828 21360 6880 21412
rect 12532 21360 12584 21412
rect 12716 21360 12768 21412
rect 13176 21360 13228 21412
rect 13820 21428 13872 21480
rect 14740 21428 14792 21480
rect 15568 21360 15620 21412
rect 16764 21403 16816 21412
rect 16764 21369 16773 21403
rect 16773 21369 16807 21403
rect 16807 21369 16816 21403
rect 16764 21360 16816 21369
rect 17040 21360 17092 21412
rect 17224 21360 17276 21412
rect 6184 21335 6236 21344
rect 6184 21301 6193 21335
rect 6193 21301 6227 21335
rect 6227 21301 6236 21335
rect 6184 21292 6236 21301
rect 6368 21335 6420 21344
rect 6368 21301 6377 21335
rect 6377 21301 6411 21335
rect 6411 21301 6420 21335
rect 6368 21292 6420 21301
rect 7104 21292 7156 21344
rect 8760 21292 8812 21344
rect 12072 21292 12124 21344
rect 12808 21335 12860 21344
rect 12808 21301 12817 21335
rect 12817 21301 12851 21335
rect 12851 21301 12860 21335
rect 12808 21292 12860 21301
rect 13728 21292 13780 21344
rect 14924 21292 14976 21344
rect 16580 21335 16632 21344
rect 16580 21301 16589 21335
rect 16589 21301 16623 21335
rect 16623 21301 16632 21335
rect 16580 21292 16632 21301
rect 7648 21190 7700 21242
rect 7712 21190 7764 21242
rect 7776 21190 7828 21242
rect 7840 21190 7892 21242
rect 14315 21190 14367 21242
rect 14379 21190 14431 21242
rect 14443 21190 14495 21242
rect 14507 21190 14559 21242
rect 1400 21088 1452 21140
rect 6184 21088 6236 21140
rect 6736 21088 6788 21140
rect 7288 21088 7340 21140
rect 12440 21088 12492 21140
rect 12716 21088 12768 21140
rect 13176 21131 13228 21140
rect 13176 21097 13185 21131
rect 13185 21097 13219 21131
rect 13219 21097 13228 21131
rect 13176 21088 13228 21097
rect 13820 21131 13872 21140
rect 13820 21097 13829 21131
rect 13829 21097 13863 21131
rect 13863 21097 13872 21131
rect 13820 21088 13872 21097
rect 14188 21131 14240 21140
rect 14188 21097 14197 21131
rect 14197 21097 14231 21131
rect 14231 21097 14240 21131
rect 14188 21088 14240 21097
rect 16672 21088 16724 21140
rect 5908 21063 5960 21072
rect 5908 21029 5917 21063
rect 5917 21029 5951 21063
rect 5951 21029 5960 21063
rect 5908 21020 5960 21029
rect 6644 21063 6696 21072
rect 6644 21029 6653 21063
rect 6653 21029 6687 21063
rect 6687 21029 6696 21063
rect 6644 21020 6696 21029
rect 1400 20995 1452 21004
rect 1400 20961 1409 20995
rect 1409 20961 1443 20995
rect 1443 20961 1452 20995
rect 1400 20952 1452 20961
rect 1676 20995 1728 21004
rect 1676 20961 1685 20995
rect 1685 20961 1719 20995
rect 1719 20961 1728 20995
rect 1676 20952 1728 20961
rect 3884 20952 3936 21004
rect 4804 20952 4856 21004
rect 5816 20995 5868 21004
rect 5816 20961 5825 20995
rect 5825 20961 5859 20995
rect 5859 20961 5868 20995
rect 5816 20952 5868 20961
rect 7104 20995 7156 21004
rect 7104 20961 7113 20995
rect 7113 20961 7147 20995
rect 7147 20961 7156 20995
rect 7104 20952 7156 20961
rect 7472 20995 7524 21004
rect 7472 20961 7481 20995
rect 7481 20961 7515 20995
rect 7515 20961 7524 20995
rect 7472 20952 7524 20961
rect 8576 21020 8628 21072
rect 15568 21020 15620 21072
rect 16764 21020 16816 21072
rect 17132 21063 17184 21072
rect 9036 20952 9088 21004
rect 13360 20952 13412 21004
rect 15108 20995 15160 21004
rect 15108 20961 15117 20995
rect 15117 20961 15151 20995
rect 15151 20961 15160 20995
rect 15108 20952 15160 20961
rect 15660 20952 15712 21004
rect 16028 20995 16080 21004
rect 16028 20961 16037 20995
rect 16037 20961 16071 20995
rect 16071 20961 16080 20995
rect 16028 20952 16080 20961
rect 16304 20952 16356 21004
rect 17132 21029 17141 21063
rect 17141 21029 17175 21063
rect 17175 21029 17184 21063
rect 17132 21020 17184 21029
rect 17500 20952 17552 21004
rect 2964 20791 3016 20800
rect 2964 20757 2973 20791
rect 2973 20757 3007 20791
rect 3007 20757 3016 20791
rect 2964 20748 3016 20757
rect 4160 20748 4212 20800
rect 12440 20748 12492 20800
rect 13176 20748 13228 20800
rect 13728 20748 13780 20800
rect 16764 20748 16816 20800
rect 17224 20748 17276 20800
rect 4315 20646 4367 20698
rect 4379 20646 4431 20698
rect 4443 20646 4495 20698
rect 4507 20646 4559 20698
rect 10982 20646 11034 20698
rect 11046 20646 11098 20698
rect 11110 20646 11162 20698
rect 11174 20646 11226 20698
rect 17648 20646 17700 20698
rect 17712 20646 17764 20698
rect 17776 20646 17828 20698
rect 17840 20646 17892 20698
rect 1676 20587 1728 20596
rect 1676 20553 1685 20587
rect 1685 20553 1719 20587
rect 1719 20553 1728 20587
rect 1676 20544 1728 20553
rect 3608 20587 3660 20596
rect 3608 20553 3617 20587
rect 3617 20553 3651 20587
rect 3651 20553 3660 20587
rect 3608 20544 3660 20553
rect 7104 20544 7156 20596
rect 8760 20587 8812 20596
rect 8760 20553 8769 20587
rect 8769 20553 8803 20587
rect 8803 20553 8812 20587
rect 8760 20544 8812 20553
rect 9036 20587 9088 20596
rect 9036 20553 9045 20587
rect 9045 20553 9079 20587
rect 9079 20553 9088 20587
rect 9036 20544 9088 20553
rect 13360 20587 13412 20596
rect 13360 20553 13369 20587
rect 13369 20553 13403 20587
rect 13403 20553 13412 20587
rect 13360 20544 13412 20553
rect 1400 20476 1452 20528
rect 6644 20476 6696 20528
rect 9404 20519 9456 20528
rect 3884 20383 3936 20392
rect 3884 20349 3893 20383
rect 3893 20349 3927 20383
rect 3927 20349 3936 20383
rect 3884 20340 3936 20349
rect 4068 20383 4120 20392
rect 4068 20349 4077 20383
rect 4077 20349 4111 20383
rect 4111 20349 4120 20383
rect 4068 20340 4120 20349
rect 7472 20408 7524 20460
rect 9404 20485 9413 20519
rect 9413 20485 9447 20519
rect 9447 20485 9456 20519
rect 9404 20476 9456 20485
rect 8208 20408 8260 20460
rect 12348 20451 12400 20460
rect 12348 20417 12357 20451
rect 12357 20417 12391 20451
rect 12391 20417 12400 20451
rect 12348 20408 12400 20417
rect 3700 20247 3752 20256
rect 3700 20213 3709 20247
rect 3709 20213 3743 20247
rect 3743 20213 3752 20247
rect 3700 20204 3752 20213
rect 5448 20247 5500 20256
rect 5448 20213 5457 20247
rect 5457 20213 5491 20247
rect 5491 20213 5500 20247
rect 5448 20204 5500 20213
rect 6920 20204 6972 20256
rect 8024 20247 8076 20256
rect 8024 20213 8033 20247
rect 8033 20213 8067 20247
rect 8067 20213 8076 20247
rect 9864 20383 9916 20392
rect 9864 20349 9873 20383
rect 9873 20349 9907 20383
rect 9907 20349 9916 20383
rect 9864 20340 9916 20349
rect 12532 20383 12584 20392
rect 12532 20349 12541 20383
rect 12541 20349 12575 20383
rect 12575 20349 12584 20383
rect 12532 20340 12584 20349
rect 11888 20315 11940 20324
rect 11888 20281 11897 20315
rect 11897 20281 11931 20315
rect 11931 20281 11940 20315
rect 12992 20340 13044 20392
rect 14832 20544 14884 20596
rect 15108 20587 15160 20596
rect 15108 20553 15117 20587
rect 15117 20553 15151 20587
rect 15151 20553 15160 20587
rect 15108 20544 15160 20553
rect 16028 20544 16080 20596
rect 16580 20476 16632 20528
rect 15200 20340 15252 20392
rect 15844 20340 15896 20392
rect 17408 20340 17460 20392
rect 17500 20383 17552 20392
rect 17500 20349 17509 20383
rect 17509 20349 17543 20383
rect 17543 20349 17552 20383
rect 17500 20340 17552 20349
rect 11888 20272 11940 20281
rect 13084 20315 13136 20324
rect 8024 20204 8076 20213
rect 12164 20204 12216 20256
rect 13084 20281 13093 20315
rect 13093 20281 13127 20315
rect 13127 20281 13136 20315
rect 13084 20272 13136 20281
rect 13820 20247 13872 20256
rect 13820 20213 13829 20247
rect 13829 20213 13863 20247
rect 13863 20213 13872 20247
rect 13820 20204 13872 20213
rect 14924 20204 14976 20256
rect 15568 20204 15620 20256
rect 7648 20102 7700 20154
rect 7712 20102 7764 20154
rect 7776 20102 7828 20154
rect 7840 20102 7892 20154
rect 14315 20102 14367 20154
rect 14379 20102 14431 20154
rect 14443 20102 14495 20154
rect 14507 20102 14559 20154
rect 1400 20000 1452 20052
rect 5816 20000 5868 20052
rect 6552 20000 6604 20052
rect 7472 20000 7524 20052
rect 12164 20043 12216 20052
rect 12164 20009 12173 20043
rect 12173 20009 12207 20043
rect 12207 20009 12216 20043
rect 12164 20000 12216 20009
rect 16304 20043 16356 20052
rect 16304 20009 16313 20043
rect 16313 20009 16347 20043
rect 16347 20009 16356 20043
rect 16304 20000 16356 20009
rect 17408 20000 17460 20052
rect 3424 19907 3476 19916
rect 3424 19873 3433 19907
rect 3433 19873 3467 19907
rect 3467 19873 3476 19907
rect 3424 19864 3476 19873
rect 6368 19864 6420 19916
rect 6920 19907 6972 19916
rect 6920 19873 6929 19907
rect 6929 19873 6963 19907
rect 6963 19873 6972 19907
rect 6920 19864 6972 19873
rect 15292 19864 15344 19916
rect 3608 19796 3660 19848
rect 6736 19796 6788 19848
rect 12624 19839 12676 19848
rect 12624 19805 12633 19839
rect 12633 19805 12667 19839
rect 12667 19805 12676 19839
rect 12624 19796 12676 19805
rect 12808 19796 12860 19848
rect 13728 19796 13780 19848
rect 15844 19907 15896 19916
rect 15844 19873 15853 19907
rect 15853 19873 15887 19907
rect 15887 19873 15896 19907
rect 15844 19864 15896 19873
rect 17500 19864 17552 19916
rect 12992 19728 13044 19780
rect 14740 19771 14792 19780
rect 14740 19737 14749 19771
rect 14749 19737 14783 19771
rect 14783 19737 14792 19771
rect 14740 19728 14792 19737
rect 15200 19771 15252 19780
rect 15200 19737 15209 19771
rect 15209 19737 15243 19771
rect 15243 19737 15252 19771
rect 15200 19728 15252 19737
rect 4712 19703 4764 19712
rect 4712 19669 4721 19703
rect 4721 19669 4755 19703
rect 4755 19669 4764 19703
rect 4712 19660 4764 19669
rect 6828 19660 6880 19712
rect 7012 19660 7064 19712
rect 9864 19703 9916 19712
rect 9864 19669 9873 19703
rect 9873 19669 9907 19703
rect 9907 19669 9916 19703
rect 9864 19660 9916 19669
rect 13820 19703 13872 19712
rect 13820 19669 13829 19703
rect 13829 19669 13863 19703
rect 13863 19669 13872 19703
rect 13820 19660 13872 19669
rect 14188 19703 14240 19712
rect 14188 19669 14197 19703
rect 14197 19669 14231 19703
rect 14231 19669 14240 19703
rect 14188 19660 14240 19669
rect 17224 19660 17276 19712
rect 17500 19660 17552 19712
rect 4315 19558 4367 19610
rect 4379 19558 4431 19610
rect 4443 19558 4495 19610
rect 4507 19558 4559 19610
rect 10982 19558 11034 19610
rect 11046 19558 11098 19610
rect 11110 19558 11162 19610
rect 11174 19558 11226 19610
rect 17648 19558 17700 19610
rect 17712 19558 17764 19610
rect 17776 19558 17828 19610
rect 17840 19558 17892 19610
rect 3424 19499 3476 19508
rect 3424 19465 3433 19499
rect 3433 19465 3467 19499
rect 3467 19465 3476 19499
rect 3424 19456 3476 19465
rect 3700 19499 3752 19508
rect 3700 19465 3709 19499
rect 3709 19465 3743 19499
rect 3743 19465 3752 19499
rect 3700 19456 3752 19465
rect 6552 19499 6604 19508
rect 6552 19465 6561 19499
rect 6561 19465 6595 19499
rect 6595 19465 6604 19499
rect 6552 19456 6604 19465
rect 6736 19456 6788 19508
rect 12164 19456 12216 19508
rect 13728 19499 13780 19508
rect 12348 19388 12400 19440
rect 12808 19388 12860 19440
rect 13176 19388 13228 19440
rect 13728 19465 13737 19499
rect 13737 19465 13771 19499
rect 13771 19465 13780 19499
rect 13728 19456 13780 19465
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 1492 19252 1544 19304
rect 5080 19295 5132 19304
rect 5080 19261 5089 19295
rect 5089 19261 5123 19295
rect 5123 19261 5132 19295
rect 5080 19252 5132 19261
rect 13084 19320 13136 19372
rect 13820 19388 13872 19440
rect 16304 19388 16356 19440
rect 5448 19295 5500 19304
rect 4068 19184 4120 19236
rect 4160 19116 4212 19168
rect 5448 19261 5457 19295
rect 5457 19261 5491 19295
rect 5491 19261 5500 19295
rect 5448 19252 5500 19261
rect 6368 19252 6420 19304
rect 8024 19184 8076 19236
rect 11612 19184 11664 19236
rect 13176 19252 13228 19304
rect 13544 19252 13596 19304
rect 15016 19295 15068 19304
rect 15016 19261 15025 19295
rect 15025 19261 15059 19295
rect 15059 19261 15068 19295
rect 15016 19252 15068 19261
rect 15844 19295 15896 19304
rect 15844 19261 15853 19295
rect 15853 19261 15887 19295
rect 15887 19261 15896 19295
rect 15844 19252 15896 19261
rect 17316 19295 17368 19304
rect 17316 19261 17325 19295
rect 17325 19261 17359 19295
rect 17359 19261 17368 19295
rect 17316 19252 17368 19261
rect 17500 19320 17552 19372
rect 13360 19184 13412 19236
rect 14740 19184 14792 19236
rect 16764 19227 16816 19236
rect 5724 19116 5776 19168
rect 7380 19116 7432 19168
rect 11796 19159 11848 19168
rect 11796 19125 11805 19159
rect 11805 19125 11839 19159
rect 11839 19125 11848 19159
rect 11796 19116 11848 19125
rect 12164 19159 12216 19168
rect 12164 19125 12173 19159
rect 12173 19125 12207 19159
rect 12207 19125 12216 19159
rect 12164 19116 12216 19125
rect 15292 19116 15344 19168
rect 16764 19193 16773 19227
rect 16773 19193 16807 19227
rect 16807 19193 16816 19227
rect 16764 19184 16816 19193
rect 7648 19014 7700 19066
rect 7712 19014 7764 19066
rect 7776 19014 7828 19066
rect 7840 19014 7892 19066
rect 14315 19014 14367 19066
rect 14379 19014 14431 19066
rect 14443 19014 14495 19066
rect 14507 19014 14559 19066
rect 1492 18912 1544 18964
rect 5080 18912 5132 18964
rect 6368 18912 6420 18964
rect 12440 18912 12492 18964
rect 13084 18912 13136 18964
rect 10784 18819 10836 18828
rect 10784 18785 10793 18819
rect 10793 18785 10827 18819
rect 10827 18785 10836 18819
rect 10784 18776 10836 18785
rect 10876 18776 10928 18828
rect 11336 18819 11388 18828
rect 11336 18785 11345 18819
rect 11345 18785 11379 18819
rect 11379 18785 11388 18819
rect 11336 18776 11388 18785
rect 11888 18776 11940 18828
rect 12532 18776 12584 18828
rect 14004 18776 14056 18828
rect 14280 18776 14332 18828
rect 14924 18776 14976 18828
rect 15752 18776 15804 18828
rect 16488 18819 16540 18828
rect 16488 18785 16497 18819
rect 16497 18785 16531 18819
rect 16531 18785 16540 18819
rect 16488 18776 16540 18785
rect 11520 18751 11572 18760
rect 11520 18717 11529 18751
rect 11529 18717 11563 18751
rect 11563 18717 11572 18751
rect 11520 18708 11572 18717
rect 14740 18708 14792 18760
rect 16120 18708 16172 18760
rect 11888 18640 11940 18692
rect 13176 18640 13228 18692
rect 15108 18640 15160 18692
rect 16580 18683 16632 18692
rect 16580 18649 16589 18683
rect 16589 18649 16623 18683
rect 16623 18649 16632 18683
rect 16580 18640 16632 18649
rect 5724 18572 5776 18624
rect 12624 18572 12676 18624
rect 12992 18572 13044 18624
rect 4315 18470 4367 18522
rect 4379 18470 4431 18522
rect 4443 18470 4495 18522
rect 4507 18470 4559 18522
rect 10982 18470 11034 18522
rect 11046 18470 11098 18522
rect 11110 18470 11162 18522
rect 11174 18470 11226 18522
rect 17648 18470 17700 18522
rect 17712 18470 17764 18522
rect 17776 18470 17828 18522
rect 17840 18470 17892 18522
rect 3792 18411 3844 18420
rect 3792 18377 3801 18411
rect 3801 18377 3835 18411
rect 3835 18377 3844 18411
rect 3792 18368 3844 18377
rect 8024 18411 8076 18420
rect 8024 18377 8033 18411
rect 8033 18377 8067 18411
rect 8067 18377 8076 18411
rect 8024 18368 8076 18377
rect 10876 18411 10928 18420
rect 10876 18377 10885 18411
rect 10885 18377 10919 18411
rect 10919 18377 10928 18411
rect 10876 18368 10928 18377
rect 14648 18411 14700 18420
rect 14648 18377 14657 18411
rect 14657 18377 14691 18411
rect 14691 18377 14700 18411
rect 14648 18368 14700 18377
rect 12164 18343 12216 18352
rect 12164 18309 12173 18343
rect 12173 18309 12207 18343
rect 12207 18309 12216 18343
rect 12164 18300 12216 18309
rect 12532 18300 12584 18352
rect 13636 18343 13688 18352
rect 13636 18309 13645 18343
rect 13645 18309 13679 18343
rect 13679 18309 13688 18343
rect 13636 18300 13688 18309
rect 13820 18300 13872 18352
rect 3700 18232 3752 18284
rect 4160 18275 4212 18284
rect 4160 18241 4169 18275
rect 4169 18241 4203 18275
rect 4203 18241 4212 18275
rect 4160 18232 4212 18241
rect 3792 18164 3844 18216
rect 11796 18207 11848 18216
rect 11796 18173 11805 18207
rect 11805 18173 11839 18207
rect 11839 18173 11848 18207
rect 11796 18164 11848 18173
rect 11888 18164 11940 18216
rect 16396 18232 16448 18284
rect 12532 18096 12584 18148
rect 14740 18164 14792 18216
rect 14924 18164 14976 18216
rect 16120 18164 16172 18216
rect 16856 18207 16908 18216
rect 16856 18173 16865 18207
rect 16865 18173 16899 18207
rect 16899 18173 16908 18207
rect 16856 18164 16908 18173
rect 14556 18096 14608 18148
rect 1676 18071 1728 18080
rect 1676 18037 1685 18071
rect 1685 18037 1719 18071
rect 1719 18037 1728 18071
rect 1676 18028 1728 18037
rect 5724 18028 5776 18080
rect 11612 18028 11664 18080
rect 12072 18028 12124 18080
rect 15752 18028 15804 18080
rect 16212 18071 16264 18080
rect 16212 18037 16221 18071
rect 16221 18037 16255 18071
rect 16255 18037 16264 18071
rect 16212 18028 16264 18037
rect 7648 17926 7700 17978
rect 7712 17926 7764 17978
rect 7776 17926 7828 17978
rect 7840 17926 7892 17978
rect 14315 17926 14367 17978
rect 14379 17926 14431 17978
rect 14443 17926 14495 17978
rect 14507 17926 14559 17978
rect 4160 17867 4212 17876
rect 4160 17833 4169 17867
rect 4169 17833 4203 17867
rect 4203 17833 4212 17867
rect 4160 17824 4212 17833
rect 10784 17867 10836 17876
rect 10784 17833 10793 17867
rect 10793 17833 10827 17867
rect 10827 17833 10836 17867
rect 10784 17824 10836 17833
rect 11796 17867 11848 17876
rect 11796 17833 11805 17867
rect 11805 17833 11839 17867
rect 11839 17833 11848 17867
rect 11796 17824 11848 17833
rect 12440 17824 12492 17876
rect 16488 17867 16540 17876
rect 9312 17756 9364 17808
rect 16488 17833 16497 17867
rect 16497 17833 16531 17867
rect 16531 17833 16540 17867
rect 16488 17824 16540 17833
rect 1584 17688 1636 17740
rect 1768 17731 1820 17740
rect 1768 17697 1777 17731
rect 1777 17697 1811 17731
rect 1811 17697 1820 17731
rect 1768 17688 1820 17697
rect 7380 17688 7432 17740
rect 8024 17688 8076 17740
rect 11336 17731 11388 17740
rect 11336 17697 11345 17731
rect 11345 17697 11379 17731
rect 11379 17697 11388 17731
rect 11336 17688 11388 17697
rect 13360 17688 13412 17740
rect 14372 17688 14424 17740
rect 15108 17731 15160 17740
rect 15108 17697 15117 17731
rect 15117 17697 15151 17731
rect 15151 17697 15160 17731
rect 15108 17688 15160 17697
rect 3148 17663 3200 17672
rect 3148 17629 3157 17663
rect 3157 17629 3191 17663
rect 3191 17629 3200 17663
rect 3148 17620 3200 17629
rect 7564 17663 7616 17672
rect 7564 17629 7573 17663
rect 7573 17629 7607 17663
rect 7607 17629 7616 17663
rect 7564 17620 7616 17629
rect 13728 17663 13780 17672
rect 13728 17629 13737 17663
rect 13737 17629 13771 17663
rect 13771 17629 13780 17663
rect 13728 17620 13780 17629
rect 14740 17552 14792 17604
rect 11888 17484 11940 17536
rect 13452 17484 13504 17536
rect 13636 17484 13688 17536
rect 14004 17484 14056 17536
rect 14924 17527 14976 17536
rect 14924 17493 14933 17527
rect 14933 17493 14967 17527
rect 14967 17493 14976 17527
rect 14924 17484 14976 17493
rect 16120 17527 16172 17536
rect 16120 17493 16129 17527
rect 16129 17493 16163 17527
rect 16163 17493 16172 17527
rect 16120 17484 16172 17493
rect 16396 17484 16448 17536
rect 4315 17382 4367 17434
rect 4379 17382 4431 17434
rect 4443 17382 4495 17434
rect 4507 17382 4559 17434
rect 10982 17382 11034 17434
rect 11046 17382 11098 17434
rect 11110 17382 11162 17434
rect 11174 17382 11226 17434
rect 17648 17382 17700 17434
rect 17712 17382 17764 17434
rect 17776 17382 17828 17434
rect 17840 17382 17892 17434
rect 1676 17280 1728 17332
rect 1860 17280 1912 17332
rect 9404 17323 9456 17332
rect 9404 17289 9413 17323
rect 9413 17289 9447 17323
rect 9447 17289 9456 17323
rect 9404 17280 9456 17289
rect 11336 17280 11388 17332
rect 1676 17144 1728 17196
rect 4160 17144 4212 17196
rect 4712 17187 4764 17196
rect 4712 17153 4721 17187
rect 4721 17153 4755 17187
rect 4755 17153 4764 17187
rect 4712 17144 4764 17153
rect 7564 17144 7616 17196
rect 12164 17212 12216 17264
rect 12440 17212 12492 17264
rect 12808 17187 12860 17196
rect 9680 17119 9732 17128
rect 9680 17085 9689 17119
rect 9689 17085 9723 17119
rect 9723 17085 9732 17119
rect 9680 17076 9732 17085
rect 8024 16940 8076 16992
rect 11060 16983 11112 16992
rect 11060 16949 11069 16983
rect 11069 16949 11103 16983
rect 11103 16949 11112 16983
rect 11060 16940 11112 16949
rect 11888 16940 11940 16992
rect 12440 17119 12492 17128
rect 12440 17085 12449 17119
rect 12449 17085 12483 17119
rect 12483 17085 12492 17119
rect 12808 17153 12817 17187
rect 12817 17153 12851 17187
rect 12851 17153 12860 17187
rect 12808 17144 12860 17153
rect 13360 17212 13412 17264
rect 15108 17212 15160 17264
rect 15568 17255 15620 17264
rect 15568 17221 15577 17255
rect 15577 17221 15611 17255
rect 15611 17221 15620 17255
rect 15568 17212 15620 17221
rect 14740 17187 14792 17196
rect 14740 17153 14749 17187
rect 14749 17153 14783 17187
rect 14783 17153 14792 17187
rect 14740 17144 14792 17153
rect 12440 17076 12492 17085
rect 15292 17076 15344 17128
rect 14372 17051 14424 17060
rect 14372 17017 14381 17051
rect 14381 17017 14415 17051
rect 14415 17017 14424 17051
rect 14372 17008 14424 17017
rect 14740 17008 14792 17060
rect 15660 17008 15712 17060
rect 16304 17076 16356 17128
rect 12256 16940 12308 16992
rect 12440 16940 12492 16992
rect 13728 16940 13780 16992
rect 7648 16838 7700 16890
rect 7712 16838 7764 16890
rect 7776 16838 7828 16890
rect 7840 16838 7892 16890
rect 14315 16838 14367 16890
rect 14379 16838 14431 16890
rect 14443 16838 14495 16890
rect 14507 16838 14559 16890
rect 1676 16779 1728 16788
rect 1676 16745 1685 16779
rect 1685 16745 1719 16779
rect 1719 16745 1728 16779
rect 1676 16736 1728 16745
rect 1768 16736 1820 16788
rect 4712 16779 4764 16788
rect 4712 16745 4721 16779
rect 4721 16745 4755 16779
rect 4755 16745 4764 16779
rect 4712 16736 4764 16745
rect 12440 16736 12492 16788
rect 12532 16736 12584 16788
rect 1584 16668 1636 16720
rect 2320 16711 2372 16720
rect 2320 16677 2329 16711
rect 2329 16677 2363 16711
rect 2363 16677 2372 16711
rect 2320 16668 2372 16677
rect 13360 16736 13412 16788
rect 16120 16779 16172 16788
rect 16120 16745 16129 16779
rect 16129 16745 16163 16779
rect 16163 16745 16172 16779
rect 16120 16736 16172 16745
rect 3056 16643 3108 16652
rect 3056 16609 3065 16643
rect 3065 16609 3099 16643
rect 3099 16609 3108 16643
rect 3056 16600 3108 16609
rect 4712 16600 4764 16652
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 13360 16600 13412 16652
rect 14188 16600 14240 16652
rect 16120 16643 16172 16652
rect 16120 16609 16129 16643
rect 16129 16609 16163 16643
rect 16163 16609 16172 16643
rect 16120 16600 16172 16609
rect 1860 16532 1912 16584
rect 2688 16532 2740 16584
rect 11796 16532 11848 16584
rect 15660 16575 15712 16584
rect 15660 16541 15669 16575
rect 15669 16541 15703 16575
rect 15703 16541 15712 16575
rect 15660 16532 15712 16541
rect 13820 16464 13872 16516
rect 15292 16507 15344 16516
rect 15292 16473 15301 16507
rect 15301 16473 15335 16507
rect 15335 16473 15344 16507
rect 15292 16464 15344 16473
rect 11612 16396 11664 16448
rect 13452 16439 13504 16448
rect 13452 16405 13461 16439
rect 13461 16405 13495 16439
rect 13495 16405 13504 16439
rect 13452 16396 13504 16405
rect 14924 16396 14976 16448
rect 4315 16294 4367 16346
rect 4379 16294 4431 16346
rect 4443 16294 4495 16346
rect 4507 16294 4559 16346
rect 10982 16294 11034 16346
rect 11046 16294 11098 16346
rect 11110 16294 11162 16346
rect 11174 16294 11226 16346
rect 17648 16294 17700 16346
rect 17712 16294 17764 16346
rect 17776 16294 17828 16346
rect 17840 16294 17892 16346
rect 3056 16192 3108 16244
rect 3976 16192 4028 16244
rect 10876 16192 10928 16244
rect 12808 16235 12860 16244
rect 12808 16201 12817 16235
rect 12817 16201 12851 16235
rect 12851 16201 12860 16235
rect 12808 16192 12860 16201
rect 13360 16192 13412 16244
rect 14188 16192 14240 16244
rect 1400 16056 1452 16108
rect 11336 16056 11388 16108
rect 1492 16031 1544 16040
rect 1492 15997 1501 16031
rect 1501 15997 1535 16031
rect 1535 15997 1544 16031
rect 1492 15988 1544 15997
rect 3148 16031 3200 16040
rect 3148 15997 3157 16031
rect 3157 15997 3191 16031
rect 3191 15997 3200 16031
rect 3148 15988 3200 15997
rect 4068 16031 4120 16040
rect 4068 15997 4077 16031
rect 4077 15997 4111 16031
rect 4111 15997 4120 16031
rect 4068 15988 4120 15997
rect 11612 15988 11664 16040
rect 15936 16124 15988 16176
rect 10876 15920 10928 15972
rect 12348 16056 12400 16108
rect 13728 16099 13780 16108
rect 13728 16065 13737 16099
rect 13737 16065 13771 16099
rect 13771 16065 13780 16099
rect 13728 16056 13780 16065
rect 15660 16056 15712 16108
rect 12808 15988 12860 16040
rect 15384 15988 15436 16040
rect 16396 16056 16448 16108
rect 5632 15895 5684 15904
rect 5632 15861 5641 15895
rect 5641 15861 5675 15895
rect 5675 15861 5684 15895
rect 5632 15852 5684 15861
rect 14924 15852 14976 15904
rect 16120 15852 16172 15904
rect 17040 15852 17092 15904
rect 7648 15750 7700 15802
rect 7712 15750 7764 15802
rect 7776 15750 7828 15802
rect 7840 15750 7892 15802
rect 14315 15750 14367 15802
rect 14379 15750 14431 15802
rect 14443 15750 14495 15802
rect 14507 15750 14559 15802
rect 1400 15648 1452 15700
rect 1492 15308 1544 15360
rect 2688 15308 2740 15360
rect 4068 15648 4120 15700
rect 10140 15648 10192 15700
rect 12532 15648 12584 15700
rect 15384 15691 15436 15700
rect 11428 15623 11480 15632
rect 11428 15589 11437 15623
rect 11437 15589 11471 15623
rect 11471 15589 11480 15623
rect 11428 15580 11480 15589
rect 3792 15555 3844 15564
rect 3792 15521 3801 15555
rect 3801 15521 3835 15555
rect 3835 15521 3844 15555
rect 3792 15512 3844 15521
rect 6920 15512 6972 15564
rect 7656 15512 7708 15564
rect 9864 15512 9916 15564
rect 12900 15512 12952 15564
rect 13820 15512 13872 15564
rect 15384 15657 15393 15691
rect 15393 15657 15427 15691
rect 15427 15657 15436 15691
rect 15384 15648 15436 15657
rect 15108 15512 15160 15564
rect 16212 15512 16264 15564
rect 16488 15555 16540 15564
rect 16488 15521 16497 15555
rect 16497 15521 16531 15555
rect 16531 15521 16540 15555
rect 16488 15512 16540 15521
rect 7564 15487 7616 15496
rect 7564 15453 7573 15487
rect 7573 15453 7607 15487
rect 7607 15453 7616 15487
rect 7564 15444 7616 15453
rect 9772 15487 9824 15496
rect 9772 15453 9781 15487
rect 9781 15453 9815 15487
rect 9815 15453 9824 15487
rect 9772 15444 9824 15453
rect 10232 15444 10284 15496
rect 14924 15487 14976 15496
rect 14924 15453 14933 15487
rect 14933 15453 14967 15487
rect 14967 15453 14976 15487
rect 14924 15444 14976 15453
rect 14280 15419 14332 15428
rect 14280 15385 14289 15419
rect 14289 15385 14323 15419
rect 14323 15385 14332 15419
rect 14280 15376 14332 15385
rect 15384 15376 15436 15428
rect 5080 15351 5132 15360
rect 5080 15317 5089 15351
rect 5089 15317 5123 15351
rect 5123 15317 5132 15351
rect 5080 15308 5132 15317
rect 11796 15351 11848 15360
rect 11796 15317 11805 15351
rect 11805 15317 11839 15351
rect 11839 15317 11848 15351
rect 11796 15308 11848 15317
rect 13452 15308 13504 15360
rect 15660 15351 15712 15360
rect 15660 15317 15669 15351
rect 15669 15317 15703 15351
rect 15703 15317 15712 15351
rect 15660 15308 15712 15317
rect 16304 15308 16356 15360
rect 16856 15351 16908 15360
rect 16856 15317 16865 15351
rect 16865 15317 16899 15351
rect 16899 15317 16908 15351
rect 16856 15308 16908 15317
rect 4315 15206 4367 15258
rect 4379 15206 4431 15258
rect 4443 15206 4495 15258
rect 4507 15206 4559 15258
rect 10982 15206 11034 15258
rect 11046 15206 11098 15258
rect 11110 15206 11162 15258
rect 11174 15206 11226 15258
rect 17648 15206 17700 15258
rect 17712 15206 17764 15258
rect 17776 15206 17828 15258
rect 17840 15206 17892 15258
rect 3792 15104 3844 15156
rect 4160 15104 4212 15156
rect 4712 15147 4764 15156
rect 4712 15113 4721 15147
rect 4721 15113 4755 15147
rect 4755 15113 4764 15147
rect 4712 15104 4764 15113
rect 7564 15104 7616 15156
rect 7656 15147 7708 15156
rect 7656 15113 7665 15147
rect 7665 15113 7699 15147
rect 7699 15113 7708 15147
rect 10876 15147 10928 15156
rect 7656 15104 7708 15113
rect 10876 15113 10885 15147
rect 10885 15113 10919 15147
rect 10919 15113 10928 15147
rect 10876 15104 10928 15113
rect 12900 15104 12952 15156
rect 13728 15147 13780 15156
rect 11704 15036 11756 15088
rect 12348 15011 12400 15020
rect 12348 14977 12357 15011
rect 12357 14977 12391 15011
rect 12391 14977 12400 15011
rect 12348 14968 12400 14977
rect 4896 14943 4948 14952
rect 4896 14909 4905 14943
rect 4905 14909 4939 14943
rect 4939 14909 4948 14943
rect 4896 14900 4948 14909
rect 10876 14900 10928 14952
rect 11796 14900 11848 14952
rect 13728 15113 13737 15147
rect 13737 15113 13771 15147
rect 13771 15113 13780 15147
rect 13728 15104 13780 15113
rect 15108 15147 15160 15156
rect 15108 15113 15117 15147
rect 15117 15113 15151 15147
rect 15151 15113 15160 15147
rect 15108 15104 15160 15113
rect 16488 15104 16540 15156
rect 16396 15079 16448 15088
rect 16396 15045 16405 15079
rect 16405 15045 16439 15079
rect 16439 15045 16448 15079
rect 16396 15036 16448 15045
rect 13728 14900 13780 14952
rect 16672 14900 16724 14952
rect 16948 14943 17000 14952
rect 9864 14807 9916 14816
rect 9864 14773 9873 14807
rect 9873 14773 9907 14807
rect 9907 14773 9916 14807
rect 9864 14764 9916 14773
rect 10232 14807 10284 14816
rect 10232 14773 10241 14807
rect 10241 14773 10275 14807
rect 10275 14773 10284 14807
rect 10232 14764 10284 14773
rect 14924 14832 14976 14884
rect 15108 14832 15160 14884
rect 16948 14909 16957 14943
rect 16957 14909 16991 14943
rect 16991 14909 17000 14943
rect 16948 14900 17000 14909
rect 16856 14832 16908 14884
rect 15292 14764 15344 14816
rect 15844 14764 15896 14816
rect 7648 14662 7700 14714
rect 7712 14662 7764 14714
rect 7776 14662 7828 14714
rect 7840 14662 7892 14714
rect 14315 14662 14367 14714
rect 14379 14662 14431 14714
rect 14443 14662 14495 14714
rect 14507 14662 14559 14714
rect 4896 14603 4948 14612
rect 4896 14569 4905 14603
rect 4905 14569 4939 14603
rect 4939 14569 4948 14603
rect 4896 14560 4948 14569
rect 12440 14560 12492 14612
rect 13360 14560 13412 14612
rect 15384 14603 15436 14612
rect 15384 14569 15393 14603
rect 15393 14569 15427 14603
rect 15427 14569 15436 14603
rect 15384 14560 15436 14569
rect 11704 14492 11756 14544
rect 12716 14535 12768 14544
rect 12716 14501 12725 14535
rect 12725 14501 12759 14535
rect 12759 14501 12768 14535
rect 12716 14492 12768 14501
rect 2320 14467 2372 14476
rect 2320 14433 2329 14467
rect 2329 14433 2363 14467
rect 2363 14433 2372 14467
rect 2320 14424 2372 14433
rect 2596 14467 2648 14476
rect 2596 14433 2605 14467
rect 2605 14433 2639 14467
rect 2639 14433 2648 14467
rect 2596 14424 2648 14433
rect 10692 14424 10744 14476
rect 13820 14424 13872 14476
rect 14464 14467 14516 14476
rect 14464 14433 14473 14467
rect 14473 14433 14507 14467
rect 14507 14433 14516 14467
rect 14464 14424 14516 14433
rect 14556 14424 14608 14476
rect 3976 14399 4028 14408
rect 3976 14365 3985 14399
rect 3985 14365 4019 14399
rect 4019 14365 4028 14399
rect 3976 14356 4028 14365
rect 14740 14356 14792 14408
rect 16488 14424 16540 14476
rect 16856 14467 16908 14476
rect 16856 14433 16865 14467
rect 16865 14433 16899 14467
rect 16899 14433 16908 14467
rect 16856 14424 16908 14433
rect 15016 14288 15068 14340
rect 16212 14331 16264 14340
rect 16212 14297 16221 14331
rect 16221 14297 16255 14331
rect 16255 14297 16264 14331
rect 16212 14288 16264 14297
rect 11704 14220 11756 14272
rect 12900 14220 12952 14272
rect 13820 14263 13872 14272
rect 13820 14229 13829 14263
rect 13829 14229 13863 14263
rect 13863 14229 13872 14263
rect 13820 14220 13872 14229
rect 4315 14118 4367 14170
rect 4379 14118 4431 14170
rect 4443 14118 4495 14170
rect 4507 14118 4559 14170
rect 10982 14118 11034 14170
rect 11046 14118 11098 14170
rect 11110 14118 11162 14170
rect 11174 14118 11226 14170
rect 17648 14118 17700 14170
rect 17712 14118 17764 14170
rect 17776 14118 17828 14170
rect 17840 14118 17892 14170
rect 2596 14016 2648 14068
rect 5632 14059 5684 14068
rect 5632 14025 5641 14059
rect 5641 14025 5675 14059
rect 5675 14025 5684 14059
rect 5632 14016 5684 14025
rect 7288 14059 7340 14068
rect 7288 14025 7297 14059
rect 7297 14025 7331 14059
rect 7331 14025 7340 14059
rect 7288 14016 7340 14025
rect 12164 14016 12216 14068
rect 14556 14016 14608 14068
rect 16304 14016 16356 14068
rect 16580 14016 16632 14068
rect 2320 13948 2372 14000
rect 12440 13948 12492 14000
rect 12716 13948 12768 14000
rect 14464 13991 14516 14000
rect 14464 13957 14473 13991
rect 14473 13957 14507 13991
rect 14507 13957 14516 13991
rect 14464 13948 14516 13957
rect 16764 13991 16816 14000
rect 16764 13957 16773 13991
rect 16773 13957 16807 13991
rect 16807 13957 16816 13991
rect 16764 13948 16816 13957
rect 5724 13855 5776 13864
rect 5724 13821 5733 13855
rect 5733 13821 5767 13855
rect 5767 13821 5776 13855
rect 5724 13812 5776 13821
rect 10692 13812 10744 13864
rect 12716 13812 12768 13864
rect 13268 13855 13320 13864
rect 13268 13821 13277 13855
rect 13277 13821 13311 13855
rect 13311 13821 13320 13855
rect 13268 13812 13320 13821
rect 13360 13855 13412 13864
rect 13360 13821 13369 13855
rect 13369 13821 13403 13855
rect 13403 13821 13412 13855
rect 13360 13812 13412 13821
rect 12624 13744 12676 13796
rect 15292 13855 15344 13864
rect 15292 13821 15301 13855
rect 15301 13821 15335 13855
rect 15335 13821 15344 13855
rect 15292 13812 15344 13821
rect 16488 13812 16540 13864
rect 16580 13812 16632 13864
rect 17408 13880 17460 13932
rect 17132 13855 17184 13864
rect 17132 13821 17141 13855
rect 17141 13821 17175 13855
rect 17175 13821 17184 13855
rect 17132 13812 17184 13821
rect 16856 13744 16908 13796
rect 10324 13719 10376 13728
rect 10324 13685 10333 13719
rect 10333 13685 10367 13719
rect 10367 13685 10376 13719
rect 10324 13676 10376 13685
rect 10876 13676 10928 13728
rect 12716 13676 12768 13728
rect 7648 13574 7700 13626
rect 7712 13574 7764 13626
rect 7776 13574 7828 13626
rect 7840 13574 7892 13626
rect 14315 13574 14367 13626
rect 14379 13574 14431 13626
rect 14443 13574 14495 13626
rect 14507 13574 14559 13626
rect 1492 13472 1544 13524
rect 2320 13472 2372 13524
rect 4896 13515 4948 13524
rect 4896 13481 4905 13515
rect 4905 13481 4939 13515
rect 4939 13481 4948 13515
rect 4896 13472 4948 13481
rect 5724 13515 5776 13524
rect 5724 13481 5733 13515
rect 5733 13481 5767 13515
rect 5767 13481 5776 13515
rect 5724 13472 5776 13481
rect 11336 13472 11388 13524
rect 12624 13472 12676 13524
rect 13176 13472 13228 13524
rect 16304 13472 16356 13524
rect 16856 13515 16908 13524
rect 16856 13481 16865 13515
rect 16865 13481 16899 13515
rect 16899 13481 16908 13515
rect 16856 13472 16908 13481
rect 12900 13404 12952 13456
rect 14924 13404 14976 13456
rect 2964 13379 3016 13388
rect 2964 13345 2973 13379
rect 2973 13345 3007 13379
rect 3007 13345 3016 13379
rect 2964 13336 3016 13345
rect 3240 13379 3292 13388
rect 3240 13345 3249 13379
rect 3249 13345 3283 13379
rect 3283 13345 3292 13379
rect 3240 13336 3292 13345
rect 7472 13336 7524 13388
rect 9496 13336 9548 13388
rect 10324 13379 10376 13388
rect 10324 13345 10333 13379
rect 10333 13345 10367 13379
rect 10367 13345 10376 13379
rect 10324 13336 10376 13345
rect 10876 13379 10928 13388
rect 10876 13345 10885 13379
rect 10885 13345 10919 13379
rect 10919 13345 10928 13379
rect 10876 13336 10928 13345
rect 11428 13336 11480 13388
rect 12808 13379 12860 13388
rect 4620 13311 4672 13320
rect 4620 13277 4629 13311
rect 4629 13277 4663 13311
rect 4663 13277 4672 13311
rect 4620 13268 4672 13277
rect 7840 13311 7892 13320
rect 7840 13277 7849 13311
rect 7849 13277 7883 13311
rect 7883 13277 7892 13311
rect 7840 13268 7892 13277
rect 12808 13345 12817 13379
rect 12817 13345 12851 13379
rect 12851 13345 12860 13379
rect 12808 13336 12860 13345
rect 13820 13336 13872 13388
rect 14372 13336 14424 13388
rect 12716 13268 12768 13320
rect 13452 13268 13504 13320
rect 14740 13311 14792 13320
rect 14740 13277 14749 13311
rect 14749 13277 14783 13311
rect 14783 13277 14792 13311
rect 14740 13268 14792 13277
rect 15844 13336 15896 13388
rect 12624 13243 12676 13252
rect 12624 13209 12633 13243
rect 12633 13209 12667 13243
rect 12667 13209 12676 13243
rect 12624 13200 12676 13209
rect 14188 13200 14240 13252
rect 15660 13200 15712 13252
rect 9772 13175 9824 13184
rect 9772 13141 9781 13175
rect 9781 13141 9815 13175
rect 9815 13141 9824 13175
rect 9772 13132 9824 13141
rect 13728 13132 13780 13184
rect 4315 13030 4367 13082
rect 4379 13030 4431 13082
rect 4443 13030 4495 13082
rect 4507 13030 4559 13082
rect 10982 13030 11034 13082
rect 11046 13030 11098 13082
rect 11110 13030 11162 13082
rect 11174 13030 11226 13082
rect 17648 13030 17700 13082
rect 17712 13030 17764 13082
rect 17776 13030 17828 13082
rect 17840 13030 17892 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 1676 12928 1728 12980
rect 2688 12928 2740 12980
rect 2964 12928 3016 12980
rect 3332 12971 3384 12980
rect 3332 12937 3341 12971
rect 3341 12937 3375 12971
rect 3375 12937 3384 12971
rect 3332 12928 3384 12937
rect 3792 12971 3844 12980
rect 3792 12937 3801 12971
rect 3801 12937 3835 12971
rect 3835 12937 3844 12971
rect 3792 12928 3844 12937
rect 5632 12971 5684 12980
rect 5632 12937 5641 12971
rect 5641 12937 5675 12971
rect 5675 12937 5684 12971
rect 5632 12928 5684 12937
rect 7472 12928 7524 12980
rect 7840 12928 7892 12980
rect 14372 12928 14424 12980
rect 15292 12928 15344 12980
rect 3240 12860 3292 12912
rect 7104 12860 7156 12912
rect 7564 12860 7616 12912
rect 12072 12860 12124 12912
rect 12256 12860 12308 12912
rect 15568 12903 15620 12912
rect 15568 12869 15577 12903
rect 15577 12869 15611 12903
rect 15611 12869 15620 12903
rect 15568 12860 15620 12869
rect 11520 12792 11572 12844
rect 11796 12835 11848 12844
rect 11796 12801 11805 12835
rect 11805 12801 11839 12835
rect 11839 12801 11848 12835
rect 11796 12792 11848 12801
rect 12808 12792 12860 12844
rect 15660 12792 15712 12844
rect 16304 12928 16356 12980
rect 16764 12928 16816 12980
rect 17132 12928 17184 12980
rect 4068 12767 4120 12776
rect 4068 12733 4077 12767
rect 4077 12733 4111 12767
rect 4111 12733 4120 12767
rect 4068 12724 4120 12733
rect 4804 12724 4856 12776
rect 9772 12724 9824 12776
rect 10876 12724 10928 12776
rect 12900 12767 12952 12776
rect 12900 12733 12909 12767
rect 12909 12733 12943 12767
rect 12943 12733 12952 12767
rect 12900 12724 12952 12733
rect 13084 12767 13136 12776
rect 13084 12733 13093 12767
rect 13093 12733 13127 12767
rect 13127 12733 13136 12767
rect 13084 12724 13136 12733
rect 13452 12767 13504 12776
rect 13452 12733 13461 12767
rect 13461 12733 13495 12767
rect 13495 12733 13504 12767
rect 13452 12724 13504 12733
rect 15384 12724 15436 12776
rect 16120 12767 16172 12776
rect 16120 12733 16129 12767
rect 16129 12733 16163 12767
rect 16163 12733 16172 12767
rect 16120 12724 16172 12733
rect 11520 12656 11572 12708
rect 13728 12699 13780 12708
rect 13728 12665 13737 12699
rect 13737 12665 13771 12699
rect 13771 12665 13780 12699
rect 13728 12656 13780 12665
rect 1952 12588 2004 12640
rect 10508 12588 10560 12640
rect 12624 12588 12676 12640
rect 16948 12631 17000 12640
rect 16948 12597 16957 12631
rect 16957 12597 16991 12631
rect 16991 12597 17000 12631
rect 16948 12588 17000 12597
rect 7648 12486 7700 12538
rect 7712 12486 7764 12538
rect 7776 12486 7828 12538
rect 7840 12486 7892 12538
rect 14315 12486 14367 12538
rect 14379 12486 14431 12538
rect 14443 12486 14495 12538
rect 14507 12486 14559 12538
rect 11336 12384 11388 12436
rect 3056 12359 3108 12368
rect 3056 12325 3065 12359
rect 3065 12325 3099 12359
rect 3099 12325 3108 12359
rect 3056 12316 3108 12325
rect 9220 12316 9272 12368
rect 10508 12359 10560 12368
rect 10508 12325 10517 12359
rect 10517 12325 10551 12359
rect 10551 12325 10560 12359
rect 10508 12316 10560 12325
rect 11704 12384 11756 12436
rect 11796 12384 11848 12436
rect 11980 12384 12032 12436
rect 12716 12384 12768 12436
rect 14924 12427 14976 12436
rect 14924 12393 14933 12427
rect 14933 12393 14967 12427
rect 14967 12393 14976 12427
rect 14924 12384 14976 12393
rect 12256 12359 12308 12368
rect 12256 12325 12265 12359
rect 12265 12325 12299 12359
rect 12299 12325 12308 12359
rect 12256 12316 12308 12325
rect 15936 12316 15988 12368
rect 1676 12291 1728 12300
rect 1676 12257 1685 12291
rect 1685 12257 1719 12291
rect 1719 12257 1728 12291
rect 1676 12248 1728 12257
rect 3792 12248 3844 12300
rect 6552 12248 6604 12300
rect 10140 12248 10192 12300
rect 11888 12248 11940 12300
rect 13268 12291 13320 12300
rect 13268 12257 13277 12291
rect 13277 12257 13311 12291
rect 13311 12257 13320 12291
rect 13268 12248 13320 12257
rect 13728 12291 13780 12300
rect 13728 12257 13737 12291
rect 13737 12257 13771 12291
rect 13771 12257 13780 12291
rect 13728 12248 13780 12257
rect 14188 12291 14240 12300
rect 14188 12257 14197 12291
rect 14197 12257 14231 12291
rect 14231 12257 14240 12291
rect 14188 12248 14240 12257
rect 1860 12180 1912 12232
rect 7012 12180 7064 12232
rect 11244 12180 11296 12232
rect 10508 12112 10560 12164
rect 13544 12180 13596 12232
rect 13820 12223 13872 12232
rect 13820 12189 13829 12223
rect 13829 12189 13863 12223
rect 13863 12189 13872 12223
rect 13820 12180 13872 12189
rect 14004 12180 14056 12232
rect 15752 12248 15804 12300
rect 16580 12291 16632 12300
rect 16580 12257 16589 12291
rect 16589 12257 16623 12291
rect 16623 12257 16632 12291
rect 16580 12248 16632 12257
rect 16764 12291 16816 12300
rect 16764 12257 16773 12291
rect 16773 12257 16807 12291
rect 16807 12257 16816 12291
rect 16764 12248 16816 12257
rect 17316 12248 17368 12300
rect 15936 12180 15988 12232
rect 16028 12180 16080 12232
rect 16396 12155 16448 12164
rect 16396 12121 16405 12155
rect 16405 12121 16439 12155
rect 16439 12121 16448 12155
rect 16396 12112 16448 12121
rect 4068 12087 4120 12096
rect 4068 12053 4077 12087
rect 4077 12053 4111 12087
rect 4111 12053 4120 12087
rect 4068 12044 4120 12053
rect 5816 12087 5868 12096
rect 5816 12053 5825 12087
rect 5825 12053 5859 12087
rect 5859 12053 5868 12087
rect 5816 12044 5868 12053
rect 11428 12044 11480 12096
rect 11612 12044 11664 12096
rect 12716 12087 12768 12096
rect 12716 12053 12725 12087
rect 12725 12053 12759 12087
rect 12759 12053 12768 12087
rect 12716 12044 12768 12053
rect 13084 12044 13136 12096
rect 14188 12044 14240 12096
rect 14740 12044 14792 12096
rect 14832 12044 14884 12096
rect 15292 12044 15344 12096
rect 15752 12044 15804 12096
rect 4315 11942 4367 11994
rect 4379 11942 4431 11994
rect 4443 11942 4495 11994
rect 4507 11942 4559 11994
rect 10982 11942 11034 11994
rect 11046 11942 11098 11994
rect 11110 11942 11162 11994
rect 11174 11942 11226 11994
rect 17648 11942 17700 11994
rect 17712 11942 17764 11994
rect 17776 11942 17828 11994
rect 17840 11942 17892 11994
rect 2964 11883 3016 11892
rect 2964 11849 2973 11883
rect 2973 11849 3007 11883
rect 3007 11849 3016 11883
rect 2964 11840 3016 11849
rect 3792 11883 3844 11892
rect 3792 11849 3801 11883
rect 3801 11849 3835 11883
rect 3835 11849 3844 11883
rect 3792 11840 3844 11849
rect 5908 11883 5960 11892
rect 5908 11849 5917 11883
rect 5917 11849 5951 11883
rect 5951 11849 5960 11883
rect 5908 11840 5960 11849
rect 8484 11883 8536 11892
rect 8484 11849 8493 11883
rect 8493 11849 8527 11883
rect 8527 11849 8536 11883
rect 8484 11840 8536 11849
rect 10508 11883 10560 11892
rect 10508 11849 10517 11883
rect 10517 11849 10551 11883
rect 10551 11849 10560 11883
rect 10508 11840 10560 11849
rect 13268 11840 13320 11892
rect 14740 11840 14792 11892
rect 16580 11840 16632 11892
rect 13636 11815 13688 11824
rect 13636 11781 13645 11815
rect 13645 11781 13679 11815
rect 13679 11781 13688 11815
rect 13636 11772 13688 11781
rect 16672 11772 16724 11824
rect 1584 11704 1636 11756
rect 9312 11704 9364 11756
rect 9588 11704 9640 11756
rect 11060 11747 11112 11756
rect 11060 11713 11069 11747
rect 11069 11713 11103 11747
rect 11103 11713 11112 11747
rect 11060 11704 11112 11713
rect 13728 11704 13780 11756
rect 15108 11704 15160 11756
rect 15660 11704 15712 11756
rect 1492 11636 1544 11688
rect 4068 11636 4120 11688
rect 3424 11543 3476 11552
rect 3424 11509 3433 11543
rect 3433 11509 3467 11543
rect 3467 11509 3476 11543
rect 7104 11679 7156 11688
rect 7104 11645 7113 11679
rect 7113 11645 7147 11679
rect 7147 11645 7156 11679
rect 7104 11636 7156 11645
rect 6552 11543 6604 11552
rect 3424 11500 3476 11509
rect 6552 11509 6561 11543
rect 6561 11509 6595 11543
rect 6595 11509 6604 11543
rect 6552 11500 6604 11509
rect 6920 11543 6972 11552
rect 6920 11509 6929 11543
rect 6929 11509 6963 11543
rect 6963 11509 6972 11543
rect 10140 11679 10192 11688
rect 10140 11645 10149 11679
rect 10149 11645 10183 11679
rect 10183 11645 10192 11679
rect 10140 11636 10192 11645
rect 6920 11500 6972 11509
rect 10692 11500 10744 11552
rect 11428 11636 11480 11688
rect 11796 11636 11848 11688
rect 13820 11679 13872 11688
rect 13820 11645 13829 11679
rect 13829 11645 13863 11679
rect 13863 11645 13872 11679
rect 13820 11636 13872 11645
rect 14188 11679 14240 11688
rect 14188 11645 14197 11679
rect 14197 11645 14231 11679
rect 14231 11645 14240 11679
rect 14188 11636 14240 11645
rect 14280 11679 14332 11688
rect 14280 11645 14289 11679
rect 14289 11645 14323 11679
rect 14323 11645 14332 11679
rect 14280 11636 14332 11645
rect 14832 11636 14884 11688
rect 15752 11679 15804 11688
rect 15752 11645 15761 11679
rect 15761 11645 15795 11679
rect 15795 11645 15804 11679
rect 15752 11636 15804 11645
rect 15936 11679 15988 11688
rect 15936 11645 15945 11679
rect 15945 11645 15979 11679
rect 15979 11645 15988 11679
rect 15936 11636 15988 11645
rect 16304 11636 16356 11688
rect 11888 11568 11940 11620
rect 11704 11500 11756 11552
rect 12716 11500 12768 11552
rect 14004 11500 14056 11552
rect 15108 11543 15160 11552
rect 15108 11509 15117 11543
rect 15117 11509 15151 11543
rect 15151 11509 15160 11543
rect 15108 11500 15160 11509
rect 17316 11543 17368 11552
rect 17316 11509 17325 11543
rect 17325 11509 17359 11543
rect 17359 11509 17368 11543
rect 17316 11500 17368 11509
rect 7648 11398 7700 11450
rect 7712 11398 7764 11450
rect 7776 11398 7828 11450
rect 7840 11398 7892 11450
rect 14315 11398 14367 11450
rect 14379 11398 14431 11450
rect 14443 11398 14495 11450
rect 14507 11398 14559 11450
rect 8116 11339 8168 11348
rect 8116 11305 8125 11339
rect 8125 11305 8159 11339
rect 8159 11305 8168 11339
rect 8116 11296 8168 11305
rect 12256 11339 12308 11348
rect 12256 11305 12265 11339
rect 12265 11305 12299 11339
rect 12299 11305 12308 11339
rect 12256 11296 12308 11305
rect 14096 11296 14148 11348
rect 6552 11228 6604 11280
rect 11796 11271 11848 11280
rect 1768 11203 1820 11212
rect 1768 11169 1777 11203
rect 1777 11169 1811 11203
rect 1811 11169 1820 11203
rect 1768 11160 1820 11169
rect 2228 11160 2280 11212
rect 3792 11160 3844 11212
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 10140 11160 10192 11212
rect 11796 11237 11805 11271
rect 11805 11237 11839 11271
rect 11839 11237 11848 11271
rect 11796 11228 11848 11237
rect 11888 11228 11940 11280
rect 14832 11296 14884 11348
rect 16764 11296 16816 11348
rect 1952 11092 2004 11144
rect 9680 11092 9732 11144
rect 11980 11160 12032 11212
rect 7104 11024 7156 11076
rect 3792 10956 3844 11008
rect 4068 10999 4120 11008
rect 4068 10965 4077 10999
rect 4077 10965 4111 10999
rect 4111 10965 4120 10999
rect 4068 10956 4120 10965
rect 10048 11024 10100 11076
rect 11244 11092 11296 11144
rect 11428 11092 11480 11144
rect 12072 11092 12124 11144
rect 12716 11092 12768 11144
rect 13544 11160 13596 11212
rect 15292 11160 15344 11212
rect 14188 11135 14240 11144
rect 14188 11101 14197 11135
rect 14197 11101 14231 11135
rect 14231 11101 14240 11135
rect 14188 11092 14240 11101
rect 15476 11092 15528 11144
rect 9772 10956 9824 11008
rect 10140 10999 10192 11008
rect 10140 10965 10149 10999
rect 10149 10965 10183 10999
rect 10183 10965 10192 10999
rect 10140 10956 10192 10965
rect 11336 11024 11388 11076
rect 13728 10956 13780 11008
rect 16396 10956 16448 11008
rect 4315 10854 4367 10906
rect 4379 10854 4431 10906
rect 4443 10854 4495 10906
rect 4507 10854 4559 10906
rect 10982 10854 11034 10906
rect 11046 10854 11098 10906
rect 11110 10854 11162 10906
rect 11174 10854 11226 10906
rect 17648 10854 17700 10906
rect 17712 10854 17764 10906
rect 17776 10854 17828 10906
rect 17840 10854 17892 10906
rect 3332 10795 3384 10804
rect 3332 10761 3341 10795
rect 3341 10761 3375 10795
rect 3375 10761 3384 10795
rect 3332 10752 3384 10761
rect 3792 10795 3844 10804
rect 3792 10761 3801 10795
rect 3801 10761 3835 10795
rect 3835 10761 3844 10795
rect 3792 10752 3844 10761
rect 6920 10752 6972 10804
rect 9680 10752 9732 10804
rect 11888 10752 11940 10804
rect 12440 10752 12492 10804
rect 13544 10752 13596 10804
rect 14740 10795 14792 10804
rect 14740 10761 14749 10795
rect 14749 10761 14783 10795
rect 14783 10761 14792 10795
rect 14740 10752 14792 10761
rect 16580 10727 16632 10736
rect 16580 10693 16589 10727
rect 16589 10693 16623 10727
rect 16623 10693 16632 10727
rect 16580 10684 16632 10693
rect 2044 10616 2096 10668
rect 2412 10616 2464 10668
rect 4252 10616 4304 10668
rect 8760 10659 8812 10668
rect 8760 10625 8769 10659
rect 8769 10625 8803 10659
rect 8803 10625 8812 10659
rect 8760 10616 8812 10625
rect 13912 10659 13964 10668
rect 13912 10625 13921 10659
rect 13921 10625 13955 10659
rect 13955 10625 13964 10659
rect 13912 10616 13964 10625
rect 16212 10616 16264 10668
rect 1492 10548 1544 10600
rect 4068 10548 4120 10600
rect 4436 10548 4488 10600
rect 8024 10591 8076 10600
rect 8024 10557 8033 10591
rect 8033 10557 8067 10591
rect 8067 10557 8076 10591
rect 8024 10548 8076 10557
rect 8116 10548 8168 10600
rect 8392 10548 8444 10600
rect 9680 10591 9732 10600
rect 9680 10557 9689 10591
rect 9689 10557 9723 10591
rect 9723 10557 9732 10591
rect 9680 10548 9732 10557
rect 9404 10523 9456 10532
rect 9404 10489 9413 10523
rect 9413 10489 9447 10523
rect 9447 10489 9456 10523
rect 11612 10548 11664 10600
rect 13268 10548 13320 10600
rect 13820 10591 13872 10600
rect 13820 10557 13829 10591
rect 13829 10557 13863 10591
rect 13863 10557 13872 10591
rect 13820 10548 13872 10557
rect 14096 10548 14148 10600
rect 9404 10480 9456 10489
rect 13728 10480 13780 10532
rect 8024 10412 8076 10464
rect 14924 10412 14976 10464
rect 15936 10548 15988 10600
rect 16304 10548 16356 10600
rect 7648 10310 7700 10362
rect 7712 10310 7764 10362
rect 7776 10310 7828 10362
rect 7840 10310 7892 10362
rect 14315 10310 14367 10362
rect 14379 10310 14431 10362
rect 14443 10310 14495 10362
rect 14507 10310 14559 10362
rect 4252 10208 4304 10260
rect 11336 10251 11388 10260
rect 11336 10217 11345 10251
rect 11345 10217 11379 10251
rect 11379 10217 11388 10251
rect 11336 10208 11388 10217
rect 11520 10208 11572 10260
rect 12256 10251 12308 10260
rect 12256 10217 12265 10251
rect 12265 10217 12299 10251
rect 12299 10217 12308 10251
rect 12256 10208 12308 10217
rect 12716 10251 12768 10260
rect 12716 10217 12725 10251
rect 12725 10217 12759 10251
rect 12759 10217 12768 10251
rect 12716 10208 12768 10217
rect 13820 10208 13872 10260
rect 16396 10251 16448 10260
rect 16396 10217 16405 10251
rect 16405 10217 16439 10251
rect 16439 10217 16448 10251
rect 16396 10208 16448 10217
rect 16580 10208 16632 10260
rect 3148 10183 3200 10192
rect 3148 10149 3157 10183
rect 3157 10149 3191 10183
rect 3191 10149 3200 10183
rect 3148 10140 3200 10149
rect 4436 10140 4488 10192
rect 8116 10140 8168 10192
rect 8484 10183 8536 10192
rect 8484 10149 8493 10183
rect 8493 10149 8527 10183
rect 8527 10149 8536 10183
rect 8484 10140 8536 10149
rect 13360 10140 13412 10192
rect 1216 10072 1268 10124
rect 2228 10072 2280 10124
rect 8208 10072 8260 10124
rect 9588 10115 9640 10124
rect 9588 10081 9597 10115
rect 9597 10081 9631 10115
rect 9631 10081 9640 10115
rect 9588 10072 9640 10081
rect 12164 10072 12216 10124
rect 12900 10115 12952 10124
rect 12900 10081 12909 10115
rect 12909 10081 12943 10115
rect 12943 10081 12952 10115
rect 12900 10072 12952 10081
rect 14004 10115 14056 10124
rect 14004 10081 14013 10115
rect 14013 10081 14047 10115
rect 14047 10081 14056 10115
rect 14004 10072 14056 10081
rect 16212 10140 16264 10192
rect 15016 10072 15068 10124
rect 15292 10115 15344 10124
rect 15292 10081 15301 10115
rect 15301 10081 15335 10115
rect 15335 10081 15344 10115
rect 15292 10072 15344 10081
rect 1492 10047 1544 10056
rect 1492 10013 1501 10047
rect 1501 10013 1535 10047
rect 1535 10013 1544 10047
rect 1492 10004 1544 10013
rect 9496 10004 9548 10056
rect 14740 10004 14792 10056
rect 15844 10072 15896 10124
rect 7840 9868 7892 9920
rect 10876 9911 10928 9920
rect 10876 9877 10885 9911
rect 10885 9877 10919 9911
rect 10919 9877 10928 9911
rect 10876 9868 10928 9877
rect 11888 9911 11940 9920
rect 11888 9877 11897 9911
rect 11897 9877 11931 9911
rect 11931 9877 11940 9911
rect 11888 9868 11940 9877
rect 12716 9868 12768 9920
rect 14096 9936 14148 9988
rect 13820 9911 13872 9920
rect 13820 9877 13829 9911
rect 13829 9877 13863 9911
rect 13863 9877 13872 9911
rect 13820 9868 13872 9877
rect 15200 9868 15252 9920
rect 16304 9868 16356 9920
rect 4315 9766 4367 9818
rect 4379 9766 4431 9818
rect 4443 9766 4495 9818
rect 4507 9766 4559 9818
rect 10982 9766 11034 9818
rect 11046 9766 11098 9818
rect 11110 9766 11162 9818
rect 11174 9766 11226 9818
rect 17648 9766 17700 9818
rect 17712 9766 17764 9818
rect 17776 9766 17828 9818
rect 17840 9766 17892 9818
rect 2044 9707 2096 9716
rect 2044 9673 2053 9707
rect 2053 9673 2087 9707
rect 2087 9673 2096 9707
rect 2044 9664 2096 9673
rect 2228 9664 2280 9716
rect 8116 9707 8168 9716
rect 8116 9673 8125 9707
rect 8125 9673 8159 9707
rect 8159 9673 8168 9707
rect 8116 9664 8168 9673
rect 8392 9664 8444 9716
rect 11428 9664 11480 9716
rect 11980 9664 12032 9716
rect 12900 9707 12952 9716
rect 12900 9673 12909 9707
rect 12909 9673 12943 9707
rect 12943 9673 12952 9707
rect 12900 9664 12952 9673
rect 1768 9596 1820 9648
rect 9588 9596 9640 9648
rect 11336 9596 11388 9648
rect 12440 9596 12492 9648
rect 15292 9664 15344 9716
rect 15568 9596 15620 9648
rect 17040 9596 17092 9648
rect 9496 9528 9548 9580
rect 7840 9503 7892 9512
rect 7840 9469 7849 9503
rect 7849 9469 7883 9503
rect 7883 9469 7892 9503
rect 7840 9460 7892 9469
rect 11428 9503 11480 9512
rect 11428 9469 11437 9503
rect 11437 9469 11471 9503
rect 11471 9469 11480 9503
rect 11428 9460 11480 9469
rect 11520 9503 11572 9512
rect 11520 9469 11529 9503
rect 11529 9469 11563 9503
rect 11563 9469 11572 9503
rect 11520 9460 11572 9469
rect 12348 9460 12400 9512
rect 15108 9528 15160 9580
rect 16304 9528 16356 9580
rect 13268 9460 13320 9512
rect 14096 9460 14148 9512
rect 14740 9460 14792 9512
rect 15016 9460 15068 9512
rect 16580 9460 16632 9512
rect 13820 9392 13872 9444
rect 15200 9392 15252 9444
rect 16396 9392 16448 9444
rect 16672 9392 16724 9444
rect 8208 9324 8260 9376
rect 8576 9367 8628 9376
rect 8576 9333 8585 9367
rect 8585 9333 8619 9367
rect 8619 9333 8628 9367
rect 8576 9324 8628 9333
rect 10048 9367 10100 9376
rect 10048 9333 10057 9367
rect 10057 9333 10091 9367
rect 10091 9333 10100 9367
rect 10048 9324 10100 9333
rect 11336 9324 11388 9376
rect 16304 9367 16356 9376
rect 16304 9333 16313 9367
rect 16313 9333 16347 9367
rect 16347 9333 16356 9367
rect 16304 9324 16356 9333
rect 7648 9222 7700 9274
rect 7712 9222 7764 9274
rect 7776 9222 7828 9274
rect 7840 9222 7892 9274
rect 14315 9222 14367 9274
rect 14379 9222 14431 9274
rect 14443 9222 14495 9274
rect 14507 9222 14559 9274
rect 1492 9120 1544 9172
rect 1676 9120 1728 9172
rect 1952 9163 2004 9172
rect 1952 9129 1961 9163
rect 1961 9129 1995 9163
rect 1995 9129 2004 9163
rect 1952 9120 2004 9129
rect 11428 9120 11480 9172
rect 13820 9163 13872 9172
rect 13820 9129 13829 9163
rect 13829 9129 13863 9163
rect 13863 9129 13872 9163
rect 13820 9120 13872 9129
rect 14096 9120 14148 9172
rect 11152 9095 11204 9104
rect 11152 9061 11161 9095
rect 11161 9061 11195 9095
rect 11195 9061 11204 9095
rect 11152 9052 11204 9061
rect 12348 9052 12400 9104
rect 9496 9027 9548 9036
rect 9496 8993 9505 9027
rect 9505 8993 9539 9027
rect 9539 8993 9548 9027
rect 9496 8984 9548 8993
rect 9772 9027 9824 9036
rect 9772 8993 9781 9027
rect 9781 8993 9815 9027
rect 9815 8993 9824 9027
rect 9772 8984 9824 8993
rect 12624 9027 12676 9036
rect 12624 8993 12633 9027
rect 12633 8993 12667 9027
rect 12667 8993 12676 9027
rect 12624 8984 12676 8993
rect 12992 9027 13044 9036
rect 12992 8993 13001 9027
rect 13001 8993 13035 9027
rect 13035 8993 13044 9027
rect 12992 8984 13044 8993
rect 13268 9027 13320 9036
rect 13268 8993 13277 9027
rect 13277 8993 13311 9027
rect 13311 8993 13320 9027
rect 13268 8984 13320 8993
rect 13912 8984 13964 9036
rect 16212 9095 16264 9104
rect 16212 9061 16221 9095
rect 16221 9061 16255 9095
rect 16255 9061 16264 9095
rect 16212 9052 16264 9061
rect 15200 9027 15252 9036
rect 15200 8993 15209 9027
rect 15209 8993 15243 9027
rect 15243 8993 15252 9027
rect 15200 8984 15252 8993
rect 16304 9027 16356 9036
rect 16304 8993 16313 9027
rect 16313 8993 16347 9027
rect 16347 8993 16356 9027
rect 16304 8984 16356 8993
rect 15108 8916 15160 8968
rect 15660 8916 15712 8968
rect 13176 8848 13228 8900
rect 15200 8848 15252 8900
rect 15844 8780 15896 8832
rect 4315 8678 4367 8730
rect 4379 8678 4431 8730
rect 4443 8678 4495 8730
rect 4507 8678 4559 8730
rect 10982 8678 11034 8730
rect 11046 8678 11098 8730
rect 11110 8678 11162 8730
rect 11174 8678 11226 8730
rect 17648 8678 17700 8730
rect 17712 8678 17764 8730
rect 17776 8678 17828 8730
rect 17840 8678 17892 8730
rect 9772 8576 9824 8628
rect 11336 8619 11388 8628
rect 11336 8585 11345 8619
rect 11345 8585 11379 8619
rect 11379 8585 11388 8619
rect 11336 8576 11388 8585
rect 11520 8619 11572 8628
rect 11520 8585 11529 8619
rect 11529 8585 11563 8619
rect 11563 8585 11572 8619
rect 11520 8576 11572 8585
rect 12440 8576 12492 8628
rect 13268 8576 13320 8628
rect 14004 8576 14056 8628
rect 15108 8619 15160 8628
rect 15108 8585 15117 8619
rect 15117 8585 15151 8619
rect 15151 8585 15160 8619
rect 15108 8576 15160 8585
rect 16396 8576 16448 8628
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 9496 8440 9548 8492
rect 10600 8483 10652 8492
rect 10600 8449 10609 8483
rect 10609 8449 10643 8483
rect 10643 8449 10652 8483
rect 10600 8440 10652 8449
rect 10508 8415 10560 8424
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 11612 8440 11664 8492
rect 12072 8415 12124 8424
rect 12072 8381 12081 8415
rect 12081 8381 12115 8415
rect 12115 8381 12124 8415
rect 12072 8372 12124 8381
rect 12348 8415 12400 8424
rect 12348 8381 12357 8415
rect 12357 8381 12391 8415
rect 12391 8381 12400 8415
rect 12348 8372 12400 8381
rect 12992 8508 13044 8560
rect 15568 8551 15620 8560
rect 15568 8517 15577 8551
rect 15577 8517 15611 8551
rect 15611 8517 15620 8551
rect 15568 8508 15620 8517
rect 15660 8440 15712 8492
rect 14832 8372 14884 8424
rect 15844 8372 15896 8424
rect 12624 8304 12676 8356
rect 13360 8304 13412 8356
rect 15660 8304 15712 8356
rect 7648 8134 7700 8186
rect 7712 8134 7764 8186
rect 7776 8134 7828 8186
rect 7840 8134 7892 8186
rect 14315 8134 14367 8186
rect 14379 8134 14431 8186
rect 14443 8134 14495 8186
rect 14507 8134 14559 8186
rect 12072 8032 12124 8084
rect 14740 8032 14792 8084
rect 15384 8032 15436 8084
rect 11336 7964 11388 8016
rect 11796 7964 11848 8016
rect 12808 7964 12860 8016
rect 8760 7939 8812 7948
rect 8760 7905 8769 7939
rect 8769 7905 8803 7939
rect 8803 7905 8812 7939
rect 8760 7896 8812 7905
rect 8852 7896 8904 7948
rect 11980 7896 12032 7948
rect 14188 7896 14240 7948
rect 14740 7896 14792 7948
rect 15016 7964 15068 8016
rect 15292 7896 15344 7948
rect 12440 7871 12492 7880
rect 12440 7837 12449 7871
rect 12449 7837 12483 7871
rect 12483 7837 12492 7871
rect 12440 7828 12492 7837
rect 12716 7828 12768 7880
rect 15016 7871 15068 7880
rect 15016 7837 15025 7871
rect 15025 7837 15059 7871
rect 15059 7837 15068 7871
rect 15016 7828 15068 7837
rect 15660 7828 15712 7880
rect 16304 7828 16356 7880
rect 13820 7760 13872 7812
rect 10324 7735 10376 7744
rect 10324 7701 10333 7735
rect 10333 7701 10367 7735
rect 10367 7701 10376 7735
rect 10324 7692 10376 7701
rect 4315 7590 4367 7642
rect 4379 7590 4431 7642
rect 4443 7590 4495 7642
rect 4507 7590 4559 7642
rect 10982 7590 11034 7642
rect 11046 7590 11098 7642
rect 11110 7590 11162 7642
rect 11174 7590 11226 7642
rect 17648 7590 17700 7642
rect 17712 7590 17764 7642
rect 17776 7590 17828 7642
rect 17840 7590 17892 7642
rect 8668 7488 8720 7540
rect 9588 7488 9640 7540
rect 10692 7488 10744 7540
rect 12808 7531 12860 7540
rect 8760 7463 8812 7472
rect 8760 7429 8769 7463
rect 8769 7429 8803 7463
rect 8803 7429 8812 7463
rect 8760 7420 8812 7429
rect 12808 7497 12817 7531
rect 12817 7497 12851 7531
rect 12851 7497 12860 7531
rect 12808 7488 12860 7497
rect 11520 7420 11572 7472
rect 10324 7352 10376 7404
rect 13176 7352 13228 7404
rect 14924 7352 14976 7404
rect 16488 7395 16540 7404
rect 5632 7327 5684 7336
rect 5632 7293 5641 7327
rect 5641 7293 5675 7327
rect 5675 7293 5684 7327
rect 5632 7284 5684 7293
rect 5540 7191 5592 7200
rect 5540 7157 5549 7191
rect 5549 7157 5583 7191
rect 5583 7157 5592 7191
rect 11336 7284 11388 7336
rect 11428 7284 11480 7336
rect 13360 7327 13412 7336
rect 13360 7293 13369 7327
rect 13369 7293 13403 7327
rect 13403 7293 13412 7327
rect 13360 7284 13412 7293
rect 13820 7327 13872 7336
rect 13820 7293 13829 7327
rect 13829 7293 13863 7327
rect 13863 7293 13872 7327
rect 13820 7284 13872 7293
rect 15108 7284 15160 7336
rect 16488 7361 16497 7395
rect 16497 7361 16531 7395
rect 16531 7361 16540 7395
rect 16488 7352 16540 7361
rect 16212 7327 16264 7336
rect 7288 7259 7340 7268
rect 7288 7225 7297 7259
rect 7297 7225 7331 7259
rect 7331 7225 7340 7259
rect 7288 7216 7340 7225
rect 11796 7216 11848 7268
rect 15292 7216 15344 7268
rect 16212 7293 16221 7327
rect 16221 7293 16255 7327
rect 16255 7293 16264 7327
rect 16212 7284 16264 7293
rect 5540 7148 5592 7157
rect 7648 7046 7700 7098
rect 7712 7046 7764 7098
rect 7776 7046 7828 7098
rect 7840 7046 7892 7098
rect 14315 7046 14367 7098
rect 14379 7046 14431 7098
rect 14443 7046 14495 7098
rect 14507 7046 14559 7098
rect 5724 6987 5776 6996
rect 5724 6953 5733 6987
rect 5733 6953 5767 6987
rect 5767 6953 5776 6987
rect 5724 6944 5776 6953
rect 12716 6987 12768 6996
rect 12716 6953 12725 6987
rect 12725 6953 12759 6987
rect 12759 6953 12768 6987
rect 12716 6944 12768 6953
rect 13360 6944 13412 6996
rect 13268 6876 13320 6928
rect 10140 6851 10192 6860
rect 10140 6817 10149 6851
rect 10149 6817 10183 6851
rect 10183 6817 10192 6851
rect 10140 6808 10192 6817
rect 12164 6808 12216 6860
rect 14924 6876 14976 6928
rect 15384 6876 15436 6928
rect 9680 6740 9732 6792
rect 10232 6740 10284 6792
rect 11980 6672 12032 6724
rect 15844 6808 15896 6860
rect 16948 6851 17000 6860
rect 16948 6817 16957 6851
rect 16957 6817 16991 6851
rect 16991 6817 17000 6851
rect 16948 6808 17000 6817
rect 17408 6808 17460 6860
rect 13912 6783 13964 6792
rect 13912 6749 13921 6783
rect 13921 6749 13955 6783
rect 13955 6749 13964 6783
rect 13912 6740 13964 6749
rect 17040 6783 17092 6792
rect 17040 6749 17049 6783
rect 17049 6749 17083 6783
rect 17083 6749 17092 6783
rect 17040 6740 17092 6749
rect 13820 6672 13872 6724
rect 14740 6672 14792 6724
rect 15200 6672 15252 6724
rect 16212 6672 16264 6724
rect 16488 6672 16540 6724
rect 17408 6715 17460 6724
rect 17408 6681 17417 6715
rect 17417 6681 17451 6715
rect 17451 6681 17460 6715
rect 17408 6672 17460 6681
rect 15292 6604 15344 6656
rect 4315 6502 4367 6554
rect 4379 6502 4431 6554
rect 4443 6502 4495 6554
rect 4507 6502 4559 6554
rect 10982 6502 11034 6554
rect 11046 6502 11098 6554
rect 11110 6502 11162 6554
rect 11174 6502 11226 6554
rect 17648 6502 17700 6554
rect 17712 6502 17764 6554
rect 17776 6502 17828 6554
rect 17840 6502 17892 6554
rect 10140 6400 10192 6452
rect 10232 6443 10284 6452
rect 10232 6409 10241 6443
rect 10241 6409 10275 6443
rect 10275 6409 10284 6443
rect 10232 6400 10284 6409
rect 10784 6400 10836 6452
rect 11520 6400 11572 6452
rect 13176 6443 13228 6452
rect 13176 6409 13185 6443
rect 13185 6409 13219 6443
rect 13219 6409 13228 6443
rect 13176 6400 13228 6409
rect 14188 6400 14240 6452
rect 15844 6443 15896 6452
rect 15844 6409 15853 6443
rect 15853 6409 15887 6443
rect 15887 6409 15896 6443
rect 15844 6400 15896 6409
rect 16948 6400 17000 6452
rect 13636 6375 13688 6384
rect 11612 6307 11664 6316
rect 11612 6273 11621 6307
rect 11621 6273 11655 6307
rect 11655 6273 11664 6307
rect 11612 6264 11664 6273
rect 13636 6341 13645 6375
rect 13645 6341 13679 6375
rect 13679 6341 13688 6375
rect 13636 6332 13688 6341
rect 14740 6375 14792 6384
rect 14740 6341 14749 6375
rect 14749 6341 14783 6375
rect 14783 6341 14792 6375
rect 14740 6332 14792 6341
rect 17040 6375 17092 6384
rect 17040 6341 17049 6375
rect 17049 6341 17083 6375
rect 17083 6341 17092 6375
rect 17040 6332 17092 6341
rect 11704 6196 11756 6248
rect 14648 6264 14700 6316
rect 17132 6264 17184 6316
rect 14004 6239 14056 6248
rect 14004 6205 14013 6239
rect 14013 6205 14047 6239
rect 14047 6205 14056 6239
rect 14004 6196 14056 6205
rect 13268 6128 13320 6180
rect 16764 6196 16816 6248
rect 17316 6196 17368 6248
rect 17500 6196 17552 6248
rect 14004 6060 14056 6112
rect 7648 5958 7700 6010
rect 7712 5958 7764 6010
rect 7776 5958 7828 6010
rect 7840 5958 7892 6010
rect 14315 5958 14367 6010
rect 14379 5958 14431 6010
rect 14443 5958 14495 6010
rect 14507 5958 14559 6010
rect 11704 5899 11756 5908
rect 11704 5865 11713 5899
rect 11713 5865 11747 5899
rect 11747 5865 11756 5899
rect 11704 5856 11756 5865
rect 12164 5899 12216 5908
rect 12164 5865 12173 5899
rect 12173 5865 12207 5899
rect 12207 5865 12216 5899
rect 12164 5856 12216 5865
rect 13268 5856 13320 5908
rect 13820 5899 13872 5908
rect 13820 5865 13829 5899
rect 13829 5865 13863 5899
rect 13863 5865 13872 5899
rect 13820 5856 13872 5865
rect 14004 5856 14056 5908
rect 14648 5856 14700 5908
rect 16028 5899 16080 5908
rect 16028 5865 16037 5899
rect 16037 5865 16071 5899
rect 16071 5865 16080 5899
rect 16028 5856 16080 5865
rect 16856 5856 16908 5908
rect 17316 5856 17368 5908
rect 8944 5831 8996 5840
rect 8944 5797 8953 5831
rect 8953 5797 8987 5831
rect 8987 5797 8996 5831
rect 8944 5788 8996 5797
rect 13176 5831 13228 5840
rect 13176 5797 13185 5831
rect 13185 5797 13219 5831
rect 13219 5797 13228 5831
rect 13176 5788 13228 5797
rect 14924 5788 14976 5840
rect 15292 5831 15344 5840
rect 15292 5797 15301 5831
rect 15301 5797 15335 5831
rect 15335 5797 15344 5831
rect 15292 5788 15344 5797
rect 1676 5720 1728 5772
rect 2228 5720 2280 5772
rect 3792 5763 3844 5772
rect 3792 5729 3801 5763
rect 3801 5729 3835 5763
rect 3835 5729 3844 5763
rect 3792 5720 3844 5729
rect 7380 5720 7432 5772
rect 9680 5720 9732 5772
rect 9864 5720 9916 5772
rect 12532 5763 12584 5772
rect 12532 5729 12541 5763
rect 12541 5729 12575 5763
rect 12575 5729 12584 5763
rect 12532 5720 12584 5729
rect 14648 5763 14700 5772
rect 14648 5729 14657 5763
rect 14657 5729 14691 5763
rect 14691 5729 14700 5763
rect 14648 5720 14700 5729
rect 16580 5763 16632 5772
rect 16580 5729 16589 5763
rect 16589 5729 16623 5763
rect 16623 5729 16632 5763
rect 16580 5720 16632 5729
rect 16948 5763 17000 5772
rect 16948 5729 16957 5763
rect 16957 5729 16991 5763
rect 16991 5729 17000 5763
rect 16948 5720 17000 5729
rect 17132 5720 17184 5772
rect 7748 5652 7800 5704
rect 11428 5695 11480 5704
rect 11428 5661 11437 5695
rect 11437 5661 11471 5695
rect 11471 5661 11480 5695
rect 11428 5652 11480 5661
rect 16396 5627 16448 5636
rect 16396 5593 16405 5627
rect 16405 5593 16439 5627
rect 16439 5593 16448 5627
rect 16396 5584 16448 5593
rect 4315 5414 4367 5466
rect 4379 5414 4431 5466
rect 4443 5414 4495 5466
rect 4507 5414 4559 5466
rect 10982 5414 11034 5466
rect 11046 5414 11098 5466
rect 11110 5414 11162 5466
rect 11174 5414 11226 5466
rect 17648 5414 17700 5466
rect 17712 5414 17764 5466
rect 17776 5414 17828 5466
rect 17840 5414 17892 5466
rect 1676 5312 1728 5364
rect 7748 5355 7800 5364
rect 7748 5321 7757 5355
rect 7757 5321 7791 5355
rect 7791 5321 7800 5355
rect 7748 5312 7800 5321
rect 9680 5312 9732 5364
rect 10232 5355 10284 5364
rect 10232 5321 10241 5355
rect 10241 5321 10275 5355
rect 10275 5321 10284 5355
rect 10232 5312 10284 5321
rect 12532 5355 12584 5364
rect 12532 5321 12541 5355
rect 12541 5321 12575 5355
rect 12575 5321 12584 5355
rect 12532 5312 12584 5321
rect 13268 5312 13320 5364
rect 16580 5312 16632 5364
rect 12440 5244 12492 5296
rect 15568 5287 15620 5296
rect 14004 5219 14056 5228
rect 14004 5185 14013 5219
rect 14013 5185 14047 5219
rect 14047 5185 14056 5219
rect 14004 5176 14056 5185
rect 2136 5151 2188 5160
rect 2136 5117 2145 5151
rect 2145 5117 2179 5151
rect 2179 5117 2188 5151
rect 2136 5108 2188 5117
rect 13912 5151 13964 5160
rect 13912 5117 13921 5151
rect 13921 5117 13955 5151
rect 13955 5117 13964 5151
rect 13912 5108 13964 5117
rect 15568 5253 15577 5287
rect 15577 5253 15611 5287
rect 15611 5253 15620 5287
rect 15568 5244 15620 5253
rect 17132 5244 17184 5296
rect 14188 5151 14240 5160
rect 14188 5117 14197 5151
rect 14197 5117 14231 5151
rect 14231 5117 14240 5151
rect 14188 5108 14240 5117
rect 15476 5108 15528 5160
rect 7288 5015 7340 5024
rect 7288 4981 7297 5015
rect 7297 4981 7331 5015
rect 7331 4981 7340 5015
rect 7288 4972 7340 4981
rect 9864 5015 9916 5024
rect 9864 4981 9873 5015
rect 9873 4981 9907 5015
rect 9907 4981 9916 5015
rect 9864 4972 9916 4981
rect 14648 5015 14700 5024
rect 14648 4981 14657 5015
rect 14657 4981 14691 5015
rect 14691 4981 14700 5015
rect 14648 4972 14700 4981
rect 7648 4870 7700 4922
rect 7712 4870 7764 4922
rect 7776 4870 7828 4922
rect 7840 4870 7892 4922
rect 14315 4870 14367 4922
rect 14379 4870 14431 4922
rect 14443 4870 14495 4922
rect 14507 4870 14559 4922
rect 1400 4768 1452 4820
rect 1676 4811 1728 4820
rect 1676 4777 1685 4811
rect 1685 4777 1719 4811
rect 1719 4777 1728 4811
rect 1676 4768 1728 4777
rect 13912 4768 13964 4820
rect 14096 4811 14148 4820
rect 14096 4777 14105 4811
rect 14105 4777 14139 4811
rect 14139 4777 14148 4811
rect 14096 4768 14148 4777
rect 16948 4768 17000 4820
rect 14556 4700 14608 4752
rect 15016 4700 15068 4752
rect 15476 4700 15528 4752
rect 15752 4743 15804 4752
rect 15752 4709 15761 4743
rect 15761 4709 15795 4743
rect 15795 4709 15804 4743
rect 15752 4700 15804 4709
rect 14188 4564 14240 4616
rect 15200 4632 15252 4684
rect 15936 4675 15988 4684
rect 15936 4641 15945 4675
rect 15945 4641 15979 4675
rect 15979 4641 15988 4675
rect 15936 4632 15988 4641
rect 14832 4496 14884 4548
rect 4315 4326 4367 4378
rect 4379 4326 4431 4378
rect 4443 4326 4495 4378
rect 4507 4326 4559 4378
rect 10982 4326 11034 4378
rect 11046 4326 11098 4378
rect 11110 4326 11162 4378
rect 11174 4326 11226 4378
rect 17648 4326 17700 4378
rect 17712 4326 17764 4378
rect 17776 4326 17828 4378
rect 17840 4326 17892 4378
rect 14188 4267 14240 4276
rect 14188 4233 14197 4267
rect 14197 4233 14231 4267
rect 14231 4233 14240 4267
rect 14188 4224 14240 4233
rect 14556 4267 14608 4276
rect 14556 4233 14565 4267
rect 14565 4233 14599 4267
rect 14599 4233 14608 4267
rect 14556 4224 14608 4233
rect 15936 4224 15988 4276
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 1676 4131 1728 4140
rect 1676 4097 1685 4131
rect 1685 4097 1719 4131
rect 1719 4097 1728 4131
rect 1676 4088 1728 4097
rect 3056 4131 3108 4140
rect 3056 4097 3065 4131
rect 3065 4097 3099 4131
rect 3099 4097 3108 4131
rect 3056 4088 3108 4097
rect 10232 4131 10284 4140
rect 10232 4097 10241 4131
rect 10241 4097 10275 4131
rect 10275 4097 10284 4131
rect 10232 4088 10284 4097
rect 12348 4088 12400 4140
rect 10048 3927 10100 3936
rect 10048 3893 10057 3927
rect 10057 3893 10091 3927
rect 10091 3893 10100 3927
rect 10048 3884 10100 3893
rect 7648 3782 7700 3834
rect 7712 3782 7764 3834
rect 7776 3782 7828 3834
rect 7840 3782 7892 3834
rect 14315 3782 14367 3834
rect 14379 3782 14431 3834
rect 14443 3782 14495 3834
rect 14507 3782 14559 3834
rect 1676 3723 1728 3732
rect 1676 3689 1685 3723
rect 1685 3689 1719 3723
rect 1719 3689 1728 3723
rect 1676 3680 1728 3689
rect 10232 3723 10284 3732
rect 10232 3689 10241 3723
rect 10241 3689 10275 3723
rect 10275 3689 10284 3723
rect 10232 3680 10284 3689
rect 4315 3238 4367 3290
rect 4379 3238 4431 3290
rect 4443 3238 4495 3290
rect 4507 3238 4559 3290
rect 10982 3238 11034 3290
rect 11046 3238 11098 3290
rect 11110 3238 11162 3290
rect 11174 3238 11226 3290
rect 17648 3238 17700 3290
rect 17712 3238 17764 3290
rect 17776 3238 17828 3290
rect 17840 3238 17892 3290
rect 7648 2694 7700 2746
rect 7712 2694 7764 2746
rect 7776 2694 7828 2746
rect 7840 2694 7892 2746
rect 14315 2694 14367 2746
rect 14379 2694 14431 2746
rect 14443 2694 14495 2746
rect 14507 2694 14559 2746
rect 9772 2592 9824 2644
rect 10140 2592 10192 2644
rect 9496 2456 9548 2508
rect 9772 2431 9824 2440
rect 9772 2397 9781 2431
rect 9781 2397 9815 2431
rect 9815 2397 9824 2431
rect 9772 2388 9824 2397
rect 9496 2295 9548 2304
rect 9496 2261 9505 2295
rect 9505 2261 9539 2295
rect 9539 2261 9548 2295
rect 9496 2252 9548 2261
rect 11336 2295 11388 2304
rect 11336 2261 11345 2295
rect 11345 2261 11379 2295
rect 11379 2261 11388 2295
rect 11336 2252 11388 2261
rect 12256 2252 12308 2304
rect 4315 2150 4367 2202
rect 4379 2150 4431 2202
rect 4443 2150 4495 2202
rect 4507 2150 4559 2202
rect 10982 2150 11034 2202
rect 11046 2150 11098 2202
rect 11110 2150 11162 2202
rect 11174 2150 11226 2202
rect 17648 2150 17700 2202
rect 17712 2150 17764 2202
rect 17776 2150 17828 2202
rect 17840 2150 17892 2202
<< metal2 >>
rect 3606 79520 3662 79529
rect 3606 79455 3662 79464
rect 2870 77888 2926 77897
rect 2870 77823 2926 77832
rect 2134 77072 2190 77081
rect 2134 77007 2190 77016
rect 2148 74866 2176 77007
rect 2136 74860 2188 74866
rect 2136 74802 2188 74808
rect 2228 74792 2280 74798
rect 2228 74734 2280 74740
rect 2136 74248 2188 74254
rect 2136 74190 2188 74196
rect 2148 73914 2176 74190
rect 2240 74118 2268 74734
rect 2780 74316 2832 74322
rect 2780 74258 2832 74264
rect 2688 74248 2740 74254
rect 2688 74190 2740 74196
rect 2228 74112 2280 74118
rect 2228 74054 2280 74060
rect 2240 73914 2268 74054
rect 2136 73908 2188 73914
rect 2136 73850 2188 73856
rect 2228 73908 2280 73914
rect 2228 73850 2280 73856
rect 2700 73250 2728 74190
rect 2792 73710 2820 74258
rect 2780 73704 2832 73710
rect 2780 73646 2832 73652
rect 2792 73370 2820 73646
rect 2780 73364 2832 73370
rect 2780 73306 2832 73312
rect 2884 73302 2912 77823
rect 3240 77512 3292 77518
rect 3240 77454 3292 77460
rect 2964 75200 3016 75206
rect 2964 75142 3016 75148
rect 2976 74798 3004 75142
rect 2964 74792 3016 74798
rect 2964 74734 3016 74740
rect 2872 73296 2924 73302
rect 2700 73222 2820 73250
rect 2872 73238 2924 73244
rect 2688 73160 2740 73166
rect 2688 73102 2740 73108
rect 2700 72826 2728 73102
rect 2688 72820 2740 72826
rect 2688 72762 2740 72768
rect 2792 72146 2820 73222
rect 3056 73092 3108 73098
rect 3056 73034 3108 73040
rect 3068 72826 3096 73034
rect 3056 72820 3108 72826
rect 3056 72762 3108 72768
rect 3252 72604 3280 77454
rect 3332 77444 3384 77450
rect 3332 77386 3384 77392
rect 3160 72576 3280 72604
rect 2870 72312 2926 72321
rect 2870 72247 2926 72256
rect 2780 72140 2832 72146
rect 2780 72082 2832 72088
rect 2792 70650 2820 72082
rect 1492 70644 1544 70650
rect 1492 70586 1544 70592
rect 2780 70644 2832 70650
rect 2780 70586 2832 70592
rect 1504 69970 1532 70586
rect 1768 70304 1820 70310
rect 1768 70246 1820 70252
rect 1492 69964 1544 69970
rect 1492 69906 1544 69912
rect 1504 68338 1532 69906
rect 1780 69902 1808 70246
rect 1768 69896 1820 69902
rect 1768 69838 1820 69844
rect 1780 69290 1808 69838
rect 2504 69760 2556 69766
rect 2504 69702 2556 69708
rect 2516 69426 2544 69702
rect 2884 69465 2912 72247
rect 2870 69456 2926 69465
rect 2504 69420 2556 69426
rect 2870 69391 2926 69400
rect 2504 69362 2556 69368
rect 1768 69284 1820 69290
rect 1768 69226 1820 69232
rect 2228 69216 2280 69222
rect 2228 69158 2280 69164
rect 2042 69048 2098 69057
rect 2042 68983 2098 68992
rect 1676 68808 1728 68814
rect 1676 68750 1728 68756
rect 1492 68332 1544 68338
rect 1492 68274 1544 68280
rect 1504 67862 1532 68274
rect 1492 67856 1544 67862
rect 1492 67798 1544 67804
rect 1306 67416 1362 67425
rect 1306 67351 1362 67360
rect 1216 61260 1268 61266
rect 1216 61202 1268 61208
rect 1228 58546 1256 61202
rect 1216 58540 1268 58546
rect 1216 58482 1268 58488
rect 1320 58138 1348 67351
rect 1688 66745 1716 68750
rect 1768 68672 1820 68678
rect 1768 68614 1820 68620
rect 1780 68338 1808 68614
rect 1768 68332 1820 68338
rect 1768 68274 1820 68280
rect 1768 67720 1820 67726
rect 1768 67662 1820 67668
rect 1674 66736 1730 66745
rect 1674 66671 1730 66680
rect 1780 65113 1808 67662
rect 1860 67176 1912 67182
rect 1860 67118 1912 67124
rect 1872 66502 1900 67118
rect 1860 66496 1912 66502
rect 1860 66438 1912 66444
rect 1872 65958 1900 66438
rect 1860 65952 1912 65958
rect 1860 65894 1912 65900
rect 1766 65104 1822 65113
rect 1766 65039 1822 65048
rect 1768 65000 1820 65006
rect 1768 64942 1820 64948
rect 1780 64326 1808 64942
rect 1768 64320 1820 64326
rect 1768 64262 1820 64268
rect 1676 63776 1728 63782
rect 1676 63718 1728 63724
rect 1688 63238 1716 63718
rect 1780 63374 1808 64262
rect 1768 63368 1820 63374
rect 1768 63310 1820 63316
rect 1676 63232 1728 63238
rect 1676 63174 1728 63180
rect 1492 62756 1544 62762
rect 1492 62698 1544 62704
rect 1504 62665 1532 62698
rect 1490 62656 1546 62665
rect 1490 62591 1546 62600
rect 1676 62348 1728 62354
rect 1676 62290 1728 62296
rect 1688 62234 1716 62290
rect 1688 62206 1808 62234
rect 1676 61736 1728 61742
rect 1676 61678 1728 61684
rect 1492 61668 1544 61674
rect 1492 61610 1544 61616
rect 1504 61033 1532 61610
rect 1490 61024 1546 61033
rect 1490 60959 1546 60968
rect 1688 60518 1716 61678
rect 1780 61198 1808 62206
rect 1768 61192 1820 61198
rect 1768 61134 1820 61140
rect 1676 60512 1728 60518
rect 1676 60454 1728 60460
rect 1582 60344 1638 60353
rect 1582 60279 1638 60288
rect 1492 59696 1544 59702
rect 1492 59638 1544 59644
rect 1398 59528 1454 59537
rect 1398 59463 1454 59472
rect 1308 58132 1360 58138
rect 1308 58074 1360 58080
rect 1412 58070 1440 59463
rect 1504 59090 1532 59638
rect 1596 59158 1624 60279
rect 1584 59152 1636 59158
rect 1584 59094 1636 59100
rect 1492 59084 1544 59090
rect 1492 59026 1544 59032
rect 1688 59022 1716 60454
rect 1780 59974 1808 61134
rect 1768 59968 1820 59974
rect 1768 59910 1820 59916
rect 1768 59152 1820 59158
rect 1768 59094 1820 59100
rect 1676 59016 1728 59022
rect 1676 58958 1728 58964
rect 1780 58546 1808 59094
rect 1768 58540 1820 58546
rect 1768 58482 1820 58488
rect 1768 58336 1820 58342
rect 1768 58278 1820 58284
rect 1400 58064 1452 58070
rect 1400 58006 1452 58012
rect 1492 57928 1544 57934
rect 1492 57870 1544 57876
rect 1400 57860 1452 57866
rect 1400 57802 1452 57808
rect 1306 47424 1362 47433
rect 1306 47359 1362 47368
rect 1320 44946 1348 47359
rect 1308 44940 1360 44946
rect 1308 44882 1360 44888
rect 1412 33561 1440 57802
rect 1504 56506 1532 57870
rect 1582 57080 1638 57089
rect 1582 57015 1638 57024
rect 1492 56500 1544 56506
rect 1492 56442 1544 56448
rect 1492 54596 1544 54602
rect 1492 54538 1544 54544
rect 1504 54126 1532 54538
rect 1596 54194 1624 57015
rect 1676 56908 1728 56914
rect 1676 56850 1728 56856
rect 1688 55962 1716 56850
rect 1780 56846 1808 58278
rect 1768 56840 1820 56846
rect 1768 56782 1820 56788
rect 1676 55956 1728 55962
rect 1676 55898 1728 55904
rect 1780 55894 1808 56782
rect 1768 55888 1820 55894
rect 1768 55830 1820 55836
rect 1780 55418 1808 55830
rect 1768 55412 1820 55418
rect 1768 55354 1820 55360
rect 1768 54528 1820 54534
rect 1768 54470 1820 54476
rect 1584 54188 1636 54194
rect 1584 54130 1636 54136
rect 1676 54188 1728 54194
rect 1676 54130 1728 54136
rect 1492 54120 1544 54126
rect 1492 54062 1544 54068
rect 1688 53786 1716 54130
rect 1780 54126 1808 54470
rect 1768 54120 1820 54126
rect 1768 54062 1820 54068
rect 1676 53780 1728 53786
rect 1676 53722 1728 53728
rect 1780 53666 1808 54062
rect 1872 53825 1900 65894
rect 1950 61840 2006 61849
rect 1950 61775 2006 61784
rect 1964 60722 1992 61775
rect 1952 60716 2004 60722
rect 1952 60658 2004 60664
rect 1952 59968 2004 59974
rect 1952 59910 2004 59916
rect 1964 57866 1992 59910
rect 1952 57860 2004 57866
rect 1952 57802 2004 57808
rect 2056 57458 2084 68983
rect 2240 68882 2268 69158
rect 2516 68882 2544 69362
rect 2596 69352 2648 69358
rect 2596 69294 2648 69300
rect 2962 69320 3018 69329
rect 2608 69222 2636 69294
rect 2962 69255 3018 69264
rect 2596 69216 2648 69222
rect 2596 69158 2648 69164
rect 2228 68876 2280 68882
rect 2228 68818 2280 68824
rect 2504 68876 2556 68882
rect 2504 68818 2556 68824
rect 2136 68672 2188 68678
rect 2136 68614 2188 68620
rect 2148 66774 2176 68614
rect 2240 67930 2268 68818
rect 2228 67924 2280 67930
rect 2228 67866 2280 67872
rect 2504 67856 2556 67862
rect 2504 67798 2556 67804
rect 2320 67720 2372 67726
rect 2320 67662 2372 67668
rect 2332 66842 2360 67662
rect 2320 66836 2372 66842
rect 2320 66778 2372 66784
rect 2136 66768 2188 66774
rect 2136 66710 2188 66716
rect 2148 65754 2176 66710
rect 2136 65748 2188 65754
rect 2136 65690 2188 65696
rect 2320 65748 2372 65754
rect 2320 65690 2372 65696
rect 2228 65408 2280 65414
rect 2228 65350 2280 65356
rect 2240 65006 2268 65350
rect 2228 65000 2280 65006
rect 2228 64942 2280 64948
rect 2136 63844 2188 63850
rect 2136 63786 2188 63792
rect 2148 63481 2176 63786
rect 2134 63472 2190 63481
rect 2134 63407 2190 63416
rect 2136 63368 2188 63374
rect 2136 63310 2188 63316
rect 2148 62676 2176 63310
rect 2228 63232 2280 63238
rect 2228 63174 2280 63180
rect 2240 62830 2268 63174
rect 2228 62824 2280 62830
rect 2228 62766 2280 62772
rect 2148 62648 2268 62676
rect 2136 62280 2188 62286
rect 2136 62222 2188 62228
rect 2148 61810 2176 62222
rect 2136 61804 2188 61810
rect 2136 61746 2188 61752
rect 2240 61690 2268 62648
rect 2148 61662 2268 61690
rect 2044 57452 2096 57458
rect 2044 57394 2096 57400
rect 1858 53816 1914 53825
rect 1858 53751 1914 53760
rect 1688 53638 1808 53666
rect 1688 53106 1716 53638
rect 1676 53100 1728 53106
rect 1676 53042 1728 53048
rect 1688 52630 1716 53042
rect 1676 52624 1728 52630
rect 1674 52592 1676 52601
rect 1728 52592 1730 52601
rect 1674 52527 1730 52536
rect 1858 52320 1914 52329
rect 1858 52255 1914 52264
rect 1584 51604 1636 51610
rect 1584 51546 1636 51552
rect 1490 51504 1546 51513
rect 1490 51439 1546 51448
rect 1504 46594 1532 51439
rect 1596 50862 1624 51546
rect 1584 50856 1636 50862
rect 1584 50798 1636 50804
rect 1768 50856 1820 50862
rect 1768 50798 1820 50804
rect 1596 49094 1624 50798
rect 1780 50182 1808 50798
rect 1768 50176 1820 50182
rect 1768 50118 1820 50124
rect 1584 49088 1636 49094
rect 1584 49030 1636 49036
rect 1596 48770 1624 49030
rect 1596 48754 1716 48770
rect 1596 48748 1728 48754
rect 1596 48742 1676 48748
rect 1676 48690 1728 48696
rect 1584 48680 1636 48686
rect 1584 48622 1636 48628
rect 1596 48006 1624 48622
rect 1584 48000 1636 48006
rect 1584 47942 1636 47948
rect 1596 47025 1624 47942
rect 1676 47660 1728 47666
rect 1676 47602 1728 47608
rect 1688 47054 1716 47602
rect 1676 47048 1728 47054
rect 1582 47016 1638 47025
rect 1676 46990 1728 46996
rect 1582 46951 1638 46960
rect 1504 46566 1624 46594
rect 1492 46436 1544 46442
rect 1492 46378 1544 46384
rect 1504 45830 1532 46378
rect 1492 45824 1544 45830
rect 1492 45766 1544 45772
rect 1504 44305 1532 45766
rect 1596 45506 1624 46566
rect 1676 46572 1728 46578
rect 1676 46514 1728 46520
rect 1688 46170 1716 46514
rect 1676 46164 1728 46170
rect 1676 46106 1728 46112
rect 1780 45937 1808 50118
rect 1766 45928 1822 45937
rect 1766 45863 1822 45872
rect 1596 45478 1808 45506
rect 1584 45416 1636 45422
rect 1584 45358 1636 45364
rect 1596 44742 1624 45358
rect 1584 44736 1636 44742
rect 1584 44678 1636 44684
rect 1490 44296 1546 44305
rect 1490 44231 1546 44240
rect 1596 43489 1624 44678
rect 1676 44532 1728 44538
rect 1676 44474 1728 44480
rect 1688 43790 1716 44474
rect 1676 43784 1728 43790
rect 1676 43726 1728 43732
rect 1582 43480 1638 43489
rect 1582 43415 1638 43424
rect 1688 43314 1716 43726
rect 1676 43308 1728 43314
rect 1676 43250 1728 43256
rect 1584 43240 1636 43246
rect 1504 43188 1584 43194
rect 1504 43182 1636 43188
rect 1504 43166 1624 43182
rect 1504 42566 1532 43166
rect 1688 42906 1716 43250
rect 1676 42900 1728 42906
rect 1676 42842 1728 42848
rect 1492 42560 1544 42566
rect 1492 42502 1544 42508
rect 1504 41857 1532 42502
rect 1688 42226 1716 42842
rect 1676 42220 1728 42226
rect 1676 42162 1728 42168
rect 1584 42152 1636 42158
rect 1584 42094 1636 42100
rect 1490 41848 1546 41857
rect 1490 41783 1546 41792
rect 1596 41478 1624 42094
rect 1688 41818 1716 42162
rect 1676 41812 1728 41818
rect 1676 41754 1728 41760
rect 1584 41472 1636 41478
rect 1582 41440 1584 41449
rect 1636 41440 1638 41449
rect 1582 41375 1638 41384
rect 1780 41274 1808 45478
rect 1768 41268 1820 41274
rect 1768 41210 1820 41216
rect 1676 41132 1728 41138
rect 1676 41074 1728 41080
rect 1584 41064 1636 41070
rect 1584 41006 1636 41012
rect 1596 40390 1624 41006
rect 1688 40390 1716 41074
rect 1584 40384 1636 40390
rect 1582 40352 1584 40361
rect 1676 40384 1728 40390
rect 1636 40352 1638 40361
rect 1676 40326 1728 40332
rect 1582 40287 1638 40296
rect 1584 38412 1636 38418
rect 1584 38354 1636 38360
rect 1596 38298 1624 38354
rect 1688 38350 1716 40326
rect 1504 38270 1624 38298
rect 1676 38344 1728 38350
rect 1676 38286 1728 38292
rect 1504 37330 1532 38270
rect 1688 38010 1716 38286
rect 1676 38004 1728 38010
rect 1676 37946 1728 37952
rect 1872 37890 1900 52255
rect 1950 49056 2006 49065
rect 1950 48991 2006 49000
rect 1964 45014 1992 48991
rect 2044 48680 2096 48686
rect 2148 48657 2176 61662
rect 2228 59016 2280 59022
rect 2228 58958 2280 58964
rect 2240 57934 2268 58958
rect 2332 58177 2360 65690
rect 2516 65686 2544 67798
rect 2608 66706 2636 69158
rect 2780 68808 2832 68814
rect 2780 68750 2832 68756
rect 2792 68202 2820 68750
rect 2780 68196 2832 68202
rect 2780 68138 2832 68144
rect 2792 67726 2820 68138
rect 2872 68128 2924 68134
rect 2872 68070 2924 68076
rect 2884 67794 2912 68070
rect 2872 67788 2924 67794
rect 2872 67730 2924 67736
rect 2780 67720 2832 67726
rect 2780 67662 2832 67668
rect 2792 67046 2820 67662
rect 2884 67386 2912 67730
rect 2872 67380 2924 67386
rect 2872 67322 2924 67328
rect 2780 67040 2832 67046
rect 2780 66982 2832 66988
rect 2596 66700 2648 66706
rect 2596 66642 2648 66648
rect 2608 66298 2636 66642
rect 2596 66292 2648 66298
rect 2596 66234 2648 66240
rect 2792 65958 2820 66982
rect 2872 66836 2924 66842
rect 2872 66778 2924 66784
rect 2884 66298 2912 66778
rect 2872 66292 2924 66298
rect 2872 66234 2924 66240
rect 2884 66094 2912 66234
rect 2872 66088 2924 66094
rect 2872 66030 2924 66036
rect 2780 65952 2832 65958
rect 2780 65894 2832 65900
rect 2504 65680 2556 65686
rect 2504 65622 2556 65628
rect 2596 65068 2648 65074
rect 2596 65010 2648 65016
rect 2504 64932 2556 64938
rect 2504 64874 2556 64880
rect 2412 64320 2464 64326
rect 2412 64262 2464 64268
rect 2424 63850 2452 64262
rect 2412 63844 2464 63850
rect 2412 63786 2464 63792
rect 2516 63481 2544 64874
rect 2502 63472 2558 63481
rect 2424 63430 2502 63458
rect 2424 62490 2452 63430
rect 2502 63407 2558 63416
rect 2502 63336 2558 63345
rect 2502 63271 2558 63280
rect 2516 62914 2544 63271
rect 2608 63034 2636 65010
rect 2688 64388 2740 64394
rect 2688 64330 2740 64336
rect 2700 63918 2728 64330
rect 2792 64054 2820 65894
rect 2872 65680 2924 65686
rect 2872 65622 2924 65628
rect 2884 64870 2912 65622
rect 2872 64864 2924 64870
rect 2872 64806 2924 64812
rect 2884 64530 2912 64806
rect 2872 64524 2924 64530
rect 2872 64466 2924 64472
rect 2870 64288 2926 64297
rect 2870 64223 2926 64232
rect 2780 64048 2832 64054
rect 2780 63990 2832 63996
rect 2688 63912 2740 63918
rect 2686 63880 2688 63889
rect 2740 63880 2742 63889
rect 2686 63815 2742 63824
rect 2688 63300 2740 63306
rect 2688 63242 2740 63248
rect 2596 63028 2648 63034
rect 2596 62970 2648 62976
rect 2516 62886 2636 62914
rect 2504 62824 2556 62830
rect 2504 62766 2556 62772
rect 2412 62484 2464 62490
rect 2412 62426 2464 62432
rect 2516 61810 2544 62766
rect 2504 61804 2556 61810
rect 2504 61746 2556 61752
rect 2608 60330 2636 62886
rect 2700 62234 2728 63242
rect 2884 62422 2912 64223
rect 2872 62416 2924 62422
rect 2872 62358 2924 62364
rect 2700 62206 2820 62234
rect 2976 62218 3004 69255
rect 3056 69216 3108 69222
rect 3054 69184 3056 69193
rect 3108 69184 3110 69193
rect 3054 69119 3110 69128
rect 3056 64456 3108 64462
rect 3056 64398 3108 64404
rect 3068 63850 3096 64398
rect 3056 63844 3108 63850
rect 3056 63786 3108 63792
rect 2688 61804 2740 61810
rect 2688 61746 2740 61752
rect 2700 61266 2728 61746
rect 2688 61260 2740 61266
rect 2688 61202 2740 61208
rect 2688 60648 2740 60654
rect 2688 60590 2740 60596
rect 2700 60489 2728 60590
rect 2686 60480 2742 60489
rect 2686 60415 2742 60424
rect 2424 60302 2636 60330
rect 2700 60314 2728 60415
rect 2688 60308 2740 60314
rect 2318 58168 2374 58177
rect 2318 58103 2374 58112
rect 2228 57928 2280 57934
rect 2228 57870 2280 57876
rect 2240 57254 2268 57870
rect 2228 57248 2280 57254
rect 2228 57190 2280 57196
rect 2240 55078 2268 57190
rect 2424 55826 2452 60302
rect 2688 60250 2740 60256
rect 2502 60208 2558 60217
rect 2792 60178 2820 62206
rect 2964 62212 3016 62218
rect 2964 62154 3016 62160
rect 3160 61792 3188 72576
rect 3240 72140 3292 72146
rect 3240 72082 3292 72088
rect 3252 71738 3280 72082
rect 3240 71732 3292 71738
rect 3240 71674 3292 71680
rect 3344 71618 3372 77386
rect 3422 75440 3478 75449
rect 3422 75375 3478 75384
rect 2976 61764 3188 61792
rect 3252 71590 3372 71618
rect 2872 60648 2924 60654
rect 2872 60590 2924 60596
rect 2502 60143 2558 60152
rect 2780 60172 2832 60178
rect 2412 55820 2464 55826
rect 2412 55762 2464 55768
rect 2228 55072 2280 55078
rect 2228 55014 2280 55020
rect 2240 54194 2268 55014
rect 2412 54732 2464 54738
rect 2412 54674 2464 54680
rect 2318 54632 2374 54641
rect 2318 54567 2374 54576
rect 2228 54188 2280 54194
rect 2228 54130 2280 54136
rect 2228 53712 2280 53718
rect 2228 53654 2280 53660
rect 2240 50862 2268 53654
rect 2228 50856 2280 50862
rect 2228 50798 2280 50804
rect 2240 49978 2268 50798
rect 2228 49972 2280 49978
rect 2228 49914 2280 49920
rect 2226 49736 2282 49745
rect 2226 49671 2282 49680
rect 2044 48622 2096 48628
rect 2134 48648 2190 48657
rect 2056 47598 2084 48622
rect 2134 48583 2190 48592
rect 2044 47592 2096 47598
rect 2044 47534 2096 47540
rect 2056 46986 2084 47534
rect 2044 46980 2096 46986
rect 2044 46922 2096 46928
rect 2240 45608 2268 49671
rect 2332 49638 2360 54567
rect 2424 53446 2452 54674
rect 2412 53440 2464 53446
rect 2412 53382 2464 53388
rect 2424 53242 2452 53382
rect 2412 53236 2464 53242
rect 2412 53178 2464 53184
rect 2412 53032 2464 53038
rect 2412 52974 2464 52980
rect 2424 52358 2452 52974
rect 2412 52352 2464 52358
rect 2412 52294 2464 52300
rect 2424 50726 2452 52294
rect 2412 50720 2464 50726
rect 2412 50662 2464 50668
rect 2320 49632 2372 49638
rect 2320 49574 2372 49580
rect 2424 49230 2452 50662
rect 2516 50017 2544 60143
rect 2780 60114 2832 60120
rect 2884 60110 2912 60590
rect 2872 60104 2924 60110
rect 2872 60046 2924 60052
rect 2688 59968 2740 59974
rect 2688 59910 2740 59916
rect 2594 59664 2650 59673
rect 2594 59599 2650 59608
rect 2502 50008 2558 50017
rect 2502 49943 2558 49952
rect 2504 49768 2556 49774
rect 2504 49710 2556 49716
rect 2516 49434 2544 49710
rect 2504 49428 2556 49434
rect 2504 49370 2556 49376
rect 2412 49224 2464 49230
rect 2412 49166 2464 49172
rect 2424 48550 2452 49166
rect 2412 48544 2464 48550
rect 2332 48504 2412 48532
rect 2332 46170 2360 48504
rect 2412 48486 2464 48492
rect 2412 47048 2464 47054
rect 2412 46990 2464 46996
rect 2320 46164 2372 46170
rect 2320 46106 2372 46112
rect 2148 45580 2268 45608
rect 2148 45370 2176 45580
rect 2332 45506 2360 46106
rect 2240 45490 2360 45506
rect 2228 45484 2360 45490
rect 2280 45478 2360 45484
rect 2228 45426 2280 45432
rect 2148 45342 2268 45370
rect 2240 45098 2268 45342
rect 2148 45070 2268 45098
rect 2332 45082 2360 45478
rect 2424 45121 2452 46990
rect 2504 46980 2556 46986
rect 2504 46922 2556 46928
rect 2516 46034 2544 46922
rect 2504 46028 2556 46034
rect 2504 45970 2556 45976
rect 2502 45928 2558 45937
rect 2502 45863 2558 45872
rect 2410 45112 2466 45121
rect 2320 45076 2372 45082
rect 1952 45008 2004 45014
rect 1952 44950 2004 44956
rect 1952 43784 2004 43790
rect 1952 43726 2004 43732
rect 1964 42702 1992 43726
rect 1952 42696 2004 42702
rect 1950 42664 1952 42673
rect 2004 42664 2006 42673
rect 1950 42599 2006 42608
rect 2148 39642 2176 45070
rect 2410 45047 2466 45056
rect 2320 45018 2372 45024
rect 2228 45008 2280 45014
rect 2228 44950 2280 44956
rect 2136 39636 2188 39642
rect 2136 39578 2188 39584
rect 2134 39536 2190 39545
rect 2134 39471 2190 39480
rect 1596 37862 1900 37890
rect 1492 37324 1544 37330
rect 1492 37266 1544 37272
rect 1504 35465 1532 37266
rect 1596 35986 1624 37862
rect 1860 37800 1912 37806
rect 1860 37742 1912 37748
rect 1768 37664 1820 37670
rect 1768 37606 1820 37612
rect 1780 37126 1808 37606
rect 1872 37330 1900 37742
rect 1860 37324 1912 37330
rect 1860 37266 1912 37272
rect 1768 37120 1820 37126
rect 1768 37062 1820 37068
rect 1780 36582 1808 37062
rect 1768 36576 1820 36582
rect 1768 36518 1820 36524
rect 1780 36122 1808 36518
rect 1872 36281 1900 37266
rect 1858 36272 1914 36281
rect 1858 36207 1914 36216
rect 1780 36094 1900 36122
rect 1872 36038 1900 36094
rect 1860 36032 1912 36038
rect 1596 35958 1808 35986
rect 1860 35974 1912 35980
rect 2044 36032 2096 36038
rect 2044 35974 2096 35980
rect 1584 35624 1636 35630
rect 1584 35566 1636 35572
rect 1490 35456 1546 35465
rect 1490 35391 1546 35400
rect 1596 34950 1624 35566
rect 1584 34944 1636 34950
rect 1584 34886 1636 34892
rect 1492 34536 1544 34542
rect 1492 34478 1544 34484
rect 1398 33552 1454 33561
rect 1398 33487 1454 33496
rect 1400 32904 1452 32910
rect 1400 32846 1452 32852
rect 1412 32366 1440 32846
rect 1400 32360 1452 32366
rect 1400 32302 1452 32308
rect 1504 31822 1532 34478
rect 1596 33833 1624 34886
rect 1582 33824 1638 33833
rect 1582 33759 1638 33768
rect 1780 33674 1808 35958
rect 1872 35698 1900 35974
rect 1860 35692 1912 35698
rect 1860 35634 1912 35640
rect 1596 33646 1808 33674
rect 1596 32065 1624 33646
rect 1676 33584 1728 33590
rect 1676 33526 1728 33532
rect 1582 32056 1638 32065
rect 1582 31991 1638 32000
rect 1584 31884 1636 31890
rect 1584 31826 1636 31832
rect 1492 31816 1544 31822
rect 1492 31758 1544 31764
rect 1504 31414 1532 31758
rect 1492 31408 1544 31414
rect 1492 31350 1544 31356
rect 1504 29714 1532 31350
rect 1596 31210 1624 31826
rect 1688 31362 1716 33526
rect 1768 33312 1820 33318
rect 1768 33254 1820 33260
rect 1780 32434 1808 33254
rect 1860 32904 1912 32910
rect 1860 32846 1912 32852
rect 1768 32428 1820 32434
rect 1768 32370 1820 32376
rect 1780 31793 1808 32370
rect 1872 32337 1900 32846
rect 1858 32328 1914 32337
rect 1858 32263 1914 32272
rect 1766 31784 1822 31793
rect 1766 31719 1822 31728
rect 1872 31482 1900 32263
rect 1950 31920 2006 31929
rect 1950 31855 2006 31864
rect 1860 31476 1912 31482
rect 1860 31418 1912 31424
rect 1688 31334 1900 31362
rect 1584 31204 1636 31210
rect 1584 31146 1636 31152
rect 1596 30705 1624 31146
rect 1768 30796 1820 30802
rect 1768 30738 1820 30744
rect 1582 30696 1638 30705
rect 1780 30682 1808 30738
rect 1582 30631 1638 30640
rect 1688 30654 1808 30682
rect 1688 30054 1716 30654
rect 1676 30048 1728 30054
rect 1676 29990 1728 29996
rect 1688 29889 1716 29990
rect 1674 29880 1730 29889
rect 1674 29815 1730 29824
rect 1492 29708 1544 29714
rect 1492 29650 1544 29656
rect 1504 29170 1532 29650
rect 1492 29164 1544 29170
rect 1492 29106 1544 29112
rect 1676 28688 1728 28694
rect 1676 28630 1728 28636
rect 1584 28620 1636 28626
rect 1584 28562 1636 28568
rect 1596 28257 1624 28562
rect 1582 28248 1638 28257
rect 1582 28183 1584 28192
rect 1636 28183 1638 28192
rect 1584 28154 1636 28160
rect 1596 28123 1624 28154
rect 1688 28121 1716 28630
rect 1674 28112 1730 28121
rect 1596 28056 1674 28064
rect 1596 28036 1676 28056
rect 1596 26761 1624 28036
rect 1728 28047 1730 28056
rect 1676 28018 1728 28024
rect 1676 27464 1728 27470
rect 1676 27406 1728 27412
rect 1582 26752 1638 26761
rect 1582 26687 1638 26696
rect 1688 26602 1716 27406
rect 1596 26574 1716 26602
rect 1596 26450 1624 26574
rect 1584 26444 1636 26450
rect 1584 26386 1636 26392
rect 1676 26444 1728 26450
rect 1676 26386 1728 26392
rect 1688 26042 1716 26386
rect 1676 26036 1728 26042
rect 1676 25978 1728 25984
rect 1400 25152 1452 25158
rect 1400 25094 1452 25100
rect 1412 24750 1440 25094
rect 1766 24848 1822 24857
rect 1872 24818 1900 31334
rect 1964 28642 1992 31855
rect 2056 29850 2084 35974
rect 2148 31278 2176 39471
rect 2136 31272 2188 31278
rect 2136 31214 2188 31220
rect 2136 30728 2188 30734
rect 2136 30670 2188 30676
rect 2148 30054 2176 30670
rect 2136 30048 2188 30054
rect 2134 30016 2136 30025
rect 2188 30016 2190 30025
rect 2134 29951 2190 29960
rect 2044 29844 2096 29850
rect 2044 29786 2096 29792
rect 2056 29102 2084 29786
rect 2136 29708 2188 29714
rect 2136 29650 2188 29656
rect 2044 29096 2096 29102
rect 2148 29073 2176 29650
rect 2044 29038 2096 29044
rect 2134 29064 2190 29073
rect 2134 28999 2190 29008
rect 2148 28762 2176 28999
rect 2136 28756 2188 28762
rect 2136 28698 2188 28704
rect 1964 28614 2084 28642
rect 1952 28552 2004 28558
rect 1950 28520 1952 28529
rect 2004 28520 2006 28529
rect 1950 28455 2006 28464
rect 2056 27538 2084 28614
rect 2044 27532 2096 27538
rect 2044 27474 2096 27480
rect 2056 27130 2084 27474
rect 2044 27124 2096 27130
rect 2044 27066 2096 27072
rect 2044 26376 2096 26382
rect 2044 26318 2096 26324
rect 2056 26042 2084 26318
rect 2044 26036 2096 26042
rect 2044 25978 2096 25984
rect 1766 24783 1822 24792
rect 1860 24812 1912 24818
rect 1400 24744 1452 24750
rect 1400 24686 1452 24692
rect 1412 21146 1440 24686
rect 1780 23730 1808 24783
rect 1860 24754 1912 24760
rect 1872 24410 1900 24754
rect 1860 24404 1912 24410
rect 1860 24346 1912 24352
rect 2134 24304 2190 24313
rect 2134 24239 2190 24248
rect 1860 24200 1912 24206
rect 1860 24142 1912 24148
rect 1768 23724 1820 23730
rect 1768 23666 1820 23672
rect 1780 23322 1808 23666
rect 1872 23662 1900 24142
rect 1860 23656 1912 23662
rect 1860 23598 1912 23604
rect 1768 23316 1820 23322
rect 1768 23258 1820 23264
rect 1872 23050 1900 23598
rect 1860 23044 1912 23050
rect 1860 22986 1912 22992
rect 1674 22672 1730 22681
rect 1674 22607 1730 22616
rect 1490 21856 1546 21865
rect 1490 21791 1546 21800
rect 1400 21140 1452 21146
rect 1400 21082 1452 21088
rect 1412 21010 1440 21082
rect 1400 21004 1452 21010
rect 1400 20946 1452 20952
rect 1412 20534 1440 20946
rect 1400 20528 1452 20534
rect 1400 20470 1452 20476
rect 1412 20058 1440 20470
rect 1400 20052 1452 20058
rect 1400 19994 1452 20000
rect 1412 19378 1440 19994
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1412 18850 1440 19314
rect 1504 19310 1532 21791
rect 1688 21010 1716 22607
rect 1872 22098 1900 22986
rect 2148 22098 2176 24239
rect 1860 22092 1912 22098
rect 1860 22034 1912 22040
rect 2136 22092 2188 22098
rect 2136 22034 2188 22040
rect 1872 21622 1900 22034
rect 2148 21690 2176 22034
rect 2136 21684 2188 21690
rect 2136 21626 2188 21632
rect 1860 21616 1912 21622
rect 1860 21558 1912 21564
rect 1676 21004 1728 21010
rect 1676 20946 1728 20952
rect 1688 20602 1716 20946
rect 1676 20596 1728 20602
rect 1676 20538 1728 20544
rect 1766 19544 1822 19553
rect 1766 19479 1822 19488
rect 1492 19304 1544 19310
rect 1492 19246 1544 19252
rect 1504 18970 1532 19246
rect 1492 18964 1544 18970
rect 1492 18906 1544 18912
rect 1412 18822 1624 18850
rect 1398 18728 1454 18737
rect 1398 18663 1454 18672
rect 1412 16114 1440 18663
rect 1596 17746 1624 18822
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1584 17740 1636 17746
rect 1584 17682 1636 17688
rect 1596 16726 1624 17682
rect 1688 17338 1716 18022
rect 1780 17746 1808 19479
rect 1768 17740 1820 17746
rect 1768 17682 1820 17688
rect 1676 17332 1728 17338
rect 1676 17274 1728 17280
rect 1674 17232 1730 17241
rect 1674 17167 1676 17176
rect 1728 17167 1730 17176
rect 1676 17138 1728 17144
rect 1688 16794 1716 17138
rect 1780 16794 1808 17682
rect 1860 17332 1912 17338
rect 1860 17274 1912 17280
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 1584 16720 1636 16726
rect 1584 16662 1636 16668
rect 1872 16590 1900 17274
rect 1860 16584 1912 16590
rect 1860 16526 1912 16532
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1412 15706 1440 16050
rect 1492 16040 1544 16046
rect 1492 15982 1544 15988
rect 1400 15700 1452 15706
rect 1400 15642 1452 15648
rect 1214 15464 1270 15473
rect 1214 15399 1270 15408
rect 1228 10130 1256 15399
rect 1504 15366 1532 15982
rect 1492 15360 1544 15366
rect 1492 15302 1544 15308
rect 1492 13524 1544 13530
rect 1492 13466 1544 13472
rect 1504 11694 1532 13466
rect 1582 13152 1638 13161
rect 1582 13087 1638 13096
rect 1596 12986 1624 13087
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1596 11762 1624 12922
rect 1688 12306 1716 12922
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 1860 12232 1912 12238
rect 1964 12186 1992 12582
rect 1912 12180 1992 12186
rect 1860 12174 1992 12180
rect 1872 12158 1992 12174
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 1492 11688 1544 11694
rect 1492 11630 1544 11636
rect 1504 10606 1532 11630
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1216 10124 1268 10130
rect 1216 10066 1268 10072
rect 1504 10062 1532 10542
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1504 9178 1532 9998
rect 1780 9654 1808 11154
rect 1964 11150 1992 12158
rect 2240 11218 2268 44950
rect 2332 44538 2360 45018
rect 2412 44940 2464 44946
rect 2412 44882 2464 44888
rect 2320 44532 2372 44538
rect 2320 44474 2372 44480
rect 2320 39636 2372 39642
rect 2320 39578 2372 39584
rect 2332 36038 2360 39578
rect 2320 36032 2372 36038
rect 2320 35974 2372 35980
rect 2320 35216 2372 35222
rect 2320 35158 2372 35164
rect 2332 34678 2360 35158
rect 2320 34672 2372 34678
rect 2318 34640 2320 34649
rect 2372 34640 2374 34649
rect 2318 34575 2374 34584
rect 2320 31272 2372 31278
rect 2320 31214 2372 31220
rect 2332 26450 2360 31214
rect 2320 26444 2372 26450
rect 2320 26386 2372 26392
rect 2320 16720 2372 16726
rect 2320 16662 2372 16668
rect 2332 14482 2360 16662
rect 2320 14476 2372 14482
rect 2320 14418 2372 14424
rect 2332 14006 2360 14418
rect 2320 14000 2372 14006
rect 2320 13942 2372 13948
rect 2332 13530 2360 13942
rect 2320 13524 2372 13530
rect 2320 13466 2372 13472
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 1768 9648 1820 9654
rect 1768 9590 1820 9596
rect 1964 9178 1992 11086
rect 2424 10674 2452 44882
rect 2516 44033 2544 45863
rect 2502 44024 2558 44033
rect 2502 43959 2558 43968
rect 2504 41268 2556 41274
rect 2504 41210 2556 41216
rect 2516 35816 2544 41210
rect 2608 38457 2636 59599
rect 2700 59566 2728 59910
rect 2688 59560 2740 59566
rect 2740 59508 2820 59514
rect 2688 59502 2820 59508
rect 2700 59486 2820 59502
rect 2792 58682 2820 59486
rect 2872 59424 2924 59430
rect 2872 59366 2924 59372
rect 2884 59226 2912 59366
rect 2872 59220 2924 59226
rect 2872 59162 2924 59168
rect 2780 58676 2832 58682
rect 2780 58618 2832 58624
rect 2688 56704 2740 56710
rect 2688 56646 2740 56652
rect 2700 56370 2728 56646
rect 2688 56364 2740 56370
rect 2688 56306 2740 56312
rect 2700 55962 2728 56306
rect 2884 56302 2912 59162
rect 2872 56296 2924 56302
rect 2872 56238 2924 56244
rect 2688 55956 2740 55962
rect 2688 55898 2740 55904
rect 2688 55820 2740 55826
rect 2688 55762 2740 55768
rect 2700 40633 2728 55762
rect 2884 54738 2912 56238
rect 2872 54732 2924 54738
rect 2872 54674 2924 54680
rect 2884 54330 2912 54674
rect 2872 54324 2924 54330
rect 2872 54266 2924 54272
rect 2884 53718 2912 54266
rect 2872 53712 2924 53718
rect 2872 53654 2924 53660
rect 2780 53440 2832 53446
rect 2780 53382 2832 53388
rect 2792 51814 2820 53382
rect 2870 53136 2926 53145
rect 2870 53071 2926 53080
rect 2780 51808 2832 51814
rect 2778 51776 2780 51785
rect 2832 51776 2834 51785
rect 2778 51711 2834 51720
rect 2884 49745 2912 53071
rect 2870 49736 2926 49745
rect 2870 49671 2926 49680
rect 2872 49632 2924 49638
rect 2872 49574 2924 49580
rect 2778 48240 2834 48249
rect 2778 48175 2834 48184
rect 2686 40624 2742 40633
rect 2686 40559 2742 40568
rect 2686 39400 2742 39409
rect 2686 39335 2742 39344
rect 2700 39098 2728 39335
rect 2688 39092 2740 39098
rect 2688 39034 2740 39040
rect 2594 38448 2650 38457
rect 2594 38383 2650 38392
rect 2516 35788 2636 35816
rect 2504 35692 2556 35698
rect 2504 35634 2556 35640
rect 2516 35086 2544 35634
rect 2504 35080 2556 35086
rect 2504 35022 2556 35028
rect 2516 34542 2544 35022
rect 2504 34536 2556 34542
rect 2504 34478 2556 34484
rect 2608 33658 2636 35788
rect 2596 33652 2648 33658
rect 2596 33594 2648 33600
rect 2792 33454 2820 48175
rect 2884 47297 2912 49574
rect 2976 47802 3004 61764
rect 3056 61668 3108 61674
rect 3056 61610 3108 61616
rect 3068 61402 3096 61610
rect 3148 61600 3200 61606
rect 3148 61542 3200 61548
rect 3056 61396 3108 61402
rect 3056 61338 3108 61344
rect 3160 61282 3188 61542
rect 3068 61254 3188 61282
rect 3068 60654 3096 61254
rect 3146 61160 3202 61169
rect 3146 61095 3202 61104
rect 3056 60648 3108 60654
rect 3056 60590 3108 60596
rect 3068 58342 3096 60590
rect 3056 58336 3108 58342
rect 3056 58278 3108 58284
rect 3056 57792 3108 57798
rect 3056 57734 3108 57740
rect 3068 57390 3096 57734
rect 3056 57384 3108 57390
rect 3054 57352 3056 57361
rect 3108 57352 3110 57361
rect 3054 57287 3110 57296
rect 3056 56976 3108 56982
rect 3056 56918 3108 56924
rect 3068 55026 3096 56918
rect 3160 55418 3188 61095
rect 3148 55412 3200 55418
rect 3148 55354 3200 55360
rect 3160 55214 3188 55354
rect 3148 55208 3200 55214
rect 3148 55150 3200 55156
rect 3068 54998 3188 55026
rect 3056 53644 3108 53650
rect 3056 53586 3108 53592
rect 3068 52698 3096 53586
rect 3160 53446 3188 54998
rect 3148 53440 3200 53446
rect 3148 53382 3200 53388
rect 3160 52902 3188 53382
rect 3148 52896 3200 52902
rect 3148 52838 3200 52844
rect 3146 52728 3202 52737
rect 3056 52692 3108 52698
rect 3146 52663 3202 52672
rect 3056 52634 3108 52640
rect 3160 52562 3188 52663
rect 3148 52556 3200 52562
rect 3148 52498 3200 52504
rect 3056 52488 3108 52494
rect 3056 52430 3108 52436
rect 3068 51338 3096 52430
rect 3160 51610 3188 52498
rect 3148 51604 3200 51610
rect 3148 51546 3200 51552
rect 3148 51468 3200 51474
rect 3148 51410 3200 51416
rect 3056 51332 3108 51338
rect 3056 51274 3108 51280
rect 3054 49872 3110 49881
rect 3054 49807 3110 49816
rect 2964 47796 3016 47802
rect 2964 47738 3016 47744
rect 2870 47288 2926 47297
rect 2870 47223 2926 47232
rect 2964 45280 3016 45286
rect 2964 45222 3016 45228
rect 2870 42800 2926 42809
rect 2870 42735 2926 42744
rect 2884 42362 2912 42735
rect 2872 42356 2924 42362
rect 2872 42298 2924 42304
rect 2976 42242 3004 45222
rect 2884 42214 3004 42242
rect 2884 41585 2912 42214
rect 2870 41576 2926 41585
rect 2870 41511 2926 41520
rect 2964 39568 3016 39574
rect 2964 39510 3016 39516
rect 2780 33448 2832 33454
rect 2780 33390 2832 33396
rect 2688 33380 2740 33386
rect 2688 33322 2740 33328
rect 2700 32366 2728 33322
rect 2870 33144 2926 33153
rect 2976 33114 3004 39510
rect 2870 33079 2926 33088
rect 2964 33108 3016 33114
rect 2884 32570 2912 33079
rect 2964 33050 3016 33056
rect 2872 32564 2924 32570
rect 2872 32506 2924 32512
rect 2688 32360 2740 32366
rect 2688 32302 2740 32308
rect 2700 32230 2728 32302
rect 2688 32224 2740 32230
rect 2688 32166 2740 32172
rect 2700 30734 2728 32166
rect 2688 30728 2740 30734
rect 2688 30670 2740 30676
rect 2596 29164 2648 29170
rect 2596 29106 2648 29112
rect 2608 28762 2636 29106
rect 2596 28756 2648 28762
rect 2596 28698 2648 28704
rect 2608 28218 2636 28698
rect 2596 28212 2648 28218
rect 2596 28154 2648 28160
rect 2608 27470 2636 28154
rect 2596 27464 2648 27470
rect 2596 27406 2648 27412
rect 2780 27464 2832 27470
rect 2780 27406 2832 27412
rect 2792 26994 2820 27406
rect 2780 26988 2832 26994
rect 2780 26930 2832 26936
rect 2872 26920 2924 26926
rect 2872 26862 2924 26868
rect 2884 26042 2912 26862
rect 2872 26036 2924 26042
rect 2872 25978 2924 25984
rect 2778 25936 2834 25945
rect 2778 25871 2834 25880
rect 2792 24274 2820 25871
rect 2780 24268 2832 24274
rect 2700 24228 2780 24256
rect 2700 23322 2728 24228
rect 2780 24210 2832 24216
rect 2792 24145 2820 24210
rect 2688 23316 2740 23322
rect 2688 23258 2740 23264
rect 2964 20800 3016 20806
rect 2964 20742 3016 20748
rect 2976 19825 3004 20742
rect 2962 19816 3018 19825
rect 2962 19751 3018 19760
rect 2778 17096 2834 17105
rect 2778 17031 2834 17040
rect 2688 16584 2740 16590
rect 2688 16526 2740 16532
rect 2594 16280 2650 16289
rect 2594 16215 2650 16224
rect 2608 14482 2636 16215
rect 2700 15366 2728 16526
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2596 14476 2648 14482
rect 2596 14418 2648 14424
rect 2608 14074 2636 14418
rect 2596 14068 2648 14074
rect 2596 14010 2648 14016
rect 2792 13002 2820 17031
rect 3068 16658 3096 49807
rect 3160 31958 3188 51410
rect 3252 51066 3280 71590
rect 3332 67788 3384 67794
rect 3332 67730 3384 67736
rect 3344 67046 3372 67730
rect 3332 67040 3384 67046
rect 3332 66982 3384 66988
rect 3344 66706 3372 66982
rect 3332 66700 3384 66706
rect 3332 66642 3384 66648
rect 3344 65958 3372 66642
rect 3436 66230 3464 75375
rect 3516 73160 3568 73166
rect 3516 73102 3568 73108
rect 3528 72486 3556 73102
rect 3516 72480 3568 72486
rect 3516 72422 3568 72428
rect 3620 72298 3648 79455
rect 16026 78840 16082 78849
rect 16026 78775 16082 78784
rect 3790 78704 3846 78713
rect 3790 78639 3792 78648
rect 3844 78639 3846 78648
rect 4804 78668 4856 78674
rect 3792 78610 3844 78616
rect 4804 78610 4856 78616
rect 4289 77276 4585 77296
rect 4345 77274 4369 77276
rect 4425 77274 4449 77276
rect 4505 77274 4529 77276
rect 4367 77222 4369 77274
rect 4431 77222 4443 77274
rect 4505 77222 4507 77274
rect 4345 77220 4369 77222
rect 4425 77220 4449 77222
rect 4505 77220 4529 77222
rect 4289 77200 4585 77220
rect 4066 76256 4122 76265
rect 4122 76214 4200 76242
rect 4066 76191 4122 76200
rect 4172 75478 4200 76214
rect 4289 76188 4585 76208
rect 4345 76186 4369 76188
rect 4425 76186 4449 76188
rect 4505 76186 4529 76188
rect 4367 76134 4369 76186
rect 4431 76134 4443 76186
rect 4505 76134 4507 76186
rect 4345 76132 4369 76134
rect 4425 76132 4449 76134
rect 4505 76132 4529 76134
rect 4289 76112 4585 76132
rect 4160 75472 4212 75478
rect 4160 75414 4212 75420
rect 3976 75268 4028 75274
rect 3976 75210 4028 75216
rect 3988 74798 4016 75210
rect 4160 75200 4212 75206
rect 4160 75142 4212 75148
rect 4172 74798 4200 75142
rect 4289 75100 4585 75120
rect 4345 75098 4369 75100
rect 4425 75098 4449 75100
rect 4505 75098 4529 75100
rect 4367 75046 4369 75098
rect 4431 75046 4443 75098
rect 4505 75046 4507 75098
rect 4345 75044 4369 75046
rect 4425 75044 4449 75046
rect 4505 75044 4529 75046
rect 4289 75024 4585 75044
rect 3976 74792 4028 74798
rect 3976 74734 4028 74740
rect 4160 74792 4212 74798
rect 4160 74734 4212 74740
rect 4816 74746 4844 78610
rect 15934 78160 15990 78169
rect 15934 78095 15990 78104
rect 7622 77820 7918 77840
rect 7678 77818 7702 77820
rect 7758 77818 7782 77820
rect 7838 77818 7862 77820
rect 7700 77766 7702 77818
rect 7764 77766 7776 77818
rect 7838 77766 7840 77818
rect 7678 77764 7702 77766
rect 7758 77764 7782 77766
rect 7838 77764 7862 77766
rect 7622 77744 7918 77764
rect 14289 77820 14585 77840
rect 14345 77818 14369 77820
rect 14425 77818 14449 77820
rect 14505 77818 14529 77820
rect 14367 77766 14369 77818
rect 14431 77766 14443 77818
rect 14505 77766 14507 77818
rect 14345 77764 14369 77766
rect 14425 77764 14449 77766
rect 14505 77764 14529 77766
rect 14289 77744 14585 77764
rect 15948 77518 15976 78095
rect 15936 77512 15988 77518
rect 15936 77454 15988 77460
rect 16040 77450 16068 78775
rect 16028 77444 16080 77450
rect 16028 77386 16080 77392
rect 10956 77276 11252 77296
rect 11012 77274 11036 77276
rect 11092 77274 11116 77276
rect 11172 77274 11196 77276
rect 11034 77222 11036 77274
rect 11098 77222 11110 77274
rect 11172 77222 11174 77274
rect 11012 77220 11036 77222
rect 11092 77220 11116 77222
rect 11172 77220 11196 77222
rect 10956 77200 11252 77220
rect 17622 77276 17918 77296
rect 17678 77274 17702 77276
rect 17758 77274 17782 77276
rect 17838 77274 17862 77276
rect 17700 77222 17702 77274
rect 17764 77222 17776 77274
rect 17838 77222 17840 77274
rect 17678 77220 17702 77222
rect 17758 77220 17782 77222
rect 17838 77220 17862 77222
rect 17622 77200 17918 77220
rect 7622 76732 7918 76752
rect 7678 76730 7702 76732
rect 7758 76730 7782 76732
rect 7838 76730 7862 76732
rect 7700 76678 7702 76730
rect 7764 76678 7776 76730
rect 7838 76678 7840 76730
rect 7678 76676 7702 76678
rect 7758 76676 7782 76678
rect 7838 76676 7862 76678
rect 7622 76656 7918 76676
rect 14289 76732 14585 76752
rect 14345 76730 14369 76732
rect 14425 76730 14449 76732
rect 14505 76730 14529 76732
rect 14367 76678 14369 76730
rect 14431 76678 14443 76730
rect 14505 76678 14507 76730
rect 14345 76676 14369 76678
rect 14425 76676 14449 76678
rect 14505 76676 14529 76678
rect 14289 76656 14585 76676
rect 10956 76188 11252 76208
rect 11012 76186 11036 76188
rect 11092 76186 11116 76188
rect 11172 76186 11196 76188
rect 11034 76134 11036 76186
rect 11098 76134 11110 76186
rect 11172 76134 11174 76186
rect 11012 76132 11036 76134
rect 11092 76132 11116 76134
rect 11172 76132 11196 76134
rect 10956 76112 11252 76132
rect 17622 76188 17918 76208
rect 17678 76186 17702 76188
rect 17758 76186 17782 76188
rect 17838 76186 17862 76188
rect 17700 76134 17702 76186
rect 17764 76134 17776 76186
rect 17838 76134 17840 76186
rect 17678 76132 17702 76134
rect 17758 76132 17782 76134
rect 17838 76132 17862 76134
rect 17622 76112 17918 76132
rect 7622 75644 7918 75664
rect 7678 75642 7702 75644
rect 7758 75642 7782 75644
rect 7838 75642 7862 75644
rect 7700 75590 7702 75642
rect 7764 75590 7776 75642
rect 7838 75590 7840 75642
rect 7678 75588 7702 75590
rect 7758 75588 7782 75590
rect 7838 75588 7862 75590
rect 7622 75568 7918 75588
rect 14289 75644 14585 75664
rect 14345 75642 14369 75644
rect 14425 75642 14449 75644
rect 14505 75642 14529 75644
rect 14367 75590 14369 75642
rect 14431 75590 14443 75642
rect 14505 75590 14507 75642
rect 14345 75588 14369 75590
rect 14425 75588 14449 75590
rect 14505 75588 14529 75590
rect 14289 75568 14585 75588
rect 5172 75404 5224 75410
rect 5172 75346 5224 75352
rect 7104 75404 7156 75410
rect 7104 75346 7156 75352
rect 4896 75336 4948 75342
rect 4894 75304 4896 75313
rect 4948 75304 4950 75313
rect 4894 75239 4950 75248
rect 4908 74866 4936 75239
rect 5184 75002 5212 75346
rect 7010 75304 7066 75313
rect 7010 75239 7066 75248
rect 7024 75002 7052 75239
rect 5172 74996 5224 75002
rect 5172 74938 5224 74944
rect 7012 74996 7064 75002
rect 7012 74938 7064 74944
rect 4896 74860 4948 74866
rect 4896 74802 4948 74808
rect 4988 74792 5040 74798
rect 3988 74662 4016 74734
rect 4068 74724 4120 74730
rect 4816 74718 4936 74746
rect 4988 74734 5040 74740
rect 6736 74792 6788 74798
rect 6736 74734 6788 74740
rect 4068 74666 4120 74672
rect 3976 74656 4028 74662
rect 3976 74598 4028 74604
rect 4080 74610 4108 74666
rect 4618 74624 4674 74633
rect 3882 73400 3938 73409
rect 3882 73335 3938 73344
rect 3896 72826 3924 73335
rect 3988 73166 4016 74598
rect 4080 74582 4200 74610
rect 4172 74458 4200 74582
rect 4618 74559 4674 74568
rect 4160 74452 4212 74458
rect 4160 74394 4212 74400
rect 4289 74012 4585 74032
rect 4345 74010 4369 74012
rect 4425 74010 4449 74012
rect 4505 74010 4529 74012
rect 4367 73958 4369 74010
rect 4431 73958 4443 74010
rect 4505 73958 4507 74010
rect 4345 73956 4369 73958
rect 4425 73956 4449 73958
rect 4505 73956 4529 73958
rect 4289 73936 4585 73956
rect 4344 73704 4396 73710
rect 4344 73646 4396 73652
rect 4252 73636 4304 73642
rect 4252 73578 4304 73584
rect 3976 73160 4028 73166
rect 4264 73137 4292 73578
rect 4356 73273 4384 73646
rect 4342 73264 4398 73273
rect 4342 73199 4344 73208
rect 4396 73199 4398 73208
rect 4344 73170 4396 73176
rect 3976 73102 4028 73108
rect 4250 73128 4306 73137
rect 4250 73063 4306 73072
rect 4289 72924 4585 72944
rect 4345 72922 4369 72924
rect 4425 72922 4449 72924
rect 4505 72922 4529 72924
rect 4367 72870 4369 72922
rect 4431 72870 4443 72922
rect 4505 72870 4507 72922
rect 4345 72868 4369 72870
rect 4425 72868 4449 72870
rect 4505 72868 4529 72870
rect 4289 72848 4585 72868
rect 3884 72820 3936 72826
rect 3884 72762 3936 72768
rect 4632 72690 4660 74559
rect 4802 73808 4858 73817
rect 4802 73743 4858 73752
rect 4816 73302 4844 73743
rect 4804 73296 4856 73302
rect 4804 73238 4856 73244
rect 4712 73024 4764 73030
rect 4712 72966 4764 72972
rect 4724 72690 4752 72966
rect 4620 72684 4672 72690
rect 4620 72626 4672 72632
rect 4712 72684 4764 72690
rect 4712 72626 4764 72632
rect 4068 72480 4120 72486
rect 4120 72440 4200 72468
rect 4068 72422 4120 72428
rect 3528 72270 3648 72298
rect 3528 68950 3556 72270
rect 3700 72140 3752 72146
rect 3700 72082 3752 72088
rect 3712 71398 3740 72082
rect 3700 71392 3752 71398
rect 3698 71360 3700 71369
rect 3752 71360 3754 71369
rect 3698 71295 3754 71304
rect 4172 70922 4200 72440
rect 4289 71836 4585 71856
rect 4345 71834 4369 71836
rect 4425 71834 4449 71836
rect 4505 71834 4529 71836
rect 4367 71782 4369 71834
rect 4431 71782 4443 71834
rect 4505 71782 4507 71834
rect 4345 71780 4369 71782
rect 4425 71780 4449 71782
rect 4505 71780 4529 71782
rect 4289 71760 4585 71780
rect 4528 71052 4580 71058
rect 4528 70994 4580 71000
rect 4712 71052 4764 71058
rect 4712 70994 4764 71000
rect 4540 70938 4568 70994
rect 4160 70916 4212 70922
rect 4540 70910 4660 70938
rect 4160 70858 4212 70864
rect 4289 70748 4585 70768
rect 4345 70746 4369 70748
rect 4425 70746 4449 70748
rect 4505 70746 4529 70748
rect 4367 70694 4369 70746
rect 4431 70694 4443 70746
rect 4505 70694 4507 70746
rect 4345 70692 4369 70694
rect 4425 70692 4449 70694
rect 4505 70692 4529 70694
rect 4289 70672 4585 70692
rect 4632 70310 4660 70910
rect 4724 70650 4752 70994
rect 4712 70644 4764 70650
rect 4712 70586 4764 70592
rect 4724 70417 4752 70586
rect 4710 70408 4766 70417
rect 4710 70343 4766 70352
rect 4068 70304 4120 70310
rect 4068 70246 4120 70252
rect 4620 70304 4672 70310
rect 4620 70246 4672 70252
rect 3974 69864 4030 69873
rect 3974 69799 4030 69808
rect 3608 69216 3660 69222
rect 3608 69158 3660 69164
rect 3700 69216 3752 69222
rect 3700 69158 3752 69164
rect 3620 69057 3648 69158
rect 3606 69048 3662 69057
rect 3606 68983 3662 68992
rect 3516 68944 3568 68950
rect 3516 68886 3568 68892
rect 3608 68672 3660 68678
rect 3608 68614 3660 68620
rect 3620 68116 3648 68614
rect 3712 68218 3740 69158
rect 3884 68876 3936 68882
rect 3884 68818 3936 68824
rect 3712 68190 3832 68218
rect 3700 68128 3752 68134
rect 3620 68088 3700 68116
rect 3700 68070 3752 68076
rect 3712 67794 3740 68070
rect 3700 67788 3752 67794
rect 3700 67730 3752 67736
rect 3804 67658 3832 68190
rect 3896 68134 3924 68818
rect 3884 68128 3936 68134
rect 3884 68070 3936 68076
rect 3896 67930 3924 68070
rect 3884 67924 3936 67930
rect 3884 67866 3936 67872
rect 3792 67652 3844 67658
rect 3792 67594 3844 67600
rect 3424 66224 3476 66230
rect 3424 66166 3476 66172
rect 3608 66088 3660 66094
rect 3608 66030 3660 66036
rect 3332 65952 3384 65958
rect 3332 65894 3384 65900
rect 3514 65920 3570 65929
rect 3344 65618 3372 65894
rect 3514 65855 3570 65864
rect 3332 65612 3384 65618
rect 3332 65554 3384 65560
rect 3344 65210 3372 65554
rect 3332 65204 3384 65210
rect 3332 65146 3384 65152
rect 3424 64660 3476 64666
rect 3424 64602 3476 64608
rect 3436 63306 3464 64602
rect 3424 63300 3476 63306
rect 3424 63242 3476 63248
rect 3424 62280 3476 62286
rect 3424 62222 3476 62228
rect 3436 61606 3464 62222
rect 3424 61600 3476 61606
rect 3424 61542 3476 61548
rect 3436 61402 3464 61542
rect 3424 61396 3476 61402
rect 3424 61338 3476 61344
rect 3424 61124 3476 61130
rect 3424 61066 3476 61072
rect 3436 60858 3464 61066
rect 3424 60852 3476 60858
rect 3424 60794 3476 60800
rect 3330 60616 3386 60625
rect 3330 60551 3386 60560
rect 3240 51060 3292 51066
rect 3240 51002 3292 51008
rect 3240 50312 3292 50318
rect 3240 50254 3292 50260
rect 3252 49842 3280 50254
rect 3240 49836 3292 49842
rect 3240 49778 3292 49784
rect 3238 49192 3294 49201
rect 3238 49127 3294 49136
rect 3252 48890 3280 49127
rect 3240 48884 3292 48890
rect 3240 48826 3292 48832
rect 3240 47048 3292 47054
rect 3240 46990 3292 46996
rect 3252 46753 3280 46990
rect 3238 46744 3294 46753
rect 3238 46679 3294 46688
rect 3252 46646 3280 46679
rect 3240 46640 3292 46646
rect 3240 46582 3292 46588
rect 3238 45928 3294 45937
rect 3238 45863 3294 45872
rect 3252 43926 3280 45863
rect 3240 43920 3292 43926
rect 3240 43862 3292 43868
rect 3238 43344 3294 43353
rect 3238 43279 3294 43288
rect 3252 41274 3280 43279
rect 3240 41268 3292 41274
rect 3240 41210 3292 41216
rect 3344 39574 3372 60551
rect 3424 60104 3476 60110
rect 3424 60046 3476 60052
rect 3436 59430 3464 60046
rect 3424 59424 3476 59430
rect 3422 59392 3424 59401
rect 3476 59392 3478 59401
rect 3422 59327 3478 59336
rect 3528 59072 3556 65855
rect 3620 64002 3648 66030
rect 3700 65408 3752 65414
rect 3700 65350 3752 65356
rect 3712 65074 3740 65350
rect 3700 65068 3752 65074
rect 3700 65010 3752 65016
rect 3620 63974 3740 64002
rect 3608 63912 3660 63918
rect 3608 63854 3660 63860
rect 3620 59242 3648 63854
rect 3712 61266 3740 63974
rect 3700 61260 3752 61266
rect 3700 61202 3752 61208
rect 3712 60858 3740 61202
rect 3804 61169 3832 67594
rect 3988 67250 4016 69799
rect 4080 69358 4108 70246
rect 4804 69964 4856 69970
rect 4804 69906 4856 69912
rect 4620 69760 4672 69766
rect 4620 69702 4672 69708
rect 4289 69660 4585 69680
rect 4345 69658 4369 69660
rect 4425 69658 4449 69660
rect 4505 69658 4529 69660
rect 4367 69606 4369 69658
rect 4431 69606 4443 69658
rect 4505 69606 4507 69658
rect 4345 69604 4369 69606
rect 4425 69604 4449 69606
rect 4505 69604 4529 69606
rect 4289 69584 4585 69604
rect 4160 69488 4212 69494
rect 4160 69430 4212 69436
rect 4068 69352 4120 69358
rect 4068 69294 4120 69300
rect 4068 68808 4120 68814
rect 4172 68796 4200 69430
rect 4632 69358 4660 69702
rect 4710 69592 4766 69601
rect 4710 69527 4766 69536
rect 4620 69352 4672 69358
rect 4620 69294 4672 69300
rect 4120 68768 4200 68796
rect 4068 68750 4120 68756
rect 4080 67930 4108 68750
rect 4289 68572 4585 68592
rect 4345 68570 4369 68572
rect 4425 68570 4449 68572
rect 4505 68570 4529 68572
rect 4367 68518 4369 68570
rect 4431 68518 4443 68570
rect 4505 68518 4507 68570
rect 4345 68516 4369 68518
rect 4425 68516 4449 68518
rect 4505 68516 4529 68518
rect 4289 68496 4585 68516
rect 4158 68232 4214 68241
rect 4158 68167 4214 68176
rect 4068 67924 4120 67930
rect 4068 67866 4120 67872
rect 4068 67788 4120 67794
rect 4068 67730 4120 67736
rect 3976 67244 4028 67250
rect 3976 67186 4028 67192
rect 3976 65476 4028 65482
rect 3976 65418 4028 65424
rect 3988 64530 4016 65418
rect 4080 65142 4108 67730
rect 4068 65136 4120 65142
rect 4068 65078 4120 65084
rect 4080 64666 4108 65078
rect 4068 64660 4120 64666
rect 4068 64602 4120 64608
rect 3884 64524 3936 64530
rect 3884 64466 3936 64472
rect 3976 64524 4028 64530
rect 3976 64466 4028 64472
rect 3896 63442 3924 64466
rect 4068 64048 4120 64054
rect 4066 64016 4068 64025
rect 4120 64016 4122 64025
rect 4172 63986 4200 68167
rect 4289 67484 4585 67504
rect 4345 67482 4369 67484
rect 4425 67482 4449 67484
rect 4505 67482 4529 67484
rect 4367 67430 4369 67482
rect 4431 67430 4443 67482
rect 4505 67430 4507 67482
rect 4345 67428 4369 67430
rect 4425 67428 4449 67430
rect 4505 67428 4529 67430
rect 4289 67408 4585 67428
rect 4252 67176 4304 67182
rect 4252 67118 4304 67124
rect 4264 66842 4292 67118
rect 4252 66836 4304 66842
rect 4252 66778 4304 66784
rect 4289 66396 4585 66416
rect 4345 66394 4369 66396
rect 4425 66394 4449 66396
rect 4505 66394 4529 66396
rect 4367 66342 4369 66394
rect 4431 66342 4443 66394
rect 4505 66342 4507 66394
rect 4345 66340 4369 66342
rect 4425 66340 4449 66342
rect 4505 66340 4529 66342
rect 4289 66320 4585 66340
rect 4632 65958 4660 69294
rect 4724 68785 4752 69527
rect 4816 69222 4844 69906
rect 4804 69216 4856 69222
rect 4804 69158 4856 69164
rect 4710 68776 4766 68785
rect 4710 68711 4766 68720
rect 4712 67652 4764 67658
rect 4712 67594 4764 67600
rect 4620 65952 4672 65958
rect 4620 65894 4672 65900
rect 4289 65308 4585 65328
rect 4345 65306 4369 65308
rect 4425 65306 4449 65308
rect 4505 65306 4529 65308
rect 4367 65254 4369 65306
rect 4431 65254 4443 65306
rect 4505 65254 4507 65306
rect 4345 65252 4369 65254
rect 4425 65252 4449 65254
rect 4505 65252 4529 65254
rect 4289 65232 4585 65252
rect 4724 65006 4752 67594
rect 4816 65618 4844 69158
rect 4908 67930 4936 74718
rect 5000 74254 5028 74734
rect 5448 74656 5500 74662
rect 5448 74598 5500 74604
rect 5460 74474 5488 74598
rect 5460 74458 5580 74474
rect 5460 74452 5592 74458
rect 5460 74446 5540 74452
rect 5540 74394 5592 74400
rect 6092 74452 6144 74458
rect 6092 74394 6144 74400
rect 5908 74384 5960 74390
rect 5908 74326 5960 74332
rect 5356 74316 5408 74322
rect 5356 74258 5408 74264
rect 4988 74248 5040 74254
rect 4988 74190 5040 74196
rect 5080 74180 5132 74186
rect 5080 74122 5132 74128
rect 5092 73710 5120 74122
rect 5368 73710 5396 74258
rect 5448 74112 5500 74118
rect 5448 74054 5500 74060
rect 5080 73704 5132 73710
rect 5078 73672 5080 73681
rect 5264 73704 5316 73710
rect 5132 73672 5134 73681
rect 5264 73646 5316 73652
rect 5356 73704 5408 73710
rect 5356 73646 5408 73652
rect 5078 73607 5134 73616
rect 5276 73166 5304 73646
rect 5460 73250 5488 74054
rect 5920 73846 5948 74326
rect 5908 73840 5960 73846
rect 5908 73782 5960 73788
rect 5920 73574 5948 73782
rect 6104 73778 6132 74394
rect 6460 74180 6512 74186
rect 6460 74122 6512 74128
rect 6092 73772 6144 73778
rect 6092 73714 6144 73720
rect 5908 73568 5960 73574
rect 5908 73510 5960 73516
rect 6000 73568 6052 73574
rect 6000 73510 6052 73516
rect 5460 73234 5580 73250
rect 5448 73228 5580 73234
rect 5500 73222 5580 73228
rect 5448 73170 5500 73176
rect 4988 73160 5040 73166
rect 4988 73102 5040 73108
rect 5264 73160 5316 73166
rect 5264 73102 5316 73108
rect 5000 72282 5028 73102
rect 5080 73092 5132 73098
rect 5080 73034 5132 73040
rect 4988 72276 5040 72282
rect 4988 72218 5040 72224
rect 5092 72162 5120 73034
rect 5448 72684 5500 72690
rect 5448 72626 5500 72632
rect 5264 72616 5316 72622
rect 5264 72558 5316 72564
rect 5000 72134 5120 72162
rect 5000 68814 5028 72134
rect 5276 71738 5304 72558
rect 5460 72162 5488 72626
rect 5552 72282 5580 73222
rect 5816 73160 5868 73166
rect 5816 73102 5868 73108
rect 5920 73114 5948 73510
rect 6012 73409 6040 73510
rect 5998 73400 6054 73409
rect 5998 73335 6054 73344
rect 6012 73234 6040 73335
rect 6000 73228 6052 73234
rect 6000 73170 6052 73176
rect 5828 72486 5856 73102
rect 5920 73086 6040 73114
rect 5816 72480 5868 72486
rect 5816 72422 5868 72428
rect 5540 72276 5592 72282
rect 5540 72218 5592 72224
rect 5460 72134 5580 72162
rect 5264 71732 5316 71738
rect 5264 71674 5316 71680
rect 5448 71596 5500 71602
rect 5448 71538 5500 71544
rect 5080 71528 5132 71534
rect 5080 71470 5132 71476
rect 5092 71058 5120 71470
rect 5460 71194 5488 71538
rect 5448 71188 5500 71194
rect 5448 71130 5500 71136
rect 5080 71052 5132 71058
rect 5080 70994 5132 71000
rect 5552 70650 5580 72134
rect 5540 70644 5592 70650
rect 5540 70586 5592 70592
rect 5724 70508 5776 70514
rect 5724 70450 5776 70456
rect 5264 69760 5316 69766
rect 5264 69702 5316 69708
rect 4988 68808 5040 68814
rect 4988 68750 5040 68756
rect 5078 68776 5134 68785
rect 5000 68338 5028 68750
rect 5078 68711 5080 68720
rect 5132 68711 5134 68720
rect 5080 68682 5132 68688
rect 4988 68332 5040 68338
rect 4988 68274 5040 68280
rect 4896 67924 4948 67930
rect 4896 67866 4948 67872
rect 4896 67788 4948 67794
rect 4896 67730 4948 67736
rect 4908 67386 4936 67730
rect 4896 67380 4948 67386
rect 4896 67322 4948 67328
rect 4896 65952 4948 65958
rect 4896 65894 4948 65900
rect 4804 65612 4856 65618
rect 4804 65554 4856 65560
rect 4908 65056 4936 65894
rect 4816 65028 4936 65056
rect 4712 65000 4764 65006
rect 4712 64942 4764 64948
rect 4620 64524 4672 64530
rect 4620 64466 4672 64472
rect 4289 64220 4585 64240
rect 4345 64218 4369 64220
rect 4425 64218 4449 64220
rect 4505 64218 4529 64220
rect 4367 64166 4369 64218
rect 4431 64166 4443 64218
rect 4505 64166 4507 64218
rect 4345 64164 4369 64166
rect 4425 64164 4449 64166
rect 4505 64164 4529 64166
rect 4289 64144 4585 64164
rect 4066 63951 4122 63960
rect 4160 63980 4212 63986
rect 4160 63922 4212 63928
rect 4158 63880 4214 63889
rect 4068 63844 4120 63850
rect 4158 63815 4214 63824
rect 4068 63786 4120 63792
rect 3884 63436 3936 63442
rect 3884 63378 3936 63384
rect 3896 62490 3924 63378
rect 3976 63368 4028 63374
rect 3976 63310 4028 63316
rect 3988 63034 4016 63310
rect 4080 63238 4108 63786
rect 4068 63232 4120 63238
rect 4068 63174 4120 63180
rect 3976 63028 4028 63034
rect 3976 62970 4028 62976
rect 4080 62762 4108 63174
rect 4172 63034 4200 63815
rect 4632 63782 4660 64466
rect 4712 63980 4764 63986
rect 4712 63922 4764 63928
rect 4620 63776 4672 63782
rect 4620 63718 4672 63724
rect 4528 63368 4580 63374
rect 4526 63336 4528 63345
rect 4580 63336 4582 63345
rect 4526 63271 4582 63280
rect 4289 63132 4585 63152
rect 4345 63130 4369 63132
rect 4425 63130 4449 63132
rect 4505 63130 4529 63132
rect 4367 63078 4369 63130
rect 4431 63078 4443 63130
rect 4505 63078 4507 63130
rect 4345 63076 4369 63078
rect 4425 63076 4449 63078
rect 4505 63076 4529 63078
rect 4289 63056 4585 63076
rect 4160 63028 4212 63034
rect 4160 62970 4212 62976
rect 4068 62756 4120 62762
rect 4068 62698 4120 62704
rect 4160 62688 4212 62694
rect 4160 62630 4212 62636
rect 3884 62484 3936 62490
rect 3884 62426 3936 62432
rect 3896 61810 3924 62426
rect 3976 62280 4028 62286
rect 3976 62222 4028 62228
rect 3988 61946 4016 62222
rect 4068 62212 4120 62218
rect 4068 62154 4120 62160
rect 3976 61940 4028 61946
rect 3976 61882 4028 61888
rect 3884 61804 3936 61810
rect 3884 61746 3936 61752
rect 4080 61418 4108 62154
rect 3988 61390 4108 61418
rect 3790 61160 3846 61169
rect 3790 61095 3846 61104
rect 3988 60874 4016 61390
rect 4068 61056 4120 61062
rect 4068 60998 4120 61004
rect 3700 60852 3752 60858
rect 3700 60794 3752 60800
rect 3896 60846 4016 60874
rect 3790 60616 3846 60625
rect 3790 60551 3846 60560
rect 3712 60110 3740 60141
rect 3700 60104 3752 60110
rect 3698 60072 3700 60081
rect 3752 60072 3754 60081
rect 3698 60007 3754 60016
rect 3712 59770 3740 60007
rect 3700 59764 3752 59770
rect 3700 59706 3752 59712
rect 3620 59214 3740 59242
rect 3528 59044 3648 59072
rect 3424 58336 3476 58342
rect 3424 58278 3476 58284
rect 3436 56982 3464 58278
rect 3516 57860 3568 57866
rect 3516 57802 3568 57808
rect 3424 56976 3476 56982
rect 3424 56918 3476 56924
rect 3528 56914 3556 57802
rect 3516 56908 3568 56914
rect 3516 56850 3568 56856
rect 3528 56710 3556 56850
rect 3516 56704 3568 56710
rect 3516 56646 3568 56652
rect 3516 56432 3568 56438
rect 3516 56374 3568 56380
rect 3528 55418 3556 56374
rect 3424 55412 3476 55418
rect 3424 55354 3476 55360
rect 3516 55412 3568 55418
rect 3516 55354 3568 55360
rect 3436 48346 3464 55354
rect 3528 54126 3556 55354
rect 3516 54120 3568 54126
rect 3516 54062 3568 54068
rect 3620 53582 3648 59044
rect 3712 57934 3740 59214
rect 3700 57928 3752 57934
rect 3700 57870 3752 57876
rect 3712 57458 3740 57870
rect 3700 57452 3752 57458
rect 3700 57394 3752 57400
rect 3700 57248 3752 57254
rect 3700 57190 3752 57196
rect 3712 56370 3740 57190
rect 3700 56364 3752 56370
rect 3700 56306 3752 56312
rect 3698 56264 3754 56273
rect 3698 56199 3754 56208
rect 3608 53576 3660 53582
rect 3608 53518 3660 53524
rect 3516 52896 3568 52902
rect 3516 52838 3568 52844
rect 3528 52698 3556 52838
rect 3516 52692 3568 52698
rect 3516 52634 3568 52640
rect 3516 52488 3568 52494
rect 3516 52430 3568 52436
rect 3528 51785 3556 52430
rect 3514 51776 3570 51785
rect 3514 51711 3570 51720
rect 3606 51368 3662 51377
rect 3606 51303 3662 51312
rect 3516 51264 3568 51270
rect 3516 51206 3568 51212
rect 3528 50318 3556 51206
rect 3516 50312 3568 50318
rect 3516 50254 3568 50260
rect 3516 49292 3568 49298
rect 3516 49234 3568 49240
rect 3528 48890 3556 49234
rect 3516 48884 3568 48890
rect 3516 48826 3568 48832
rect 3424 48340 3476 48346
rect 3424 48282 3476 48288
rect 3422 48240 3478 48249
rect 3422 48175 3478 48184
rect 3436 45490 3464 48175
rect 3620 47122 3648 51303
rect 3712 50454 3740 56199
rect 3804 51474 3832 60551
rect 3792 51468 3844 51474
rect 3792 51410 3844 51416
rect 3792 51332 3844 51338
rect 3792 51274 3844 51280
rect 3700 50448 3752 50454
rect 3700 50390 3752 50396
rect 3700 50312 3752 50318
rect 3700 50254 3752 50260
rect 3712 48754 3740 50254
rect 3700 48748 3752 48754
rect 3700 48690 3752 48696
rect 3700 48340 3752 48346
rect 3700 48282 3752 48288
rect 3516 47116 3568 47122
rect 3516 47058 3568 47064
rect 3608 47116 3660 47122
rect 3608 47058 3660 47064
rect 3528 46374 3556 47058
rect 3620 46714 3648 47058
rect 3608 46708 3660 46714
rect 3608 46650 3660 46656
rect 3516 46368 3568 46374
rect 3516 46310 3568 46316
rect 3606 46064 3662 46073
rect 3606 45999 3662 46008
rect 3516 45960 3568 45966
rect 3516 45902 3568 45908
rect 3528 45626 3556 45902
rect 3516 45620 3568 45626
rect 3516 45562 3568 45568
rect 3424 45484 3476 45490
rect 3424 45426 3476 45432
rect 3528 45234 3556 45562
rect 3436 45206 3556 45234
rect 3436 42702 3464 45206
rect 3516 43648 3568 43654
rect 3516 43590 3568 43596
rect 3528 42770 3556 43590
rect 3620 43314 3648 45999
rect 3712 43450 3740 48282
rect 3700 43444 3752 43450
rect 3700 43386 3752 43392
rect 3608 43308 3660 43314
rect 3608 43250 3660 43256
rect 3712 43246 3740 43386
rect 3700 43240 3752 43246
rect 3700 43182 3752 43188
rect 3712 42820 3740 43182
rect 3804 42906 3832 51274
rect 3792 42900 3844 42906
rect 3792 42842 3844 42848
rect 3620 42792 3740 42820
rect 3790 42800 3846 42809
rect 3516 42764 3568 42770
rect 3516 42706 3568 42712
rect 3424 42696 3476 42702
rect 3424 42638 3476 42644
rect 3436 41818 3464 42638
rect 3528 42362 3556 42706
rect 3516 42356 3568 42362
rect 3516 42298 3568 42304
rect 3424 41812 3476 41818
rect 3424 41754 3476 41760
rect 3620 39574 3648 42792
rect 3790 42735 3846 42744
rect 3698 40216 3754 40225
rect 3698 40151 3700 40160
rect 3752 40151 3754 40160
rect 3700 40122 3752 40128
rect 3332 39568 3384 39574
rect 3332 39510 3384 39516
rect 3608 39568 3660 39574
rect 3608 39510 3660 39516
rect 3240 39500 3292 39506
rect 3240 39442 3292 39448
rect 3700 39500 3752 39506
rect 3700 39442 3752 39448
rect 3252 39098 3280 39442
rect 3332 39432 3384 39438
rect 3332 39374 3384 39380
rect 3344 39098 3372 39374
rect 3240 39092 3292 39098
rect 3240 39034 3292 39040
rect 3332 39092 3384 39098
rect 3332 39034 3384 39040
rect 3332 38888 3384 38894
rect 3332 38830 3384 38836
rect 3238 38312 3294 38321
rect 3238 38247 3294 38256
rect 3252 38010 3280 38247
rect 3240 38004 3292 38010
rect 3240 37946 3292 37952
rect 3240 37120 3292 37126
rect 3240 37062 3292 37068
rect 3252 36582 3280 37062
rect 3240 36576 3292 36582
rect 3240 36518 3292 36524
rect 3252 33998 3280 36518
rect 3240 33992 3292 33998
rect 3240 33934 3292 33940
rect 3252 33386 3280 33934
rect 3240 33380 3292 33386
rect 3240 33322 3292 33328
rect 3344 32026 3372 38830
rect 3712 38826 3740 39442
rect 3804 39098 3832 42735
rect 3792 39092 3844 39098
rect 3792 39034 3844 39040
rect 3804 38894 3832 39034
rect 3792 38888 3844 38894
rect 3792 38830 3844 38836
rect 3700 38820 3752 38826
rect 3700 38762 3752 38768
rect 3516 38412 3568 38418
rect 3516 38354 3568 38360
rect 3528 38010 3556 38354
rect 3516 38004 3568 38010
rect 3516 37946 3568 37952
rect 3514 37904 3570 37913
rect 3514 37839 3570 37848
rect 3422 36816 3478 36825
rect 3422 36751 3478 36760
rect 3332 32020 3384 32026
rect 3332 31962 3384 31968
rect 3148 31952 3200 31958
rect 3148 31894 3200 31900
rect 3332 31748 3384 31754
rect 3332 31690 3384 31696
rect 3148 29028 3200 29034
rect 3148 28970 3200 28976
rect 3160 25265 3188 28970
rect 3344 27062 3372 31690
rect 3436 30870 3464 36751
rect 3528 34066 3556 37839
rect 3608 37800 3660 37806
rect 3608 37742 3660 37748
rect 3620 37262 3648 37742
rect 3712 37330 3740 38762
rect 3792 37664 3844 37670
rect 3792 37606 3844 37612
rect 3700 37324 3752 37330
rect 3700 37266 3752 37272
rect 3608 37256 3660 37262
rect 3608 37198 3660 37204
rect 3804 37097 3832 37606
rect 3790 37088 3846 37097
rect 3790 37023 3846 37032
rect 3896 35834 3924 60846
rect 4080 60738 4108 60998
rect 3988 60710 4108 60738
rect 3988 58460 4016 60710
rect 4068 58948 4120 58954
rect 4068 58890 4120 58896
rect 4080 58614 4108 58890
rect 4068 58608 4120 58614
rect 4068 58550 4120 58556
rect 3988 58432 4108 58460
rect 3974 57896 4030 57905
rect 3974 57831 4030 57840
rect 3988 47410 4016 57831
rect 4080 56438 4108 58432
rect 4068 56432 4120 56438
rect 4068 56374 4120 56380
rect 4068 56160 4120 56166
rect 4068 56102 4120 56108
rect 4080 54534 4108 56102
rect 4068 54528 4120 54534
rect 4068 54470 4120 54476
rect 4080 53038 4108 54470
rect 4068 53032 4120 53038
rect 4068 52974 4120 52980
rect 4068 52896 4120 52902
rect 4068 52838 4120 52844
rect 4080 51406 4108 52838
rect 4172 52018 4200 62630
rect 4289 62044 4585 62064
rect 4345 62042 4369 62044
rect 4425 62042 4449 62044
rect 4505 62042 4529 62044
rect 4367 61990 4369 62042
rect 4431 61990 4443 62042
rect 4505 61990 4507 62042
rect 4345 61988 4369 61990
rect 4425 61988 4449 61990
rect 4505 61988 4529 61990
rect 4289 61968 4585 61988
rect 4632 61062 4660 63718
rect 4724 62694 4752 63922
rect 4816 62830 4844 65028
rect 4896 64932 4948 64938
rect 4896 64874 4948 64880
rect 4908 64326 4936 64874
rect 4896 64320 4948 64326
rect 4896 64262 4948 64268
rect 4908 63850 4936 64262
rect 4896 63844 4948 63850
rect 4896 63786 4948 63792
rect 4804 62824 4856 62830
rect 4804 62766 4856 62772
rect 4712 62688 4764 62694
rect 4712 62630 4764 62636
rect 4804 62688 4856 62694
rect 4804 62630 4856 62636
rect 4816 62490 4844 62630
rect 4804 62484 4856 62490
rect 4804 62426 4856 62432
rect 4712 62212 4764 62218
rect 4712 62154 4764 62160
rect 4724 61742 4752 62154
rect 4712 61736 4764 61742
rect 4712 61678 4764 61684
rect 4724 61334 4752 61678
rect 4816 61402 4844 62426
rect 4804 61396 4856 61402
rect 4804 61338 4856 61344
rect 4712 61328 4764 61334
rect 4712 61270 4764 61276
rect 4620 61056 4672 61062
rect 4620 60998 4672 61004
rect 4289 60956 4585 60976
rect 4345 60954 4369 60956
rect 4425 60954 4449 60956
rect 4505 60954 4529 60956
rect 4367 60902 4369 60954
rect 4431 60902 4443 60954
rect 4505 60902 4507 60954
rect 4345 60900 4369 60902
rect 4425 60900 4449 60902
rect 4505 60900 4529 60902
rect 4289 60880 4585 60900
rect 4620 60648 4672 60654
rect 4620 60590 4672 60596
rect 4344 60512 4396 60518
rect 4342 60480 4344 60489
rect 4396 60480 4398 60489
rect 4342 60415 4398 60424
rect 4632 60314 4660 60590
rect 4620 60308 4672 60314
rect 4620 60250 4672 60256
rect 4289 59868 4585 59888
rect 4345 59866 4369 59868
rect 4425 59866 4449 59868
rect 4505 59866 4529 59868
rect 4367 59814 4369 59866
rect 4431 59814 4443 59866
rect 4505 59814 4507 59866
rect 4345 59812 4369 59814
rect 4425 59812 4449 59814
rect 4505 59812 4529 59814
rect 4289 59792 4585 59812
rect 4618 59256 4674 59265
rect 4618 59191 4674 59200
rect 4632 59090 4660 59191
rect 4620 59084 4672 59090
rect 4620 59026 4672 59032
rect 4289 58780 4585 58800
rect 4345 58778 4369 58780
rect 4425 58778 4449 58780
rect 4505 58778 4529 58780
rect 4367 58726 4369 58778
rect 4431 58726 4443 58778
rect 4505 58726 4507 58778
rect 4345 58724 4369 58726
rect 4425 58724 4449 58726
rect 4505 58724 4529 58726
rect 4289 58704 4585 58724
rect 4632 58682 4660 59026
rect 4620 58676 4672 58682
rect 4620 58618 4672 58624
rect 4632 58478 4660 58618
rect 4620 58472 4672 58478
rect 4620 58414 4672 58420
rect 4620 57928 4672 57934
rect 4620 57870 4672 57876
rect 4289 57692 4585 57712
rect 4345 57690 4369 57692
rect 4425 57690 4449 57692
rect 4505 57690 4529 57692
rect 4367 57638 4369 57690
rect 4431 57638 4443 57690
rect 4505 57638 4507 57690
rect 4345 57636 4369 57638
rect 4425 57636 4449 57638
rect 4505 57636 4529 57638
rect 4289 57616 4585 57636
rect 4632 57254 4660 57870
rect 4620 57248 4672 57254
rect 4620 57190 4672 57196
rect 4289 56604 4585 56624
rect 4345 56602 4369 56604
rect 4425 56602 4449 56604
rect 4505 56602 4529 56604
rect 4367 56550 4369 56602
rect 4431 56550 4443 56602
rect 4505 56550 4507 56602
rect 4345 56548 4369 56550
rect 4425 56548 4449 56550
rect 4505 56548 4529 56550
rect 4289 56528 4585 56548
rect 4344 56296 4396 56302
rect 4344 56238 4396 56244
rect 4356 55690 4384 56238
rect 4724 55876 4752 61270
rect 4816 59770 4844 61338
rect 4804 59764 4856 59770
rect 4804 59706 4856 59712
rect 4816 59226 4844 59706
rect 4804 59220 4856 59226
rect 4804 59162 4856 59168
rect 4804 57996 4856 58002
rect 4804 57938 4856 57944
rect 4816 57050 4844 57938
rect 4804 57044 4856 57050
rect 4804 56986 4856 56992
rect 4804 56908 4856 56914
rect 4804 56850 4856 56856
rect 4816 56506 4844 56850
rect 4804 56500 4856 56506
rect 4804 56442 4856 56448
rect 4816 56273 4844 56442
rect 4802 56264 4858 56273
rect 4802 56199 4858 56208
rect 4804 56160 4856 56166
rect 4804 56102 4856 56108
rect 4632 55848 4752 55876
rect 4344 55684 4396 55690
rect 4344 55626 4396 55632
rect 4289 55516 4585 55536
rect 4345 55514 4369 55516
rect 4425 55514 4449 55516
rect 4505 55514 4529 55516
rect 4367 55462 4369 55514
rect 4431 55462 4443 55514
rect 4505 55462 4507 55514
rect 4345 55460 4369 55462
rect 4425 55460 4449 55462
rect 4505 55460 4529 55462
rect 4289 55440 4585 55460
rect 4436 55072 4488 55078
rect 4434 55040 4436 55049
rect 4488 55040 4490 55049
rect 4434 54975 4490 54984
rect 4289 54428 4585 54448
rect 4345 54426 4369 54428
rect 4425 54426 4449 54428
rect 4505 54426 4529 54428
rect 4367 54374 4369 54426
rect 4431 54374 4443 54426
rect 4505 54374 4507 54426
rect 4345 54372 4369 54374
rect 4425 54372 4449 54374
rect 4505 54372 4529 54374
rect 4289 54352 4585 54372
rect 4528 54052 4580 54058
rect 4528 53994 4580 54000
rect 4252 53984 4304 53990
rect 4252 53926 4304 53932
rect 4264 53718 4292 53926
rect 4540 53718 4568 53994
rect 4252 53712 4304 53718
rect 4252 53654 4304 53660
rect 4528 53712 4580 53718
rect 4528 53654 4580 53660
rect 4342 53544 4398 53553
rect 4342 53479 4344 53488
rect 4396 53479 4398 53488
rect 4344 53450 4396 53456
rect 4289 53340 4585 53360
rect 4345 53338 4369 53340
rect 4425 53338 4449 53340
rect 4505 53338 4529 53340
rect 4367 53286 4369 53338
rect 4431 53286 4443 53338
rect 4505 53286 4507 53338
rect 4345 53284 4369 53286
rect 4425 53284 4449 53286
rect 4505 53284 4529 53286
rect 4289 53264 4585 53284
rect 4526 53136 4582 53145
rect 4526 53071 4582 53080
rect 4540 53038 4568 53071
rect 4528 53032 4580 53038
rect 4528 52974 4580 52980
rect 4540 52630 4568 52974
rect 4528 52624 4580 52630
rect 4528 52566 4580 52572
rect 4289 52252 4585 52272
rect 4345 52250 4369 52252
rect 4425 52250 4449 52252
rect 4505 52250 4529 52252
rect 4367 52198 4369 52250
rect 4431 52198 4443 52250
rect 4505 52198 4507 52250
rect 4345 52196 4369 52198
rect 4425 52196 4449 52198
rect 4505 52196 4529 52198
rect 4289 52176 4585 52196
rect 4160 52012 4212 52018
rect 4160 51954 4212 51960
rect 4528 51944 4580 51950
rect 4528 51886 4580 51892
rect 4160 51876 4212 51882
rect 4160 51818 4212 51824
rect 4068 51400 4120 51406
rect 4068 51342 4120 51348
rect 4080 51066 4108 51342
rect 4068 51060 4120 51066
rect 4068 51002 4120 51008
rect 4172 50386 4200 51818
rect 4540 51338 4568 51886
rect 4528 51332 4580 51338
rect 4528 51274 4580 51280
rect 4289 51164 4585 51184
rect 4345 51162 4369 51164
rect 4425 51162 4449 51164
rect 4505 51162 4529 51164
rect 4367 51110 4369 51162
rect 4431 51110 4443 51162
rect 4505 51110 4507 51162
rect 4345 51108 4369 51110
rect 4425 51108 4449 51110
rect 4505 51108 4529 51110
rect 4289 51088 4585 51108
rect 4528 50992 4580 50998
rect 4528 50934 4580 50940
rect 4252 50720 4304 50726
rect 4540 50708 4568 50934
rect 4632 50810 4660 55848
rect 4712 55616 4764 55622
rect 4712 55558 4764 55564
rect 4724 55146 4752 55558
rect 4712 55140 4764 55146
rect 4712 55082 4764 55088
rect 4816 55078 4844 56102
rect 4908 55894 4936 63786
rect 5000 62880 5028 68274
rect 5092 68270 5120 68682
rect 5080 68264 5132 68270
rect 5080 68206 5132 68212
rect 5092 66570 5120 68206
rect 5172 67584 5224 67590
rect 5172 67526 5224 67532
rect 5184 67046 5212 67526
rect 5276 67153 5304 69702
rect 5354 69184 5410 69193
rect 5354 69119 5410 69128
rect 5368 68882 5396 69119
rect 5540 69012 5592 69018
rect 5540 68954 5592 68960
rect 5356 68876 5408 68882
rect 5356 68818 5408 68824
rect 5368 68202 5396 68818
rect 5356 68196 5408 68202
rect 5356 68138 5408 68144
rect 5262 67144 5318 67153
rect 5262 67079 5318 67088
rect 5172 67040 5224 67046
rect 5172 66982 5224 66988
rect 5080 66564 5132 66570
rect 5080 66506 5132 66512
rect 5184 66502 5212 66982
rect 5276 66706 5304 67079
rect 5264 66700 5316 66706
rect 5264 66642 5316 66648
rect 5172 66496 5224 66502
rect 5172 66438 5224 66444
rect 5184 66298 5212 66438
rect 5172 66292 5224 66298
rect 5172 66234 5224 66240
rect 5080 66088 5132 66094
rect 5080 66030 5132 66036
rect 5092 65414 5120 66030
rect 5080 65408 5132 65414
rect 5080 65350 5132 65356
rect 5092 63782 5120 65350
rect 5080 63776 5132 63782
rect 5080 63718 5132 63724
rect 5000 62852 5120 62880
rect 4988 62756 5040 62762
rect 4988 62698 5040 62704
rect 5000 60625 5028 62698
rect 4986 60616 5042 60625
rect 4986 60551 5042 60560
rect 4988 59084 5040 59090
rect 4988 59026 5040 59032
rect 5000 58857 5028 59026
rect 4986 58848 5042 58857
rect 4986 58783 5042 58792
rect 5000 58682 5028 58783
rect 4988 58676 5040 58682
rect 4988 58618 5040 58624
rect 5092 58562 5120 62852
rect 5000 58534 5120 58562
rect 5000 56506 5028 58534
rect 5080 58336 5132 58342
rect 5080 58278 5132 58284
rect 4988 56500 5040 56506
rect 4988 56442 5040 56448
rect 4988 56364 5040 56370
rect 4988 56306 5040 56312
rect 4896 55888 4948 55894
rect 4896 55830 4948 55836
rect 4804 55072 4856 55078
rect 4804 55014 4856 55020
rect 4908 54874 4936 55830
rect 5000 55826 5028 56306
rect 5092 56137 5120 58278
rect 5078 56128 5134 56137
rect 5078 56063 5134 56072
rect 5184 55944 5212 66234
rect 5276 65210 5304 66642
rect 5264 65204 5316 65210
rect 5264 65146 5316 65152
rect 5264 63912 5316 63918
rect 5264 63854 5316 63860
rect 5276 63578 5304 63854
rect 5264 63572 5316 63578
rect 5264 63514 5316 63520
rect 5368 63458 5396 68138
rect 5446 66192 5502 66201
rect 5446 66127 5502 66136
rect 5460 65550 5488 66127
rect 5448 65544 5500 65550
rect 5448 65486 5500 65492
rect 5552 65498 5580 68954
rect 5632 68264 5684 68270
rect 5632 68206 5684 68212
rect 5644 67182 5672 68206
rect 5632 67176 5684 67182
rect 5632 67118 5684 67124
rect 5632 66700 5684 66706
rect 5632 66642 5684 66648
rect 5644 66162 5672 66642
rect 5632 66156 5684 66162
rect 5632 66098 5684 66104
rect 5460 64025 5488 65486
rect 5552 65470 5672 65498
rect 5540 65408 5592 65414
rect 5540 65350 5592 65356
rect 5552 65074 5580 65350
rect 5540 65068 5592 65074
rect 5540 65010 5592 65016
rect 5446 64016 5502 64025
rect 5446 63951 5502 63960
rect 5276 63430 5396 63458
rect 5276 61010 5304 63430
rect 5460 63322 5488 63951
rect 5644 63481 5672 65470
rect 5630 63472 5686 63481
rect 5630 63407 5686 63416
rect 5368 63294 5488 63322
rect 5368 61690 5396 63294
rect 5644 63050 5672 63407
rect 5460 63034 5672 63050
rect 5448 63028 5672 63034
rect 5500 63022 5672 63028
rect 5448 62970 5500 62976
rect 5632 62824 5684 62830
rect 5632 62766 5684 62772
rect 5368 61662 5580 61690
rect 5448 61600 5500 61606
rect 5448 61542 5500 61548
rect 5460 61266 5488 61542
rect 5448 61260 5500 61266
rect 5448 61202 5500 61208
rect 5276 60982 5396 61010
rect 5264 60852 5316 60858
rect 5264 60794 5316 60800
rect 5092 55916 5212 55944
rect 4988 55820 5040 55826
rect 4988 55762 5040 55768
rect 4896 54868 4948 54874
rect 4816 54828 4896 54856
rect 4712 54120 4764 54126
rect 4712 54062 4764 54068
rect 4724 52698 4752 54062
rect 4712 52692 4764 52698
rect 4712 52634 4764 52640
rect 4816 51898 4844 54828
rect 4896 54810 4948 54816
rect 4896 53644 4948 53650
rect 4896 53586 4948 53592
rect 4908 53242 4936 53586
rect 4988 53440 5040 53446
rect 4988 53382 5040 53388
rect 4896 53236 4948 53242
rect 4896 53178 4948 53184
rect 5000 52018 5028 53382
rect 4988 52012 5040 52018
rect 4988 51954 5040 51960
rect 4816 51870 5028 51898
rect 5092 51882 5120 55916
rect 5172 55820 5224 55826
rect 5172 55762 5224 55768
rect 5184 55282 5212 55762
rect 5172 55276 5224 55282
rect 5172 55218 5224 55224
rect 5172 53712 5224 53718
rect 5172 53654 5224 53660
rect 5184 52698 5212 53654
rect 5172 52692 5224 52698
rect 5172 52634 5224 52640
rect 5170 52184 5226 52193
rect 5170 52119 5226 52128
rect 4712 51808 4764 51814
rect 4712 51750 4764 51756
rect 4804 51808 4856 51814
rect 4804 51750 4856 51756
rect 4724 51105 4752 51750
rect 4710 51096 4766 51105
rect 4710 51031 4766 51040
rect 4632 50782 4752 50810
rect 4540 50680 4660 50708
rect 4252 50662 4304 50668
rect 4068 50380 4120 50386
rect 4068 50322 4120 50328
rect 4160 50380 4212 50386
rect 4160 50322 4212 50328
rect 4080 50289 4108 50322
rect 4066 50280 4122 50289
rect 4066 50215 4122 50224
rect 4080 49298 4108 50215
rect 4172 49978 4200 50322
rect 4264 50318 4292 50662
rect 4252 50312 4304 50318
rect 4252 50254 4304 50260
rect 4289 50076 4585 50096
rect 4345 50074 4369 50076
rect 4425 50074 4449 50076
rect 4505 50074 4529 50076
rect 4367 50022 4369 50074
rect 4431 50022 4443 50074
rect 4505 50022 4507 50074
rect 4345 50020 4369 50022
rect 4425 50020 4449 50022
rect 4505 50020 4529 50022
rect 4289 50000 4585 50020
rect 4160 49972 4212 49978
rect 4160 49914 4212 49920
rect 4068 49292 4120 49298
rect 4068 49234 4120 49240
rect 4172 47569 4200 49914
rect 4289 48988 4585 49008
rect 4345 48986 4369 48988
rect 4425 48986 4449 48988
rect 4505 48986 4529 48988
rect 4367 48934 4369 48986
rect 4431 48934 4443 48986
rect 4505 48934 4507 48986
rect 4345 48932 4369 48934
rect 4425 48932 4449 48934
rect 4505 48932 4529 48934
rect 4289 48912 4585 48932
rect 4289 47900 4585 47920
rect 4345 47898 4369 47900
rect 4425 47898 4449 47900
rect 4505 47898 4529 47900
rect 4367 47846 4369 47898
rect 4431 47846 4443 47898
rect 4505 47846 4507 47898
rect 4345 47844 4369 47846
rect 4425 47844 4449 47846
rect 4505 47844 4529 47846
rect 4289 47824 4585 47844
rect 4158 47560 4214 47569
rect 4158 47495 4214 47504
rect 3988 47382 4200 47410
rect 3976 47048 4028 47054
rect 3976 46990 4028 46996
rect 4068 47048 4120 47054
rect 4068 46990 4120 46996
rect 3988 44946 4016 46990
rect 4080 46714 4108 46990
rect 4068 46708 4120 46714
rect 4068 46650 4120 46656
rect 4068 46368 4120 46374
rect 4068 46310 4120 46316
rect 4080 46170 4108 46310
rect 4068 46164 4120 46170
rect 4068 46106 4120 46112
rect 4068 45960 4120 45966
rect 4068 45902 4120 45908
rect 4080 45286 4108 45902
rect 4068 45280 4120 45286
rect 4068 45222 4120 45228
rect 3976 44940 4028 44946
rect 3976 44882 4028 44888
rect 3988 44538 4016 44882
rect 4068 44872 4120 44878
rect 4068 44814 4120 44820
rect 3976 44532 4028 44538
rect 3976 44474 4028 44480
rect 4080 44470 4108 44814
rect 4068 44464 4120 44470
rect 3974 44432 4030 44441
rect 4068 44406 4120 44412
rect 3974 44367 4030 44376
rect 3988 44334 4016 44367
rect 3976 44328 4028 44334
rect 3976 44270 4028 44276
rect 4172 43926 4200 47382
rect 4289 46812 4585 46832
rect 4345 46810 4369 46812
rect 4425 46810 4449 46812
rect 4505 46810 4529 46812
rect 4367 46758 4369 46810
rect 4431 46758 4443 46810
rect 4505 46758 4507 46810
rect 4345 46756 4369 46758
rect 4425 46756 4449 46758
rect 4505 46756 4529 46758
rect 4289 46736 4585 46756
rect 4526 46608 4582 46617
rect 4526 46543 4528 46552
rect 4580 46543 4582 46552
rect 4528 46514 4580 46520
rect 4289 45724 4585 45744
rect 4345 45722 4369 45724
rect 4425 45722 4449 45724
rect 4505 45722 4529 45724
rect 4367 45670 4369 45722
rect 4431 45670 4443 45722
rect 4505 45670 4507 45722
rect 4345 45668 4369 45670
rect 4425 45668 4449 45670
rect 4505 45668 4529 45670
rect 4289 45648 4585 45668
rect 4250 45112 4306 45121
rect 4250 45047 4252 45056
rect 4304 45047 4306 45056
rect 4252 45018 4304 45024
rect 4289 44636 4585 44656
rect 4345 44634 4369 44636
rect 4425 44634 4449 44636
rect 4505 44634 4529 44636
rect 4367 44582 4369 44634
rect 4431 44582 4443 44634
rect 4505 44582 4507 44634
rect 4345 44580 4369 44582
rect 4425 44580 4449 44582
rect 4505 44580 4529 44582
rect 4289 44560 4585 44580
rect 4252 44464 4304 44470
rect 4252 44406 4304 44412
rect 4160 43920 4212 43926
rect 4160 43862 4212 43868
rect 3976 43852 4028 43858
rect 3976 43794 4028 43800
rect 3988 43450 4016 43794
rect 4068 43784 4120 43790
rect 4264 43738 4292 44406
rect 4068 43726 4120 43732
rect 4080 43450 4108 43726
rect 4172 43710 4292 43738
rect 3976 43444 4028 43450
rect 3976 43386 4028 43392
rect 4068 43444 4120 43450
rect 4068 43386 4120 43392
rect 3988 43081 4016 43386
rect 3974 43072 4030 43081
rect 3974 43007 4030 43016
rect 3974 42936 4030 42945
rect 3974 42871 4030 42880
rect 4068 42900 4120 42906
rect 3988 38486 4016 42871
rect 4068 42842 4120 42848
rect 3976 38480 4028 38486
rect 3976 38422 4028 38428
rect 3976 38344 4028 38350
rect 3976 38286 4028 38292
rect 3988 37806 4016 38286
rect 3976 37800 4028 37806
rect 3976 37742 4028 37748
rect 3976 37256 4028 37262
rect 3976 37198 4028 37204
rect 3988 36854 4016 37198
rect 3976 36848 4028 36854
rect 3976 36790 4028 36796
rect 3884 35828 3936 35834
rect 3884 35770 3936 35776
rect 3976 35080 4028 35086
rect 3974 35048 3976 35057
rect 4028 35048 4030 35057
rect 3974 34983 4030 34992
rect 3516 34060 3568 34066
rect 3516 34002 3568 34008
rect 3528 33658 3556 34002
rect 3516 33652 3568 33658
rect 3516 33594 3568 33600
rect 3976 33448 4028 33454
rect 3976 33390 4028 33396
rect 3792 33312 3844 33318
rect 3792 33254 3844 33260
rect 3804 33017 3832 33254
rect 3790 33008 3846 33017
rect 3790 32943 3846 32952
rect 3516 32768 3568 32774
rect 3516 32710 3568 32716
rect 3528 32570 3556 32710
rect 3516 32564 3568 32570
rect 3516 32506 3568 32512
rect 3528 32230 3556 32506
rect 3516 32224 3568 32230
rect 3516 32166 3568 32172
rect 3516 32020 3568 32026
rect 3516 31962 3568 31968
rect 3424 30864 3476 30870
rect 3424 30806 3476 30812
rect 3424 28960 3476 28966
rect 3424 28902 3476 28908
rect 3436 28762 3464 28902
rect 3424 28756 3476 28762
rect 3424 28698 3476 28704
rect 3528 27538 3556 31962
rect 3698 30696 3754 30705
rect 3698 30631 3754 30640
rect 3712 29782 3740 30631
rect 3700 29776 3752 29782
rect 3700 29718 3752 29724
rect 3608 28620 3660 28626
rect 3608 28562 3660 28568
rect 3620 28218 3648 28562
rect 3608 28212 3660 28218
rect 3608 28154 3660 28160
rect 3516 27532 3568 27538
rect 3516 27474 3568 27480
rect 3424 27328 3476 27334
rect 3424 27270 3476 27276
rect 3332 27056 3384 27062
rect 3332 26998 3384 27004
rect 3240 26376 3292 26382
rect 3240 26318 3292 26324
rect 3252 25809 3280 26318
rect 3344 26042 3372 26998
rect 3436 26353 3464 27270
rect 3528 27130 3556 27474
rect 3516 27124 3568 27130
rect 3516 27066 3568 27072
rect 3528 26450 3556 27066
rect 3608 26920 3660 26926
rect 3608 26862 3660 26868
rect 3620 26518 3648 26862
rect 3608 26512 3660 26518
rect 3608 26454 3660 26460
rect 3516 26444 3568 26450
rect 3516 26386 3568 26392
rect 3422 26344 3478 26353
rect 3422 26279 3478 26288
rect 3332 26036 3384 26042
rect 3332 25978 3384 25984
rect 3436 25922 3464 26279
rect 3528 26042 3556 26386
rect 3516 26036 3568 26042
rect 3516 25978 3568 25984
rect 3436 25894 3648 25922
rect 3238 25800 3294 25809
rect 3238 25735 3294 25744
rect 3146 25256 3202 25265
rect 3146 25191 3202 25200
rect 3516 24676 3568 24682
rect 3516 24618 3568 24624
rect 3148 23588 3200 23594
rect 3148 23530 3200 23536
rect 3160 23089 3188 23530
rect 3330 23488 3386 23497
rect 3330 23423 3386 23432
rect 3146 23080 3202 23089
rect 3146 23015 3202 23024
rect 3344 20505 3372 23423
rect 3424 21888 3476 21894
rect 3424 21830 3476 21836
rect 3436 21593 3464 21830
rect 3422 21584 3478 21593
rect 3422 21519 3478 21528
rect 3422 21040 3478 21049
rect 3422 20975 3478 20984
rect 3330 20496 3386 20505
rect 3330 20431 3386 20440
rect 3436 19922 3464 20975
rect 3528 20482 3556 24618
rect 3620 20602 3648 25894
rect 3700 25832 3752 25838
rect 3700 25774 3752 25780
rect 3712 25158 3740 25774
rect 3884 25356 3936 25362
rect 3884 25298 3936 25304
rect 3792 25220 3844 25226
rect 3792 25162 3844 25168
rect 3700 25152 3752 25158
rect 3700 25094 3752 25100
rect 3712 24954 3740 25094
rect 3700 24948 3752 24954
rect 3700 24890 3752 24896
rect 3804 24698 3832 25162
rect 3896 24886 3924 25298
rect 3884 24880 3936 24886
rect 3884 24822 3936 24828
rect 3884 24744 3936 24750
rect 3804 24692 3884 24698
rect 3804 24686 3936 24692
rect 3804 24670 3924 24686
rect 3896 23322 3924 24670
rect 3884 23316 3936 23322
rect 3884 23258 3936 23264
rect 3792 23180 3844 23186
rect 3792 23122 3844 23128
rect 3804 22438 3832 23122
rect 3792 22432 3844 22438
rect 3792 22374 3844 22380
rect 3804 22234 3832 22374
rect 3792 22228 3844 22234
rect 3792 22170 3844 22176
rect 3896 22166 3924 23258
rect 3884 22160 3936 22166
rect 3884 22102 3936 22108
rect 3884 21004 3936 21010
rect 3884 20946 3936 20952
rect 3608 20596 3660 20602
rect 3608 20538 3660 20544
rect 3528 20454 3832 20482
rect 3514 20360 3570 20369
rect 3514 20295 3570 20304
rect 3424 19916 3476 19922
rect 3424 19858 3476 19864
rect 3436 19514 3464 19858
rect 3424 19508 3476 19514
rect 3424 19450 3476 19456
rect 3528 17785 3556 20295
rect 3700 20256 3752 20262
rect 3700 20198 3752 20204
rect 3608 19848 3660 19854
rect 3712 19836 3740 20198
rect 3660 19808 3740 19836
rect 3608 19790 3660 19796
rect 3712 19514 3740 19808
rect 3700 19508 3752 19514
rect 3700 19450 3752 19456
rect 3712 18290 3740 19450
rect 3804 18873 3832 20454
rect 3896 20398 3924 20946
rect 3884 20392 3936 20398
rect 3884 20334 3936 20340
rect 3790 18864 3846 18873
rect 3790 18799 3846 18808
rect 3804 18426 3832 18799
rect 3792 18420 3844 18426
rect 3792 18362 3844 18368
rect 3700 18284 3752 18290
rect 3700 18226 3752 18232
rect 3804 18222 3832 18362
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 3790 17912 3846 17921
rect 3790 17847 3846 17856
rect 3514 17776 3570 17785
rect 3514 17711 3570 17720
rect 3148 17672 3200 17678
rect 3146 17640 3148 17649
rect 3200 17640 3202 17649
rect 3146 17575 3202 17584
rect 3056 16652 3108 16658
rect 3056 16594 3108 16600
rect 3068 16250 3096 16594
rect 3056 16244 3108 16250
rect 3056 16186 3108 16192
rect 3148 16040 3200 16046
rect 3146 16008 3148 16017
rect 3200 16008 3202 16017
rect 3146 15943 3202 15952
rect 3804 15570 3832 17847
rect 3988 16250 4016 33390
rect 4080 31754 4108 42842
rect 4172 42362 4200 43710
rect 4289 43548 4585 43568
rect 4345 43546 4369 43548
rect 4425 43546 4449 43548
rect 4505 43546 4529 43548
rect 4367 43494 4369 43546
rect 4431 43494 4443 43546
rect 4505 43494 4507 43546
rect 4345 43492 4369 43494
rect 4425 43492 4449 43494
rect 4505 43492 4529 43494
rect 4289 43472 4585 43492
rect 4289 42460 4585 42480
rect 4345 42458 4369 42460
rect 4425 42458 4449 42460
rect 4505 42458 4529 42460
rect 4367 42406 4369 42458
rect 4431 42406 4443 42458
rect 4505 42406 4507 42458
rect 4345 42404 4369 42406
rect 4425 42404 4449 42406
rect 4505 42404 4529 42406
rect 4289 42384 4585 42404
rect 4160 42356 4212 42362
rect 4160 42298 4212 42304
rect 4172 41750 4200 42298
rect 4252 42016 4304 42022
rect 4252 41958 4304 41964
rect 4160 41744 4212 41750
rect 4160 41686 4212 41692
rect 4264 41596 4292 41958
rect 4172 41568 4292 41596
rect 4172 32910 4200 41568
rect 4289 41372 4585 41392
rect 4345 41370 4369 41372
rect 4425 41370 4449 41372
rect 4505 41370 4529 41372
rect 4367 41318 4369 41370
rect 4431 41318 4443 41370
rect 4505 41318 4507 41370
rect 4345 41316 4369 41318
rect 4425 41316 4449 41318
rect 4505 41316 4529 41318
rect 4289 41296 4585 41316
rect 4250 41168 4306 41177
rect 4250 41103 4306 41112
rect 4264 40594 4292 41103
rect 4632 41070 4660 50680
rect 4724 47462 4752 50782
rect 4712 47456 4764 47462
rect 4712 47398 4764 47404
rect 4710 47288 4766 47297
rect 4710 47223 4766 47232
rect 4724 46578 4752 47223
rect 4712 46572 4764 46578
rect 4712 46514 4764 46520
rect 4712 46436 4764 46442
rect 4712 46378 4764 46384
rect 4620 41064 4672 41070
rect 4620 41006 4672 41012
rect 4252 40588 4304 40594
rect 4252 40530 4304 40536
rect 4289 40284 4585 40304
rect 4345 40282 4369 40284
rect 4425 40282 4449 40284
rect 4505 40282 4529 40284
rect 4367 40230 4369 40282
rect 4431 40230 4443 40282
rect 4505 40230 4507 40282
rect 4345 40228 4369 40230
rect 4425 40228 4449 40230
rect 4505 40228 4529 40230
rect 4289 40208 4585 40228
rect 4620 39976 4672 39982
rect 4342 39944 4398 39953
rect 4620 39918 4672 39924
rect 4342 39879 4398 39888
rect 4436 39908 4488 39914
rect 4356 39846 4384 39879
rect 4436 39850 4488 39856
rect 4344 39840 4396 39846
rect 4344 39782 4396 39788
rect 4448 39642 4476 39850
rect 4632 39642 4660 39918
rect 4436 39636 4488 39642
rect 4436 39578 4488 39584
rect 4620 39636 4672 39642
rect 4620 39578 4672 39584
rect 4620 39500 4672 39506
rect 4620 39442 4672 39448
rect 4289 39196 4585 39216
rect 4345 39194 4369 39196
rect 4425 39194 4449 39196
rect 4505 39194 4529 39196
rect 4367 39142 4369 39194
rect 4431 39142 4443 39194
rect 4505 39142 4507 39194
rect 4345 39140 4369 39142
rect 4425 39140 4449 39142
rect 4505 39140 4529 39142
rect 4289 39120 4585 39140
rect 4632 38554 4660 39442
rect 4724 38962 4752 46378
rect 4712 38956 4764 38962
rect 4712 38898 4764 38904
rect 4620 38548 4672 38554
rect 4620 38490 4672 38496
rect 4289 38108 4585 38128
rect 4345 38106 4369 38108
rect 4425 38106 4449 38108
rect 4505 38106 4529 38108
rect 4367 38054 4369 38106
rect 4431 38054 4443 38106
rect 4505 38054 4507 38106
rect 4345 38052 4369 38054
rect 4425 38052 4449 38054
rect 4505 38052 4529 38054
rect 4289 38032 4585 38052
rect 4289 37020 4585 37040
rect 4345 37018 4369 37020
rect 4425 37018 4449 37020
rect 4505 37018 4529 37020
rect 4367 36966 4369 37018
rect 4431 36966 4443 37018
rect 4505 36966 4507 37018
rect 4345 36964 4369 36966
rect 4425 36964 4449 36966
rect 4505 36964 4529 36966
rect 4289 36944 4585 36964
rect 4289 35932 4585 35952
rect 4345 35930 4369 35932
rect 4425 35930 4449 35932
rect 4505 35930 4529 35932
rect 4367 35878 4369 35930
rect 4431 35878 4443 35930
rect 4505 35878 4507 35930
rect 4345 35876 4369 35878
rect 4425 35876 4449 35878
rect 4505 35876 4529 35878
rect 4289 35856 4585 35876
rect 4816 35714 4844 51750
rect 4894 51096 4950 51105
rect 4894 51031 4950 51040
rect 4908 50522 4936 51031
rect 4896 50516 4948 50522
rect 4896 50458 4948 50464
rect 5000 49858 5028 51870
rect 5080 51876 5132 51882
rect 5080 51818 5132 51824
rect 5184 51474 5212 52119
rect 5276 51814 5304 60794
rect 5368 60636 5396 60982
rect 5552 60858 5580 61662
rect 5540 60852 5592 60858
rect 5540 60794 5592 60800
rect 5368 60608 5488 60636
rect 5354 60480 5410 60489
rect 5354 60415 5410 60424
rect 5264 51808 5316 51814
rect 5264 51750 5316 51756
rect 5262 51640 5318 51649
rect 5262 51575 5318 51584
rect 5172 51468 5224 51474
rect 5172 51410 5224 51416
rect 5080 51332 5132 51338
rect 5080 51274 5132 51280
rect 4908 49830 5028 49858
rect 4908 48686 4936 49830
rect 4988 49768 5040 49774
rect 4988 49710 5040 49716
rect 4896 48680 4948 48686
rect 4896 48622 4948 48628
rect 4908 48006 4936 48622
rect 4896 48000 4948 48006
rect 4896 47942 4948 47948
rect 4896 47456 4948 47462
rect 4896 47398 4948 47404
rect 4908 43382 4936 47398
rect 5000 47161 5028 49710
rect 5092 48890 5120 51274
rect 5184 51066 5212 51410
rect 5172 51060 5224 51066
rect 5172 51002 5224 51008
rect 5172 50856 5224 50862
rect 5172 50798 5224 50804
rect 5184 50522 5212 50798
rect 5172 50516 5224 50522
rect 5172 50458 5224 50464
rect 5184 49910 5212 50458
rect 5172 49904 5224 49910
rect 5172 49846 5224 49852
rect 5172 49768 5224 49774
rect 5172 49710 5224 49716
rect 5184 49094 5212 49710
rect 5172 49088 5224 49094
rect 5172 49030 5224 49036
rect 5080 48884 5132 48890
rect 5080 48826 5132 48832
rect 5184 48754 5212 49030
rect 5080 48748 5132 48754
rect 5080 48690 5132 48696
rect 5172 48748 5224 48754
rect 5172 48690 5224 48696
rect 4986 47152 5042 47161
rect 4986 47087 5042 47096
rect 5092 46968 5120 48690
rect 5172 48204 5224 48210
rect 5172 48146 5224 48152
rect 5184 47802 5212 48146
rect 5172 47796 5224 47802
rect 5172 47738 5224 47744
rect 5172 47456 5224 47462
rect 5172 47398 5224 47404
rect 5000 46940 5120 46968
rect 5000 43926 5028 46940
rect 5078 46880 5134 46889
rect 5078 46815 5134 46824
rect 4988 43920 5040 43926
rect 4988 43862 5040 43868
rect 4988 43784 5040 43790
rect 4988 43726 5040 43732
rect 4896 43376 4948 43382
rect 4896 43318 4948 43324
rect 4896 43240 4948 43246
rect 4896 43182 4948 43188
rect 4908 42770 4936 43182
rect 5000 42906 5028 43726
rect 4988 42900 5040 42906
rect 4988 42842 5040 42848
rect 4896 42764 4948 42770
rect 4896 42706 4948 42712
rect 4908 42294 4936 42706
rect 4896 42288 4948 42294
rect 4896 42230 4948 42236
rect 5092 41970 5120 46815
rect 5184 46578 5212 47398
rect 5172 46572 5224 46578
rect 5172 46514 5224 46520
rect 5276 46442 5304 51575
rect 5368 49065 5396 60415
rect 5460 59265 5488 60608
rect 5644 59770 5672 62766
rect 5736 60738 5764 70450
rect 5828 69562 5856 72422
rect 5908 72004 5960 72010
rect 5908 71946 5960 71952
rect 5920 70446 5948 71946
rect 5908 70440 5960 70446
rect 5908 70382 5960 70388
rect 5920 69766 5948 70382
rect 5908 69760 5960 69766
rect 5908 69702 5960 69708
rect 5816 69556 5868 69562
rect 5816 69498 5868 69504
rect 5814 69456 5870 69465
rect 5814 69391 5816 69400
rect 5868 69391 5870 69400
rect 5816 69362 5868 69368
rect 6012 69018 6040 73086
rect 6104 72690 6132 73714
rect 6184 73296 6236 73302
rect 6184 73238 6236 73244
rect 6092 72684 6144 72690
rect 6092 72626 6144 72632
rect 6104 72282 6132 72626
rect 6196 72486 6224 73238
rect 6472 73030 6500 74122
rect 6552 74112 6604 74118
rect 6552 74054 6604 74060
rect 6564 73778 6592 74054
rect 6552 73772 6604 73778
rect 6552 73714 6604 73720
rect 6460 73024 6512 73030
rect 6460 72966 6512 72972
rect 6472 72622 6500 72966
rect 6460 72616 6512 72622
rect 6460 72558 6512 72564
rect 6184 72480 6236 72486
rect 6184 72422 6236 72428
rect 6092 72276 6144 72282
rect 6092 72218 6144 72224
rect 6104 71602 6132 72218
rect 6092 71596 6144 71602
rect 6092 71538 6144 71544
rect 6196 70292 6224 72422
rect 6564 72146 6592 73714
rect 6748 73166 6776 74734
rect 7116 74186 7144 75346
rect 7288 75200 7340 75206
rect 7288 75142 7340 75148
rect 7104 74180 7156 74186
rect 7104 74122 7156 74128
rect 7196 73704 7248 73710
rect 7010 73672 7066 73681
rect 7196 73646 7248 73652
rect 7010 73607 7066 73616
rect 6918 73264 6974 73273
rect 6918 73199 6974 73208
rect 6736 73160 6788 73166
rect 6736 73102 6788 73108
rect 6552 72140 6604 72146
rect 6552 72082 6604 72088
rect 6748 72010 6776 73102
rect 6932 73098 6960 73199
rect 6920 73092 6972 73098
rect 6920 73034 6972 73040
rect 7024 72826 7052 73607
rect 7012 72820 7064 72826
rect 7012 72762 7064 72768
rect 7102 72176 7158 72185
rect 6828 72140 6880 72146
rect 7102 72111 7104 72120
rect 6828 72082 6880 72088
rect 7156 72111 7158 72120
rect 7104 72082 7156 72088
rect 6736 72004 6788 72010
rect 6736 71946 6788 71952
rect 6840 71738 6868 72082
rect 7208 72010 7236 73646
rect 7300 73302 7328 75142
rect 10956 75100 11252 75120
rect 11012 75098 11036 75100
rect 11092 75098 11116 75100
rect 11172 75098 11196 75100
rect 11034 75046 11036 75098
rect 11098 75046 11110 75098
rect 11172 75046 11174 75098
rect 11012 75044 11036 75046
rect 11092 75044 11116 75046
rect 11172 75044 11196 75046
rect 10956 75024 11252 75044
rect 17622 75100 17918 75120
rect 17678 75098 17702 75100
rect 17758 75098 17782 75100
rect 17838 75098 17862 75100
rect 17700 75046 17702 75098
rect 17764 75046 17776 75098
rect 17838 75046 17840 75098
rect 17678 75044 17702 75046
rect 17758 75044 17782 75046
rect 17838 75044 17862 75046
rect 17622 75024 17918 75044
rect 7380 74724 7432 74730
rect 7380 74666 7432 74672
rect 7392 74390 7420 74666
rect 7622 74556 7918 74576
rect 7678 74554 7702 74556
rect 7758 74554 7782 74556
rect 7838 74554 7862 74556
rect 7700 74502 7702 74554
rect 7764 74502 7776 74554
rect 7838 74502 7840 74554
rect 7678 74500 7702 74502
rect 7758 74500 7782 74502
rect 7838 74500 7862 74502
rect 7622 74480 7918 74500
rect 14289 74556 14585 74576
rect 14345 74554 14369 74556
rect 14425 74554 14449 74556
rect 14505 74554 14529 74556
rect 14367 74502 14369 74554
rect 14431 74502 14443 74554
rect 14505 74502 14507 74554
rect 14345 74500 14369 74502
rect 14425 74500 14449 74502
rect 14505 74500 14529 74502
rect 14289 74480 14585 74500
rect 7380 74384 7432 74390
rect 7380 74326 7432 74332
rect 8300 74384 8352 74390
rect 8300 74326 8352 74332
rect 7748 74316 7800 74322
rect 7748 74258 7800 74264
rect 7760 73642 7788 74258
rect 7380 73636 7432 73642
rect 7380 73578 7432 73584
rect 7748 73636 7800 73642
rect 7748 73578 7800 73584
rect 7288 73296 7340 73302
rect 7288 73238 7340 73244
rect 7392 73148 7420 73578
rect 7622 73468 7918 73488
rect 7678 73466 7702 73468
rect 7758 73466 7782 73468
rect 7838 73466 7862 73468
rect 7700 73414 7702 73466
rect 7764 73414 7776 73466
rect 7838 73414 7840 73466
rect 7678 73412 7702 73414
rect 7758 73412 7782 73414
rect 7838 73412 7862 73414
rect 7622 73392 7918 73412
rect 7300 73120 7420 73148
rect 7196 72004 7248 72010
rect 7196 71946 7248 71952
rect 6828 71732 6880 71738
rect 6828 71674 6880 71680
rect 6552 71596 6604 71602
rect 6552 71538 6604 71544
rect 6196 70264 6316 70292
rect 6000 69012 6052 69018
rect 6000 68954 6052 68960
rect 6092 68672 6144 68678
rect 6092 68614 6144 68620
rect 5908 67176 5960 67182
rect 5908 67118 5960 67124
rect 5920 66638 5948 67118
rect 5908 66632 5960 66638
rect 5908 66574 5960 66580
rect 6000 66564 6052 66570
rect 6000 66506 6052 66512
rect 5816 65068 5868 65074
rect 5816 65010 5868 65016
rect 5828 64326 5856 65010
rect 5816 64320 5868 64326
rect 5816 64262 5868 64268
rect 5828 62830 5856 64262
rect 5816 62824 5868 62830
rect 5816 62766 5868 62772
rect 5736 60710 5948 60738
rect 5632 59764 5684 59770
rect 5632 59706 5684 59712
rect 5816 59560 5868 59566
rect 5816 59502 5868 59508
rect 5446 59256 5502 59265
rect 5446 59191 5502 59200
rect 5448 59152 5500 59158
rect 5448 59094 5500 59100
rect 5460 57594 5488 59094
rect 5724 59084 5776 59090
rect 5724 59026 5776 59032
rect 5538 58168 5594 58177
rect 5538 58103 5594 58112
rect 5448 57588 5500 57594
rect 5448 57530 5500 57536
rect 5448 57248 5500 57254
rect 5448 57190 5500 57196
rect 5460 51474 5488 57190
rect 5552 55350 5580 58103
rect 5736 58070 5764 59026
rect 5724 58064 5776 58070
rect 5724 58006 5776 58012
rect 5630 57352 5686 57361
rect 5630 57287 5686 57296
rect 5644 56506 5672 57287
rect 5724 57248 5776 57254
rect 5724 57190 5776 57196
rect 5736 56710 5764 57190
rect 5724 56704 5776 56710
rect 5724 56646 5776 56652
rect 5632 56500 5684 56506
rect 5632 56442 5684 56448
rect 5828 56386 5856 59502
rect 5644 56358 5856 56386
rect 5540 55344 5592 55350
rect 5540 55286 5592 55292
rect 5540 55140 5592 55146
rect 5540 55082 5592 55088
rect 5552 54738 5580 55082
rect 5540 54732 5592 54738
rect 5540 54674 5592 54680
rect 5552 54330 5580 54674
rect 5540 54324 5592 54330
rect 5540 54266 5592 54272
rect 5552 53718 5580 54266
rect 5540 53712 5592 53718
rect 5540 53654 5592 53660
rect 5540 53576 5592 53582
rect 5540 53518 5592 53524
rect 5552 52902 5580 53518
rect 5644 53009 5672 56358
rect 5724 55616 5776 55622
rect 5724 55558 5776 55564
rect 5736 55282 5764 55558
rect 5724 55276 5776 55282
rect 5724 55218 5776 55224
rect 5724 55140 5776 55146
rect 5724 55082 5776 55088
rect 5736 54534 5764 55082
rect 5816 54596 5868 54602
rect 5816 54538 5868 54544
rect 5724 54528 5776 54534
rect 5724 54470 5776 54476
rect 5630 53000 5686 53009
rect 5630 52935 5686 52944
rect 5540 52896 5592 52902
rect 5540 52838 5592 52844
rect 5632 52896 5684 52902
rect 5632 52838 5684 52844
rect 5540 52692 5592 52698
rect 5540 52634 5592 52640
rect 5552 52018 5580 52634
rect 5540 52012 5592 52018
rect 5540 51954 5592 51960
rect 5538 51776 5594 51785
rect 5538 51711 5594 51720
rect 5448 51468 5500 51474
rect 5448 51410 5500 51416
rect 5552 51354 5580 51711
rect 5460 51338 5580 51354
rect 5448 51332 5580 51338
rect 5500 51326 5580 51332
rect 5448 51274 5500 51280
rect 5540 51264 5592 51270
rect 5446 51232 5502 51241
rect 5540 51206 5592 51212
rect 5446 51167 5502 51176
rect 5354 49056 5410 49065
rect 5354 48991 5410 49000
rect 5356 48680 5408 48686
rect 5356 48622 5408 48628
rect 5368 48142 5396 48622
rect 5356 48136 5408 48142
rect 5356 48078 5408 48084
rect 5356 48000 5408 48006
rect 5356 47942 5408 47948
rect 5264 46436 5316 46442
rect 5264 46378 5316 46384
rect 5172 46368 5224 46374
rect 5172 46310 5224 46316
rect 5184 42401 5212 46310
rect 5264 44872 5316 44878
rect 5264 44814 5316 44820
rect 5276 44334 5304 44814
rect 5264 44328 5316 44334
rect 5264 44270 5316 44276
rect 5262 43888 5318 43897
rect 5262 43823 5318 43832
rect 5170 42392 5226 42401
rect 5170 42327 5226 42336
rect 5170 42256 5226 42265
rect 5170 42191 5226 42200
rect 5184 42158 5212 42191
rect 5172 42152 5224 42158
rect 5172 42094 5224 42100
rect 5000 41942 5120 41970
rect 5000 41834 5028 41942
rect 4908 41806 5028 41834
rect 5078 41848 5134 41857
rect 4908 40118 4936 41806
rect 5184 41818 5212 42094
rect 5276 42022 5304 43823
rect 5264 42016 5316 42022
rect 5264 41958 5316 41964
rect 5078 41783 5134 41792
rect 5172 41812 5224 41818
rect 4988 41744 5040 41750
rect 4988 41686 5040 41692
rect 5092 41698 5120 41783
rect 5172 41754 5224 41760
rect 5000 40730 5028 41686
rect 5092 41670 5212 41698
rect 5080 41064 5132 41070
rect 5080 41006 5132 41012
rect 4988 40724 5040 40730
rect 4988 40666 5040 40672
rect 5092 40610 5120 41006
rect 5000 40582 5120 40610
rect 4896 40112 4948 40118
rect 4896 40054 4948 40060
rect 4896 39908 4948 39914
rect 4896 39850 4948 39856
rect 4908 36922 4936 39850
rect 4896 36916 4948 36922
rect 4896 36858 4948 36864
rect 4908 36582 4936 36858
rect 4896 36576 4948 36582
rect 4896 36518 4948 36524
rect 4908 36310 4936 36518
rect 4896 36304 4948 36310
rect 4896 36246 4948 36252
rect 4724 35686 4844 35714
rect 4620 35012 4672 35018
rect 4620 34954 4672 34960
rect 4289 34844 4585 34864
rect 4345 34842 4369 34844
rect 4425 34842 4449 34844
rect 4505 34842 4529 34844
rect 4367 34790 4369 34842
rect 4431 34790 4443 34842
rect 4505 34790 4507 34842
rect 4345 34788 4369 34790
rect 4425 34788 4449 34790
rect 4505 34788 4529 34790
rect 4289 34768 4585 34788
rect 4632 34610 4660 34954
rect 4620 34604 4672 34610
rect 4620 34546 4672 34552
rect 4289 33756 4585 33776
rect 4345 33754 4369 33756
rect 4425 33754 4449 33756
rect 4505 33754 4529 33756
rect 4367 33702 4369 33754
rect 4431 33702 4443 33754
rect 4505 33702 4507 33754
rect 4345 33700 4369 33702
rect 4425 33700 4449 33702
rect 4505 33700 4529 33702
rect 4289 33680 4585 33700
rect 4724 32978 4752 35686
rect 5000 34610 5028 40582
rect 5080 38888 5132 38894
rect 5080 38830 5132 38836
rect 5092 38214 5120 38830
rect 5080 38208 5132 38214
rect 5080 38150 5132 38156
rect 5092 37466 5120 38150
rect 5080 37460 5132 37466
rect 5080 37402 5132 37408
rect 5080 34944 5132 34950
rect 5080 34886 5132 34892
rect 4988 34604 5040 34610
rect 4988 34546 5040 34552
rect 5092 34542 5120 34886
rect 5080 34536 5132 34542
rect 5080 34478 5132 34484
rect 4896 33992 4948 33998
rect 4894 33960 4896 33969
rect 4948 33960 4950 33969
rect 4894 33895 4950 33904
rect 4712 32972 4764 32978
rect 4712 32914 4764 32920
rect 4160 32904 4212 32910
rect 4160 32846 4212 32852
rect 4289 32668 4585 32688
rect 4345 32666 4369 32668
rect 4425 32666 4449 32668
rect 4505 32666 4529 32668
rect 4367 32614 4369 32666
rect 4431 32614 4443 32666
rect 4505 32614 4507 32666
rect 4345 32612 4369 32614
rect 4425 32612 4449 32614
rect 4505 32612 4529 32614
rect 4289 32592 4585 32612
rect 5092 32570 5120 34478
rect 5080 32564 5132 32570
rect 5080 32506 5132 32512
rect 4988 32360 5040 32366
rect 4988 32302 5040 32308
rect 5000 31890 5028 32302
rect 4988 31884 5040 31890
rect 4988 31826 5040 31832
rect 4068 31748 4120 31754
rect 4068 31690 4120 31696
rect 4289 31580 4585 31600
rect 4345 31578 4369 31580
rect 4425 31578 4449 31580
rect 4505 31578 4529 31580
rect 4367 31526 4369 31578
rect 4431 31526 4443 31578
rect 4505 31526 4507 31578
rect 4345 31524 4369 31526
rect 4425 31524 4449 31526
rect 4505 31524 4529 31526
rect 4289 31504 4585 31524
rect 4066 30832 4122 30841
rect 4066 30767 4122 30776
rect 4080 27441 4108 30767
rect 4988 30728 5040 30734
rect 4988 30670 5040 30676
rect 5000 30569 5028 30670
rect 4986 30560 5042 30569
rect 4289 30492 4585 30512
rect 4986 30495 5042 30504
rect 4345 30490 4369 30492
rect 4425 30490 4449 30492
rect 4505 30490 4529 30492
rect 4367 30438 4369 30490
rect 4431 30438 4443 30490
rect 4505 30438 4507 30490
rect 4345 30436 4369 30438
rect 4425 30436 4449 30438
rect 4505 30436 4529 30438
rect 4289 30416 4585 30436
rect 5000 30394 5028 30495
rect 4988 30388 5040 30394
rect 4988 30330 5040 30336
rect 4436 30252 4488 30258
rect 4436 30194 4488 30200
rect 4448 29782 4476 30194
rect 4896 30184 4948 30190
rect 4896 30126 4948 30132
rect 4526 30016 4582 30025
rect 4526 29951 4582 29960
rect 4540 29850 4568 29951
rect 4528 29844 4580 29850
rect 4528 29786 4580 29792
rect 4436 29776 4488 29782
rect 4436 29718 4488 29724
rect 4712 29708 4764 29714
rect 4712 29650 4764 29656
rect 4289 29404 4585 29424
rect 4345 29402 4369 29404
rect 4425 29402 4449 29404
rect 4505 29402 4529 29404
rect 4367 29350 4369 29402
rect 4431 29350 4443 29402
rect 4505 29350 4507 29402
rect 4345 29348 4369 29350
rect 4425 29348 4449 29350
rect 4505 29348 4529 29350
rect 4289 29328 4585 29348
rect 4724 28626 4752 29650
rect 4908 29034 4936 30126
rect 4896 29028 4948 29034
rect 4896 28970 4948 28976
rect 4712 28620 4764 28626
rect 4712 28562 4764 28568
rect 4289 28316 4585 28336
rect 4345 28314 4369 28316
rect 4425 28314 4449 28316
rect 4505 28314 4529 28316
rect 4367 28262 4369 28314
rect 4431 28262 4443 28314
rect 4505 28262 4507 28314
rect 4345 28260 4369 28262
rect 4425 28260 4449 28262
rect 4505 28260 4529 28262
rect 4289 28240 4585 28260
rect 4712 28008 4764 28014
rect 4712 27950 4764 27956
rect 4344 27872 4396 27878
rect 4344 27814 4396 27820
rect 4356 27606 4384 27814
rect 4160 27600 4212 27606
rect 4160 27542 4212 27548
rect 4344 27600 4396 27606
rect 4344 27542 4396 27548
rect 4066 27432 4122 27441
rect 4066 27367 4122 27376
rect 4172 26926 4200 27542
rect 4724 27538 4752 27950
rect 5184 27606 5212 41670
rect 5264 41676 5316 41682
rect 5264 41618 5316 41624
rect 5276 40662 5304 41618
rect 5264 40656 5316 40662
rect 5264 40598 5316 40604
rect 5264 40520 5316 40526
rect 5264 40462 5316 40468
rect 5276 39642 5304 40462
rect 5264 39636 5316 39642
rect 5264 39578 5316 39584
rect 5368 39506 5396 47942
rect 5356 39500 5408 39506
rect 5356 39442 5408 39448
rect 5368 39098 5396 39442
rect 5356 39092 5408 39098
rect 5356 39034 5408 39040
rect 5356 38412 5408 38418
rect 5356 38354 5408 38360
rect 5262 37360 5318 37369
rect 5262 37295 5318 37304
rect 5276 36718 5304 37295
rect 5264 36712 5316 36718
rect 5264 36654 5316 36660
rect 5276 36378 5304 36654
rect 5264 36372 5316 36378
rect 5264 36314 5316 36320
rect 5368 36242 5396 38354
rect 5356 36236 5408 36242
rect 5356 36178 5408 36184
rect 5368 35834 5396 36178
rect 5356 35828 5408 35834
rect 5356 35770 5408 35776
rect 5460 34610 5488 51167
rect 5552 50998 5580 51206
rect 5540 50992 5592 50998
rect 5540 50934 5592 50940
rect 5552 50522 5580 50934
rect 5644 50862 5672 52838
rect 5736 51066 5764 54470
rect 5828 53650 5856 54538
rect 5816 53644 5868 53650
rect 5816 53586 5868 53592
rect 5724 51060 5776 51066
rect 5724 51002 5776 51008
rect 5722 50960 5778 50969
rect 5828 50930 5856 53586
rect 5722 50895 5778 50904
rect 5816 50924 5868 50930
rect 5632 50856 5684 50862
rect 5632 50798 5684 50804
rect 5632 50720 5684 50726
rect 5632 50662 5684 50668
rect 5540 50516 5592 50522
rect 5540 50458 5592 50464
rect 5538 49192 5594 49201
rect 5538 49127 5540 49136
rect 5592 49127 5594 49136
rect 5540 49098 5592 49104
rect 5538 49056 5594 49065
rect 5538 48991 5594 49000
rect 5552 46986 5580 48991
rect 5644 48929 5672 50662
rect 5630 48920 5686 48929
rect 5630 48855 5686 48864
rect 5632 47116 5684 47122
rect 5632 47058 5684 47064
rect 5540 46980 5592 46986
rect 5540 46922 5592 46928
rect 5644 46714 5672 47058
rect 5632 46708 5684 46714
rect 5632 46650 5684 46656
rect 5540 46640 5592 46646
rect 5540 46582 5592 46588
rect 5552 44316 5580 46582
rect 5644 46510 5672 46541
rect 5632 46504 5684 46510
rect 5630 46472 5632 46481
rect 5684 46472 5686 46481
rect 5630 46407 5686 46416
rect 5644 46170 5672 46407
rect 5632 46164 5684 46170
rect 5632 46106 5684 46112
rect 5632 45824 5684 45830
rect 5632 45766 5684 45772
rect 5644 45626 5672 45766
rect 5632 45620 5684 45626
rect 5632 45562 5684 45568
rect 5632 45416 5684 45422
rect 5632 45358 5684 45364
rect 5644 44441 5672 45358
rect 5630 44432 5686 44441
rect 5630 44367 5686 44376
rect 5632 44328 5684 44334
rect 5552 44288 5632 44316
rect 5632 44270 5684 44276
rect 5540 43376 5592 43382
rect 5540 43318 5592 43324
rect 5552 41206 5580 43318
rect 5644 41546 5672 44270
rect 5736 41993 5764 50895
rect 5816 50866 5868 50872
rect 5814 50824 5870 50833
rect 5814 50759 5870 50768
rect 5828 49978 5856 50759
rect 5816 49972 5868 49978
rect 5816 49914 5868 49920
rect 5828 49774 5856 49914
rect 5816 49768 5868 49774
rect 5816 49710 5868 49716
rect 5814 48240 5870 48249
rect 5814 48175 5816 48184
rect 5868 48175 5870 48184
rect 5816 48146 5868 48152
rect 5816 47728 5868 47734
rect 5814 47696 5816 47705
rect 5868 47696 5870 47705
rect 5814 47631 5870 47640
rect 5816 47456 5868 47462
rect 5816 47398 5868 47404
rect 5828 46374 5856 47398
rect 5816 46368 5868 46374
rect 5816 46310 5868 46316
rect 5828 45286 5856 46310
rect 5816 45280 5868 45286
rect 5816 45222 5868 45228
rect 5828 43110 5856 45222
rect 5816 43104 5868 43110
rect 5816 43046 5868 43052
rect 5722 41984 5778 41993
rect 5722 41919 5778 41928
rect 5724 41744 5776 41750
rect 5724 41686 5776 41692
rect 5632 41540 5684 41546
rect 5632 41482 5684 41488
rect 5630 41440 5686 41449
rect 5630 41375 5686 41384
rect 5540 41200 5592 41206
rect 5644 41177 5672 41375
rect 5540 41142 5592 41148
rect 5630 41168 5686 41177
rect 5630 41103 5686 41112
rect 5632 41064 5684 41070
rect 5630 41032 5632 41041
rect 5684 41032 5686 41041
rect 5630 40967 5686 40976
rect 5538 40896 5594 40905
rect 5538 40831 5594 40840
rect 5552 38554 5580 40831
rect 5644 40458 5672 40967
rect 5632 40452 5684 40458
rect 5632 40394 5684 40400
rect 5736 39930 5764 41686
rect 5644 39902 5764 39930
rect 5644 39030 5672 39902
rect 5724 39840 5776 39846
rect 5724 39782 5776 39788
rect 5736 39098 5764 39782
rect 5724 39092 5776 39098
rect 5724 39034 5776 39040
rect 5632 39024 5684 39030
rect 5632 38966 5684 38972
rect 5540 38548 5592 38554
rect 5540 38490 5592 38496
rect 5540 37868 5592 37874
rect 5540 37810 5592 37816
rect 5552 36666 5580 37810
rect 5644 37210 5672 38966
rect 5644 37182 5764 37210
rect 5632 37120 5684 37126
rect 5632 37062 5684 37068
rect 5644 36854 5672 37062
rect 5632 36848 5684 36854
rect 5632 36790 5684 36796
rect 5552 36638 5672 36666
rect 5540 36576 5592 36582
rect 5540 36518 5592 36524
rect 5448 34604 5500 34610
rect 5448 34546 5500 34552
rect 5356 32904 5408 32910
rect 5356 32846 5408 32852
rect 5368 32366 5396 32846
rect 5356 32360 5408 32366
rect 5356 32302 5408 32308
rect 5368 32026 5396 32302
rect 5356 32020 5408 32026
rect 5356 31962 5408 31968
rect 5368 30190 5396 31962
rect 5356 30184 5408 30190
rect 5356 30126 5408 30132
rect 5448 30184 5500 30190
rect 5448 30126 5500 30132
rect 5460 29209 5488 30126
rect 5446 29200 5502 29209
rect 5446 29135 5502 29144
rect 5264 28620 5316 28626
rect 5264 28562 5316 28568
rect 5276 27878 5304 28562
rect 5264 27872 5316 27878
rect 5264 27814 5316 27820
rect 5172 27600 5224 27606
rect 5172 27542 5224 27548
rect 4712 27532 4764 27538
rect 4712 27474 4764 27480
rect 4289 27228 4585 27248
rect 4345 27226 4369 27228
rect 4425 27226 4449 27228
rect 4505 27226 4529 27228
rect 4367 27174 4369 27226
rect 4431 27174 4443 27226
rect 4505 27174 4507 27226
rect 4345 27172 4369 27174
rect 4425 27172 4449 27174
rect 4505 27172 4529 27174
rect 4289 27152 4585 27172
rect 4724 27130 4752 27474
rect 4712 27124 4764 27130
rect 4712 27066 4764 27072
rect 4160 26920 4212 26926
rect 4160 26862 4212 26868
rect 4620 26580 4672 26586
rect 4620 26522 4672 26528
rect 4160 26240 4212 26246
rect 4160 26182 4212 26188
rect 4172 26042 4200 26182
rect 4289 26140 4585 26160
rect 4345 26138 4369 26140
rect 4425 26138 4449 26140
rect 4505 26138 4529 26140
rect 4367 26086 4369 26138
rect 4431 26086 4443 26138
rect 4505 26086 4507 26138
rect 4345 26084 4369 26086
rect 4425 26084 4449 26086
rect 4505 26084 4529 26086
rect 4289 26064 4585 26084
rect 4160 26036 4212 26042
rect 4160 25978 4212 25984
rect 4632 25362 4660 26522
rect 4724 25974 4752 27066
rect 4988 26920 5040 26926
rect 4988 26862 5040 26868
rect 4712 25968 4764 25974
rect 4712 25910 4764 25916
rect 4620 25356 4672 25362
rect 4620 25298 4672 25304
rect 4158 25256 4214 25265
rect 4158 25191 4214 25200
rect 4068 24064 4120 24070
rect 4068 24006 4120 24012
rect 4080 23225 4108 24006
rect 4066 23216 4122 23225
rect 4066 23151 4122 23160
rect 4172 23118 4200 25191
rect 4620 25152 4672 25158
rect 4620 25094 4672 25100
rect 4289 25052 4585 25072
rect 4345 25050 4369 25052
rect 4425 25050 4449 25052
rect 4505 25050 4529 25052
rect 4367 24998 4369 25050
rect 4431 24998 4443 25050
rect 4505 24998 4507 25050
rect 4345 24996 4369 24998
rect 4425 24996 4449 24998
rect 4505 24996 4529 24998
rect 4289 24976 4585 24996
rect 4632 24750 4660 25094
rect 4620 24744 4672 24750
rect 4620 24686 4672 24692
rect 5000 24410 5028 26862
rect 5170 26616 5226 26625
rect 5170 26551 5226 26560
rect 5184 26518 5212 26551
rect 5172 26512 5224 26518
rect 5172 26454 5224 26460
rect 5170 24440 5226 24449
rect 4988 24404 5040 24410
rect 5170 24375 5226 24384
rect 4988 24346 5040 24352
rect 4289 23964 4585 23984
rect 4345 23962 4369 23964
rect 4425 23962 4449 23964
rect 4505 23962 4529 23964
rect 4367 23910 4369 23962
rect 4431 23910 4443 23962
rect 4505 23910 4507 23962
rect 4345 23908 4369 23910
rect 4425 23908 4449 23910
rect 4505 23908 4529 23910
rect 4289 23888 4585 23908
rect 4712 23180 4764 23186
rect 4712 23122 4764 23128
rect 4160 23112 4212 23118
rect 4160 23054 4212 23060
rect 4172 22794 4200 23054
rect 4724 22953 4752 23122
rect 4710 22944 4766 22953
rect 4289 22876 4585 22896
rect 4710 22879 4766 22888
rect 4345 22874 4369 22876
rect 4425 22874 4449 22876
rect 4505 22874 4529 22876
rect 4367 22822 4369 22874
rect 4431 22822 4443 22874
rect 4505 22822 4507 22874
rect 4345 22820 4369 22822
rect 4425 22820 4449 22822
rect 4505 22820 4529 22822
rect 4289 22800 4585 22820
rect 4080 22778 4200 22794
rect 4068 22772 4200 22778
rect 4120 22766 4200 22772
rect 4068 22714 4120 22720
rect 4724 22234 4752 22879
rect 5000 22574 5028 24346
rect 5080 24064 5132 24070
rect 5080 24006 5132 24012
rect 5092 23526 5120 24006
rect 5184 23594 5212 24375
rect 5172 23588 5224 23594
rect 5172 23530 5224 23536
rect 5080 23520 5132 23526
rect 5078 23488 5080 23497
rect 5132 23488 5134 23497
rect 5078 23423 5134 23432
rect 5276 23254 5304 27814
rect 5552 24410 5580 36518
rect 5644 33658 5672 36638
rect 5736 35494 5764 37182
rect 5828 36582 5856 43046
rect 5920 36854 5948 60710
rect 6012 59566 6040 66506
rect 6104 65414 6132 68614
rect 6184 67584 6236 67590
rect 6184 67526 6236 67532
rect 6196 67182 6224 67526
rect 6184 67176 6236 67182
rect 6184 67118 6236 67124
rect 6092 65408 6144 65414
rect 6092 65350 6144 65356
rect 6104 65210 6132 65350
rect 6092 65204 6144 65210
rect 6092 65146 6144 65152
rect 6288 64104 6316 70264
rect 6564 69902 6592 71538
rect 7194 71360 7250 71369
rect 7194 71295 7250 71304
rect 6736 71052 6788 71058
rect 6736 70994 6788 71000
rect 6748 70106 6776 70994
rect 6828 70984 6880 70990
rect 6828 70926 6880 70932
rect 6840 70446 6868 70926
rect 6828 70440 6880 70446
rect 6828 70382 6880 70388
rect 6736 70100 6788 70106
rect 6736 70042 6788 70048
rect 6552 69896 6604 69902
rect 6552 69838 6604 69844
rect 6368 69352 6420 69358
rect 6368 69294 6420 69300
rect 6380 68746 6408 69294
rect 6368 68740 6420 68746
rect 6368 68682 6420 68688
rect 6564 68678 6592 69838
rect 6736 69488 6788 69494
rect 6642 69456 6698 69465
rect 6736 69430 6788 69436
rect 6642 69391 6698 69400
rect 6656 69358 6684 69391
rect 6644 69352 6696 69358
rect 6644 69294 6696 69300
rect 6656 69018 6684 69294
rect 6644 69012 6696 69018
rect 6644 68954 6696 68960
rect 6552 68672 6604 68678
rect 6552 68614 6604 68620
rect 6748 68474 6776 69430
rect 7208 69358 7236 71295
rect 7196 69352 7248 69358
rect 7196 69294 7248 69300
rect 7102 69048 7158 69057
rect 7102 68983 7158 68992
rect 7012 68808 7064 68814
rect 7012 68750 7064 68756
rect 6920 68740 6972 68746
rect 6920 68682 6972 68688
rect 6736 68468 6788 68474
rect 6736 68410 6788 68416
rect 6748 67386 6776 68410
rect 6932 67386 6960 68682
rect 6736 67380 6788 67386
rect 6736 67322 6788 67328
rect 6920 67380 6972 67386
rect 6920 67322 6972 67328
rect 6828 67108 6880 67114
rect 6880 67068 6960 67096
rect 6828 67050 6880 67056
rect 6552 66700 6604 66706
rect 6552 66642 6604 66648
rect 6736 66700 6788 66706
rect 6736 66642 6788 66648
rect 6368 64456 6420 64462
rect 6368 64398 6420 64404
rect 6380 64122 6408 64398
rect 6104 64076 6316 64104
rect 6368 64116 6420 64122
rect 6104 63986 6132 64076
rect 6368 64058 6420 64064
rect 6092 63980 6144 63986
rect 6092 63922 6144 63928
rect 6104 63578 6132 63922
rect 6092 63572 6144 63578
rect 6092 63514 6144 63520
rect 6368 63572 6420 63578
rect 6368 63514 6420 63520
rect 6090 63336 6146 63345
rect 6090 63271 6146 63280
rect 6000 59560 6052 59566
rect 6000 59502 6052 59508
rect 6000 58948 6052 58954
rect 6000 58890 6052 58896
rect 6012 58478 6040 58890
rect 6000 58472 6052 58478
rect 6000 58414 6052 58420
rect 6104 55876 6132 63271
rect 6274 60616 6330 60625
rect 6274 60551 6330 60560
rect 6182 60072 6238 60081
rect 6182 60007 6184 60016
rect 6236 60007 6238 60016
rect 6184 59978 6236 59984
rect 6288 59770 6316 60551
rect 6276 59764 6328 59770
rect 6276 59706 6328 59712
rect 6184 59696 6236 59702
rect 6184 59638 6236 59644
rect 6196 57934 6224 59638
rect 6288 59401 6316 59706
rect 6274 59392 6330 59401
rect 6274 59327 6330 59336
rect 6380 58478 6408 63514
rect 6564 62694 6592 66642
rect 6748 64852 6776 66642
rect 6828 66496 6880 66502
rect 6828 66438 6880 66444
rect 6840 66026 6868 66438
rect 6828 66020 6880 66026
rect 6828 65962 6880 65968
rect 6840 64920 6868 65962
rect 6932 65210 6960 67068
rect 6920 65204 6972 65210
rect 6920 65146 6972 65152
rect 6840 64892 6960 64920
rect 6748 64824 6868 64852
rect 6644 64660 6696 64666
rect 6644 64602 6696 64608
rect 6656 63578 6684 64602
rect 6644 63572 6696 63578
rect 6696 63532 6776 63560
rect 6644 63514 6696 63520
rect 6644 62824 6696 62830
rect 6644 62766 6696 62772
rect 6552 62688 6604 62694
rect 6552 62630 6604 62636
rect 6460 60172 6512 60178
rect 6460 60114 6512 60120
rect 6472 59634 6500 60114
rect 6460 59628 6512 59634
rect 6460 59570 6512 59576
rect 6368 58472 6420 58478
rect 6368 58414 6420 58420
rect 6276 58132 6328 58138
rect 6380 58120 6408 58414
rect 6472 58138 6500 59570
rect 6328 58092 6408 58120
rect 6460 58132 6512 58138
rect 6276 58074 6328 58080
rect 6460 58074 6512 58080
rect 6460 57996 6512 58002
rect 6460 57938 6512 57944
rect 6184 57928 6236 57934
rect 6184 57870 6236 57876
rect 6196 57050 6224 57870
rect 6276 57792 6328 57798
rect 6276 57734 6328 57740
rect 6184 57044 6236 57050
rect 6184 56986 6236 56992
rect 6184 56908 6236 56914
rect 6184 56850 6236 56856
rect 6196 56166 6224 56850
rect 6288 56846 6316 57734
rect 6368 57520 6420 57526
rect 6368 57462 6420 57468
rect 6276 56840 6328 56846
rect 6276 56782 6328 56788
rect 6380 56302 6408 57462
rect 6368 56296 6420 56302
rect 6368 56238 6420 56244
rect 6184 56160 6236 56166
rect 6184 56102 6236 56108
rect 6012 55848 6132 55876
rect 6012 50810 6040 55848
rect 6196 55808 6224 56102
rect 6276 55956 6328 55962
rect 6380 55944 6408 56238
rect 6472 55962 6500 57938
rect 6328 55916 6408 55944
rect 6460 55956 6512 55962
rect 6276 55898 6328 55904
rect 6460 55898 6512 55904
rect 6104 55780 6224 55808
rect 6104 55418 6132 55780
rect 6288 55729 6316 55898
rect 6274 55720 6330 55729
rect 6184 55684 6236 55690
rect 6274 55655 6330 55664
rect 6184 55626 6236 55632
rect 6092 55412 6144 55418
rect 6092 55354 6144 55360
rect 6104 55214 6132 55354
rect 6092 55208 6144 55214
rect 6092 55150 6144 55156
rect 6104 53530 6132 55150
rect 6196 54330 6224 55626
rect 6276 55616 6328 55622
rect 6276 55558 6328 55564
rect 6288 55214 6316 55558
rect 6276 55208 6328 55214
rect 6276 55150 6328 55156
rect 6184 54324 6236 54330
rect 6184 54266 6236 54272
rect 6184 54120 6236 54126
rect 6182 54088 6184 54097
rect 6236 54088 6238 54097
rect 6182 54023 6238 54032
rect 6184 53984 6236 53990
rect 6184 53926 6236 53932
rect 6196 53650 6224 53926
rect 6184 53644 6236 53650
rect 6184 53586 6236 53592
rect 6104 53502 6224 53530
rect 6092 53440 6144 53446
rect 6092 53382 6144 53388
rect 6104 52737 6132 53382
rect 6090 52728 6146 52737
rect 6090 52663 6146 52672
rect 6092 52352 6144 52358
rect 6092 52294 6144 52300
rect 6104 51950 6132 52294
rect 6196 52193 6224 53502
rect 6182 52184 6238 52193
rect 6182 52119 6238 52128
rect 6184 52080 6236 52086
rect 6184 52022 6236 52028
rect 6092 51944 6144 51950
rect 6092 51886 6144 51892
rect 6196 51610 6224 52022
rect 6184 51604 6236 51610
rect 6184 51546 6236 51552
rect 6288 51490 6316 55150
rect 6368 54528 6420 54534
rect 6368 54470 6420 54476
rect 6380 53961 6408 54470
rect 6472 54126 6500 55898
rect 6460 54120 6512 54126
rect 6460 54062 6512 54068
rect 6366 53952 6422 53961
rect 6366 53887 6422 53896
rect 6472 53786 6500 54062
rect 6460 53780 6512 53786
rect 6460 53722 6512 53728
rect 6564 53666 6592 62630
rect 6656 59809 6684 62766
rect 6642 59800 6698 59809
rect 6748 59770 6776 63532
rect 6840 62830 6868 64824
rect 6828 62824 6880 62830
rect 6828 62766 6880 62772
rect 6932 61946 6960 64892
rect 7024 63730 7052 68750
rect 7116 66706 7144 68983
rect 7196 67176 7248 67182
rect 7194 67144 7196 67153
rect 7248 67144 7250 67153
rect 7194 67079 7250 67088
rect 7104 66700 7156 66706
rect 7104 66642 7156 66648
rect 7300 66586 7328 73120
rect 8312 73098 8340 74326
rect 10600 74112 10652 74118
rect 10600 74054 10652 74060
rect 10612 73710 10640 74054
rect 10956 74012 11252 74032
rect 11012 74010 11036 74012
rect 11092 74010 11116 74012
rect 11172 74010 11196 74012
rect 11034 73958 11036 74010
rect 11098 73958 11110 74010
rect 11172 73958 11174 74010
rect 11012 73956 11036 73958
rect 11092 73956 11116 73958
rect 11172 73956 11196 73958
rect 10956 73936 11252 73956
rect 17622 74012 17918 74032
rect 17678 74010 17702 74012
rect 17758 74010 17782 74012
rect 17838 74010 17862 74012
rect 17700 73958 17702 74010
rect 17764 73958 17776 74010
rect 17838 73958 17840 74010
rect 17678 73956 17702 73958
rect 17758 73956 17782 73958
rect 17838 73956 17862 73958
rect 17622 73936 17918 73956
rect 10692 73772 10744 73778
rect 10692 73714 10744 73720
rect 9312 73704 9364 73710
rect 9312 73646 9364 73652
rect 10600 73704 10652 73710
rect 10600 73646 10652 73652
rect 8482 73400 8538 73409
rect 9324 73370 9352 73646
rect 8482 73335 8538 73344
rect 9312 73364 9364 73370
rect 8300 73092 8352 73098
rect 8300 73034 8352 73040
rect 8312 72826 8340 73034
rect 8300 72820 8352 72826
rect 8300 72762 8352 72768
rect 8024 72616 8076 72622
rect 8024 72558 8076 72564
rect 7622 72380 7918 72400
rect 7678 72378 7702 72380
rect 7758 72378 7782 72380
rect 7838 72378 7862 72380
rect 7700 72326 7702 72378
rect 7764 72326 7776 72378
rect 7838 72326 7840 72378
rect 7678 72324 7702 72326
rect 7758 72324 7782 72326
rect 7838 72324 7862 72326
rect 7622 72304 7918 72324
rect 7472 71392 7524 71398
rect 7472 71334 7524 71340
rect 7484 70417 7512 71334
rect 7622 71292 7918 71312
rect 7678 71290 7702 71292
rect 7758 71290 7782 71292
rect 7838 71290 7862 71292
rect 7700 71238 7702 71290
rect 7764 71238 7776 71290
rect 7838 71238 7840 71290
rect 7678 71236 7702 71238
rect 7758 71236 7782 71238
rect 7838 71236 7862 71238
rect 7622 71216 7918 71236
rect 7840 70508 7892 70514
rect 7840 70450 7892 70456
rect 7852 70417 7880 70450
rect 7470 70408 7526 70417
rect 7470 70343 7526 70352
rect 7838 70408 7894 70417
rect 7838 70343 7894 70352
rect 7484 70310 7512 70343
rect 8036 70310 8064 72558
rect 8116 72072 8168 72078
rect 8116 72014 8168 72020
rect 8128 71058 8156 72014
rect 8208 71936 8260 71942
rect 8208 71878 8260 71884
rect 8220 71534 8248 71878
rect 8208 71528 8260 71534
rect 8208 71470 8260 71476
rect 8392 71528 8444 71534
rect 8392 71470 8444 71476
rect 8116 71052 8168 71058
rect 8116 70994 8168 71000
rect 8404 70854 8432 71470
rect 8392 70848 8444 70854
rect 8392 70790 8444 70796
rect 8116 70508 8168 70514
rect 8116 70450 8168 70456
rect 7472 70304 7524 70310
rect 7472 70246 7524 70252
rect 8024 70304 8076 70310
rect 8024 70246 8076 70252
rect 7380 69964 7432 69970
rect 7380 69906 7432 69912
rect 7392 69222 7420 69906
rect 7484 69426 7512 70246
rect 7622 70204 7918 70224
rect 7678 70202 7702 70204
rect 7758 70202 7782 70204
rect 7838 70202 7862 70204
rect 7700 70150 7702 70202
rect 7764 70150 7776 70202
rect 7838 70150 7840 70202
rect 7678 70148 7702 70150
rect 7758 70148 7782 70150
rect 7838 70148 7862 70150
rect 7622 70128 7918 70148
rect 7472 69420 7524 69426
rect 7472 69362 7524 69368
rect 7380 69216 7432 69222
rect 7380 69158 7432 69164
rect 7392 68678 7420 69158
rect 7622 69116 7918 69136
rect 7678 69114 7702 69116
rect 7758 69114 7782 69116
rect 7838 69114 7862 69116
rect 7700 69062 7702 69114
rect 7764 69062 7776 69114
rect 7838 69062 7840 69114
rect 7678 69060 7702 69062
rect 7758 69060 7782 69062
rect 7838 69060 7862 69062
rect 7622 69040 7918 69060
rect 8022 68912 8078 68921
rect 7944 68856 8022 68864
rect 7944 68836 8024 68856
rect 7380 68672 7432 68678
rect 7380 68614 7432 68620
rect 7392 68270 7420 68614
rect 7944 68406 7972 68836
rect 8076 68847 8078 68856
rect 8024 68818 8076 68824
rect 8024 68740 8076 68746
rect 8024 68682 8076 68688
rect 7932 68400 7984 68406
rect 7932 68342 7984 68348
rect 7380 68264 7432 68270
rect 7380 68206 7432 68212
rect 7208 66558 7328 66586
rect 7208 64569 7236 66558
rect 7288 66496 7340 66502
rect 7288 66438 7340 66444
rect 7300 66094 7328 66438
rect 7288 66088 7340 66094
rect 7288 66030 7340 66036
rect 7194 64560 7250 64569
rect 7300 64530 7328 66030
rect 7194 64495 7250 64504
rect 7288 64524 7340 64530
rect 7288 64466 7340 64472
rect 7104 64388 7156 64394
rect 7104 64330 7156 64336
rect 7116 63918 7144 64330
rect 7104 63912 7156 63918
rect 7104 63854 7156 63860
rect 7196 63844 7248 63850
rect 7196 63786 7248 63792
rect 7024 63702 7144 63730
rect 7116 62121 7144 63702
rect 7208 63617 7236 63786
rect 7194 63608 7250 63617
rect 7194 63543 7250 63552
rect 7300 62694 7328 64466
rect 7288 62688 7340 62694
rect 7288 62630 7340 62636
rect 7194 62384 7250 62393
rect 7194 62319 7250 62328
rect 7102 62112 7158 62121
rect 7102 62047 7158 62056
rect 6920 61940 6972 61946
rect 6920 61882 6972 61888
rect 7104 61940 7156 61946
rect 7104 61882 7156 61888
rect 6642 59735 6698 59744
rect 6736 59764 6788 59770
rect 6736 59706 6788 59712
rect 6644 58880 6696 58886
rect 6644 58822 6696 58828
rect 6656 58585 6684 58822
rect 6642 58576 6698 58585
rect 6642 58511 6698 58520
rect 6748 58138 6776 59706
rect 6920 59628 6972 59634
rect 6920 59570 6972 59576
rect 6828 59084 6880 59090
rect 6932 59072 6960 59570
rect 6880 59044 6960 59072
rect 6828 59026 6880 59032
rect 6840 58546 7052 58562
rect 6828 58540 7052 58546
rect 6880 58534 7052 58540
rect 6828 58482 6880 58488
rect 6920 58404 6972 58410
rect 6920 58346 6972 58352
rect 6736 58132 6788 58138
rect 6736 58074 6788 58080
rect 6736 57860 6788 57866
rect 6736 57802 6788 57808
rect 6748 57458 6776 57802
rect 6736 57452 6788 57458
rect 6736 57394 6788 57400
rect 6644 57316 6696 57322
rect 6644 57258 6696 57264
rect 6380 53638 6592 53666
rect 6380 52902 6408 53638
rect 6656 53530 6684 57258
rect 6748 57202 6776 57394
rect 6828 57384 6880 57390
rect 6932 57372 6960 58346
rect 6880 57344 6960 57372
rect 6828 57326 6880 57332
rect 6748 57174 6960 57202
rect 6828 56976 6880 56982
rect 6828 56918 6880 56924
rect 6736 56704 6788 56710
rect 6736 56646 6788 56652
rect 6748 56302 6776 56646
rect 6736 56296 6788 56302
rect 6736 56238 6788 56244
rect 6736 56160 6788 56166
rect 6736 56102 6788 56108
rect 6748 54534 6776 56102
rect 6736 54528 6788 54534
rect 6736 54470 6788 54476
rect 6748 54369 6776 54470
rect 6734 54360 6790 54369
rect 6734 54295 6790 54304
rect 6736 54256 6788 54262
rect 6734 54224 6736 54233
rect 6788 54224 6790 54233
rect 6734 54159 6790 54168
rect 6734 54088 6790 54097
rect 6734 54023 6790 54032
rect 6472 53502 6684 53530
rect 6368 52896 6420 52902
rect 6368 52838 6420 52844
rect 6368 52692 6420 52698
rect 6368 52634 6420 52640
rect 6092 51468 6144 51474
rect 6092 51410 6144 51416
rect 6196 51462 6316 51490
rect 6104 51066 6132 51410
rect 6092 51060 6144 51066
rect 6092 51002 6144 51008
rect 6012 50782 6132 50810
rect 6104 50402 6132 50782
rect 6012 50374 6132 50402
rect 6012 48822 6040 50374
rect 6090 50280 6146 50289
rect 6090 50215 6146 50224
rect 6104 49910 6132 50215
rect 6092 49904 6144 49910
rect 6092 49846 6144 49852
rect 6092 49700 6144 49706
rect 6092 49642 6144 49648
rect 6104 49337 6132 49642
rect 6090 49328 6146 49337
rect 6090 49263 6146 49272
rect 6000 48816 6052 48822
rect 6000 48758 6052 48764
rect 5998 48648 6054 48657
rect 5998 48583 6054 48592
rect 6012 44470 6040 48583
rect 6104 48385 6132 49263
rect 6090 48376 6146 48385
rect 6090 48311 6146 48320
rect 6092 48136 6144 48142
rect 6092 48078 6144 48084
rect 6104 47977 6132 48078
rect 6090 47968 6146 47977
rect 6090 47903 6146 47912
rect 6092 47592 6144 47598
rect 6092 47534 6144 47540
rect 6104 46510 6132 47534
rect 6092 46504 6144 46510
rect 6092 46446 6144 46452
rect 6104 45422 6132 46446
rect 6196 45626 6224 51462
rect 6380 51354 6408 52634
rect 6472 51814 6500 53502
rect 6644 53440 6696 53446
rect 6644 53382 6696 53388
rect 6656 53106 6684 53382
rect 6644 53100 6696 53106
rect 6644 53042 6696 53048
rect 6644 52964 6696 52970
rect 6644 52906 6696 52912
rect 6552 52896 6604 52902
rect 6552 52838 6604 52844
rect 6564 52154 6592 52838
rect 6552 52148 6604 52154
rect 6552 52090 6604 52096
rect 6564 51950 6592 52090
rect 6552 51944 6604 51950
rect 6552 51886 6604 51892
rect 6460 51808 6512 51814
rect 6460 51750 6512 51756
rect 6550 51776 6606 51785
rect 6288 51326 6408 51354
rect 6288 49706 6316 51326
rect 6368 51264 6420 51270
rect 6472 51241 6500 51750
rect 6550 51711 6606 51720
rect 6368 51206 6420 51212
rect 6458 51232 6514 51241
rect 6380 50318 6408 51206
rect 6458 51167 6514 51176
rect 6460 50856 6512 50862
rect 6460 50798 6512 50804
rect 6368 50312 6420 50318
rect 6368 50254 6420 50260
rect 6472 50153 6500 50798
rect 6458 50144 6514 50153
rect 6458 50079 6514 50088
rect 6460 49972 6512 49978
rect 6460 49914 6512 49920
rect 6368 49768 6420 49774
rect 6368 49710 6420 49716
rect 6276 49700 6328 49706
rect 6276 49642 6328 49648
rect 6274 49600 6330 49609
rect 6274 49535 6330 49544
rect 6288 49434 6316 49535
rect 6276 49428 6328 49434
rect 6276 49370 6328 49376
rect 6276 48816 6328 48822
rect 6276 48758 6328 48764
rect 6184 45620 6236 45626
rect 6184 45562 6236 45568
rect 6182 45520 6238 45529
rect 6182 45455 6238 45464
rect 6092 45416 6144 45422
rect 6092 45358 6144 45364
rect 6104 44810 6132 45358
rect 6196 44946 6224 45455
rect 6184 44940 6236 44946
rect 6184 44882 6236 44888
rect 6288 44826 6316 48758
rect 6092 44804 6144 44810
rect 6092 44746 6144 44752
rect 6196 44798 6316 44826
rect 6000 44464 6052 44470
rect 6000 44406 6052 44412
rect 6000 44260 6052 44266
rect 6000 44202 6052 44208
rect 6012 42362 6040 44202
rect 6104 43246 6132 44746
rect 6196 43382 6224 44798
rect 6276 44736 6328 44742
rect 6276 44678 6328 44684
rect 6288 44334 6316 44678
rect 6276 44328 6328 44334
rect 6276 44270 6328 44276
rect 6184 43376 6236 43382
rect 6184 43318 6236 43324
rect 6092 43240 6144 43246
rect 6092 43182 6144 43188
rect 6104 42634 6132 43182
rect 6196 43081 6224 43318
rect 6288 43314 6316 44270
rect 6276 43308 6328 43314
rect 6276 43250 6328 43256
rect 6182 43072 6238 43081
rect 6182 43007 6238 43016
rect 6196 42906 6224 43007
rect 6184 42900 6236 42906
rect 6184 42842 6236 42848
rect 6182 42800 6238 42809
rect 6182 42735 6238 42744
rect 6092 42628 6144 42634
rect 6092 42570 6144 42576
rect 6000 42356 6052 42362
rect 6000 42298 6052 42304
rect 6012 42158 6040 42298
rect 6000 42152 6052 42158
rect 6000 42094 6052 42100
rect 5998 41712 6054 41721
rect 5998 41647 6000 41656
rect 6052 41647 6054 41656
rect 6000 41618 6052 41624
rect 6000 41540 6052 41546
rect 6000 41482 6052 41488
rect 6012 39982 6040 41482
rect 6000 39976 6052 39982
rect 6000 39918 6052 39924
rect 5998 39536 6054 39545
rect 5998 39471 6054 39480
rect 6012 37874 6040 39471
rect 6000 37868 6052 37874
rect 6000 37810 6052 37816
rect 6000 37732 6052 37738
rect 6000 37674 6052 37680
rect 5908 36848 5960 36854
rect 5908 36790 5960 36796
rect 5816 36576 5868 36582
rect 5816 36518 5868 36524
rect 5814 36408 5870 36417
rect 5814 36343 5870 36352
rect 5724 35488 5776 35494
rect 5724 35430 5776 35436
rect 5828 34542 5856 36343
rect 6012 36281 6040 37674
rect 5998 36272 6054 36281
rect 5998 36207 6054 36216
rect 5908 36032 5960 36038
rect 5908 35974 5960 35980
rect 5816 34536 5868 34542
rect 5816 34478 5868 34484
rect 5632 33652 5684 33658
rect 5632 33594 5684 33600
rect 5632 33516 5684 33522
rect 5632 33458 5684 33464
rect 5644 32910 5672 33458
rect 5722 33416 5778 33425
rect 5722 33351 5724 33360
rect 5776 33351 5778 33360
rect 5816 33380 5868 33386
rect 5724 33322 5776 33328
rect 5816 33322 5868 33328
rect 5828 33046 5856 33322
rect 5816 33040 5868 33046
rect 5816 32982 5868 32988
rect 5632 32904 5684 32910
rect 5632 32846 5684 32852
rect 5632 32428 5684 32434
rect 5632 32370 5684 32376
rect 5644 30954 5672 32370
rect 5828 32366 5856 32982
rect 5816 32360 5868 32366
rect 5816 32302 5868 32308
rect 5814 31920 5870 31929
rect 5814 31855 5816 31864
rect 5868 31855 5870 31864
rect 5816 31826 5868 31832
rect 5920 31770 5948 35974
rect 6000 35488 6052 35494
rect 6000 35430 6052 35436
rect 6012 35154 6040 35430
rect 6000 35148 6052 35154
rect 6000 35090 6052 35096
rect 6012 34746 6040 35090
rect 6000 34740 6052 34746
rect 6000 34682 6052 34688
rect 6000 33652 6052 33658
rect 6000 33594 6052 33600
rect 6012 31890 6040 33594
rect 6000 31884 6052 31890
rect 6000 31826 6052 31832
rect 5828 31742 5948 31770
rect 5644 30926 5764 30954
rect 5632 30796 5684 30802
rect 5632 30738 5684 30744
rect 5644 30258 5672 30738
rect 5632 30252 5684 30258
rect 5632 30194 5684 30200
rect 5736 30190 5764 30926
rect 5724 30184 5776 30190
rect 5724 30126 5776 30132
rect 5736 29850 5764 30126
rect 5724 29844 5776 29850
rect 5724 29786 5776 29792
rect 5632 29776 5684 29782
rect 5632 29718 5684 29724
rect 5644 29034 5672 29718
rect 5736 29170 5764 29786
rect 5724 29164 5776 29170
rect 5724 29106 5776 29112
rect 5632 29028 5684 29034
rect 5632 28970 5684 28976
rect 5828 28626 5856 31742
rect 6012 31482 6040 31826
rect 6000 31476 6052 31482
rect 6000 31418 6052 31424
rect 6000 31136 6052 31142
rect 6000 31078 6052 31084
rect 5908 30184 5960 30190
rect 5908 30126 5960 30132
rect 5920 29782 5948 30126
rect 5908 29776 5960 29782
rect 5908 29718 5960 29724
rect 5908 29028 5960 29034
rect 5908 28970 5960 28976
rect 5816 28620 5868 28626
rect 5816 28562 5868 28568
rect 5724 28484 5776 28490
rect 5724 28426 5776 28432
rect 5632 27872 5684 27878
rect 5632 27814 5684 27820
rect 5644 26586 5672 27814
rect 5736 26858 5764 28426
rect 5920 28014 5948 28970
rect 5908 28008 5960 28014
rect 5908 27950 5960 27956
rect 5920 27674 5948 27950
rect 5908 27668 5960 27674
rect 5908 27610 5960 27616
rect 5724 26852 5776 26858
rect 5724 26794 5776 26800
rect 5632 26580 5684 26586
rect 5632 26522 5684 26528
rect 5920 25838 5948 27610
rect 5908 25832 5960 25838
rect 5908 25774 5960 25780
rect 5908 25356 5960 25362
rect 5908 25298 5960 25304
rect 5920 24614 5948 25298
rect 5908 24608 5960 24614
rect 5908 24550 5960 24556
rect 5540 24404 5592 24410
rect 5540 24346 5592 24352
rect 5920 24274 5948 24550
rect 5908 24268 5960 24274
rect 5908 24210 5960 24216
rect 5356 24132 5408 24138
rect 5356 24074 5408 24080
rect 5264 23248 5316 23254
rect 5264 23190 5316 23196
rect 5368 23186 5396 24074
rect 6012 23730 6040 31078
rect 6104 29152 6132 42570
rect 6196 41818 6224 42735
rect 6276 42152 6328 42158
rect 6276 42094 6328 42100
rect 6184 41812 6236 41818
rect 6184 41754 6236 41760
rect 6184 41608 6236 41614
rect 6184 41550 6236 41556
rect 6196 41274 6224 41550
rect 6288 41449 6316 42094
rect 6274 41440 6330 41449
rect 6274 41375 6330 41384
rect 6274 41304 6330 41313
rect 6184 41268 6236 41274
rect 6274 41239 6330 41248
rect 6184 41210 6236 41216
rect 6184 41064 6236 41070
rect 6184 41006 6236 41012
rect 6196 40730 6224 41006
rect 6184 40724 6236 40730
rect 6184 40666 6236 40672
rect 6196 40497 6224 40666
rect 6182 40488 6238 40497
rect 6182 40423 6238 40432
rect 6182 39944 6238 39953
rect 6182 39879 6184 39888
rect 6236 39879 6238 39888
rect 6184 39850 6236 39856
rect 6182 39808 6238 39817
rect 6182 39743 6238 39752
rect 6196 38894 6224 39743
rect 6184 38888 6236 38894
rect 6184 38830 6236 38836
rect 6196 38214 6224 38830
rect 6184 38208 6236 38214
rect 6184 38150 6236 38156
rect 6196 37330 6224 38150
rect 6184 37324 6236 37330
rect 6184 37266 6236 37272
rect 6288 37194 6316 41239
rect 6276 37188 6328 37194
rect 6276 37130 6328 37136
rect 6288 36922 6316 37130
rect 6276 36916 6328 36922
rect 6276 36858 6328 36864
rect 6184 36848 6236 36854
rect 6184 36790 6236 36796
rect 6196 35290 6224 36790
rect 6288 36718 6316 36858
rect 6276 36712 6328 36718
rect 6274 36680 6276 36689
rect 6328 36680 6330 36689
rect 6274 36615 6330 36624
rect 6276 36576 6328 36582
rect 6276 36518 6328 36524
rect 6184 35284 6236 35290
rect 6184 35226 6236 35232
rect 6196 34610 6224 35226
rect 6184 34604 6236 34610
rect 6184 34546 6236 34552
rect 6182 33552 6238 33561
rect 6182 33487 6238 33496
rect 6196 30870 6224 33487
rect 6288 31278 6316 36518
rect 6380 35834 6408 49710
rect 6472 44146 6500 49914
rect 6564 46050 6592 51711
rect 6656 47802 6684 52906
rect 6748 51105 6776 54023
rect 6840 52970 6868 56918
rect 6932 55894 6960 57174
rect 7024 56438 7052 58534
rect 7116 56506 7144 61882
rect 7208 61198 7236 62319
rect 7196 61192 7248 61198
rect 7196 61134 7248 61140
rect 7300 59673 7328 62630
rect 7392 61334 7420 68206
rect 8036 68134 8064 68682
rect 8024 68128 8076 68134
rect 8024 68070 8076 68076
rect 7622 68028 7918 68048
rect 7678 68026 7702 68028
rect 7758 68026 7782 68028
rect 7838 68026 7862 68028
rect 7700 67974 7702 68026
rect 7764 67974 7776 68026
rect 7838 67974 7840 68026
rect 7678 67972 7702 67974
rect 7758 67972 7782 67974
rect 7838 67972 7862 67974
rect 7622 67952 7918 67972
rect 7472 67788 7524 67794
rect 7472 67730 7524 67736
rect 7484 67046 7512 67730
rect 8036 67590 8064 68070
rect 8128 67862 8156 70450
rect 8404 70446 8432 70790
rect 8392 70440 8444 70446
rect 8390 70408 8392 70417
rect 8444 70408 8446 70417
rect 8390 70343 8446 70352
rect 8206 70272 8262 70281
rect 8206 70207 8262 70216
rect 8220 69970 8248 70207
rect 8208 69964 8260 69970
rect 8208 69906 8260 69912
rect 8392 69760 8444 69766
rect 8496 69737 8524 73335
rect 9312 73306 9364 73312
rect 9508 73234 9720 73250
rect 9220 73228 9272 73234
rect 9220 73170 9272 73176
rect 9496 73228 9720 73234
rect 9548 73222 9720 73228
rect 9496 73170 9548 73176
rect 8576 73024 8628 73030
rect 8576 72966 8628 72972
rect 8588 72758 8616 72966
rect 8576 72752 8628 72758
rect 8576 72694 8628 72700
rect 8588 72078 8616 72694
rect 9232 72486 9260 73170
rect 9312 73092 9364 73098
rect 9312 73034 9364 73040
rect 9220 72480 9272 72486
rect 9220 72422 9272 72428
rect 9232 72146 9260 72422
rect 9324 72146 9352 73034
rect 9692 72486 9720 73222
rect 10048 73228 10100 73234
rect 10048 73170 10100 73176
rect 10060 72554 10088 73170
rect 10324 72684 10376 72690
rect 10324 72626 10376 72632
rect 10048 72548 10100 72554
rect 10048 72490 10100 72496
rect 9680 72480 9732 72486
rect 9680 72422 9732 72428
rect 9220 72140 9272 72146
rect 9220 72082 9272 72088
rect 9312 72140 9364 72146
rect 9312 72082 9364 72088
rect 9680 72140 9732 72146
rect 9680 72082 9732 72088
rect 8576 72072 8628 72078
rect 8576 72014 8628 72020
rect 8852 72072 8904 72078
rect 8852 72014 8904 72020
rect 8668 71732 8720 71738
rect 8668 71674 8720 71680
rect 8576 71188 8628 71194
rect 8576 71130 8628 71136
rect 8588 70650 8616 71130
rect 8576 70644 8628 70650
rect 8576 70586 8628 70592
rect 8588 70446 8616 70586
rect 8576 70440 8628 70446
rect 8576 70382 8628 70388
rect 8392 69702 8444 69708
rect 8482 69728 8538 69737
rect 8404 69465 8432 69702
rect 8482 69663 8538 69672
rect 8390 69456 8446 69465
rect 8390 69391 8446 69400
rect 8208 69352 8260 69358
rect 8208 69294 8260 69300
rect 8220 69193 8248 69294
rect 8206 69184 8262 69193
rect 8206 69119 8262 69128
rect 8588 68882 8616 70382
rect 8576 68876 8628 68882
rect 8576 68818 8628 68824
rect 8300 68808 8352 68814
rect 8300 68750 8352 68756
rect 8312 67930 8340 68750
rect 8588 68474 8616 68818
rect 8576 68468 8628 68474
rect 8576 68410 8628 68416
rect 8484 68196 8536 68202
rect 8484 68138 8536 68144
rect 8392 68128 8444 68134
rect 8392 68070 8444 68076
rect 8404 67930 8432 68070
rect 8300 67924 8352 67930
rect 8300 67866 8352 67872
rect 8392 67924 8444 67930
rect 8392 67866 8444 67872
rect 8116 67856 8168 67862
rect 8116 67798 8168 67804
rect 8312 67674 8340 67866
rect 8128 67646 8340 67674
rect 8024 67584 8076 67590
rect 8024 67526 8076 67532
rect 8036 67182 8064 67526
rect 8024 67176 8076 67182
rect 8024 67118 8076 67124
rect 7472 67040 7524 67046
rect 7472 66982 7524 66988
rect 7484 66824 7512 66982
rect 7622 66940 7918 66960
rect 7678 66938 7702 66940
rect 7758 66938 7782 66940
rect 7838 66938 7862 66940
rect 7700 66886 7702 66938
rect 7764 66886 7776 66938
rect 7838 66886 7840 66938
rect 7678 66884 7702 66886
rect 7758 66884 7782 66886
rect 7838 66884 7862 66886
rect 7622 66864 7918 66884
rect 7484 66796 7604 66824
rect 7472 66700 7524 66706
rect 7472 66642 7524 66648
rect 7484 66298 7512 66642
rect 7472 66292 7524 66298
rect 7472 66234 7524 66240
rect 7576 66201 7604 66796
rect 7562 66192 7618 66201
rect 7562 66127 7618 66136
rect 7472 65952 7524 65958
rect 7472 65894 7524 65900
rect 7484 65618 7512 65894
rect 7622 65852 7918 65872
rect 7678 65850 7702 65852
rect 7758 65850 7782 65852
rect 7838 65850 7862 65852
rect 7700 65798 7702 65850
rect 7764 65798 7776 65850
rect 7838 65798 7840 65850
rect 7678 65796 7702 65798
rect 7758 65796 7782 65798
rect 7838 65796 7862 65798
rect 7622 65776 7918 65796
rect 8036 65736 8064 67118
rect 8128 66094 8156 67646
rect 8404 67538 8432 67866
rect 8220 67510 8432 67538
rect 8220 66706 8248 67510
rect 8208 66700 8260 66706
rect 8208 66642 8260 66648
rect 8208 66496 8260 66502
rect 8260 66456 8340 66484
rect 8208 66438 8260 66444
rect 8116 66088 8168 66094
rect 8116 66030 8168 66036
rect 7944 65708 8064 65736
rect 7944 65618 7972 65708
rect 8128 65634 8156 66030
rect 8208 66020 8260 66026
rect 8208 65962 8260 65968
rect 7472 65612 7524 65618
rect 7472 65554 7524 65560
rect 7932 65612 7984 65618
rect 7932 65554 7984 65560
rect 8036 65606 8156 65634
rect 7472 65476 7524 65482
rect 7472 65418 7524 65424
rect 7484 64870 7512 65418
rect 7944 65210 7972 65554
rect 7932 65204 7984 65210
rect 7932 65146 7984 65152
rect 7472 64864 7524 64870
rect 7472 64806 7524 64812
rect 7484 63782 7512 64806
rect 7622 64764 7918 64784
rect 7678 64762 7702 64764
rect 7758 64762 7782 64764
rect 7838 64762 7862 64764
rect 7700 64710 7702 64762
rect 7764 64710 7776 64762
rect 7838 64710 7840 64762
rect 7678 64708 7702 64710
rect 7758 64708 7782 64710
rect 7838 64708 7862 64710
rect 7622 64688 7918 64708
rect 7932 63912 7984 63918
rect 7930 63880 7932 63889
rect 7984 63880 7986 63889
rect 7930 63815 7986 63824
rect 7472 63776 7524 63782
rect 7472 63718 7524 63724
rect 7622 63676 7918 63696
rect 7678 63674 7702 63676
rect 7758 63674 7782 63676
rect 7838 63674 7862 63676
rect 7700 63622 7702 63674
rect 7764 63622 7776 63674
rect 7838 63622 7840 63674
rect 7678 63620 7702 63622
rect 7758 63620 7782 63622
rect 7838 63620 7862 63622
rect 7622 63600 7918 63620
rect 8036 63442 8064 65606
rect 8116 65544 8168 65550
rect 8220 65521 8248 65962
rect 8116 65486 8168 65492
rect 8206 65512 8262 65521
rect 8024 63436 8076 63442
rect 8024 63378 8076 63384
rect 7748 63368 7800 63374
rect 7746 63336 7748 63345
rect 7800 63336 7802 63345
rect 7746 63271 7802 63280
rect 7472 62824 7524 62830
rect 7760 62801 7788 63271
rect 7472 62766 7524 62772
rect 7746 62792 7802 62801
rect 7380 61328 7432 61334
rect 7380 61270 7432 61276
rect 7380 61192 7432 61198
rect 7380 61134 7432 61140
rect 7392 60314 7420 61134
rect 7380 60308 7432 60314
rect 7380 60250 7432 60256
rect 7286 59664 7342 59673
rect 7286 59599 7342 59608
rect 7288 59560 7340 59566
rect 7392 59548 7420 60250
rect 7340 59520 7420 59548
rect 7288 59502 7340 59508
rect 7196 59492 7248 59498
rect 7196 59434 7248 59440
rect 7208 58886 7236 59434
rect 7286 59392 7342 59401
rect 7286 59327 7342 59336
rect 7196 58880 7248 58886
rect 7196 58822 7248 58828
rect 7104 56500 7156 56506
rect 7104 56442 7156 56448
rect 7012 56432 7064 56438
rect 7012 56374 7064 56380
rect 7012 56296 7064 56302
rect 7012 56238 7064 56244
rect 7024 56001 7052 56238
rect 7010 55992 7066 56001
rect 7010 55927 7066 55936
rect 6920 55888 6972 55894
rect 6920 55830 6972 55836
rect 7012 55820 7064 55826
rect 7012 55762 7064 55768
rect 6920 55752 6972 55758
rect 6920 55694 6972 55700
rect 6932 54602 6960 55694
rect 7024 55282 7052 55762
rect 7012 55276 7064 55282
rect 7012 55218 7064 55224
rect 6920 54596 6972 54602
rect 6920 54538 6972 54544
rect 6920 54188 6972 54194
rect 6920 54130 6972 54136
rect 6932 53582 6960 54130
rect 6920 53576 6972 53582
rect 6920 53518 6972 53524
rect 6920 53168 6972 53174
rect 6920 53110 6972 53116
rect 6828 52964 6880 52970
rect 6828 52906 6880 52912
rect 6932 52170 6960 53110
rect 7024 53038 7052 55218
rect 7012 53032 7064 53038
rect 7012 52974 7064 52980
rect 7104 53032 7156 53038
rect 7104 52974 7156 52980
rect 7010 52592 7066 52601
rect 7010 52527 7066 52536
rect 6840 52142 6960 52170
rect 6840 52086 6868 52142
rect 7024 52086 7052 52527
rect 7116 52494 7144 52974
rect 7104 52488 7156 52494
rect 7104 52430 7156 52436
rect 6828 52080 6880 52086
rect 6828 52022 6880 52028
rect 7012 52080 7064 52086
rect 7012 52022 7064 52028
rect 6828 51876 6880 51882
rect 6880 51836 6960 51864
rect 6828 51818 6880 51824
rect 6826 51640 6882 51649
rect 6826 51575 6882 51584
rect 6840 51406 6868 51575
rect 6828 51400 6880 51406
rect 6828 51342 6880 51348
rect 6734 51096 6790 51105
rect 6734 51031 6790 51040
rect 6826 50960 6882 50969
rect 6826 50895 6882 50904
rect 6736 50788 6788 50794
rect 6736 50730 6788 50736
rect 6644 47796 6696 47802
rect 6644 47738 6696 47744
rect 6642 47696 6698 47705
rect 6642 47631 6698 47640
rect 6656 47258 6684 47631
rect 6644 47252 6696 47258
rect 6644 47194 6696 47200
rect 6656 46986 6684 47194
rect 6644 46980 6696 46986
rect 6644 46922 6696 46928
rect 6748 46170 6776 50730
rect 6840 50454 6868 50895
rect 6828 50448 6880 50454
rect 6828 50390 6880 50396
rect 6828 49700 6880 49706
rect 6828 49642 6880 49648
rect 6840 49434 6868 49642
rect 6828 49428 6880 49434
rect 6828 49370 6880 49376
rect 6932 49298 6960 51836
rect 7012 51536 7064 51542
rect 7010 51504 7012 51513
rect 7064 51504 7066 51513
rect 7010 51439 7066 51448
rect 7012 51400 7064 51406
rect 7012 51342 7064 51348
rect 7024 50862 7052 51342
rect 7012 50856 7064 50862
rect 7010 50824 7012 50833
rect 7064 50824 7066 50833
rect 7010 50759 7066 50768
rect 7012 50720 7064 50726
rect 7012 50662 7064 50668
rect 7024 49910 7052 50662
rect 7012 49904 7064 49910
rect 7012 49846 7064 49852
rect 7012 49768 7064 49774
rect 7012 49710 7064 49716
rect 7024 49298 7052 49710
rect 6920 49292 6972 49298
rect 6920 49234 6972 49240
rect 7012 49292 7064 49298
rect 7012 49234 7064 49240
rect 6920 48748 6972 48754
rect 6920 48690 6972 48696
rect 6828 48680 6880 48686
rect 6828 48622 6880 48628
rect 6736 46164 6788 46170
rect 6736 46106 6788 46112
rect 6564 46022 6776 46050
rect 6552 45960 6604 45966
rect 6552 45902 6604 45908
rect 6564 44266 6592 45902
rect 6644 45824 6696 45830
rect 6644 45766 6696 45772
rect 6656 45422 6684 45766
rect 6644 45416 6696 45422
rect 6644 45358 6696 45364
rect 6552 44260 6604 44266
rect 6552 44202 6604 44208
rect 6472 44118 6592 44146
rect 6460 43648 6512 43654
rect 6460 43590 6512 43596
rect 6472 36038 6500 43590
rect 6460 36032 6512 36038
rect 6460 35974 6512 35980
rect 6368 35828 6420 35834
rect 6420 35788 6500 35816
rect 6368 35770 6420 35776
rect 6368 34536 6420 34542
rect 6368 34478 6420 34484
rect 6380 34134 6408 34478
rect 6368 34128 6420 34134
rect 6368 34070 6420 34076
rect 6380 33153 6408 34070
rect 6366 33144 6422 33153
rect 6366 33079 6422 33088
rect 6368 32972 6420 32978
rect 6368 32914 6420 32920
rect 6380 32366 6408 32914
rect 6368 32360 6420 32366
rect 6368 32302 6420 32308
rect 6380 31958 6408 32302
rect 6368 31952 6420 31958
rect 6368 31894 6420 31900
rect 6366 31784 6422 31793
rect 6366 31719 6422 31728
rect 6276 31272 6328 31278
rect 6276 31214 6328 31220
rect 6184 30864 6236 30870
rect 6184 30806 6236 30812
rect 6184 29164 6236 29170
rect 6104 29124 6184 29152
rect 6184 29106 6236 29112
rect 6092 28008 6144 28014
rect 6092 27950 6144 27956
rect 6104 27334 6132 27950
rect 6092 27328 6144 27334
rect 6092 27270 6144 27276
rect 6104 27062 6132 27270
rect 6092 27056 6144 27062
rect 6092 26998 6144 27004
rect 6000 23724 6052 23730
rect 6000 23666 6052 23672
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5356 23180 5408 23186
rect 5356 23122 5408 23128
rect 5356 22976 5408 22982
rect 5170 22944 5226 22953
rect 5356 22918 5408 22924
rect 5170 22879 5226 22888
rect 5184 22574 5212 22879
rect 5368 22642 5396 22918
rect 5356 22636 5408 22642
rect 5356 22578 5408 22584
rect 4988 22568 5040 22574
rect 4988 22510 5040 22516
rect 5172 22568 5224 22574
rect 5172 22510 5224 22516
rect 4804 22432 4856 22438
rect 4804 22374 4856 22380
rect 4712 22228 4764 22234
rect 4712 22170 4764 22176
rect 4289 21788 4585 21808
rect 4345 21786 4369 21788
rect 4425 21786 4449 21788
rect 4505 21786 4529 21788
rect 4367 21734 4369 21786
rect 4431 21734 4443 21786
rect 4505 21734 4507 21786
rect 4345 21732 4369 21734
rect 4425 21732 4449 21734
rect 4505 21732 4529 21734
rect 4289 21712 4585 21732
rect 4816 21010 4844 22374
rect 5000 22234 5028 22510
rect 4988 22228 5040 22234
rect 4988 22170 5040 22176
rect 5080 21956 5132 21962
rect 5080 21898 5132 21904
rect 4804 21004 4856 21010
rect 4804 20946 4856 20952
rect 4160 20800 4212 20806
rect 4160 20742 4212 20748
rect 4068 20392 4120 20398
rect 4172 20380 4200 20742
rect 4289 20700 4585 20720
rect 4345 20698 4369 20700
rect 4425 20698 4449 20700
rect 4505 20698 4529 20700
rect 4367 20646 4369 20698
rect 4431 20646 4443 20698
rect 4505 20646 4507 20698
rect 4345 20644 4369 20646
rect 4425 20644 4449 20646
rect 4505 20644 4529 20646
rect 4289 20624 4585 20644
rect 4120 20352 4200 20380
rect 4068 20334 4120 20340
rect 4066 19272 4122 19281
rect 4066 19207 4068 19216
rect 4120 19207 4122 19216
rect 4068 19178 4120 19184
rect 4172 19174 4200 20352
rect 4712 19712 4764 19718
rect 4712 19654 4764 19660
rect 4289 19612 4585 19632
rect 4345 19610 4369 19612
rect 4425 19610 4449 19612
rect 4505 19610 4529 19612
rect 4367 19558 4369 19610
rect 4431 19558 4443 19610
rect 4505 19558 4507 19610
rect 4345 19556 4369 19558
rect 4425 19556 4449 19558
rect 4505 19556 4529 19558
rect 4289 19536 4585 19556
rect 4724 19417 4752 19654
rect 4710 19408 4766 19417
rect 4710 19343 4766 19352
rect 5092 19310 5120 21898
rect 5460 21570 5488 23598
rect 5906 23488 5962 23497
rect 5906 23423 5962 23432
rect 5920 23118 5948 23423
rect 5908 23112 5960 23118
rect 5908 23054 5960 23060
rect 5724 22092 5776 22098
rect 5724 22034 5776 22040
rect 5460 21554 5580 21570
rect 5460 21548 5592 21554
rect 5460 21542 5540 21548
rect 5540 21490 5592 21496
rect 5736 21418 5764 22034
rect 5724 21412 5776 21418
rect 5724 21354 5776 21360
rect 5920 21078 5948 23054
rect 6196 22234 6224 29106
rect 6380 29102 6408 31719
rect 6368 29096 6420 29102
rect 6368 29038 6420 29044
rect 6472 26586 6500 35788
rect 6564 33454 6592 44118
rect 6656 43722 6684 45358
rect 6644 43716 6696 43722
rect 6644 43658 6696 43664
rect 6656 43246 6684 43658
rect 6644 43240 6696 43246
rect 6644 43182 6696 43188
rect 6656 39930 6684 43182
rect 6748 41052 6776 46022
rect 6840 44962 6868 48622
rect 6932 48550 6960 48690
rect 6920 48544 6972 48550
rect 6920 48486 6972 48492
rect 6932 48142 6960 48486
rect 7024 48278 7052 49234
rect 7012 48272 7064 48278
rect 7012 48214 7064 48220
rect 6920 48136 6972 48142
rect 6972 48096 7052 48124
rect 6920 48078 6972 48084
rect 6920 48000 6972 48006
rect 6920 47942 6972 47948
rect 6932 47841 6960 47942
rect 6918 47832 6974 47841
rect 6918 47767 6974 47776
rect 6920 47592 6972 47598
rect 6920 47534 6972 47540
rect 6932 46510 6960 47534
rect 6920 46504 6972 46510
rect 6920 46446 6972 46452
rect 6932 45830 6960 46446
rect 7024 46170 7052 48096
rect 7012 46164 7064 46170
rect 7012 46106 7064 46112
rect 6920 45824 6972 45830
rect 6920 45766 6972 45772
rect 7024 45121 7052 46106
rect 7010 45112 7066 45121
rect 7010 45047 7066 45056
rect 7116 45014 7144 52430
rect 7208 50930 7236 58822
rect 7300 57390 7328 59327
rect 7380 59084 7432 59090
rect 7380 59026 7432 59032
rect 7392 58993 7420 59026
rect 7378 58984 7434 58993
rect 7378 58919 7434 58928
rect 7288 57384 7340 57390
rect 7288 57326 7340 57332
rect 7380 57248 7432 57254
rect 7380 57190 7432 57196
rect 7288 56500 7340 56506
rect 7288 56442 7340 56448
rect 7300 55758 7328 56442
rect 7288 55752 7340 55758
rect 7288 55694 7340 55700
rect 7392 55706 7420 57190
rect 7484 56778 7512 62766
rect 7746 62727 7748 62736
rect 7800 62727 7802 62736
rect 7748 62698 7800 62704
rect 7622 62588 7918 62608
rect 7678 62586 7702 62588
rect 7758 62586 7782 62588
rect 7838 62586 7862 62588
rect 7700 62534 7702 62586
rect 7764 62534 7776 62586
rect 7838 62534 7840 62586
rect 7678 62532 7702 62534
rect 7758 62532 7782 62534
rect 7838 62532 7862 62534
rect 7622 62512 7918 62532
rect 7622 61500 7918 61520
rect 7678 61498 7702 61500
rect 7758 61498 7782 61500
rect 7838 61498 7862 61500
rect 7700 61446 7702 61498
rect 7764 61446 7776 61498
rect 7838 61446 7840 61498
rect 7678 61444 7702 61446
rect 7758 61444 7782 61446
rect 7838 61444 7862 61446
rect 7622 61424 7918 61444
rect 7564 61328 7616 61334
rect 7564 61270 7616 61276
rect 8024 61328 8076 61334
rect 8024 61270 8076 61276
rect 7576 60625 7604 61270
rect 7562 60616 7618 60625
rect 7562 60551 7618 60560
rect 8036 60518 8064 61270
rect 8024 60512 8076 60518
rect 8024 60454 8076 60460
rect 7622 60412 7918 60432
rect 7678 60410 7702 60412
rect 7758 60410 7782 60412
rect 7838 60410 7862 60412
rect 7700 60358 7702 60410
rect 7764 60358 7776 60410
rect 7838 60358 7840 60410
rect 7678 60356 7702 60358
rect 7758 60356 7782 60358
rect 7838 60356 7862 60358
rect 7622 60336 7918 60356
rect 7622 59324 7918 59344
rect 7678 59322 7702 59324
rect 7758 59322 7782 59324
rect 7838 59322 7862 59324
rect 7700 59270 7702 59322
rect 7764 59270 7776 59322
rect 7838 59270 7840 59322
rect 7678 59268 7702 59270
rect 7758 59268 7782 59270
rect 7838 59268 7862 59270
rect 7622 59248 7918 59268
rect 8036 58682 8064 60454
rect 8024 58676 8076 58682
rect 8024 58618 8076 58624
rect 8024 58336 8076 58342
rect 8024 58278 8076 58284
rect 7622 58236 7918 58256
rect 7678 58234 7702 58236
rect 7758 58234 7782 58236
rect 7838 58234 7862 58236
rect 7700 58182 7702 58234
rect 7764 58182 7776 58234
rect 7838 58182 7840 58234
rect 7678 58180 7702 58182
rect 7758 58180 7782 58182
rect 7838 58180 7862 58182
rect 7622 58160 7918 58180
rect 7932 58064 7984 58070
rect 7562 58032 7618 58041
rect 7932 58006 7984 58012
rect 7562 57967 7618 57976
rect 7656 57996 7708 58002
rect 7576 57526 7604 57967
rect 7656 57938 7708 57944
rect 7840 57996 7892 58002
rect 7840 57938 7892 57944
rect 7564 57520 7616 57526
rect 7564 57462 7616 57468
rect 7668 57322 7696 57938
rect 7852 57905 7880 57938
rect 7838 57896 7894 57905
rect 7838 57831 7894 57840
rect 7852 57798 7880 57831
rect 7840 57792 7892 57798
rect 7840 57734 7892 57740
rect 7944 57361 7972 58006
rect 7930 57352 7986 57361
rect 7656 57316 7708 57322
rect 7930 57287 7986 57296
rect 7656 57258 7708 57264
rect 7622 57148 7918 57168
rect 7678 57146 7702 57148
rect 7758 57146 7782 57148
rect 7838 57146 7862 57148
rect 7700 57094 7702 57146
rect 7764 57094 7776 57146
rect 7838 57094 7840 57146
rect 7678 57092 7702 57094
rect 7758 57092 7782 57094
rect 7838 57092 7862 57094
rect 7622 57072 7918 57092
rect 7840 56840 7892 56846
rect 7840 56782 7892 56788
rect 7472 56772 7524 56778
rect 7472 56714 7524 56720
rect 7852 56506 7880 56782
rect 7840 56500 7892 56506
rect 7840 56442 7892 56448
rect 7472 56228 7524 56234
rect 7472 56170 7524 56176
rect 7484 55826 7512 56170
rect 7622 56060 7918 56080
rect 7678 56058 7702 56060
rect 7758 56058 7782 56060
rect 7838 56058 7862 56060
rect 7700 56006 7702 56058
rect 7764 56006 7776 56058
rect 7838 56006 7840 56058
rect 7678 56004 7702 56006
rect 7758 56004 7782 56006
rect 7838 56004 7862 56006
rect 7622 55984 7918 56004
rect 7472 55820 7524 55826
rect 7472 55762 7524 55768
rect 7392 55678 7512 55706
rect 7380 55140 7432 55146
rect 7380 55082 7432 55088
rect 7288 55072 7340 55078
rect 7286 55040 7288 55049
rect 7340 55040 7342 55049
rect 7286 54975 7342 54984
rect 7288 54664 7340 54670
rect 7288 54606 7340 54612
rect 7196 50924 7248 50930
rect 7196 50866 7248 50872
rect 7300 50810 7328 54606
rect 7392 53961 7420 55082
rect 7378 53952 7434 53961
rect 7378 53887 7434 53896
rect 7484 53514 7512 55678
rect 7622 54972 7918 54992
rect 7678 54970 7702 54972
rect 7758 54970 7782 54972
rect 7838 54970 7862 54972
rect 7700 54918 7702 54970
rect 7764 54918 7776 54970
rect 7838 54918 7840 54970
rect 7678 54916 7702 54918
rect 7758 54916 7782 54918
rect 7838 54916 7862 54918
rect 7622 54896 7918 54916
rect 7838 54768 7894 54777
rect 7838 54703 7894 54712
rect 7852 54126 7880 54703
rect 7840 54120 7892 54126
rect 7840 54062 7892 54068
rect 7622 53884 7918 53904
rect 7678 53882 7702 53884
rect 7758 53882 7782 53884
rect 7838 53882 7862 53884
rect 7700 53830 7702 53882
rect 7764 53830 7776 53882
rect 7838 53830 7840 53882
rect 7678 53828 7702 53830
rect 7758 53828 7782 53830
rect 7838 53828 7862 53830
rect 7622 53808 7918 53828
rect 7472 53508 7524 53514
rect 7472 53450 7524 53456
rect 7380 53440 7432 53446
rect 7380 53382 7432 53388
rect 7392 53174 7420 53382
rect 7380 53168 7432 53174
rect 7380 53110 7432 53116
rect 7472 53100 7524 53106
rect 7472 53042 7524 53048
rect 7380 52896 7432 52902
rect 7380 52838 7432 52844
rect 7208 50782 7328 50810
rect 7392 50794 7420 52838
rect 7484 52698 7512 53042
rect 7622 52796 7918 52816
rect 7678 52794 7702 52796
rect 7758 52794 7782 52796
rect 7838 52794 7862 52796
rect 7700 52742 7702 52794
rect 7764 52742 7776 52794
rect 7838 52742 7840 52794
rect 7678 52740 7702 52742
rect 7758 52740 7782 52742
rect 7838 52740 7862 52742
rect 7622 52720 7918 52740
rect 7472 52692 7524 52698
rect 7472 52634 7524 52640
rect 7472 52488 7524 52494
rect 7472 52430 7524 52436
rect 7484 51338 7512 52430
rect 7622 51708 7918 51728
rect 7678 51706 7702 51708
rect 7758 51706 7782 51708
rect 7838 51706 7862 51708
rect 7700 51654 7702 51706
rect 7764 51654 7776 51706
rect 7838 51654 7840 51706
rect 7678 51652 7702 51654
rect 7758 51652 7782 51654
rect 7838 51652 7862 51654
rect 7622 51632 7918 51652
rect 7564 51536 7616 51542
rect 7564 51478 7616 51484
rect 7930 51504 7986 51513
rect 7472 51332 7524 51338
rect 7472 51274 7524 51280
rect 7484 50998 7512 51274
rect 7576 51066 7604 51478
rect 7748 51468 7800 51474
rect 7930 51439 7932 51448
rect 7748 51410 7800 51416
rect 7984 51439 7986 51448
rect 7932 51410 7984 51416
rect 7760 51377 7788 51410
rect 7746 51368 7802 51377
rect 7802 51326 7880 51354
rect 7746 51303 7802 51312
rect 7748 51264 7800 51270
rect 7748 51206 7800 51212
rect 7564 51060 7616 51066
rect 7564 51002 7616 51008
rect 7472 50992 7524 50998
rect 7472 50934 7524 50940
rect 7760 50862 7788 51206
rect 7852 51066 7880 51326
rect 7840 51060 7892 51066
rect 7840 51002 7892 51008
rect 7944 50998 7972 51410
rect 7932 50992 7984 50998
rect 7932 50934 7984 50940
rect 7472 50856 7524 50862
rect 7472 50798 7524 50804
rect 7748 50856 7800 50862
rect 7748 50798 7800 50804
rect 7380 50788 7432 50794
rect 7208 50454 7236 50782
rect 7380 50730 7432 50736
rect 7288 50720 7340 50726
rect 7288 50662 7340 50668
rect 7196 50448 7248 50454
rect 7196 50390 7248 50396
rect 7196 50312 7248 50318
rect 7196 50254 7248 50260
rect 7208 48278 7236 50254
rect 7300 48890 7328 50662
rect 7392 50522 7420 50730
rect 7380 50516 7432 50522
rect 7380 50458 7432 50464
rect 7484 50402 7512 50798
rect 7622 50620 7918 50640
rect 7678 50618 7702 50620
rect 7758 50618 7782 50620
rect 7838 50618 7862 50620
rect 7700 50566 7702 50618
rect 7764 50566 7776 50618
rect 7838 50566 7840 50618
rect 7678 50564 7702 50566
rect 7758 50564 7782 50566
rect 7838 50564 7862 50566
rect 7622 50544 7918 50564
rect 8036 50504 8064 58278
rect 8128 53666 8156 65486
rect 8206 65447 8262 65456
rect 8312 65006 8340 66456
rect 8392 65612 8444 65618
rect 8392 65554 8444 65560
rect 8300 65000 8352 65006
rect 8300 64942 8352 64948
rect 8298 64832 8354 64841
rect 8298 64767 8354 64776
rect 8312 64530 8340 64767
rect 8404 64666 8432 65554
rect 8496 64954 8524 68138
rect 8576 67040 8628 67046
rect 8576 66982 8628 66988
rect 8588 66842 8616 66982
rect 8576 66836 8628 66842
rect 8576 66778 8628 66784
rect 8576 66088 8628 66094
rect 8576 66030 8628 66036
rect 8588 65754 8616 66030
rect 8576 65748 8628 65754
rect 8576 65690 8628 65696
rect 8496 64926 8616 64954
rect 8484 64864 8536 64870
rect 8484 64806 8536 64812
rect 8392 64660 8444 64666
rect 8392 64602 8444 64608
rect 8300 64524 8352 64530
rect 8300 64466 8352 64472
rect 8208 64456 8260 64462
rect 8260 64404 8340 64410
rect 8208 64398 8340 64404
rect 8220 64382 8340 64398
rect 8208 63912 8260 63918
rect 8208 63854 8260 63860
rect 8220 60058 8248 63854
rect 8312 63238 8340 64382
rect 8404 63986 8432 64602
rect 8496 64598 8524 64806
rect 8588 64682 8616 64926
rect 8680 64841 8708 71674
rect 8864 71534 8892 72014
rect 8944 72004 8996 72010
rect 8944 71946 8996 71952
rect 8852 71528 8904 71534
rect 8852 71470 8904 71476
rect 8760 71460 8812 71466
rect 8760 71402 8812 71408
rect 8772 71058 8800 71402
rect 8850 71088 8906 71097
rect 8760 71052 8812 71058
rect 8850 71023 8906 71032
rect 8760 70994 8812 71000
rect 8772 70106 8800 70994
rect 8760 70100 8812 70106
rect 8760 70042 8812 70048
rect 8864 68202 8892 71023
rect 8852 68196 8904 68202
rect 8852 68138 8904 68144
rect 8956 67946 8984 71946
rect 9232 71398 9260 72082
rect 9324 71738 9352 72082
rect 9402 72040 9458 72049
rect 9402 71975 9458 71984
rect 9312 71732 9364 71738
rect 9312 71674 9364 71680
rect 9220 71392 9272 71398
rect 9220 71334 9272 71340
rect 9232 68762 9260 71334
rect 9416 69329 9444 71975
rect 9692 71210 9720 72082
rect 9600 71194 9720 71210
rect 9588 71188 9720 71194
rect 9640 71182 9720 71188
rect 9588 71130 9640 71136
rect 9600 71074 9628 71130
rect 9508 71046 9628 71074
rect 9508 69562 9536 71046
rect 9588 70984 9640 70990
rect 9588 70926 9640 70932
rect 9600 70689 9628 70926
rect 9586 70680 9642 70689
rect 9586 70615 9642 70624
rect 9772 70440 9824 70446
rect 9678 70408 9734 70417
rect 9772 70382 9824 70388
rect 9678 70343 9734 70352
rect 9588 70304 9640 70310
rect 9588 70246 9640 70252
rect 9600 70009 9628 70246
rect 9692 70122 9720 70343
rect 9784 70281 9812 70382
rect 9770 70272 9826 70281
rect 9770 70207 9826 70216
rect 9692 70094 9812 70122
rect 9586 70000 9642 70009
rect 9586 69935 9642 69944
rect 9680 69964 9732 69970
rect 9680 69906 9732 69912
rect 9496 69556 9548 69562
rect 9496 69498 9548 69504
rect 9402 69320 9458 69329
rect 9692 69290 9720 69906
rect 9784 69902 9812 70094
rect 9956 70032 10008 70038
rect 9956 69974 10008 69980
rect 9772 69896 9824 69902
rect 9772 69838 9824 69844
rect 9864 69828 9916 69834
rect 9864 69770 9916 69776
rect 9770 69320 9826 69329
rect 9402 69255 9458 69264
rect 9680 69284 9732 69290
rect 9770 69255 9826 69264
rect 9680 69226 9732 69232
rect 9496 69216 9548 69222
rect 9402 69184 9458 69193
rect 9496 69158 9548 69164
rect 9402 69119 9458 69128
rect 8772 67918 8984 67946
rect 9048 68734 9260 68762
rect 8772 65754 8800 67918
rect 8944 67788 8996 67794
rect 8944 67730 8996 67736
rect 8956 67046 8984 67730
rect 8944 67040 8996 67046
rect 8944 66982 8996 66988
rect 8760 65748 8812 65754
rect 8760 65690 8812 65696
rect 8760 65612 8812 65618
rect 8760 65554 8812 65560
rect 8772 64870 8800 65554
rect 8956 65006 8984 66982
rect 8944 65000 8996 65006
rect 8944 64942 8996 64948
rect 8852 64932 8904 64938
rect 8852 64874 8904 64880
rect 8760 64864 8812 64870
rect 8666 64832 8722 64841
rect 8760 64806 8812 64812
rect 8666 64767 8722 64776
rect 8588 64654 8800 64682
rect 8484 64592 8536 64598
rect 8484 64534 8536 64540
rect 8392 63980 8444 63986
rect 8392 63922 8444 63928
rect 8496 63918 8524 64534
rect 8576 64524 8628 64530
rect 8576 64466 8628 64472
rect 8484 63912 8536 63918
rect 8484 63854 8536 63860
rect 8484 63776 8536 63782
rect 8484 63718 8536 63724
rect 8390 63472 8446 63481
rect 8390 63407 8446 63416
rect 8300 63232 8352 63238
rect 8300 63174 8352 63180
rect 8404 62762 8432 63407
rect 8392 62756 8444 62762
rect 8392 62698 8444 62704
rect 8496 61810 8524 63718
rect 8588 63578 8616 64466
rect 8668 64456 8720 64462
rect 8668 64398 8720 64404
rect 8576 63572 8628 63578
rect 8576 63514 8628 63520
rect 8574 63472 8630 63481
rect 8574 63407 8630 63416
rect 8484 61804 8536 61810
rect 8484 61746 8536 61752
rect 8484 61600 8536 61606
rect 8484 61542 8536 61548
rect 8298 61296 8354 61305
rect 8298 61231 8300 61240
rect 8352 61231 8354 61240
rect 8300 61202 8352 61208
rect 8300 61056 8352 61062
rect 8300 60998 8352 61004
rect 8312 60654 8340 60998
rect 8496 60858 8524 61542
rect 8484 60852 8536 60858
rect 8484 60794 8536 60800
rect 8300 60648 8352 60654
rect 8300 60590 8352 60596
rect 8312 60314 8340 60590
rect 8392 60512 8444 60518
rect 8588 60466 8616 63407
rect 8680 61146 8708 64398
rect 8772 62937 8800 64654
rect 8758 62928 8814 62937
rect 8758 62863 8814 62872
rect 8760 62688 8812 62694
rect 8760 62630 8812 62636
rect 8772 61946 8800 62630
rect 8760 61940 8812 61946
rect 8760 61882 8812 61888
rect 8772 61266 8800 61882
rect 8760 61260 8812 61266
rect 8760 61202 8812 61208
rect 8680 61118 8800 61146
rect 8668 61056 8720 61062
rect 8668 60998 8720 61004
rect 8392 60454 8444 60460
rect 8300 60308 8352 60314
rect 8300 60250 8352 60256
rect 8404 60217 8432 60454
rect 8496 60438 8616 60466
rect 8390 60208 8446 60217
rect 8390 60143 8446 60152
rect 8220 60030 8432 60058
rect 8300 59968 8352 59974
rect 8220 59928 8300 59956
rect 8220 58342 8248 59928
rect 8300 59910 8352 59916
rect 8404 59158 8432 60030
rect 8496 59650 8524 60438
rect 8680 60296 8708 60998
rect 8588 60268 8708 60296
rect 8588 59974 8616 60268
rect 8668 60172 8720 60178
rect 8668 60114 8720 60120
rect 8576 59968 8628 59974
rect 8576 59910 8628 59916
rect 8496 59622 8616 59650
rect 8484 59492 8536 59498
rect 8484 59434 8536 59440
rect 8392 59152 8444 59158
rect 8392 59094 8444 59100
rect 8496 59090 8524 59434
rect 8484 59084 8536 59090
rect 8484 59026 8536 59032
rect 8300 58880 8352 58886
rect 8298 58848 8300 58857
rect 8352 58848 8354 58857
rect 8298 58783 8354 58792
rect 8312 58478 8340 58783
rect 8300 58472 8352 58478
rect 8300 58414 8352 58420
rect 8208 58336 8260 58342
rect 8208 58278 8260 58284
rect 8312 58154 8340 58414
rect 8220 58126 8340 58154
rect 8220 56930 8248 58126
rect 8392 57928 8444 57934
rect 8392 57870 8444 57876
rect 8404 57254 8432 57870
rect 8392 57248 8444 57254
rect 8392 57190 8444 57196
rect 8220 56902 8340 56930
rect 8208 56840 8260 56846
rect 8208 56782 8260 56788
rect 8220 54738 8248 56782
rect 8312 56302 8340 56902
rect 8300 56296 8352 56302
rect 8300 56238 8352 56244
rect 8298 55992 8354 56001
rect 8298 55927 8300 55936
rect 8352 55927 8354 55936
rect 8300 55898 8352 55904
rect 8312 55282 8340 55898
rect 8300 55276 8352 55282
rect 8300 55218 8352 55224
rect 8404 55214 8432 57190
rect 8392 55208 8444 55214
rect 8392 55150 8444 55156
rect 8208 54732 8260 54738
rect 8208 54674 8260 54680
rect 8392 54732 8444 54738
rect 8392 54674 8444 54680
rect 8300 54528 8352 54534
rect 8404 54505 8432 54674
rect 8300 54470 8352 54476
rect 8390 54496 8446 54505
rect 8312 54194 8340 54470
rect 8390 54431 8446 54440
rect 8300 54188 8352 54194
rect 8300 54130 8352 54136
rect 8392 54120 8444 54126
rect 8392 54062 8444 54068
rect 8300 54052 8352 54058
rect 8300 53994 8352 54000
rect 8128 53638 8248 53666
rect 8116 53576 8168 53582
rect 8116 53518 8168 53524
rect 8128 53242 8156 53518
rect 8116 53236 8168 53242
rect 8116 53178 8168 53184
rect 8128 52873 8156 53178
rect 8220 52902 8248 53638
rect 8208 52896 8260 52902
rect 8114 52864 8170 52873
rect 8208 52838 8260 52844
rect 8114 52799 8170 52808
rect 8206 52728 8262 52737
rect 8206 52663 8262 52672
rect 8220 52630 8248 52663
rect 8208 52624 8260 52630
rect 8208 52566 8260 52572
rect 8208 52488 8260 52494
rect 8114 52456 8170 52465
rect 8208 52430 8260 52436
rect 8114 52391 8170 52400
rect 8128 51542 8156 52391
rect 8220 51814 8248 52430
rect 8208 51808 8260 51814
rect 8312 51796 8340 53994
rect 8404 53446 8432 54062
rect 8392 53440 8444 53446
rect 8392 53382 8444 53388
rect 8404 52562 8432 53382
rect 8392 52556 8444 52562
rect 8392 52498 8444 52504
rect 8392 52420 8444 52426
rect 8392 52362 8444 52368
rect 8404 52154 8432 52362
rect 8392 52148 8444 52154
rect 8392 52090 8444 52096
rect 8392 51808 8444 51814
rect 8312 51768 8392 51796
rect 8208 51750 8260 51756
rect 8392 51750 8444 51756
rect 8116 51536 8168 51542
rect 8116 51478 8168 51484
rect 8116 51400 8168 51406
rect 8116 51342 8168 51348
rect 7392 50374 7512 50402
rect 7944 50476 8064 50504
rect 7288 48884 7340 48890
rect 7288 48826 7340 48832
rect 7300 48686 7328 48826
rect 7288 48680 7340 48686
rect 7288 48622 7340 48628
rect 7392 48532 7420 50374
rect 7472 50244 7524 50250
rect 7472 50186 7524 50192
rect 7484 50153 7512 50186
rect 7748 50176 7800 50182
rect 7470 50144 7526 50153
rect 7748 50118 7800 50124
rect 7470 50079 7526 50088
rect 7760 49774 7788 50118
rect 7944 49978 7972 50476
rect 8022 50416 8078 50425
rect 8022 50351 8078 50360
rect 7932 49972 7984 49978
rect 7932 49914 7984 49920
rect 7838 49872 7894 49881
rect 7838 49807 7894 49816
rect 7852 49774 7880 49807
rect 7472 49768 7524 49774
rect 7472 49710 7524 49716
rect 7748 49768 7800 49774
rect 7748 49710 7800 49716
rect 7840 49768 7892 49774
rect 7840 49710 7892 49716
rect 7300 48504 7420 48532
rect 7196 48272 7248 48278
rect 7196 48214 7248 48220
rect 7196 48136 7248 48142
rect 7196 48078 7248 48084
rect 7208 47462 7236 48078
rect 7196 47456 7248 47462
rect 7196 47398 7248 47404
rect 7104 45008 7156 45014
rect 6840 44934 7052 44962
rect 7104 44950 7156 44956
rect 6920 44872 6972 44878
rect 6840 44820 6920 44826
rect 6840 44814 6972 44820
rect 6840 44798 6960 44814
rect 6840 43654 6868 44798
rect 7024 44266 7052 44934
rect 7104 44804 7156 44810
rect 7104 44746 7156 44752
rect 7012 44260 7064 44266
rect 7012 44202 7064 44208
rect 6918 44024 6974 44033
rect 7116 43994 7144 44746
rect 7208 44538 7236 47398
rect 7300 47274 7328 48504
rect 7378 48376 7434 48385
rect 7378 48311 7380 48320
rect 7432 48311 7434 48320
rect 7380 48282 7432 48288
rect 7380 48204 7432 48210
rect 7380 48146 7432 48152
rect 7392 47462 7420 48146
rect 7484 48074 7512 49710
rect 7622 49532 7918 49552
rect 7678 49530 7702 49532
rect 7758 49530 7782 49532
rect 7838 49530 7862 49532
rect 7700 49478 7702 49530
rect 7764 49478 7776 49530
rect 7838 49478 7840 49530
rect 7678 49476 7702 49478
rect 7758 49476 7782 49478
rect 7838 49476 7862 49478
rect 7622 49456 7918 49476
rect 7564 49224 7616 49230
rect 7564 49166 7616 49172
rect 7932 49224 7984 49230
rect 7932 49166 7984 49172
rect 7576 48822 7604 49166
rect 7564 48816 7616 48822
rect 7564 48758 7616 48764
rect 7944 48686 7972 49166
rect 7748 48680 7800 48686
rect 7746 48648 7748 48657
rect 7932 48680 7984 48686
rect 7800 48648 7802 48657
rect 7932 48622 7984 48628
rect 7746 48583 7802 48592
rect 7622 48444 7918 48464
rect 7678 48442 7702 48444
rect 7758 48442 7782 48444
rect 7838 48442 7862 48444
rect 7700 48390 7702 48442
rect 7764 48390 7776 48442
rect 7838 48390 7840 48442
rect 7678 48388 7702 48390
rect 7758 48388 7782 48390
rect 7838 48388 7862 48390
rect 7622 48368 7918 48388
rect 7930 48240 7986 48249
rect 7930 48175 7986 48184
rect 7472 48068 7524 48074
rect 7472 48010 7524 48016
rect 7564 48000 7616 48006
rect 7564 47942 7616 47948
rect 7380 47456 7432 47462
rect 7576 47444 7604 47942
rect 7944 47818 7972 48175
rect 8036 48006 8064 50351
rect 8128 49842 8156 51342
rect 8220 51066 8248 51750
rect 8298 51232 8354 51241
rect 8298 51167 8354 51176
rect 8208 51060 8260 51066
rect 8208 51002 8260 51008
rect 8208 50788 8260 50794
rect 8208 50730 8260 50736
rect 8220 50522 8248 50730
rect 8312 50522 8340 51167
rect 8208 50516 8260 50522
rect 8208 50458 8260 50464
rect 8300 50516 8352 50522
rect 8300 50458 8352 50464
rect 8300 50244 8352 50250
rect 8300 50186 8352 50192
rect 8116 49836 8168 49842
rect 8116 49778 8168 49784
rect 8208 49768 8260 49774
rect 8208 49710 8260 49716
rect 8116 49292 8168 49298
rect 8116 49234 8168 49240
rect 8128 48521 8156 49234
rect 8220 49076 8248 49710
rect 8312 49201 8340 50186
rect 8298 49192 8354 49201
rect 8298 49127 8354 49136
rect 8300 49088 8352 49094
rect 8220 49048 8300 49076
rect 8114 48512 8170 48521
rect 8114 48447 8170 48456
rect 8116 48340 8168 48346
rect 8116 48282 8168 48288
rect 8128 48113 8156 48282
rect 8220 48142 8248 49048
rect 8300 49030 8352 49036
rect 8404 48346 8432 51750
rect 8496 50810 8524 59026
rect 8588 58698 8616 59622
rect 8680 59430 8708 60114
rect 8668 59424 8720 59430
rect 8668 59366 8720 59372
rect 8680 59022 8708 59366
rect 8668 59016 8720 59022
rect 8668 58958 8720 58964
rect 8588 58670 8708 58698
rect 8574 58576 8630 58585
rect 8574 58511 8630 58520
rect 8588 58478 8616 58511
rect 8576 58472 8628 58478
rect 8576 58414 8628 58420
rect 8588 58070 8616 58414
rect 8576 58064 8628 58070
rect 8576 58006 8628 58012
rect 8576 57792 8628 57798
rect 8576 57734 8628 57740
rect 8588 56982 8616 57734
rect 8576 56976 8628 56982
rect 8576 56918 8628 56924
rect 8576 56704 8628 56710
rect 8576 56646 8628 56652
rect 8588 54534 8616 56646
rect 8680 56506 8708 58670
rect 8668 56500 8720 56506
rect 8668 56442 8720 56448
rect 8668 55276 8720 55282
rect 8668 55218 8720 55224
rect 8576 54528 8628 54534
rect 8576 54470 8628 54476
rect 8576 53984 8628 53990
rect 8576 53926 8628 53932
rect 8588 50930 8616 53926
rect 8680 53786 8708 55218
rect 8668 53780 8720 53786
rect 8668 53722 8720 53728
rect 8668 53644 8720 53650
rect 8668 53586 8720 53592
rect 8680 53242 8708 53586
rect 8668 53236 8720 53242
rect 8668 53178 8720 53184
rect 8680 51542 8708 53178
rect 8772 52426 8800 61118
rect 8864 57882 8892 64874
rect 8956 62354 8984 64942
rect 9048 63374 9076 68734
rect 9220 68672 9272 68678
rect 9220 68614 9272 68620
rect 9128 66700 9180 66706
rect 9128 66642 9180 66648
rect 9140 65958 9168 66642
rect 9232 66570 9260 68614
rect 9220 66564 9272 66570
rect 9220 66506 9272 66512
rect 9220 66224 9272 66230
rect 9220 66166 9272 66172
rect 9232 65958 9260 66166
rect 9128 65952 9180 65958
rect 9128 65894 9180 65900
rect 9220 65952 9272 65958
rect 9220 65894 9272 65900
rect 9140 65793 9168 65894
rect 9126 65784 9182 65793
rect 9126 65719 9182 65728
rect 9128 65680 9180 65686
rect 9128 65622 9180 65628
rect 9140 64025 9168 65622
rect 9126 64016 9182 64025
rect 9126 63951 9182 63960
rect 9126 63880 9182 63889
rect 9126 63815 9182 63824
rect 9036 63368 9088 63374
rect 9036 63310 9088 63316
rect 9048 62966 9076 63310
rect 9036 62960 9088 62966
rect 9036 62902 9088 62908
rect 8944 62348 8996 62354
rect 8944 62290 8996 62296
rect 8956 61878 8984 62290
rect 9140 62098 9168 63815
rect 9232 63481 9260 65894
rect 9416 65657 9444 69119
rect 9508 68950 9536 69158
rect 9496 68944 9548 68950
rect 9496 68886 9548 68892
rect 9508 68134 9536 68886
rect 9496 68128 9548 68134
rect 9692 68116 9720 69226
rect 9784 68218 9812 69255
rect 9876 68678 9904 69770
rect 9968 69358 9996 69974
rect 9956 69352 10008 69358
rect 9956 69294 10008 69300
rect 9968 68746 9996 69294
rect 10060 68921 10088 72490
rect 10336 72185 10364 72626
rect 10508 72480 10560 72486
rect 10508 72422 10560 72428
rect 10322 72176 10378 72185
rect 10322 72111 10378 72120
rect 10520 71482 10548 72422
rect 10612 71602 10640 73646
rect 10704 73273 10732 73714
rect 11336 73704 11388 73710
rect 11336 73646 11388 73652
rect 10690 73264 10746 73273
rect 10690 73199 10746 73208
rect 10876 73024 10928 73030
rect 10876 72966 10928 72972
rect 10888 72758 10916 72966
rect 10956 72924 11252 72944
rect 11012 72922 11036 72924
rect 11092 72922 11116 72924
rect 11172 72922 11196 72924
rect 11034 72870 11036 72922
rect 11098 72870 11110 72922
rect 11172 72870 11174 72922
rect 11012 72868 11036 72870
rect 11092 72868 11116 72870
rect 11172 72868 11196 72870
rect 10956 72848 11252 72868
rect 11348 72758 11376 73646
rect 14289 73468 14585 73488
rect 14345 73466 14369 73468
rect 14425 73466 14449 73468
rect 14505 73466 14529 73468
rect 14367 73414 14369 73466
rect 14431 73414 14443 73466
rect 14505 73414 14507 73466
rect 14345 73412 14369 73414
rect 14425 73412 14449 73414
rect 14505 73412 14529 73414
rect 14289 73392 14585 73412
rect 11612 73160 11664 73166
rect 11612 73102 11664 73108
rect 10876 72752 10928 72758
rect 10876 72694 10928 72700
rect 11336 72752 11388 72758
rect 11336 72694 11388 72700
rect 10888 72622 10916 72694
rect 11624 72622 11652 73102
rect 17622 72924 17918 72944
rect 17678 72922 17702 72924
rect 17758 72922 17782 72924
rect 17838 72922 17862 72924
rect 17700 72870 17702 72922
rect 17764 72870 17776 72922
rect 17838 72870 17840 72922
rect 17678 72868 17702 72870
rect 17758 72868 17782 72870
rect 17838 72868 17862 72870
rect 17622 72848 17918 72868
rect 16302 72720 16358 72729
rect 16302 72655 16358 72664
rect 10876 72616 10928 72622
rect 10876 72558 10928 72564
rect 11612 72616 11664 72622
rect 11796 72616 11848 72622
rect 11612 72558 11664 72564
rect 11794 72584 11796 72593
rect 11980 72616 12032 72622
rect 11848 72584 11850 72593
rect 10600 71596 10652 71602
rect 10600 71538 10652 71544
rect 10520 71454 10640 71482
rect 10140 70848 10192 70854
rect 10140 70790 10192 70796
rect 10232 70848 10284 70854
rect 10232 70790 10284 70796
rect 10152 70446 10180 70790
rect 10244 70514 10272 70790
rect 10324 70644 10376 70650
rect 10324 70586 10376 70592
rect 10232 70508 10284 70514
rect 10232 70450 10284 70456
rect 10140 70440 10192 70446
rect 10336 70394 10364 70586
rect 10140 70382 10192 70388
rect 10244 70366 10364 70394
rect 10416 70440 10468 70446
rect 10416 70382 10468 70388
rect 10140 70304 10192 70310
rect 10140 70246 10192 70252
rect 10152 69970 10180 70246
rect 10140 69964 10192 69970
rect 10140 69906 10192 69912
rect 10140 69352 10192 69358
rect 10140 69294 10192 69300
rect 10046 68912 10102 68921
rect 10046 68847 10102 68856
rect 10060 68814 10088 68847
rect 10048 68808 10100 68814
rect 10048 68750 10100 68756
rect 9956 68740 10008 68746
rect 9956 68682 10008 68688
rect 9864 68672 9916 68678
rect 9864 68614 9916 68620
rect 9968 68406 9996 68682
rect 9956 68400 10008 68406
rect 9956 68342 10008 68348
rect 9784 68190 9996 68218
rect 10152 68202 10180 69294
rect 9772 68128 9824 68134
rect 9692 68088 9772 68116
rect 9496 68070 9548 68076
rect 9772 68070 9824 68076
rect 9508 67046 9536 68070
rect 9680 67176 9732 67182
rect 9678 67144 9680 67153
rect 9732 67144 9734 67153
rect 9678 67079 9734 67088
rect 9496 67040 9548 67046
rect 9496 66982 9548 66988
rect 9508 66298 9536 66982
rect 9692 66842 9720 67079
rect 9680 66836 9732 66842
rect 9680 66778 9732 66784
rect 9784 66722 9812 68070
rect 9864 67584 9916 67590
rect 9864 67526 9916 67532
rect 9600 66706 9812 66722
rect 9876 66706 9904 67526
rect 9588 66700 9812 66706
rect 9640 66694 9812 66700
rect 9588 66642 9640 66648
rect 9680 66632 9732 66638
rect 9680 66574 9732 66580
rect 9496 66292 9548 66298
rect 9496 66234 9548 66240
rect 9588 66088 9640 66094
rect 9692 66076 9720 66574
rect 9640 66048 9720 66076
rect 9588 66030 9640 66036
rect 9402 65648 9458 65657
rect 9402 65583 9458 65592
rect 9312 64320 9364 64326
rect 9312 64262 9364 64268
rect 9324 64054 9352 64262
rect 9312 64048 9364 64054
rect 9312 63990 9364 63996
rect 9218 63472 9274 63481
rect 9218 63407 9274 63416
rect 9220 63300 9272 63306
rect 9220 63242 9272 63248
rect 9232 62257 9260 63242
rect 9218 62248 9274 62257
rect 9218 62183 9274 62192
rect 9140 62070 9260 62098
rect 8944 61872 8996 61878
rect 8944 61814 8996 61820
rect 9128 61804 9180 61810
rect 9128 61746 9180 61752
rect 9036 61192 9088 61198
rect 9036 61134 9088 61140
rect 8944 60716 8996 60722
rect 8944 60658 8996 60664
rect 8956 59498 8984 60658
rect 9048 60602 9076 61134
rect 9140 60722 9168 61746
rect 9128 60716 9180 60722
rect 9128 60658 9180 60664
rect 9048 60574 9168 60602
rect 9140 60518 9168 60574
rect 9128 60512 9180 60518
rect 9128 60454 9180 60460
rect 9034 59800 9090 59809
rect 9034 59735 9036 59744
rect 9088 59735 9090 59744
rect 9036 59706 9088 59712
rect 8944 59492 8996 59498
rect 8944 59434 8996 59440
rect 9140 59090 9168 60454
rect 9128 59084 9180 59090
rect 9128 59026 9180 59032
rect 9140 58342 9168 59026
rect 9128 58336 9180 58342
rect 9128 58278 9180 58284
rect 8864 57854 9076 57882
rect 9048 57798 9076 57854
rect 9036 57792 9088 57798
rect 9036 57734 9088 57740
rect 8852 56908 8904 56914
rect 8852 56850 8904 56856
rect 8864 55962 8892 56850
rect 8944 56160 8996 56166
rect 8944 56102 8996 56108
rect 8852 55956 8904 55962
rect 8852 55898 8904 55904
rect 8864 55865 8892 55898
rect 8850 55856 8906 55865
rect 8850 55791 8906 55800
rect 8852 55684 8904 55690
rect 8852 55626 8904 55632
rect 8864 55418 8892 55626
rect 8852 55412 8904 55418
rect 8852 55354 8904 55360
rect 8864 55282 8892 55354
rect 8852 55276 8904 55282
rect 8852 55218 8904 55224
rect 8850 55040 8906 55049
rect 8850 54975 8906 54984
rect 8864 54738 8892 54975
rect 8852 54732 8904 54738
rect 8852 54674 8904 54680
rect 8850 53680 8906 53689
rect 8850 53615 8852 53624
rect 8904 53615 8906 53624
rect 8852 53586 8904 53592
rect 8864 53242 8892 53586
rect 8852 53236 8904 53242
rect 8852 53178 8904 53184
rect 8852 52556 8904 52562
rect 8852 52498 8904 52504
rect 8760 52420 8812 52426
rect 8760 52362 8812 52368
rect 8864 52306 8892 52498
rect 8772 52278 8892 52306
rect 8772 52086 8800 52278
rect 8852 52148 8904 52154
rect 8852 52090 8904 52096
rect 8760 52080 8812 52086
rect 8760 52022 8812 52028
rect 8668 51536 8720 51542
rect 8668 51478 8720 51484
rect 8772 51388 8800 52022
rect 8680 51360 8800 51388
rect 8576 50924 8628 50930
rect 8576 50866 8628 50872
rect 8496 50782 8616 50810
rect 8484 50720 8536 50726
rect 8484 50662 8536 50668
rect 8496 49910 8524 50662
rect 8588 50017 8616 50782
rect 8574 50008 8630 50017
rect 8574 49943 8630 49952
rect 8484 49904 8536 49910
rect 8484 49846 8536 49852
rect 8576 49904 8628 49910
rect 8576 49846 8628 49852
rect 8484 49768 8536 49774
rect 8484 49710 8536 49716
rect 8392 48340 8444 48346
rect 8392 48282 8444 48288
rect 8392 48204 8444 48210
rect 8392 48146 8444 48152
rect 8208 48136 8260 48142
rect 8114 48104 8170 48113
rect 8208 48078 8260 48084
rect 8114 48039 8170 48048
rect 8024 48000 8076 48006
rect 8300 48000 8352 48006
rect 8024 47942 8076 47948
rect 8114 47968 8170 47977
rect 8300 47942 8352 47948
rect 8114 47903 8170 47912
rect 7944 47790 8064 47818
rect 7380 47398 7432 47404
rect 7484 47416 7604 47444
rect 7300 47246 7420 47274
rect 7288 46028 7340 46034
rect 7288 45970 7340 45976
rect 7300 45830 7328 45970
rect 7288 45824 7340 45830
rect 7288 45766 7340 45772
rect 7300 44878 7328 45766
rect 7288 44872 7340 44878
rect 7288 44814 7340 44820
rect 7196 44532 7248 44538
rect 7196 44474 7248 44480
rect 7392 44470 7420 47246
rect 7380 44464 7432 44470
rect 7380 44406 7432 44412
rect 7484 44248 7512 47416
rect 7622 47356 7918 47376
rect 7678 47354 7702 47356
rect 7758 47354 7782 47356
rect 7838 47354 7862 47356
rect 7700 47302 7702 47354
rect 7764 47302 7776 47354
rect 7838 47302 7840 47354
rect 7678 47300 7702 47302
rect 7758 47300 7782 47302
rect 7838 47300 7862 47302
rect 7622 47280 7918 47300
rect 7748 46980 7800 46986
rect 7748 46922 7800 46928
rect 7760 46714 7788 46922
rect 7748 46708 7800 46714
rect 7748 46650 7800 46656
rect 7622 46268 7918 46288
rect 7678 46266 7702 46268
rect 7758 46266 7782 46268
rect 7838 46266 7862 46268
rect 7700 46214 7702 46266
rect 7764 46214 7776 46266
rect 7838 46214 7840 46266
rect 7678 46212 7702 46214
rect 7758 46212 7782 46214
rect 7838 46212 7862 46214
rect 7622 46192 7918 46212
rect 8036 46152 8064 47790
rect 7944 46124 8064 46152
rect 7944 45665 7972 46124
rect 8128 46034 8156 47903
rect 8312 47598 8340 47942
rect 8300 47592 8352 47598
rect 8300 47534 8352 47540
rect 8208 47456 8260 47462
rect 8208 47398 8260 47404
rect 8024 46028 8076 46034
rect 8024 45970 8076 45976
rect 8116 46028 8168 46034
rect 8116 45970 8168 45976
rect 7930 45656 7986 45665
rect 8036 45626 8064 45970
rect 7930 45591 7986 45600
rect 8024 45620 8076 45626
rect 8024 45562 8076 45568
rect 8024 45280 8076 45286
rect 8024 45222 8076 45228
rect 7622 45180 7918 45200
rect 7678 45178 7702 45180
rect 7758 45178 7782 45180
rect 7838 45178 7862 45180
rect 7700 45126 7702 45178
rect 7764 45126 7776 45178
rect 7838 45126 7840 45178
rect 7678 45124 7702 45126
rect 7758 45124 7782 45126
rect 7838 45124 7862 45126
rect 7622 45104 7918 45124
rect 7562 44976 7618 44985
rect 7562 44911 7618 44920
rect 7392 44220 7512 44248
rect 6918 43959 6974 43968
rect 7104 43988 7156 43994
rect 6932 43874 6960 43959
rect 7104 43930 7156 43936
rect 6932 43858 7052 43874
rect 6920 43852 7052 43858
rect 6972 43846 7052 43852
rect 6920 43794 6972 43800
rect 7024 43761 7052 43846
rect 7104 43852 7156 43858
rect 7104 43794 7156 43800
rect 7010 43752 7066 43761
rect 6920 43716 6972 43722
rect 7010 43687 7066 43696
rect 6920 43658 6972 43664
rect 6828 43648 6880 43654
rect 6828 43590 6880 43596
rect 6932 42265 6960 43658
rect 7024 43450 7052 43687
rect 7012 43444 7064 43450
rect 7012 43386 7064 43392
rect 7012 42560 7064 42566
rect 7116 42548 7144 43794
rect 7288 43376 7340 43382
rect 7288 43318 7340 43324
rect 7196 43240 7248 43246
rect 7196 43182 7248 43188
rect 7208 42838 7236 43182
rect 7196 42832 7248 42838
rect 7196 42774 7248 42780
rect 7064 42520 7144 42548
rect 7012 42502 7064 42508
rect 6918 42256 6974 42265
rect 6918 42191 6974 42200
rect 6918 42120 6974 42129
rect 6918 42055 6974 42064
rect 6828 41472 6880 41478
rect 6932 41460 6960 42055
rect 7024 41750 7052 42502
rect 7208 41818 7236 42774
rect 7196 41812 7248 41818
rect 7196 41754 7248 41760
rect 7012 41744 7064 41750
rect 7012 41686 7064 41692
rect 7104 41676 7156 41682
rect 7104 41618 7156 41624
rect 7116 41585 7144 41618
rect 7300 41596 7328 43318
rect 7102 41576 7158 41585
rect 7102 41511 7158 41520
rect 7208 41568 7328 41596
rect 6932 41432 7144 41460
rect 6828 41414 6880 41420
rect 6840 41206 6868 41414
rect 7010 41304 7066 41313
rect 7010 41239 7012 41248
rect 7064 41239 7066 41248
rect 7012 41210 7064 41216
rect 6828 41200 6880 41206
rect 6828 41142 6880 41148
rect 6920 41064 6972 41070
rect 6748 41024 6920 41052
rect 6920 41006 6972 41012
rect 6932 40730 6960 41006
rect 7012 40928 7064 40934
rect 7012 40870 7064 40876
rect 6920 40724 6972 40730
rect 6920 40666 6972 40672
rect 6932 40576 6960 40666
rect 6840 40548 6960 40576
rect 6656 39902 6776 39930
rect 6644 39840 6696 39846
rect 6644 39782 6696 39788
rect 6656 39302 6684 39782
rect 6644 39296 6696 39302
rect 6644 39238 6696 39244
rect 6552 33448 6604 33454
rect 6552 33390 6604 33396
rect 6564 33114 6592 33390
rect 6552 33108 6604 33114
rect 6552 33050 6604 33056
rect 6656 32994 6684 39238
rect 6748 38826 6776 39902
rect 6736 38820 6788 38826
rect 6736 38762 6788 38768
rect 6840 38554 6868 40548
rect 6920 40452 6972 40458
rect 6920 40394 6972 40400
rect 6932 40050 6960 40394
rect 6920 40044 6972 40050
rect 6920 39986 6972 39992
rect 6920 39908 6972 39914
rect 6920 39850 6972 39856
rect 6932 39098 6960 39850
rect 6920 39092 6972 39098
rect 6920 39034 6972 39040
rect 6828 38548 6880 38554
rect 6880 38508 6960 38536
rect 6828 38490 6880 38496
rect 6828 38412 6880 38418
rect 6828 38354 6880 38360
rect 6736 37800 6788 37806
rect 6734 37768 6736 37777
rect 6788 37768 6790 37777
rect 6840 37738 6868 38354
rect 6932 37806 6960 38508
rect 6920 37800 6972 37806
rect 6920 37742 6972 37748
rect 6734 37703 6790 37712
rect 6828 37732 6880 37738
rect 6748 37398 6776 37703
rect 6828 37674 6880 37680
rect 6736 37392 6788 37398
rect 6736 37334 6788 37340
rect 6840 37330 6868 37674
rect 6932 37466 6960 37742
rect 7024 37670 7052 40870
rect 7012 37664 7064 37670
rect 7012 37606 7064 37612
rect 6920 37460 6972 37466
rect 6920 37402 6972 37408
rect 7116 37346 7144 41432
rect 7208 39982 7236 41568
rect 7286 41032 7342 41041
rect 7286 40967 7342 40976
rect 7196 39976 7248 39982
rect 7196 39918 7248 39924
rect 7208 39642 7236 39918
rect 7196 39636 7248 39642
rect 7196 39578 7248 39584
rect 6828 37324 6880 37330
rect 6828 37266 6880 37272
rect 6920 37324 6972 37330
rect 6920 37266 6972 37272
rect 7024 37318 7144 37346
rect 7208 37330 7236 39578
rect 7300 38185 7328 40967
rect 7286 38176 7342 38185
rect 7286 38111 7342 38120
rect 7392 38026 7420 44220
rect 7576 44180 7604 44911
rect 8036 44402 8064 45222
rect 8128 45082 8156 45970
rect 8116 45076 8168 45082
rect 8116 45018 8168 45024
rect 8116 44532 8168 44538
rect 8116 44474 8168 44480
rect 8024 44396 8076 44402
rect 8024 44338 8076 44344
rect 8128 44334 8156 44474
rect 8116 44328 8168 44334
rect 8116 44270 8168 44276
rect 8024 44260 8076 44266
rect 8024 44202 8076 44208
rect 7484 44152 7604 44180
rect 7484 43858 7512 44152
rect 7622 44092 7918 44112
rect 7678 44090 7702 44092
rect 7758 44090 7782 44092
rect 7838 44090 7862 44092
rect 7700 44038 7702 44090
rect 7764 44038 7776 44090
rect 7838 44038 7840 44090
rect 7678 44036 7702 44038
rect 7758 44036 7782 44038
rect 7838 44036 7862 44038
rect 7622 44016 7918 44036
rect 7472 43852 7524 43858
rect 7472 43794 7524 43800
rect 7484 43450 7512 43794
rect 7472 43444 7524 43450
rect 7472 43386 7524 43392
rect 7622 43004 7918 43024
rect 7678 43002 7702 43004
rect 7758 43002 7782 43004
rect 7838 43002 7862 43004
rect 7700 42950 7702 43002
rect 7764 42950 7776 43002
rect 7838 42950 7840 43002
rect 7678 42948 7702 42950
rect 7758 42948 7782 42950
rect 7838 42948 7862 42950
rect 7622 42928 7918 42948
rect 7932 42832 7984 42838
rect 7932 42774 7984 42780
rect 7562 42664 7618 42673
rect 7562 42599 7618 42608
rect 7576 42294 7604 42599
rect 7748 42560 7800 42566
rect 7748 42502 7800 42508
rect 7564 42288 7616 42294
rect 7760 42265 7788 42502
rect 7564 42230 7616 42236
rect 7746 42256 7802 42265
rect 7746 42191 7748 42200
rect 7800 42191 7802 42200
rect 7748 42162 7800 42168
rect 7944 42090 7972 42774
rect 7472 42084 7524 42090
rect 7472 42026 7524 42032
rect 7932 42084 7984 42090
rect 7932 42026 7984 42032
rect 7484 41206 7512 42026
rect 7622 41916 7918 41936
rect 7678 41914 7702 41916
rect 7758 41914 7782 41916
rect 7838 41914 7862 41916
rect 7700 41862 7702 41914
rect 7764 41862 7776 41914
rect 7838 41862 7840 41914
rect 7678 41860 7702 41862
rect 7758 41860 7782 41862
rect 7838 41860 7862 41862
rect 7622 41840 7918 41860
rect 7472 41200 7524 41206
rect 7472 41142 7524 41148
rect 7470 41032 7526 41041
rect 7470 40967 7526 40976
rect 7484 40730 7512 40967
rect 7622 40828 7918 40848
rect 7678 40826 7702 40828
rect 7758 40826 7782 40828
rect 7838 40826 7862 40828
rect 7700 40774 7702 40826
rect 7764 40774 7776 40826
rect 7838 40774 7840 40826
rect 7678 40772 7702 40774
rect 7758 40772 7782 40774
rect 7838 40772 7862 40774
rect 7622 40752 7918 40772
rect 7472 40724 7524 40730
rect 7472 40666 7524 40672
rect 7472 40588 7524 40594
rect 7472 40530 7524 40536
rect 7484 40118 7512 40530
rect 7472 40112 7524 40118
rect 7472 40054 7524 40060
rect 7622 39740 7918 39760
rect 7678 39738 7702 39740
rect 7758 39738 7782 39740
rect 7838 39738 7862 39740
rect 7700 39686 7702 39738
rect 7764 39686 7776 39738
rect 7838 39686 7840 39738
rect 7678 39684 7702 39686
rect 7758 39684 7782 39686
rect 7838 39684 7862 39686
rect 7622 39664 7918 39684
rect 7656 39500 7708 39506
rect 7656 39442 7708 39448
rect 7564 39432 7616 39438
rect 7562 39400 7564 39409
rect 7616 39400 7618 39409
rect 7562 39335 7618 39344
rect 7668 39001 7696 39442
rect 7654 38992 7710 39001
rect 7654 38927 7710 38936
rect 7472 38888 7524 38894
rect 7472 38830 7524 38836
rect 7300 37998 7420 38026
rect 7196 37324 7248 37330
rect 6734 37088 6790 37097
rect 6734 37023 6790 37032
rect 6748 36378 6776 37023
rect 6840 36582 6868 37266
rect 6828 36576 6880 36582
rect 6828 36518 6880 36524
rect 6826 36408 6882 36417
rect 6736 36372 6788 36378
rect 6826 36343 6882 36352
rect 6736 36314 6788 36320
rect 6840 35630 6868 36343
rect 6828 35624 6880 35630
rect 6828 35566 6880 35572
rect 6932 35154 6960 37266
rect 7024 36666 7052 37318
rect 7196 37266 7248 37272
rect 7024 36638 7144 36666
rect 7012 36576 7064 36582
rect 7012 36518 7064 36524
rect 6920 35148 6972 35154
rect 6920 35090 6972 35096
rect 6736 34944 6788 34950
rect 6736 34886 6788 34892
rect 6748 34542 6776 34886
rect 6736 34536 6788 34542
rect 6736 34478 6788 34484
rect 6748 34105 6776 34478
rect 6828 34468 6880 34474
rect 6828 34410 6880 34416
rect 6734 34096 6790 34105
rect 6840 34066 6868 34410
rect 6932 34202 6960 35090
rect 6920 34196 6972 34202
rect 6920 34138 6972 34144
rect 6734 34031 6790 34040
rect 6828 34060 6880 34066
rect 6828 34002 6880 34008
rect 6736 33924 6788 33930
rect 6736 33866 6788 33872
rect 6564 32966 6684 32994
rect 6564 31482 6592 32966
rect 6644 32020 6696 32026
rect 6644 31962 6696 31968
rect 6552 31476 6604 31482
rect 6552 31418 6604 31424
rect 6564 30938 6592 31418
rect 6552 30932 6604 30938
rect 6552 30874 6604 30880
rect 6552 30048 6604 30054
rect 6552 29990 6604 29996
rect 6564 29034 6592 29990
rect 6552 29028 6604 29034
rect 6552 28970 6604 28976
rect 6460 26580 6512 26586
rect 6460 26522 6512 26528
rect 6472 25906 6500 26522
rect 6460 25900 6512 25906
rect 6460 25842 6512 25848
rect 6368 25832 6420 25838
rect 6368 25774 6420 25780
rect 6380 25226 6408 25774
rect 6564 25498 6592 28970
rect 6552 25492 6604 25498
rect 6552 25434 6604 25440
rect 6656 25294 6684 31962
rect 6748 28762 6776 33866
rect 6840 33833 6868 34002
rect 6826 33824 6882 33833
rect 6826 33759 6882 33768
rect 6826 33688 6882 33697
rect 6826 33623 6828 33632
rect 6880 33623 6882 33632
rect 6828 33594 6880 33600
rect 6920 33312 6972 33318
rect 6920 33254 6972 33260
rect 6932 33130 6960 33254
rect 6840 33114 6960 33130
rect 6828 33108 6960 33114
rect 6880 33102 6960 33108
rect 6828 33050 6880 33056
rect 6826 33008 6882 33017
rect 6826 32943 6882 32952
rect 6840 32337 6868 32943
rect 6826 32328 6882 32337
rect 6826 32263 6882 32272
rect 6840 31793 6868 32263
rect 6826 31784 6882 31793
rect 6826 31719 6882 31728
rect 6932 30326 6960 33102
rect 6920 30320 6972 30326
rect 6920 30262 6972 30268
rect 6932 30190 6960 30262
rect 6920 30184 6972 30190
rect 6920 30126 6972 30132
rect 6828 29708 6880 29714
rect 6828 29650 6880 29656
rect 6840 29170 6868 29650
rect 6828 29164 6880 29170
rect 6828 29106 6880 29112
rect 6736 28756 6788 28762
rect 6736 28698 6788 28704
rect 6748 28082 6776 28698
rect 7024 28626 7052 36518
rect 7116 28762 7144 36638
rect 7300 36242 7328 37998
rect 7484 37942 7512 38830
rect 7668 38826 7696 38927
rect 7656 38820 7708 38826
rect 7656 38762 7708 38768
rect 7622 38652 7918 38672
rect 7678 38650 7702 38652
rect 7758 38650 7782 38652
rect 7838 38650 7862 38652
rect 7700 38598 7702 38650
rect 7764 38598 7776 38650
rect 7838 38598 7840 38650
rect 7678 38596 7702 38598
rect 7758 38596 7782 38598
rect 7838 38596 7862 38598
rect 7622 38576 7918 38596
rect 7380 37936 7432 37942
rect 7380 37878 7432 37884
rect 7472 37936 7524 37942
rect 7472 37878 7524 37884
rect 7392 37369 7420 37878
rect 7472 37800 7524 37806
rect 7472 37742 7524 37748
rect 7484 37670 7512 37742
rect 7472 37664 7524 37670
rect 7472 37606 7524 37612
rect 7378 37360 7434 37369
rect 7378 37295 7434 37304
rect 7380 37256 7432 37262
rect 7380 37198 7432 37204
rect 7392 36258 7420 37198
rect 7484 36718 7512 37606
rect 7622 37564 7918 37584
rect 7678 37562 7702 37564
rect 7758 37562 7782 37564
rect 7838 37562 7862 37564
rect 7700 37510 7702 37562
rect 7764 37510 7776 37562
rect 7838 37510 7840 37562
rect 7678 37508 7702 37510
rect 7758 37508 7782 37510
rect 7838 37508 7862 37510
rect 7622 37488 7918 37508
rect 7930 37088 7986 37097
rect 7930 37023 7986 37032
rect 7944 36718 7972 37023
rect 7472 36712 7524 36718
rect 7472 36654 7524 36660
rect 7932 36712 7984 36718
rect 7932 36654 7984 36660
rect 7622 36476 7918 36496
rect 7678 36474 7702 36476
rect 7758 36474 7782 36476
rect 7838 36474 7862 36476
rect 7700 36422 7702 36474
rect 7764 36422 7776 36474
rect 7838 36422 7840 36474
rect 7678 36420 7702 36422
rect 7758 36420 7782 36422
rect 7838 36420 7862 36422
rect 7622 36400 7918 36420
rect 7196 36236 7248 36242
rect 7196 36178 7248 36184
rect 7288 36236 7340 36242
rect 7392 36230 7512 36258
rect 7288 36178 7340 36184
rect 7208 35494 7236 36178
rect 7300 35834 7328 36178
rect 7288 35828 7340 35834
rect 7340 35788 7420 35816
rect 7288 35770 7340 35776
rect 7196 35488 7248 35494
rect 7196 35430 7248 35436
rect 7208 30190 7236 35430
rect 7288 35080 7340 35086
rect 7288 35022 7340 35028
rect 7300 34066 7328 35022
rect 7288 34060 7340 34066
rect 7288 34002 7340 34008
rect 7300 33114 7328 34002
rect 7288 33108 7340 33114
rect 7288 33050 7340 33056
rect 7392 32745 7420 35788
rect 7484 34513 7512 36230
rect 7622 35388 7918 35408
rect 7678 35386 7702 35388
rect 7758 35386 7782 35388
rect 7838 35386 7862 35388
rect 7700 35334 7702 35386
rect 7764 35334 7776 35386
rect 7838 35334 7840 35386
rect 7678 35332 7702 35334
rect 7758 35332 7782 35334
rect 7838 35332 7862 35334
rect 7622 35312 7918 35332
rect 7932 34740 7984 34746
rect 7932 34682 7984 34688
rect 7944 34649 7972 34682
rect 7930 34640 7986 34649
rect 7930 34575 7986 34584
rect 7944 34542 7972 34575
rect 7932 34536 7984 34542
rect 7470 34504 7526 34513
rect 7932 34478 7984 34484
rect 7470 34439 7526 34448
rect 7472 34400 7524 34406
rect 7472 34342 7524 34348
rect 7484 34066 7512 34342
rect 7622 34300 7918 34320
rect 7678 34298 7702 34300
rect 7758 34298 7782 34300
rect 7838 34298 7862 34300
rect 7700 34246 7702 34298
rect 7764 34246 7776 34298
rect 7838 34246 7840 34298
rect 7678 34244 7702 34246
rect 7758 34244 7782 34246
rect 7838 34244 7862 34246
rect 7622 34224 7918 34244
rect 7472 34060 7524 34066
rect 7472 34002 7524 34008
rect 7484 33114 7512 34002
rect 7622 33212 7918 33232
rect 7678 33210 7702 33212
rect 7758 33210 7782 33212
rect 7838 33210 7862 33212
rect 7700 33158 7702 33210
rect 7764 33158 7776 33210
rect 7838 33158 7840 33210
rect 7678 33156 7702 33158
rect 7758 33156 7782 33158
rect 7838 33156 7862 33158
rect 7622 33136 7918 33156
rect 7472 33108 7524 33114
rect 7472 33050 7524 33056
rect 7378 32736 7434 32745
rect 8036 32722 8064 44202
rect 8128 42838 8156 44270
rect 8116 42832 8168 42838
rect 8116 42774 8168 42780
rect 8116 42560 8168 42566
rect 8116 42502 8168 42508
rect 8128 41682 8156 42502
rect 8116 41676 8168 41682
rect 8116 41618 8168 41624
rect 8116 40928 8168 40934
rect 8116 40870 8168 40876
rect 8128 40662 8156 40870
rect 8116 40656 8168 40662
rect 8116 40598 8168 40604
rect 8114 39672 8170 39681
rect 8114 39607 8170 39616
rect 8128 39574 8156 39607
rect 8116 39568 8168 39574
rect 8116 39510 8168 39516
rect 8116 38820 8168 38826
rect 8116 38762 8168 38768
rect 8128 38554 8156 38762
rect 8116 38548 8168 38554
rect 8116 38490 8168 38496
rect 8116 37936 8168 37942
rect 8116 37878 8168 37884
rect 8128 37126 8156 37878
rect 8116 37120 8168 37126
rect 8116 37062 8168 37068
rect 8116 36712 8168 36718
rect 8116 36654 8168 36660
rect 8128 36310 8156 36654
rect 8116 36304 8168 36310
rect 8116 36246 8168 36252
rect 8036 32694 8156 32722
rect 7378 32671 7434 32680
rect 8022 32600 8078 32609
rect 8022 32535 8024 32544
rect 8076 32535 8078 32544
rect 8024 32506 8076 32512
rect 8036 32366 8064 32506
rect 8024 32360 8076 32366
rect 8024 32302 8076 32308
rect 7622 32124 7918 32144
rect 7678 32122 7702 32124
rect 7758 32122 7782 32124
rect 7838 32122 7862 32124
rect 7700 32070 7702 32122
rect 7764 32070 7776 32122
rect 7838 32070 7840 32122
rect 7678 32068 7702 32070
rect 7758 32068 7782 32070
rect 7838 32068 7862 32070
rect 7622 32048 7918 32068
rect 7288 32020 7340 32026
rect 8036 32008 8064 32302
rect 7288 31962 7340 31968
rect 7944 31980 8064 32008
rect 7196 30184 7248 30190
rect 7196 30126 7248 30132
rect 7208 29306 7236 30126
rect 7196 29300 7248 29306
rect 7196 29242 7248 29248
rect 7194 29200 7250 29209
rect 7194 29135 7250 29144
rect 7104 28756 7156 28762
rect 7104 28698 7156 28704
rect 7012 28620 7064 28626
rect 7012 28562 7064 28568
rect 6736 28076 6788 28082
rect 6736 28018 6788 28024
rect 7024 27674 7052 28562
rect 7012 27668 7064 27674
rect 7012 27610 7064 27616
rect 7116 27606 7144 28698
rect 7104 27600 7156 27606
rect 7104 27542 7156 27548
rect 7116 26858 7144 27542
rect 7104 26852 7156 26858
rect 7104 26794 7156 26800
rect 7104 26444 7156 26450
rect 7104 26386 7156 26392
rect 7116 26042 7144 26386
rect 7104 26036 7156 26042
rect 7104 25978 7156 25984
rect 7104 25424 7156 25430
rect 7104 25366 7156 25372
rect 6644 25288 6696 25294
rect 6644 25230 6696 25236
rect 6368 25220 6420 25226
rect 6368 25162 6420 25168
rect 6656 24750 6684 25230
rect 6644 24744 6696 24750
rect 6644 24686 6696 24692
rect 6368 24608 6420 24614
rect 6368 24550 6420 24556
rect 6184 22228 6236 22234
rect 6184 22170 6236 22176
rect 6380 22030 6408 24550
rect 6552 24404 6604 24410
rect 6552 24346 6604 24352
rect 6564 23662 6592 24346
rect 6656 24342 6684 24686
rect 7012 24676 7064 24682
rect 7012 24618 7064 24624
rect 7024 24449 7052 24618
rect 7010 24440 7066 24449
rect 7116 24410 7144 25366
rect 7208 24750 7236 29135
rect 7196 24744 7248 24750
rect 7196 24686 7248 24692
rect 7010 24375 7066 24384
rect 7104 24404 7156 24410
rect 7104 24346 7156 24352
rect 6644 24336 6696 24342
rect 6644 24278 6696 24284
rect 7012 24268 7064 24274
rect 7012 24210 7064 24216
rect 6644 24064 6696 24070
rect 6642 24032 6644 24041
rect 6696 24032 6698 24041
rect 6642 23967 6698 23976
rect 7024 23730 7052 24210
rect 7300 23746 7328 31962
rect 7472 31816 7524 31822
rect 7472 31758 7524 31764
rect 7484 31482 7512 31758
rect 7472 31476 7524 31482
rect 7472 31418 7524 31424
rect 7944 31278 7972 31980
rect 8024 31884 8076 31890
rect 8024 31826 8076 31832
rect 8036 31414 8064 31826
rect 8024 31408 8076 31414
rect 8024 31350 8076 31356
rect 7932 31272 7984 31278
rect 7932 31214 7984 31220
rect 7472 31204 7524 31210
rect 7472 31146 7524 31152
rect 7484 30580 7512 31146
rect 7622 31036 7918 31056
rect 7678 31034 7702 31036
rect 7758 31034 7782 31036
rect 7838 31034 7862 31036
rect 7700 30982 7702 31034
rect 7764 30982 7776 31034
rect 7838 30982 7840 31034
rect 7678 30980 7702 30982
rect 7758 30980 7782 30982
rect 7838 30980 7862 30982
rect 7622 30960 7918 30980
rect 8036 30938 8064 31350
rect 8024 30932 8076 30938
rect 8024 30874 8076 30880
rect 7656 30592 7708 30598
rect 7484 30560 7656 30580
rect 7708 30560 7710 30569
rect 7484 30552 7654 30560
rect 7654 30495 7710 30504
rect 7622 29948 7918 29968
rect 7678 29946 7702 29948
rect 7758 29946 7782 29948
rect 7838 29946 7862 29948
rect 7700 29894 7702 29946
rect 7764 29894 7776 29946
rect 7838 29894 7840 29946
rect 7678 29892 7702 29894
rect 7758 29892 7782 29894
rect 7838 29892 7862 29894
rect 7622 29872 7918 29892
rect 8128 29073 8156 32694
rect 8114 29064 8170 29073
rect 8114 28999 8170 29008
rect 8024 28960 8076 28966
rect 8024 28902 8076 28908
rect 8116 28960 8168 28966
rect 8116 28902 8168 28908
rect 7622 28860 7918 28880
rect 7678 28858 7702 28860
rect 7758 28858 7782 28860
rect 7838 28858 7862 28860
rect 7700 28806 7702 28858
rect 7764 28806 7776 28858
rect 7838 28806 7840 28858
rect 7678 28804 7702 28806
rect 7758 28804 7782 28806
rect 7838 28804 7862 28806
rect 7622 28784 7918 28804
rect 8036 28626 8064 28902
rect 8128 28762 8156 28902
rect 8116 28756 8168 28762
rect 8116 28698 8168 28704
rect 8114 28656 8170 28665
rect 8024 28620 8076 28626
rect 8114 28591 8170 28600
rect 8024 28562 8076 28568
rect 8036 28218 8064 28562
rect 8024 28212 8076 28218
rect 8024 28154 8076 28160
rect 7472 27940 7524 27946
rect 7472 27882 7524 27888
rect 7380 27328 7432 27334
rect 7380 27270 7432 27276
rect 7392 25362 7420 27270
rect 7484 26926 7512 27882
rect 7622 27772 7918 27792
rect 7678 27770 7702 27772
rect 7758 27770 7782 27772
rect 7838 27770 7862 27772
rect 7700 27718 7702 27770
rect 7764 27718 7776 27770
rect 7838 27718 7840 27770
rect 7678 27716 7702 27718
rect 7758 27716 7782 27718
rect 7838 27716 7862 27718
rect 7622 27696 7918 27716
rect 7932 27600 7984 27606
rect 7932 27542 7984 27548
rect 7944 27062 7972 27542
rect 8024 27532 8076 27538
rect 8024 27474 8076 27480
rect 8036 27130 8064 27474
rect 8024 27124 8076 27130
rect 8024 27066 8076 27072
rect 7932 27056 7984 27062
rect 7932 26998 7984 27004
rect 7472 26920 7524 26926
rect 7472 26862 7524 26868
rect 7484 26586 7512 26862
rect 7622 26684 7918 26704
rect 7678 26682 7702 26684
rect 7758 26682 7782 26684
rect 7838 26682 7862 26684
rect 7700 26630 7702 26682
rect 7764 26630 7776 26682
rect 7838 26630 7840 26682
rect 7678 26628 7702 26630
rect 7758 26628 7782 26630
rect 7838 26628 7862 26630
rect 7622 26608 7918 26628
rect 7472 26580 7524 26586
rect 7472 26522 7524 26528
rect 7656 26512 7708 26518
rect 7656 26454 7708 26460
rect 7668 26042 7696 26454
rect 8128 26450 8156 28591
rect 8116 26444 8168 26450
rect 8116 26386 8168 26392
rect 7656 26036 7708 26042
rect 7656 25978 7708 25984
rect 7668 25838 7696 25978
rect 7656 25832 7708 25838
rect 7656 25774 7708 25780
rect 7622 25596 7918 25616
rect 7678 25594 7702 25596
rect 7758 25594 7782 25596
rect 7838 25594 7862 25596
rect 7700 25542 7702 25594
rect 7764 25542 7776 25594
rect 7838 25542 7840 25594
rect 7678 25540 7702 25542
rect 7758 25540 7782 25542
rect 7838 25540 7862 25542
rect 7622 25520 7918 25540
rect 7380 25356 7432 25362
rect 7380 25298 7432 25304
rect 7472 25356 7524 25362
rect 7472 25298 7524 25304
rect 7392 24886 7420 25298
rect 7380 24880 7432 24886
rect 7380 24822 7432 24828
rect 7380 24744 7432 24750
rect 7380 24686 7432 24692
rect 7392 24410 7420 24686
rect 7380 24404 7432 24410
rect 7380 24346 7432 24352
rect 7484 24041 7512 25298
rect 8024 24812 8076 24818
rect 8024 24754 8076 24760
rect 7622 24508 7918 24528
rect 7678 24506 7702 24508
rect 7758 24506 7782 24508
rect 7838 24506 7862 24508
rect 7700 24454 7702 24506
rect 7764 24454 7776 24506
rect 7838 24454 7840 24506
rect 7678 24452 7702 24454
rect 7758 24452 7782 24454
rect 7838 24452 7862 24454
rect 7622 24432 7918 24452
rect 8036 24138 8064 24754
rect 8024 24132 8076 24138
rect 8024 24074 8076 24080
rect 7470 24032 7526 24041
rect 7470 23967 7526 23976
rect 7012 23724 7064 23730
rect 7300 23718 7420 23746
rect 7012 23666 7064 23672
rect 6552 23656 6604 23662
rect 6472 23616 6552 23644
rect 6472 22234 6500 23616
rect 6552 23598 6604 23604
rect 6552 23180 6604 23186
rect 6552 23122 6604 23128
rect 6564 22778 6592 23122
rect 6552 22772 6604 22778
rect 6552 22714 6604 22720
rect 6736 22772 6788 22778
rect 6736 22714 6788 22720
rect 6460 22228 6512 22234
rect 6460 22170 6512 22176
rect 6748 22166 6776 22714
rect 6736 22160 6788 22166
rect 6736 22102 6788 22108
rect 6368 22024 6420 22030
rect 6368 21966 6420 21972
rect 6380 21486 6408 21966
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 6368 21480 6420 21486
rect 6368 21422 6420 21428
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 6368 21344 6420 21350
rect 6368 21286 6420 21292
rect 6196 21146 6224 21286
rect 6184 21140 6236 21146
rect 6184 21082 6236 21088
rect 5908 21072 5960 21078
rect 5908 21014 5960 21020
rect 5816 21004 5868 21010
rect 5816 20946 5868 20952
rect 5448 20256 5500 20262
rect 5448 20198 5500 20204
rect 5460 19310 5488 20198
rect 5828 20058 5856 20946
rect 5816 20052 5868 20058
rect 5816 19994 5868 20000
rect 6380 19922 6408 21286
rect 6656 21078 6684 21490
rect 6748 21146 6776 22102
rect 7024 22098 7052 23666
rect 7392 23662 7420 23718
rect 8036 23662 8064 24074
rect 7104 23656 7156 23662
rect 7104 23598 7156 23604
rect 7288 23656 7340 23662
rect 7288 23598 7340 23604
rect 7380 23656 7432 23662
rect 7380 23598 7432 23604
rect 8024 23656 8076 23662
rect 8024 23598 8076 23604
rect 7116 22438 7144 23598
rect 7300 23186 7328 23598
rect 7392 23322 7420 23598
rect 7622 23420 7918 23440
rect 7678 23418 7702 23420
rect 7758 23418 7782 23420
rect 7838 23418 7862 23420
rect 7700 23366 7702 23418
rect 7764 23366 7776 23418
rect 7838 23366 7840 23418
rect 7678 23364 7702 23366
rect 7758 23364 7782 23366
rect 7838 23364 7862 23366
rect 7622 23344 7918 23364
rect 7380 23316 7432 23322
rect 7380 23258 7432 23264
rect 7288 23180 7340 23186
rect 7288 23122 7340 23128
rect 7564 23180 7616 23186
rect 7564 23122 7616 23128
rect 7380 23112 7432 23118
rect 7380 23054 7432 23060
rect 7392 22438 7420 23054
rect 7576 22506 7604 23122
rect 8128 22778 8156 26386
rect 8116 22772 8168 22778
rect 8116 22714 8168 22720
rect 8128 22574 8156 22714
rect 8116 22568 8168 22574
rect 8116 22510 8168 22516
rect 7564 22500 7616 22506
rect 7564 22442 7616 22448
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 7380 22432 7432 22438
rect 7380 22374 7432 22380
rect 7116 22098 7144 22374
rect 7012 22092 7064 22098
rect 7012 22034 7064 22040
rect 7104 22092 7156 22098
rect 7104 22034 7156 22040
rect 6828 21412 6880 21418
rect 6880 21372 7052 21400
rect 6828 21354 6880 21360
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 6644 21072 6696 21078
rect 6644 21014 6696 21020
rect 6656 20534 6684 21014
rect 6644 20528 6696 20534
rect 6644 20470 6696 20476
rect 6552 20052 6604 20058
rect 6552 19994 6604 20000
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6380 19310 6408 19858
rect 6564 19514 6592 19994
rect 6656 19836 6684 20470
rect 6920 20256 6972 20262
rect 6920 20198 6972 20204
rect 6932 19922 6960 20198
rect 6920 19916 6972 19922
rect 6920 19858 6972 19864
rect 6736 19848 6788 19854
rect 6656 19808 6736 19836
rect 6736 19790 6788 19796
rect 6748 19514 6776 19790
rect 7024 19718 7052 21372
rect 7116 21350 7144 22034
rect 7392 21894 7420 22374
rect 7622 22332 7918 22352
rect 7678 22330 7702 22332
rect 7758 22330 7782 22332
rect 7838 22330 7862 22332
rect 7700 22278 7702 22330
rect 7764 22278 7776 22330
rect 7838 22278 7840 22330
rect 7678 22276 7702 22278
rect 7758 22276 7782 22278
rect 7838 22276 7862 22278
rect 7622 22256 7918 22276
rect 8114 22264 8170 22273
rect 8114 22199 8170 22208
rect 8128 22030 8156 22199
rect 8116 22024 8168 22030
rect 8116 21966 8168 21972
rect 7380 21888 7432 21894
rect 7380 21830 7432 21836
rect 7392 21690 7420 21830
rect 7380 21684 7432 21690
rect 7380 21626 7432 21632
rect 8220 21486 8248 47398
rect 8312 47054 8340 47534
rect 8404 47258 8432 48146
rect 8496 47802 8524 49710
rect 8484 47796 8536 47802
rect 8484 47738 8536 47744
rect 8588 47682 8616 49846
rect 8496 47654 8616 47682
rect 8392 47252 8444 47258
rect 8392 47194 8444 47200
rect 8300 47048 8352 47054
rect 8300 46990 8352 46996
rect 8404 46986 8432 47194
rect 8392 46980 8444 46986
rect 8392 46922 8444 46928
rect 8300 46912 8352 46918
rect 8300 46854 8352 46860
rect 8390 46880 8446 46889
rect 8312 44946 8340 46854
rect 8390 46815 8446 46824
rect 8404 45966 8432 46815
rect 8496 46102 8524 47654
rect 8576 47116 8628 47122
rect 8576 47058 8628 47064
rect 8588 46374 8616 47058
rect 8576 46368 8628 46374
rect 8576 46310 8628 46316
rect 8574 46200 8630 46209
rect 8574 46135 8630 46144
rect 8484 46096 8536 46102
rect 8484 46038 8536 46044
rect 8392 45960 8444 45966
rect 8392 45902 8444 45908
rect 8404 45626 8432 45902
rect 8392 45620 8444 45626
rect 8392 45562 8444 45568
rect 8300 44940 8352 44946
rect 8300 44882 8352 44888
rect 8300 44396 8352 44402
rect 8300 44338 8352 44344
rect 8312 43994 8340 44338
rect 8300 43988 8352 43994
rect 8300 43930 8352 43936
rect 8300 43852 8352 43858
rect 8300 43794 8352 43800
rect 8312 43450 8340 43794
rect 8300 43444 8352 43450
rect 8300 43386 8352 43392
rect 8312 42809 8340 43386
rect 8404 42906 8432 45562
rect 8496 43450 8524 46038
rect 8484 43444 8536 43450
rect 8484 43386 8536 43392
rect 8588 43246 8616 46135
rect 8680 45014 8708 51360
rect 8760 51264 8812 51270
rect 8760 51206 8812 51212
rect 8772 50969 8800 51206
rect 8758 50960 8814 50969
rect 8758 50895 8814 50904
rect 8760 50856 8812 50862
rect 8760 50798 8812 50804
rect 8772 50697 8800 50798
rect 8758 50688 8814 50697
rect 8758 50623 8814 50632
rect 8864 49910 8892 52090
rect 8956 51610 8984 56102
rect 9048 54738 9076 57734
rect 9036 54732 9088 54738
rect 9036 54674 9088 54680
rect 9048 54534 9076 54674
rect 9036 54528 9088 54534
rect 9036 54470 9088 54476
rect 9048 52154 9076 54470
rect 9036 52148 9088 52154
rect 9036 52090 9088 52096
rect 8944 51604 8996 51610
rect 8944 51546 8996 51552
rect 8956 51241 8984 51546
rect 9036 51536 9088 51542
rect 9036 51478 9088 51484
rect 8942 51232 8998 51241
rect 8942 51167 8998 51176
rect 8942 50960 8998 50969
rect 8942 50895 8998 50904
rect 8956 50726 8984 50895
rect 8944 50720 8996 50726
rect 8944 50662 8996 50668
rect 8956 50318 8984 50662
rect 8944 50312 8996 50318
rect 8944 50254 8996 50260
rect 8944 50176 8996 50182
rect 8944 50118 8996 50124
rect 8852 49904 8904 49910
rect 8852 49846 8904 49852
rect 8760 49700 8812 49706
rect 8760 49642 8812 49648
rect 8772 49434 8800 49642
rect 8852 49632 8904 49638
rect 8852 49574 8904 49580
rect 8760 49428 8812 49434
rect 8760 49370 8812 49376
rect 8864 49298 8892 49574
rect 8852 49292 8904 49298
rect 8852 49234 8904 49240
rect 8864 48550 8892 49234
rect 8852 48544 8904 48550
rect 8852 48486 8904 48492
rect 8852 48340 8904 48346
rect 8852 48282 8904 48288
rect 8760 48000 8812 48006
rect 8760 47942 8812 47948
rect 8772 47122 8800 47942
rect 8760 47116 8812 47122
rect 8760 47058 8812 47064
rect 8772 46442 8800 47058
rect 8760 46436 8812 46442
rect 8760 46378 8812 46384
rect 8668 45008 8720 45014
rect 8668 44950 8720 44956
rect 8680 43654 8708 44950
rect 8668 43648 8720 43654
rect 8668 43590 8720 43596
rect 8576 43240 8628 43246
rect 8576 43182 8628 43188
rect 8588 42906 8616 43182
rect 8392 42900 8444 42906
rect 8392 42842 8444 42848
rect 8576 42900 8628 42906
rect 8576 42842 8628 42848
rect 8298 42800 8354 42809
rect 8680 42786 8708 43590
rect 8298 42735 8354 42744
rect 8392 42764 8444 42770
rect 8392 42706 8444 42712
rect 8484 42764 8536 42770
rect 8484 42706 8536 42712
rect 8588 42758 8708 42786
rect 8300 42696 8352 42702
rect 8300 42638 8352 42644
rect 8312 41818 8340 42638
rect 8404 42362 8432 42706
rect 8392 42356 8444 42362
rect 8392 42298 8444 42304
rect 8300 41812 8352 41818
rect 8300 41754 8352 41760
rect 8300 41064 8352 41070
rect 8300 41006 8352 41012
rect 8312 40390 8340 41006
rect 8300 40384 8352 40390
rect 8300 40326 8352 40332
rect 8312 38593 8340 40326
rect 8404 39098 8432 42298
rect 8496 41818 8524 42706
rect 8484 41812 8536 41818
rect 8484 41754 8536 41760
rect 8484 41472 8536 41478
rect 8484 41414 8536 41420
rect 8392 39092 8444 39098
rect 8392 39034 8444 39040
rect 8496 38894 8524 41414
rect 8588 41206 8616 42758
rect 8668 42628 8720 42634
rect 8668 42570 8720 42576
rect 8576 41200 8628 41206
rect 8576 41142 8628 41148
rect 8576 40928 8628 40934
rect 8576 40870 8628 40876
rect 8588 39846 8616 40870
rect 8576 39840 8628 39846
rect 8576 39782 8628 39788
rect 8484 38888 8536 38894
rect 8484 38830 8536 38836
rect 8298 38584 8354 38593
rect 8298 38519 8354 38528
rect 8496 38486 8524 38830
rect 8484 38480 8536 38486
rect 8298 38448 8354 38457
rect 8484 38422 8536 38428
rect 8298 38383 8354 38392
rect 8312 37262 8340 38383
rect 8392 38344 8444 38350
rect 8392 38286 8444 38292
rect 8404 37670 8432 38286
rect 8588 38282 8616 39782
rect 8576 38276 8628 38282
rect 8576 38218 8628 38224
rect 8392 37664 8444 37670
rect 8392 37606 8444 37612
rect 8484 37664 8536 37670
rect 8484 37606 8536 37612
rect 8300 37256 8352 37262
rect 8300 37198 8352 37204
rect 8312 36922 8340 37198
rect 8300 36916 8352 36922
rect 8300 36858 8352 36864
rect 8300 36168 8352 36174
rect 8300 36110 8352 36116
rect 8312 35766 8340 36110
rect 8300 35760 8352 35766
rect 8300 35702 8352 35708
rect 8300 34468 8352 34474
rect 8300 34410 8352 34416
rect 8312 33833 8340 34410
rect 8298 33824 8354 33833
rect 8298 33759 8354 33768
rect 8312 33658 8340 33759
rect 8300 33652 8352 33658
rect 8300 33594 8352 33600
rect 8298 32736 8354 32745
rect 8298 32671 8354 32680
rect 8312 32570 8340 32671
rect 8300 32564 8352 32570
rect 8300 32506 8352 32512
rect 8404 30190 8432 37606
rect 8496 37210 8524 37606
rect 8588 37330 8616 38218
rect 8576 37324 8628 37330
rect 8576 37266 8628 37272
rect 8496 37182 8616 37210
rect 8484 37120 8536 37126
rect 8484 37062 8536 37068
rect 8496 35834 8524 37062
rect 8484 35828 8536 35834
rect 8484 35770 8536 35776
rect 8484 35148 8536 35154
rect 8484 35090 8536 35096
rect 8496 34542 8524 35090
rect 8484 34536 8536 34542
rect 8484 34478 8536 34484
rect 8588 34474 8616 37182
rect 8576 34468 8628 34474
rect 8576 34410 8628 34416
rect 8576 32564 8628 32570
rect 8576 32506 8628 32512
rect 8484 32496 8536 32502
rect 8484 32438 8536 32444
rect 8392 30184 8444 30190
rect 8392 30126 8444 30132
rect 8300 30048 8352 30054
rect 8300 29990 8352 29996
rect 8312 29714 8340 29990
rect 8300 29708 8352 29714
rect 8300 29650 8352 29656
rect 8392 29640 8444 29646
rect 8392 29582 8444 29588
rect 8404 29102 8432 29582
rect 8392 29096 8444 29102
rect 8392 29038 8444 29044
rect 8300 28484 8352 28490
rect 8300 28426 8352 28432
rect 8312 27674 8340 28426
rect 8392 28144 8444 28150
rect 8392 28086 8444 28092
rect 8404 27674 8432 28086
rect 8300 27668 8352 27674
rect 8300 27610 8352 27616
rect 8392 27668 8444 27674
rect 8392 27610 8444 27616
rect 8300 27328 8352 27334
rect 8300 27270 8352 27276
rect 8312 24886 8340 27270
rect 8404 26518 8432 27610
rect 8496 26586 8524 32438
rect 8588 27112 8616 32506
rect 8680 28626 8708 42570
rect 8772 41070 8800 46378
rect 8864 45966 8892 48282
rect 8852 45960 8904 45966
rect 8852 45902 8904 45908
rect 8956 45778 8984 50118
rect 9048 47190 9076 51478
rect 9140 48210 9168 58278
rect 9232 54330 9260 62070
rect 9324 57934 9352 63990
rect 9416 63782 9444 65583
rect 9600 65210 9628 66030
rect 9784 65958 9812 66694
rect 9864 66700 9916 66706
rect 9864 66642 9916 66648
rect 9876 66230 9904 66642
rect 9864 66224 9916 66230
rect 9864 66166 9916 66172
rect 9680 65952 9732 65958
rect 9680 65894 9732 65900
rect 9772 65952 9824 65958
rect 9772 65894 9824 65900
rect 9588 65204 9640 65210
rect 9588 65146 9640 65152
rect 9600 64530 9628 65146
rect 9588 64524 9640 64530
rect 9588 64466 9640 64472
rect 9692 63866 9720 65894
rect 9968 65498 9996 68190
rect 10140 68196 10192 68202
rect 10140 68138 10192 68144
rect 10140 67856 10192 67862
rect 10140 67798 10192 67804
rect 10048 66292 10100 66298
rect 10048 66234 10100 66240
rect 10060 66042 10088 66234
rect 10152 66230 10180 67798
rect 10140 66224 10192 66230
rect 10140 66166 10192 66172
rect 10060 66014 10180 66042
rect 10048 65952 10100 65958
rect 10046 65920 10048 65929
rect 10100 65920 10102 65929
rect 10046 65855 10102 65864
rect 10152 65770 10180 66014
rect 9876 65470 9996 65498
rect 10060 65754 10180 65770
rect 10060 65748 10192 65754
rect 10060 65742 10140 65748
rect 9876 64818 9904 65470
rect 9956 65408 10008 65414
rect 9956 65350 10008 65356
rect 9968 65006 9996 65350
rect 9956 65000 10008 65006
rect 9956 64942 10008 64948
rect 10060 64818 10088 65742
rect 10140 65690 10192 65696
rect 10152 65659 10180 65690
rect 10140 64864 10192 64870
rect 9876 64790 9996 64818
rect 9864 64660 9916 64666
rect 9864 64602 9916 64608
rect 9772 64320 9824 64326
rect 9772 64262 9824 64268
rect 9784 63918 9812 64262
rect 9600 63838 9720 63866
rect 9772 63912 9824 63918
rect 9772 63854 9824 63860
rect 9404 63776 9456 63782
rect 9404 63718 9456 63724
rect 9600 63594 9628 63838
rect 9680 63776 9732 63782
rect 9680 63718 9732 63724
rect 9508 63566 9628 63594
rect 9404 63436 9456 63442
rect 9404 63378 9456 63384
rect 9416 63034 9444 63378
rect 9404 63028 9456 63034
rect 9404 62970 9456 62976
rect 9402 62928 9458 62937
rect 9402 62863 9404 62872
rect 9456 62863 9458 62872
rect 9404 62834 9456 62840
rect 9508 62150 9536 63566
rect 9588 63436 9640 63442
rect 9692 63424 9720 63718
rect 9876 63510 9904 64602
rect 9968 64025 9996 64790
rect 10060 64812 10140 64818
rect 10060 64806 10192 64812
rect 10060 64790 10180 64806
rect 9954 64016 10010 64025
rect 9954 63951 10010 63960
rect 9956 63844 10008 63850
rect 9956 63786 10008 63792
rect 9864 63504 9916 63510
rect 9864 63446 9916 63452
rect 9640 63396 9720 63424
rect 9772 63436 9824 63442
rect 9588 63378 9640 63384
rect 9772 63378 9824 63384
rect 9680 63300 9732 63306
rect 9680 63242 9732 63248
rect 9588 63232 9640 63238
rect 9588 63174 9640 63180
rect 9496 62144 9548 62150
rect 9496 62086 9548 62092
rect 9508 61198 9536 62086
rect 9496 61192 9548 61198
rect 9496 61134 9548 61140
rect 9404 60104 9456 60110
rect 9404 60046 9456 60052
rect 9312 57928 9364 57934
rect 9312 57870 9364 57876
rect 9324 57594 9352 57870
rect 9312 57588 9364 57594
rect 9312 57530 9364 57536
rect 9312 56976 9364 56982
rect 9312 56918 9364 56924
rect 9324 56166 9352 56918
rect 9312 56160 9364 56166
rect 9312 56102 9364 56108
rect 9324 55282 9352 56102
rect 9312 55276 9364 55282
rect 9312 55218 9364 55224
rect 9220 54324 9272 54330
rect 9272 54284 9352 54312
rect 9220 54266 9272 54272
rect 9218 54224 9274 54233
rect 9218 54159 9274 54168
rect 9232 53514 9260 54159
rect 9220 53508 9272 53514
rect 9220 53450 9272 53456
rect 9220 52964 9272 52970
rect 9220 52906 9272 52912
rect 9232 52698 9260 52906
rect 9220 52692 9272 52698
rect 9220 52634 9272 52640
rect 9218 51776 9274 51785
rect 9218 51711 9274 51720
rect 9232 51474 9260 51711
rect 9220 51468 9272 51474
rect 9220 51410 9272 51416
rect 9232 51066 9260 51410
rect 9220 51060 9272 51066
rect 9220 51002 9272 51008
rect 9220 50380 9272 50386
rect 9220 50322 9272 50328
rect 9232 49978 9260 50322
rect 9220 49972 9272 49978
rect 9220 49914 9272 49920
rect 9218 49872 9274 49881
rect 9218 49807 9274 49816
rect 9128 48204 9180 48210
rect 9128 48146 9180 48152
rect 9140 47802 9168 48146
rect 9128 47796 9180 47802
rect 9128 47738 9180 47744
rect 9128 47524 9180 47530
rect 9128 47466 9180 47472
rect 9036 47184 9088 47190
rect 9036 47126 9088 47132
rect 9140 46322 9168 47466
rect 9232 47122 9260 49807
rect 9220 47116 9272 47122
rect 9220 47058 9272 47064
rect 9232 46714 9260 47058
rect 9220 46708 9272 46714
rect 9220 46650 9272 46656
rect 9140 46294 9260 46322
rect 9128 46164 9180 46170
rect 9128 46106 9180 46112
rect 9036 45960 9088 45966
rect 9036 45902 9088 45908
rect 8864 45750 8984 45778
rect 8760 41064 8812 41070
rect 8760 41006 8812 41012
rect 8864 40916 8892 45750
rect 8942 45656 8998 45665
rect 8942 45591 8998 45600
rect 8956 42362 8984 45591
rect 9048 44538 9076 45902
rect 9036 44532 9088 44538
rect 9036 44474 9088 44480
rect 9034 44160 9090 44169
rect 9034 44095 9090 44104
rect 8944 42356 8996 42362
rect 8944 42298 8996 42304
rect 8944 42152 8996 42158
rect 8944 42094 8996 42100
rect 8956 41721 8984 42094
rect 9048 42090 9076 44095
rect 9036 42084 9088 42090
rect 9036 42026 9088 42032
rect 8942 41712 8998 41721
rect 8942 41647 8998 41656
rect 8944 41608 8996 41614
rect 8944 41550 8996 41556
rect 9036 41608 9088 41614
rect 9036 41550 9088 41556
rect 8956 41206 8984 41550
rect 8944 41200 8996 41206
rect 8944 41142 8996 41148
rect 8944 41064 8996 41070
rect 8944 41006 8996 41012
rect 8772 40888 8892 40916
rect 8772 37330 8800 40888
rect 8852 40520 8904 40526
rect 8852 40462 8904 40468
rect 8864 38894 8892 40462
rect 8852 38888 8904 38894
rect 8852 38830 8904 38836
rect 8852 38752 8904 38758
rect 8852 38694 8904 38700
rect 8760 37324 8812 37330
rect 8760 37266 8812 37272
rect 8772 36378 8800 37266
rect 8760 36372 8812 36378
rect 8760 36314 8812 36320
rect 8760 33652 8812 33658
rect 8760 33594 8812 33600
rect 8772 31890 8800 33594
rect 8864 32502 8892 38694
rect 8956 38418 8984 41006
rect 9048 40594 9076 41550
rect 9140 40730 9168 46106
rect 9232 44810 9260 46294
rect 9324 46170 9352 54284
rect 9416 50522 9444 60046
rect 9496 59016 9548 59022
rect 9496 58958 9548 58964
rect 9508 58342 9536 58958
rect 9496 58336 9548 58342
rect 9496 58278 9548 58284
rect 9508 56914 9536 58278
rect 9600 58041 9628 63174
rect 9692 58614 9720 63242
rect 9784 62218 9812 63378
rect 9876 62490 9904 63446
rect 9968 63034 9996 63786
rect 10060 63238 10088 64790
rect 10140 64524 10192 64530
rect 10140 64466 10192 64472
rect 10152 63578 10180 64466
rect 10140 63572 10192 63578
rect 10140 63514 10192 63520
rect 10244 63306 10272 70366
rect 10428 69970 10456 70382
rect 10416 69964 10468 69970
rect 10416 69906 10468 69912
rect 10428 69766 10456 69906
rect 10416 69760 10468 69766
rect 10416 69702 10468 69708
rect 10428 68864 10456 69702
rect 10508 68876 10560 68882
rect 10428 68836 10508 68864
rect 10324 68400 10376 68406
rect 10324 68342 10376 68348
rect 10336 67862 10364 68342
rect 10428 67930 10456 68836
rect 10508 68818 10560 68824
rect 10416 67924 10468 67930
rect 10416 67866 10468 67872
rect 10324 67856 10376 67862
rect 10324 67798 10376 67804
rect 10428 67289 10456 67866
rect 10414 67280 10470 67289
rect 10414 67215 10470 67224
rect 10508 67244 10560 67250
rect 10428 67182 10456 67215
rect 10508 67186 10560 67192
rect 10416 67176 10468 67182
rect 10416 67118 10468 67124
rect 10416 66564 10468 66570
rect 10416 66506 10468 66512
rect 10324 65952 10376 65958
rect 10324 65894 10376 65900
rect 10336 64530 10364 65894
rect 10428 65482 10456 66506
rect 10416 65476 10468 65482
rect 10416 65418 10468 65424
rect 10324 64524 10376 64530
rect 10324 64466 10376 64472
rect 10336 64122 10364 64466
rect 10324 64116 10376 64122
rect 10324 64058 10376 64064
rect 10232 63300 10284 63306
rect 10232 63242 10284 63248
rect 10048 63232 10100 63238
rect 10048 63174 10100 63180
rect 9956 63028 10008 63034
rect 9956 62970 10008 62976
rect 10060 62937 10088 63174
rect 10046 62928 10102 62937
rect 10046 62863 10102 62872
rect 10048 62824 10100 62830
rect 10048 62766 10100 62772
rect 10232 62824 10284 62830
rect 10232 62766 10284 62772
rect 9864 62484 9916 62490
rect 9864 62426 9916 62432
rect 9864 62348 9916 62354
rect 9864 62290 9916 62296
rect 9772 62212 9824 62218
rect 9772 62154 9824 62160
rect 9772 61396 9824 61402
rect 9772 61338 9824 61344
rect 9784 61266 9812 61338
rect 9876 61266 9904 62290
rect 10060 61305 10088 62766
rect 10244 62490 10272 62766
rect 10232 62484 10284 62490
rect 10232 62426 10284 62432
rect 10140 62212 10192 62218
rect 10140 62154 10192 62160
rect 10152 61606 10180 62154
rect 10244 61674 10272 62426
rect 10336 61742 10364 64058
rect 10324 61736 10376 61742
rect 10324 61678 10376 61684
rect 10232 61668 10284 61674
rect 10232 61610 10284 61616
rect 10140 61600 10192 61606
rect 10140 61542 10192 61548
rect 10046 61296 10102 61305
rect 9772 61260 9824 61266
rect 9772 61202 9824 61208
rect 9864 61260 9916 61266
rect 10046 61231 10102 61240
rect 9864 61202 9916 61208
rect 9784 60314 9812 61202
rect 9876 60858 9904 61202
rect 10048 61192 10100 61198
rect 10048 61134 10100 61140
rect 10060 60858 10088 61134
rect 9864 60852 9916 60858
rect 9864 60794 9916 60800
rect 10048 60852 10100 60858
rect 10048 60794 10100 60800
rect 9772 60308 9824 60314
rect 9772 60250 9824 60256
rect 9784 59498 9812 60250
rect 9772 59492 9824 59498
rect 9772 59434 9824 59440
rect 9784 59090 9812 59434
rect 9876 59401 9904 60794
rect 9954 60752 10010 60761
rect 9954 60687 10010 60696
rect 9862 59392 9918 59401
rect 9862 59327 9918 59336
rect 9772 59084 9824 59090
rect 9772 59026 9824 59032
rect 9680 58608 9732 58614
rect 9680 58550 9732 58556
rect 9680 58472 9732 58478
rect 9680 58414 9732 58420
rect 9586 58032 9642 58041
rect 9586 57967 9642 57976
rect 9692 57798 9720 58414
rect 9772 57996 9824 58002
rect 9772 57938 9824 57944
rect 9680 57792 9732 57798
rect 9680 57734 9732 57740
rect 9784 57610 9812 57938
rect 9588 57588 9640 57594
rect 9588 57530 9640 57536
rect 9692 57582 9812 57610
rect 9496 56908 9548 56914
rect 9496 56850 9548 56856
rect 9494 56264 9550 56273
rect 9494 56199 9550 56208
rect 9508 55962 9536 56199
rect 9496 55956 9548 55962
rect 9496 55898 9548 55904
rect 9494 55720 9550 55729
rect 9494 55655 9550 55664
rect 9508 55350 9536 55655
rect 9496 55344 9548 55350
rect 9496 55286 9548 55292
rect 9600 55298 9628 57530
rect 9692 57089 9720 57582
rect 9864 57452 9916 57458
rect 9864 57394 9916 57400
rect 9772 57316 9824 57322
rect 9772 57258 9824 57264
rect 9678 57080 9734 57089
rect 9678 57015 9680 57024
rect 9732 57015 9734 57024
rect 9680 56986 9732 56992
rect 9692 56955 9720 56986
rect 9680 56908 9732 56914
rect 9680 56850 9732 56856
rect 9692 55962 9720 56850
rect 9680 55956 9732 55962
rect 9680 55898 9732 55904
rect 9680 55820 9732 55826
rect 9680 55762 9732 55768
rect 9692 55457 9720 55762
rect 9678 55448 9734 55457
rect 9678 55383 9734 55392
rect 9508 54670 9536 55286
rect 9600 55270 9720 55298
rect 9588 55072 9640 55078
rect 9588 55014 9640 55020
rect 9496 54664 9548 54670
rect 9496 54606 9548 54612
rect 9496 54528 9548 54534
rect 9496 54470 9548 54476
rect 9508 54126 9536 54470
rect 9496 54120 9548 54126
rect 9496 54062 9548 54068
rect 9508 53961 9536 54062
rect 9494 53952 9550 53961
rect 9494 53887 9550 53896
rect 9600 53718 9628 55014
rect 9692 54126 9720 55270
rect 9784 54806 9812 57258
rect 9876 57254 9904 57394
rect 9864 57248 9916 57254
rect 9864 57190 9916 57196
rect 9876 56409 9904 57190
rect 9862 56400 9918 56409
rect 9862 56335 9918 56344
rect 9864 56296 9916 56302
rect 9864 56238 9916 56244
rect 9876 55826 9904 56238
rect 9864 55820 9916 55826
rect 9864 55762 9916 55768
rect 9968 55706 9996 60687
rect 10046 59392 10102 59401
rect 10046 59327 10102 59336
rect 9876 55678 9996 55706
rect 9772 54800 9824 54806
rect 9772 54742 9824 54748
rect 9784 54534 9812 54742
rect 9772 54528 9824 54534
rect 9772 54470 9824 54476
rect 9772 54256 9824 54262
rect 9772 54198 9824 54204
rect 9680 54120 9732 54126
rect 9680 54062 9732 54068
rect 9692 53786 9720 54062
rect 9680 53780 9732 53786
rect 9680 53722 9732 53728
rect 9588 53712 9640 53718
rect 9588 53654 9640 53660
rect 9496 53644 9548 53650
rect 9496 53586 9548 53592
rect 9508 53242 9536 53586
rect 9588 53508 9640 53514
rect 9588 53450 9640 53456
rect 9496 53236 9548 53242
rect 9496 53178 9548 53184
rect 9508 51388 9536 53178
rect 9600 51950 9628 53450
rect 9678 52864 9734 52873
rect 9678 52799 9734 52808
rect 9588 51944 9640 51950
rect 9588 51886 9640 51892
rect 9586 51640 9642 51649
rect 9586 51575 9642 51584
rect 9600 51542 9628 51575
rect 9588 51536 9640 51542
rect 9588 51478 9640 51484
rect 9508 51360 9628 51388
rect 9692 51377 9720 52799
rect 9784 51542 9812 54198
rect 9772 51536 9824 51542
rect 9772 51478 9824 51484
rect 9600 51048 9628 51360
rect 9678 51368 9734 51377
rect 9678 51303 9734 51312
rect 9772 51332 9824 51338
rect 9772 51274 9824 51280
rect 9784 51066 9812 51274
rect 9508 51020 9628 51048
rect 9680 51060 9732 51066
rect 9404 50516 9456 50522
rect 9404 50458 9456 50464
rect 9404 50380 9456 50386
rect 9404 50322 9456 50328
rect 9416 49774 9444 50322
rect 9404 49768 9456 49774
rect 9404 49710 9456 49716
rect 9416 48278 9444 49710
rect 9404 48272 9456 48278
rect 9404 48214 9456 48220
rect 9404 46368 9456 46374
rect 9404 46310 9456 46316
rect 9312 46164 9364 46170
rect 9312 46106 9364 46112
rect 9416 46050 9444 46310
rect 9324 46022 9444 46050
rect 9220 44804 9272 44810
rect 9220 44746 9272 44752
rect 9232 44470 9260 44746
rect 9220 44464 9272 44470
rect 9220 44406 9272 44412
rect 9232 41682 9260 44406
rect 9220 41676 9272 41682
rect 9220 41618 9272 41624
rect 9218 41576 9274 41585
rect 9218 41511 9274 41520
rect 9232 41274 9260 41511
rect 9220 41268 9272 41274
rect 9220 41210 9272 41216
rect 9220 41132 9272 41138
rect 9220 41074 9272 41080
rect 9128 40724 9180 40730
rect 9128 40666 9180 40672
rect 9232 40610 9260 41074
rect 9036 40588 9088 40594
rect 9036 40530 9088 40536
rect 9140 40582 9260 40610
rect 9034 40488 9090 40497
rect 9034 40423 9036 40432
rect 9088 40423 9090 40432
rect 9036 40394 9088 40400
rect 9036 40112 9088 40118
rect 9036 40054 9088 40060
rect 8944 38412 8996 38418
rect 8944 38354 8996 38360
rect 9048 38321 9076 40054
rect 9034 38312 9090 38321
rect 9034 38247 9090 38256
rect 9140 37913 9168 40582
rect 9220 40452 9272 40458
rect 9220 40394 9272 40400
rect 9232 39846 9260 40394
rect 9220 39840 9272 39846
rect 9220 39782 9272 39788
rect 9218 38992 9274 39001
rect 9218 38927 9274 38936
rect 9232 38729 9260 38927
rect 9218 38720 9274 38729
rect 9218 38655 9274 38664
rect 9324 38554 9352 46022
rect 9404 45484 9456 45490
rect 9404 45426 9456 45432
rect 9416 42566 9444 45426
rect 9404 42560 9456 42566
rect 9404 42502 9456 42508
rect 9404 42356 9456 42362
rect 9404 42298 9456 42304
rect 9416 39574 9444 42298
rect 9508 42242 9536 51020
rect 9680 51002 9732 51008
rect 9772 51060 9824 51066
rect 9772 51002 9824 51008
rect 9692 50164 9720 51002
rect 9772 50720 9824 50726
rect 9772 50662 9824 50668
rect 9600 50136 9720 50164
rect 9600 49978 9628 50136
rect 9678 50008 9734 50017
rect 9588 49972 9640 49978
rect 9678 49943 9734 49952
rect 9588 49914 9640 49920
rect 9692 49774 9720 49943
rect 9680 49768 9732 49774
rect 9600 49728 9680 49756
rect 9600 49366 9628 49728
rect 9680 49710 9732 49716
rect 9680 49632 9732 49638
rect 9680 49574 9732 49580
rect 9588 49360 9640 49366
rect 9588 49302 9640 49308
rect 9692 49230 9720 49574
rect 9680 49224 9732 49230
rect 9680 49166 9732 49172
rect 9588 48680 9640 48686
rect 9586 48648 9588 48657
rect 9640 48648 9642 48657
rect 9586 48583 9642 48592
rect 9588 48544 9640 48550
rect 9640 48504 9720 48532
rect 9588 48486 9640 48492
rect 9588 48272 9640 48278
rect 9588 48214 9640 48220
rect 9600 44878 9628 48214
rect 9692 47462 9720 48504
rect 9680 47456 9732 47462
rect 9680 47398 9732 47404
rect 9784 46714 9812 50662
rect 9876 49280 9904 55678
rect 9956 55208 10008 55214
rect 9956 55150 10008 55156
rect 9968 54233 9996 55150
rect 9954 54224 10010 54233
rect 9954 54159 10010 54168
rect 9954 53136 10010 53145
rect 9954 53071 10010 53080
rect 9968 52562 9996 53071
rect 9956 52556 10008 52562
rect 9956 52498 10008 52504
rect 9956 52352 10008 52358
rect 9956 52294 10008 52300
rect 9968 51950 9996 52294
rect 9956 51944 10008 51950
rect 9956 51886 10008 51892
rect 9956 51604 10008 51610
rect 9956 51546 10008 51552
rect 9968 49434 9996 51546
rect 10060 49586 10088 59327
rect 10152 54262 10180 61542
rect 10244 61402 10272 61610
rect 10232 61396 10284 61402
rect 10232 61338 10284 61344
rect 10336 61282 10364 61678
rect 10244 61254 10364 61282
rect 10244 61062 10272 61254
rect 10428 61180 10456 65418
rect 10520 64054 10548 67186
rect 10612 65929 10640 71454
rect 10784 71120 10836 71126
rect 10784 71062 10836 71068
rect 10796 70650 10824 71062
rect 10784 70644 10836 70650
rect 10784 70586 10836 70592
rect 10796 70514 10824 70586
rect 10784 70508 10836 70514
rect 10784 70450 10836 70456
rect 10888 70394 10916 72558
rect 11336 71936 11388 71942
rect 11336 71878 11388 71884
rect 10956 71836 11252 71856
rect 11012 71834 11036 71836
rect 11092 71834 11116 71836
rect 11172 71834 11196 71836
rect 11034 71782 11036 71834
rect 11098 71782 11110 71834
rect 11172 71782 11174 71834
rect 11012 71780 11036 71782
rect 11092 71780 11116 71782
rect 11172 71780 11196 71782
rect 10956 71760 11252 71780
rect 11348 71602 11376 71878
rect 11336 71596 11388 71602
rect 11336 71538 11388 71544
rect 11428 71528 11480 71534
rect 11428 71470 11480 71476
rect 11336 71460 11388 71466
rect 11336 71402 11388 71408
rect 10956 70748 11252 70768
rect 11012 70746 11036 70748
rect 11092 70746 11116 70748
rect 11172 70746 11196 70748
rect 11034 70694 11036 70746
rect 11098 70694 11110 70746
rect 11172 70694 11174 70746
rect 11012 70692 11036 70694
rect 11092 70692 11116 70694
rect 11172 70692 11196 70694
rect 10956 70672 11252 70692
rect 10796 70366 10916 70394
rect 10692 68740 10744 68746
rect 10692 68682 10744 68688
rect 10704 68338 10732 68682
rect 10796 68406 10824 70366
rect 10956 69660 11252 69680
rect 11012 69658 11036 69660
rect 11092 69658 11116 69660
rect 11172 69658 11196 69660
rect 11034 69606 11036 69658
rect 11098 69606 11110 69658
rect 11172 69606 11174 69658
rect 11012 69604 11036 69606
rect 11092 69604 11116 69606
rect 11172 69604 11196 69606
rect 10956 69584 11252 69604
rect 11060 69216 11112 69222
rect 11060 69158 11112 69164
rect 11072 68898 11100 69158
rect 10888 68870 11100 68898
rect 10784 68400 10836 68406
rect 10784 68342 10836 68348
rect 10692 68332 10744 68338
rect 10692 68274 10744 68280
rect 10704 67794 10732 68274
rect 10784 68196 10836 68202
rect 10784 68138 10836 68144
rect 10692 67788 10744 67794
rect 10692 67730 10744 67736
rect 10704 66502 10732 67730
rect 10692 66496 10744 66502
rect 10692 66438 10744 66444
rect 10598 65920 10654 65929
rect 10598 65855 10654 65864
rect 10704 65618 10732 66438
rect 10692 65612 10744 65618
rect 10692 65554 10744 65560
rect 10600 65544 10652 65550
rect 10600 65486 10652 65492
rect 10612 65210 10640 65486
rect 10600 65204 10652 65210
rect 10600 65146 10652 65152
rect 10704 65090 10732 65554
rect 10796 65249 10824 68138
rect 10888 67590 10916 68870
rect 10956 68572 11252 68592
rect 11012 68570 11036 68572
rect 11092 68570 11116 68572
rect 11172 68570 11196 68572
rect 11034 68518 11036 68570
rect 11098 68518 11110 68570
rect 11172 68518 11174 68570
rect 11012 68516 11036 68518
rect 11092 68516 11116 68518
rect 11172 68516 11196 68518
rect 10956 68496 11252 68516
rect 11348 68406 11376 71402
rect 11440 71126 11468 71470
rect 11428 71120 11480 71126
rect 11428 71062 11480 71068
rect 11624 70417 11652 72558
rect 11980 72558 12032 72564
rect 12348 72616 12400 72622
rect 12400 72576 12756 72604
rect 12348 72558 12400 72564
rect 11794 72519 11850 72528
rect 11992 72282 12020 72558
rect 12532 72480 12584 72486
rect 12532 72422 12584 72428
rect 11980 72276 12032 72282
rect 11980 72218 12032 72224
rect 11704 71528 11756 71534
rect 11704 71470 11756 71476
rect 11888 71528 11940 71534
rect 11888 71470 11940 71476
rect 11716 71398 11744 71470
rect 11704 71392 11756 71398
rect 11704 71334 11756 71340
rect 11716 70650 11744 71334
rect 11900 71194 11928 71470
rect 11888 71188 11940 71194
rect 11888 71130 11940 71136
rect 11704 70644 11756 70650
rect 11704 70586 11756 70592
rect 11704 70440 11756 70446
rect 11610 70408 11666 70417
rect 11704 70382 11756 70388
rect 11610 70343 11666 70352
rect 11518 70136 11574 70145
rect 11518 70071 11574 70080
rect 11428 68672 11480 68678
rect 11428 68614 11480 68620
rect 11244 68400 11296 68406
rect 11244 68342 11296 68348
rect 11336 68400 11388 68406
rect 11336 68342 11388 68348
rect 11152 68264 11204 68270
rect 11152 68206 11204 68212
rect 11164 67862 11192 68206
rect 11152 67856 11204 67862
rect 11152 67798 11204 67804
rect 11256 67674 11284 68342
rect 11440 68270 11468 68614
rect 11428 68264 11480 68270
rect 11428 68206 11480 68212
rect 11336 68128 11388 68134
rect 11336 68070 11388 68076
rect 11348 67794 11376 68070
rect 11336 67788 11388 67794
rect 11336 67730 11388 67736
rect 11256 67646 11468 67674
rect 10876 67584 10928 67590
rect 10876 67526 10928 67532
rect 11336 67584 11388 67590
rect 11336 67526 11388 67532
rect 10956 67484 11252 67504
rect 11012 67482 11036 67484
rect 11092 67482 11116 67484
rect 11172 67482 11196 67484
rect 11034 67430 11036 67482
rect 11098 67430 11110 67482
rect 11172 67430 11174 67482
rect 11012 67428 11036 67430
rect 11092 67428 11116 67430
rect 11172 67428 11196 67430
rect 10956 67408 11252 67428
rect 11348 67046 11376 67526
rect 11336 67040 11388 67046
rect 11336 66982 11388 66988
rect 10956 66396 11252 66416
rect 11012 66394 11036 66396
rect 11092 66394 11116 66396
rect 11172 66394 11196 66396
rect 11034 66342 11036 66394
rect 11098 66342 11110 66394
rect 11172 66342 11174 66394
rect 11012 66340 11036 66342
rect 11092 66340 11116 66342
rect 11172 66340 11196 66342
rect 10956 66320 11252 66340
rect 11060 66224 11112 66230
rect 10888 66172 11060 66178
rect 10888 66166 11112 66172
rect 10888 66150 11100 66166
rect 10782 65240 10838 65249
rect 10782 65175 10838 65184
rect 10600 65068 10652 65074
rect 10704 65062 10824 65090
rect 10600 65010 10652 65016
rect 10508 64048 10560 64054
rect 10508 63990 10560 63996
rect 10520 63918 10548 63990
rect 10508 63912 10560 63918
rect 10508 63854 10560 63860
rect 10508 63572 10560 63578
rect 10508 63514 10560 63520
rect 10336 61152 10456 61180
rect 10232 61056 10284 61062
rect 10232 60998 10284 61004
rect 10140 54256 10192 54262
rect 10140 54198 10192 54204
rect 10140 54120 10192 54126
rect 10140 54062 10192 54068
rect 10152 53582 10180 54062
rect 10140 53576 10192 53582
rect 10140 53518 10192 53524
rect 10140 53440 10192 53446
rect 10140 53382 10192 53388
rect 10152 52578 10180 53382
rect 10244 53224 10272 60998
rect 10336 57594 10364 61152
rect 10416 60648 10468 60654
rect 10416 60590 10468 60596
rect 10428 60314 10456 60590
rect 10416 60308 10468 60314
rect 10416 60250 10468 60256
rect 10414 60208 10470 60217
rect 10414 60143 10470 60152
rect 10428 59566 10456 60143
rect 10416 59560 10468 59566
rect 10416 59502 10468 59508
rect 10414 59392 10470 59401
rect 10414 59327 10470 59336
rect 10428 58614 10456 59327
rect 10416 58608 10468 58614
rect 10416 58550 10468 58556
rect 10414 58440 10470 58449
rect 10414 58375 10470 58384
rect 10324 57588 10376 57594
rect 10324 57530 10376 57536
rect 10336 57390 10364 57530
rect 10324 57384 10376 57390
rect 10324 57326 10376 57332
rect 10336 55826 10364 57326
rect 10428 56846 10456 58375
rect 10416 56840 10468 56846
rect 10416 56782 10468 56788
rect 10428 56438 10456 56782
rect 10416 56432 10468 56438
rect 10414 56400 10416 56409
rect 10468 56400 10470 56409
rect 10414 56335 10470 56344
rect 10416 56228 10468 56234
rect 10416 56170 10468 56176
rect 10324 55820 10376 55826
rect 10324 55762 10376 55768
rect 10336 55418 10364 55762
rect 10324 55412 10376 55418
rect 10324 55354 10376 55360
rect 10324 54256 10376 54262
rect 10324 54198 10376 54204
rect 10336 53446 10364 54198
rect 10324 53440 10376 53446
rect 10324 53382 10376 53388
rect 10244 53196 10364 53224
rect 10230 53136 10286 53145
rect 10230 53071 10232 53080
rect 10284 53071 10286 53080
rect 10232 53042 10284 53048
rect 10152 52550 10272 52578
rect 10140 52488 10192 52494
rect 10138 52456 10140 52465
rect 10192 52456 10194 52465
rect 10138 52391 10194 52400
rect 10244 52034 10272 52550
rect 10152 52006 10272 52034
rect 10152 51513 10180 52006
rect 10232 51944 10284 51950
rect 10232 51886 10284 51892
rect 10138 51504 10194 51513
rect 10138 51439 10194 51448
rect 10140 51400 10192 51406
rect 10140 51342 10192 51348
rect 10152 50833 10180 51342
rect 10138 50824 10194 50833
rect 10138 50759 10194 50768
rect 10152 50454 10180 50759
rect 10140 50448 10192 50454
rect 10140 50390 10192 50396
rect 10152 49978 10180 50390
rect 10140 49972 10192 49978
rect 10140 49914 10192 49920
rect 10138 49872 10194 49881
rect 10138 49807 10140 49816
rect 10192 49807 10194 49816
rect 10140 49778 10192 49784
rect 10244 49745 10272 51886
rect 10336 51610 10364 53196
rect 10324 51604 10376 51610
rect 10324 51546 10376 51552
rect 10324 51468 10376 51474
rect 10324 51410 10376 51416
rect 10336 51105 10364 51410
rect 10322 51096 10378 51105
rect 10322 51031 10324 51040
rect 10376 51031 10378 51040
rect 10324 51002 10376 51008
rect 10336 50971 10364 51002
rect 10324 50856 10376 50862
rect 10322 50824 10324 50833
rect 10376 50824 10378 50833
rect 10322 50759 10378 50768
rect 10324 50720 10376 50726
rect 10324 50662 10376 50668
rect 10336 49774 10364 50662
rect 10324 49768 10376 49774
rect 10230 49736 10286 49745
rect 10324 49710 10376 49716
rect 10230 49671 10286 49680
rect 10060 49558 10272 49586
rect 9956 49428 10008 49434
rect 9956 49370 10008 49376
rect 10140 49428 10192 49434
rect 10140 49370 10192 49376
rect 10048 49292 10100 49298
rect 9876 49252 10048 49280
rect 10048 49234 10100 49240
rect 9954 49192 10010 49201
rect 9954 49127 10010 49136
rect 9864 48680 9916 48686
rect 9864 48622 9916 48628
rect 9876 47054 9904 48622
rect 9864 47048 9916 47054
rect 9864 46990 9916 46996
rect 9864 46912 9916 46918
rect 9864 46854 9916 46860
rect 9680 46708 9732 46714
rect 9680 46650 9732 46656
rect 9772 46708 9824 46714
rect 9772 46650 9824 46656
rect 9692 46034 9720 46650
rect 9680 46028 9732 46034
rect 9680 45970 9732 45976
rect 9876 45966 9904 46854
rect 9968 46510 9996 49127
rect 10060 48006 10088 49234
rect 10152 48686 10180 49370
rect 10140 48680 10192 48686
rect 10140 48622 10192 48628
rect 10152 48346 10180 48622
rect 10140 48340 10192 48346
rect 10140 48282 10192 48288
rect 10140 48136 10192 48142
rect 10140 48078 10192 48084
rect 10048 48000 10100 48006
rect 10048 47942 10100 47948
rect 9956 46504 10008 46510
rect 9956 46446 10008 46452
rect 9968 46170 9996 46446
rect 9956 46164 10008 46170
rect 9956 46106 10008 46112
rect 9864 45960 9916 45966
rect 9916 45920 9996 45948
rect 9864 45902 9916 45908
rect 9680 45824 9732 45830
rect 9680 45766 9732 45772
rect 9864 45824 9916 45830
rect 9864 45766 9916 45772
rect 9692 45082 9720 45766
rect 9876 45558 9904 45766
rect 9864 45552 9916 45558
rect 9862 45520 9864 45529
rect 9916 45520 9918 45529
rect 9862 45455 9918 45464
rect 9772 45416 9824 45422
rect 9772 45358 9824 45364
rect 9680 45076 9732 45082
rect 9680 45018 9732 45024
rect 9588 44872 9640 44878
rect 9588 44814 9640 44820
rect 9600 42770 9628 44814
rect 9692 44402 9720 45018
rect 9784 44946 9812 45358
rect 9968 45336 9996 45920
rect 9876 45308 9996 45336
rect 9876 45082 9904 45308
rect 9954 45248 10010 45257
rect 9954 45183 10010 45192
rect 9864 45076 9916 45082
rect 9864 45018 9916 45024
rect 9772 44940 9824 44946
rect 9772 44882 9824 44888
rect 9680 44396 9732 44402
rect 9680 44338 9732 44344
rect 9772 44260 9824 44266
rect 9772 44202 9824 44208
rect 9864 44260 9916 44266
rect 9864 44202 9916 44208
rect 9680 43852 9732 43858
rect 9680 43794 9732 43800
rect 9588 42764 9640 42770
rect 9588 42706 9640 42712
rect 9600 42673 9628 42706
rect 9586 42664 9642 42673
rect 9586 42599 9642 42608
rect 9692 42378 9720 43794
rect 9784 42702 9812 44202
rect 9876 43790 9904 44202
rect 9864 43784 9916 43790
rect 9862 43752 9864 43761
rect 9916 43752 9918 43761
rect 9862 43687 9918 43696
rect 9864 43308 9916 43314
rect 9864 43250 9916 43256
rect 9772 42696 9824 42702
rect 9772 42638 9824 42644
rect 9772 42560 9824 42566
rect 9772 42502 9824 42508
rect 9600 42362 9720 42378
rect 9588 42356 9720 42362
rect 9640 42350 9720 42356
rect 9588 42298 9640 42304
rect 9508 42214 9628 42242
rect 9496 42016 9548 42022
rect 9496 41958 9548 41964
rect 9508 41682 9536 41958
rect 9600 41698 9628 42214
rect 9600 41682 9720 41698
rect 9496 41676 9548 41682
rect 9496 41618 9548 41624
rect 9600 41676 9732 41682
rect 9600 41670 9680 41676
rect 9494 41440 9550 41449
rect 9494 41375 9550 41384
rect 9404 39568 9456 39574
rect 9402 39536 9404 39545
rect 9456 39536 9458 39545
rect 9402 39471 9458 39480
rect 9508 39386 9536 41375
rect 9600 40594 9628 41670
rect 9680 41618 9732 41624
rect 9680 41200 9732 41206
rect 9680 41142 9732 41148
rect 9588 40588 9640 40594
rect 9588 40530 9640 40536
rect 9600 39914 9628 40530
rect 9588 39908 9640 39914
rect 9588 39850 9640 39856
rect 9588 39636 9640 39642
rect 9692 39624 9720 41142
rect 9640 39596 9720 39624
rect 9588 39578 9640 39584
rect 9416 39358 9536 39386
rect 9312 38548 9364 38554
rect 9312 38490 9364 38496
rect 9220 38208 9272 38214
rect 9220 38150 9272 38156
rect 9126 37904 9182 37913
rect 8956 37862 9126 37890
rect 8956 34649 8984 37862
rect 9126 37839 9182 37848
rect 9128 37800 9180 37806
rect 9128 37742 9180 37748
rect 9036 37392 9088 37398
rect 9036 37334 9088 37340
rect 8942 34640 8998 34649
rect 8942 34575 8998 34584
rect 8944 34536 8996 34542
rect 8944 34478 8996 34484
rect 8852 32496 8904 32502
rect 8852 32438 8904 32444
rect 8760 31884 8812 31890
rect 8760 31826 8812 31832
rect 8852 31816 8904 31822
rect 8758 31784 8814 31793
rect 8814 31764 8852 31770
rect 8814 31758 8904 31764
rect 8814 31742 8892 31758
rect 8758 31719 8814 31728
rect 8772 31482 8800 31719
rect 8760 31476 8812 31482
rect 8760 31418 8812 31424
rect 8956 30258 8984 34478
rect 8944 30252 8996 30258
rect 8944 30194 8996 30200
rect 8760 30184 8812 30190
rect 8760 30126 8812 30132
rect 8668 28620 8720 28626
rect 8668 28562 8720 28568
rect 8680 28218 8708 28562
rect 8668 28212 8720 28218
rect 8668 28154 8720 28160
rect 8772 27334 8800 30126
rect 8852 28620 8904 28626
rect 8852 28562 8904 28568
rect 8864 28218 8892 28562
rect 8852 28212 8904 28218
rect 8852 28154 8904 28160
rect 8760 27328 8812 27334
rect 8760 27270 8812 27276
rect 8588 27084 8892 27112
rect 8668 26988 8720 26994
rect 8668 26930 8720 26936
rect 8680 26586 8708 26930
rect 8484 26580 8536 26586
rect 8484 26522 8536 26528
rect 8668 26580 8720 26586
rect 8668 26522 8720 26528
rect 8392 26512 8444 26518
rect 8392 26454 8444 26460
rect 8496 25838 8524 26522
rect 8760 26444 8812 26450
rect 8760 26386 8812 26392
rect 8668 26376 8720 26382
rect 8668 26318 8720 26324
rect 8576 26240 8628 26246
rect 8576 26182 8628 26188
rect 8588 25838 8616 26182
rect 8484 25832 8536 25838
rect 8484 25774 8536 25780
rect 8576 25832 8628 25838
rect 8576 25774 8628 25780
rect 8300 24880 8352 24886
rect 8300 24822 8352 24828
rect 8300 24744 8352 24750
rect 8300 24686 8352 24692
rect 8312 24410 8340 24686
rect 8300 24404 8352 24410
rect 8300 24346 8352 24352
rect 8484 23724 8536 23730
rect 8484 23666 8536 23672
rect 8496 23322 8524 23666
rect 8484 23316 8536 23322
rect 8484 23258 8536 23264
rect 8300 22568 8352 22574
rect 8300 22510 8352 22516
rect 8312 21690 8340 22510
rect 8484 22500 8536 22506
rect 8484 22442 8536 22448
rect 8496 22234 8524 22442
rect 8484 22228 8536 22234
rect 8484 22170 8536 22176
rect 8588 22030 8616 25774
rect 8680 25498 8708 26318
rect 8772 25974 8800 26386
rect 8760 25968 8812 25974
rect 8760 25910 8812 25916
rect 8772 25498 8800 25910
rect 8668 25492 8720 25498
rect 8668 25434 8720 25440
rect 8760 25492 8812 25498
rect 8760 25434 8812 25440
rect 8680 24138 8708 25434
rect 8864 24750 8892 27084
rect 8852 24744 8904 24750
rect 8852 24686 8904 24692
rect 8956 24274 8984 30194
rect 9048 28014 9076 37334
rect 9140 37330 9168 37742
rect 9128 37324 9180 37330
rect 9128 37266 9180 37272
rect 9140 36854 9168 37266
rect 9128 36848 9180 36854
rect 9128 36790 9180 36796
rect 9232 36242 9260 38150
rect 9324 38010 9352 38490
rect 9312 38004 9364 38010
rect 9312 37946 9364 37952
rect 9324 37670 9352 37946
rect 9312 37664 9364 37670
rect 9312 37606 9364 37612
rect 9324 37466 9352 37606
rect 9312 37460 9364 37466
rect 9312 37402 9364 37408
rect 9312 37324 9364 37330
rect 9312 37266 9364 37272
rect 9324 36922 9352 37266
rect 9312 36916 9364 36922
rect 9312 36858 9364 36864
rect 9324 36378 9352 36858
rect 9312 36372 9364 36378
rect 9312 36314 9364 36320
rect 9220 36236 9272 36242
rect 9220 36178 9272 36184
rect 9232 35834 9260 36178
rect 9220 35828 9272 35834
rect 9220 35770 9272 35776
rect 9416 35766 9444 39358
rect 9496 39296 9548 39302
rect 9496 39238 9548 39244
rect 9404 35760 9456 35766
rect 9404 35702 9456 35708
rect 9508 34490 9536 39238
rect 9692 38978 9720 39596
rect 9600 38950 9720 38978
rect 9600 38894 9628 38950
rect 9588 38888 9640 38894
rect 9588 38830 9640 38836
rect 9678 38720 9734 38729
rect 9678 38655 9734 38664
rect 9586 37768 9642 37777
rect 9586 37703 9642 37712
rect 9600 37330 9628 37703
rect 9588 37324 9640 37330
rect 9588 37266 9640 37272
rect 9600 35834 9628 37266
rect 9588 35828 9640 35834
rect 9588 35770 9640 35776
rect 9692 35222 9720 38655
rect 9784 38418 9812 42502
rect 9876 42226 9904 43250
rect 9864 42220 9916 42226
rect 9864 42162 9916 42168
rect 9864 40996 9916 41002
rect 9864 40938 9916 40944
rect 9876 40390 9904 40938
rect 9864 40384 9916 40390
rect 9864 40326 9916 40332
rect 9772 38412 9824 38418
rect 9772 38354 9824 38360
rect 9772 38276 9824 38282
rect 9772 38218 9824 38224
rect 9680 35216 9732 35222
rect 9680 35158 9732 35164
rect 9784 35068 9812 38218
rect 9876 37738 9904 40326
rect 9968 38894 9996 45183
rect 10060 40118 10088 47942
rect 10152 46918 10180 48078
rect 10140 46912 10192 46918
rect 10140 46854 10192 46860
rect 10140 46708 10192 46714
rect 10140 46650 10192 46656
rect 10048 40112 10100 40118
rect 10048 40054 10100 40060
rect 10048 39840 10100 39846
rect 10048 39782 10100 39788
rect 9956 38888 10008 38894
rect 9956 38830 10008 38836
rect 9954 38720 10010 38729
rect 9954 38655 10010 38664
rect 9968 38214 9996 38655
rect 9956 38208 10008 38214
rect 9956 38150 10008 38156
rect 9864 37732 9916 37738
rect 9864 37674 9916 37680
rect 9968 36718 9996 38150
rect 9956 36712 10008 36718
rect 9956 36654 10008 36660
rect 9956 35624 10008 35630
rect 9956 35566 10008 35572
rect 9968 35154 9996 35566
rect 9956 35148 10008 35154
rect 9956 35090 10008 35096
rect 9692 35040 9812 35068
rect 9416 34462 9536 34490
rect 9586 34504 9642 34513
rect 9126 34096 9182 34105
rect 9126 34031 9182 34040
rect 9140 33998 9168 34031
rect 9128 33992 9180 33998
rect 9128 33934 9180 33940
rect 9140 33658 9168 33934
rect 9128 33652 9180 33658
rect 9128 33594 9180 33600
rect 9128 33040 9180 33046
rect 9128 32982 9180 32988
rect 9140 32774 9168 32982
rect 9310 32872 9366 32881
rect 9310 32807 9312 32816
rect 9364 32807 9366 32816
rect 9312 32778 9364 32784
rect 9128 32768 9180 32774
rect 9128 32710 9180 32716
rect 9140 32366 9168 32710
rect 9324 32502 9352 32778
rect 9312 32496 9364 32502
rect 9312 32438 9364 32444
rect 9128 32360 9180 32366
rect 9128 32302 9180 32308
rect 9312 32360 9364 32366
rect 9312 32302 9364 32308
rect 9128 30184 9180 30190
rect 9128 30126 9180 30132
rect 9140 29714 9168 30126
rect 9128 29708 9180 29714
rect 9128 29650 9180 29656
rect 9036 28008 9088 28014
rect 9036 27950 9088 27956
rect 9048 27674 9076 27950
rect 9220 27872 9272 27878
rect 9220 27814 9272 27820
rect 9036 27668 9088 27674
rect 9036 27610 9088 27616
rect 9036 25356 9088 25362
rect 9036 25298 9088 25304
rect 9048 25265 9076 25298
rect 9034 25256 9090 25265
rect 9034 25191 9090 25200
rect 9048 24954 9076 25191
rect 9036 24948 9088 24954
rect 9036 24890 9088 24896
rect 8944 24268 8996 24274
rect 8944 24210 8996 24216
rect 8668 24132 8720 24138
rect 8668 24074 8720 24080
rect 8956 23322 8984 24210
rect 9036 24200 9088 24206
rect 9036 24142 9088 24148
rect 9048 23526 9076 24142
rect 9036 23520 9088 23526
rect 9036 23462 9088 23468
rect 8944 23316 8996 23322
rect 8944 23258 8996 23264
rect 8576 22024 8628 22030
rect 8576 21966 8628 21972
rect 8300 21684 8352 21690
rect 8300 21626 8352 21632
rect 7288 21480 7340 21486
rect 7288 21422 7340 21428
rect 8208 21480 8260 21486
rect 8208 21422 8260 21428
rect 7104 21344 7156 21350
rect 7104 21286 7156 21292
rect 7116 21010 7144 21286
rect 7300 21146 7328 21422
rect 7622 21244 7918 21264
rect 7678 21242 7702 21244
rect 7758 21242 7782 21244
rect 7838 21242 7862 21244
rect 7700 21190 7702 21242
rect 7764 21190 7776 21242
rect 7838 21190 7840 21242
rect 7678 21188 7702 21190
rect 7758 21188 7782 21190
rect 7838 21188 7862 21190
rect 7622 21168 7918 21188
rect 7288 21140 7340 21146
rect 7288 21082 7340 21088
rect 7104 21004 7156 21010
rect 7104 20946 7156 20952
rect 7472 21004 7524 21010
rect 7472 20946 7524 20952
rect 7116 20602 7144 20946
rect 7104 20596 7156 20602
rect 7104 20538 7156 20544
rect 7484 20466 7512 20946
rect 8220 20466 8248 21422
rect 8588 21078 8616 21966
rect 8760 21344 8812 21350
rect 8760 21286 8812 21292
rect 8576 21072 8628 21078
rect 8576 21014 8628 21020
rect 8772 20602 8800 21286
rect 9048 21010 9076 23462
rect 9036 21004 9088 21010
rect 9036 20946 9088 20952
rect 9048 20602 9076 20946
rect 8760 20596 8812 20602
rect 8760 20538 8812 20544
rect 9036 20596 9088 20602
rect 9036 20538 9088 20544
rect 7472 20460 7524 20466
rect 7472 20402 7524 20408
rect 8208 20460 8260 20466
rect 8208 20402 8260 20408
rect 7484 20058 7512 20402
rect 8024 20256 8076 20262
rect 8024 20198 8076 20204
rect 7622 20156 7918 20176
rect 7678 20154 7702 20156
rect 7758 20154 7782 20156
rect 7838 20154 7862 20156
rect 7700 20102 7702 20154
rect 7764 20102 7776 20154
rect 7838 20102 7840 20154
rect 7678 20100 7702 20102
rect 7758 20100 7782 20102
rect 7838 20100 7862 20102
rect 7622 20080 7918 20100
rect 7472 20052 7524 20058
rect 7472 19994 7524 20000
rect 6828 19712 6880 19718
rect 6828 19654 6880 19660
rect 7012 19712 7064 19718
rect 7012 19654 7064 19660
rect 6552 19508 6604 19514
rect 6552 19450 6604 19456
rect 6736 19508 6788 19514
rect 6736 19450 6788 19456
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 5448 19304 5500 19310
rect 5448 19246 5500 19252
rect 6368 19304 6420 19310
rect 6368 19246 6420 19252
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 5092 18970 5120 19246
rect 5724 19168 5776 19174
rect 5724 19110 5776 19116
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 5736 18630 5764 19110
rect 6380 18970 6408 19246
rect 6368 18964 6420 18970
rect 6368 18906 6420 18912
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 4289 18524 4585 18544
rect 4345 18522 4369 18524
rect 4425 18522 4449 18524
rect 4505 18522 4529 18524
rect 4367 18470 4369 18522
rect 4431 18470 4443 18522
rect 4505 18470 4507 18522
rect 4345 18468 4369 18470
rect 4425 18468 4449 18470
rect 4505 18468 4529 18470
rect 4289 18448 4585 18468
rect 4160 18284 4212 18290
rect 4160 18226 4212 18232
rect 4172 17882 4200 18226
rect 5736 18086 5764 18566
rect 5724 18080 5776 18086
rect 5724 18022 5776 18028
rect 4160 17876 4212 17882
rect 4160 17818 4212 17824
rect 4172 17202 4200 17818
rect 4289 17436 4585 17456
rect 4345 17434 4369 17436
rect 4425 17434 4449 17436
rect 4505 17434 4529 17436
rect 4367 17382 4369 17434
rect 4431 17382 4443 17434
rect 4505 17382 4507 17434
rect 4345 17380 4369 17382
rect 4425 17380 4449 17382
rect 4505 17380 4529 17382
rect 4289 17360 4585 17380
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 4172 16130 4200 17138
rect 4724 16794 4752 17138
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4289 16348 4585 16368
rect 4345 16346 4369 16348
rect 4425 16346 4449 16348
rect 4505 16346 4529 16348
rect 4367 16294 4369 16346
rect 4431 16294 4443 16346
rect 4505 16294 4507 16346
rect 4345 16292 4369 16294
rect 4425 16292 4449 16294
rect 4505 16292 4529 16294
rect 4289 16272 4585 16292
rect 4080 16102 4200 16130
rect 4080 16046 4108 16102
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 4080 15706 4108 15982
rect 4068 15700 4120 15706
rect 4120 15660 4200 15688
rect 4068 15642 4120 15648
rect 3792 15564 3844 15570
rect 3792 15506 3844 15512
rect 3804 15162 3832 15506
rect 4172 15162 4200 15660
rect 4289 15260 4585 15280
rect 4345 15258 4369 15260
rect 4425 15258 4449 15260
rect 4505 15258 4529 15260
rect 4367 15206 4369 15258
rect 4431 15206 4443 15258
rect 4505 15206 4507 15258
rect 4345 15204 4369 15206
rect 4425 15204 4449 15206
rect 4505 15204 4529 15206
rect 4289 15184 4585 15204
rect 4724 15162 4752 16594
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5080 15360 5132 15366
rect 5080 15302 5132 15308
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 4896 14952 4948 14958
rect 5092 14929 5120 15302
rect 4896 14894 4948 14900
rect 5078 14920 5134 14929
rect 3238 14648 3294 14657
rect 4908 14618 4936 14894
rect 5078 14855 5134 14864
rect 3238 14583 3294 14592
rect 4896 14612 4948 14618
rect 3252 13394 3280 14583
rect 4896 14554 4948 14560
rect 3976 14408 4028 14414
rect 3974 14376 3976 14385
rect 4028 14376 4030 14385
rect 3974 14311 4030 14320
rect 4289 14172 4585 14192
rect 4345 14170 4369 14172
rect 4425 14170 4449 14172
rect 4505 14170 4529 14172
rect 4367 14118 4369 14170
rect 4431 14118 4443 14170
rect 4505 14118 4507 14170
rect 4345 14116 4369 14118
rect 4425 14116 4449 14118
rect 4505 14116 4529 14118
rect 4289 14096 4585 14116
rect 3790 13832 3846 13841
rect 3790 13767 3846 13776
rect 2964 13388 3016 13394
rect 2964 13330 3016 13336
rect 3240 13388 3292 13394
rect 3240 13330 3292 13336
rect 2700 12986 2820 13002
rect 2976 12986 3004 13330
rect 2688 12980 2820 12986
rect 2740 12974 2820 12980
rect 2964 12980 3016 12986
rect 2688 12922 2740 12928
rect 2964 12922 3016 12928
rect 3252 12918 3280 13330
rect 3804 12986 3832 13767
rect 4908 13530 4936 14554
rect 5644 14074 5672 15846
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5736 13870 5764 18022
rect 6840 16674 6868 19654
rect 8036 19242 8064 20198
rect 8482 19544 8538 19553
rect 8482 19479 8538 19488
rect 8024 19236 8076 19242
rect 8024 19178 8076 19184
rect 7380 19168 7432 19174
rect 7380 19110 7432 19116
rect 7392 17746 7420 19110
rect 7622 19068 7918 19088
rect 7678 19066 7702 19068
rect 7758 19066 7782 19068
rect 7838 19066 7862 19068
rect 7700 19014 7702 19066
rect 7764 19014 7776 19066
rect 7838 19014 7840 19066
rect 7678 19012 7702 19014
rect 7758 19012 7782 19014
rect 7838 19012 7862 19014
rect 7622 18992 7918 19012
rect 8036 18426 8064 19178
rect 8024 18420 8076 18426
rect 8024 18362 8076 18368
rect 7622 17980 7918 18000
rect 7678 17978 7702 17980
rect 7758 17978 7782 17980
rect 7838 17978 7862 17980
rect 7700 17926 7702 17978
rect 7764 17926 7776 17978
rect 7838 17926 7840 17978
rect 7678 17924 7702 17926
rect 7758 17924 7782 17926
rect 7838 17924 7862 17926
rect 7622 17904 7918 17924
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 8024 17740 8076 17746
rect 8024 17682 8076 17688
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7576 17202 7604 17614
rect 7564 17196 7616 17202
rect 7564 17138 7616 17144
rect 8036 16998 8064 17682
rect 8024 16992 8076 16998
rect 8022 16960 8024 16969
rect 8076 16960 8078 16969
rect 7622 16892 7918 16912
rect 8022 16895 8078 16904
rect 7678 16890 7702 16892
rect 7758 16890 7782 16892
rect 7838 16890 7862 16892
rect 7700 16838 7702 16890
rect 7764 16838 7776 16890
rect 7838 16838 7840 16890
rect 7678 16836 7702 16838
rect 7758 16836 7782 16838
rect 7838 16836 7862 16838
rect 7622 16816 7918 16836
rect 6918 16688 6974 16697
rect 6840 16646 6918 16674
rect 6918 16623 6974 16632
rect 5906 16144 5962 16153
rect 5906 16079 5962 16088
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5736 13530 5764 13806
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 4620 13320 4672 13326
rect 4618 13288 4620 13297
rect 4672 13288 4674 13297
rect 4618 13223 4674 13232
rect 4289 13084 4585 13104
rect 4345 13082 4369 13084
rect 4425 13082 4449 13084
rect 4505 13082 4529 13084
rect 4367 13030 4369 13082
rect 4431 13030 4443 13082
rect 4505 13030 4507 13082
rect 4345 13028 4369 13030
rect 4425 13028 4449 13030
rect 4505 13028 4529 13030
rect 4289 13008 4585 13028
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3240 12912 3292 12918
rect 3054 12880 3110 12889
rect 3240 12854 3292 12860
rect 3054 12815 3110 12824
rect 2962 12744 3018 12753
rect 2962 12679 3018 12688
rect 2976 11898 3004 12679
rect 3068 12374 3096 12815
rect 3056 12368 3108 12374
rect 3056 12310 3108 12316
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 3344 10810 3372 12922
rect 4908 12866 4936 13466
rect 5630 13152 5686 13161
rect 5630 13087 5686 13096
rect 5644 12986 5672 13087
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 4816 12838 4936 12866
rect 4816 12782 4844 12838
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 3790 12336 3846 12345
rect 3790 12271 3792 12280
rect 3844 12271 3846 12280
rect 3792 12242 3844 12248
rect 3804 11898 3832 12242
rect 4080 12102 4108 12718
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 4080 11694 4108 12038
rect 4289 11996 4585 12016
rect 4345 11994 4369 11996
rect 4425 11994 4449 11996
rect 4505 11994 4529 11996
rect 4367 11942 4369 11994
rect 4431 11942 4443 11994
rect 4505 11942 4507 11994
rect 4345 11940 4369 11942
rect 4425 11940 4449 11942
rect 4505 11940 4529 11942
rect 4289 11920 4585 11940
rect 5828 11801 5856 12038
rect 5920 11898 5948 16079
rect 6932 15570 6960 16623
rect 7622 15804 7918 15824
rect 7678 15802 7702 15804
rect 7758 15802 7782 15804
rect 7838 15802 7862 15804
rect 7700 15750 7702 15802
rect 7764 15750 7776 15802
rect 7838 15750 7840 15802
rect 7678 15748 7702 15750
rect 7758 15748 7782 15750
rect 7838 15748 7862 15750
rect 7622 15728 7918 15748
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 7576 15162 7604 15438
rect 7668 15162 7696 15506
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7668 15042 7696 15098
rect 7484 15014 7696 15042
rect 7286 14512 7342 14521
rect 7286 14447 7342 14456
rect 7300 14074 7328 14447
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7484 13394 7512 15014
rect 7622 14716 7918 14736
rect 7678 14714 7702 14716
rect 7758 14714 7782 14716
rect 7838 14714 7862 14716
rect 7700 14662 7702 14714
rect 7764 14662 7776 14714
rect 7838 14662 7840 14714
rect 7678 14660 7702 14662
rect 7758 14660 7782 14662
rect 7838 14660 7862 14662
rect 7622 14640 7918 14660
rect 8298 13968 8354 13977
rect 8298 13903 8354 13912
rect 7622 13628 7918 13648
rect 7678 13626 7702 13628
rect 7758 13626 7782 13628
rect 7838 13626 7862 13628
rect 7700 13574 7702 13626
rect 7764 13574 7776 13626
rect 7838 13574 7840 13626
rect 7678 13572 7702 13574
rect 7758 13572 7782 13574
rect 7838 13572 7862 13574
rect 7622 13552 7918 13572
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 7484 13138 7512 13330
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 7484 13110 7604 13138
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 5814 11792 5870 11801
rect 5814 11727 5870 11736
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2056 9722 2084 10610
rect 3148 10192 3200 10198
rect 3146 10160 3148 10169
rect 3200 10160 3202 10169
rect 2228 10124 2280 10130
rect 3146 10095 3202 10104
rect 2228 10066 2280 10072
rect 2240 9722 2268 10066
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 2228 9716 2280 9722
rect 2228 9658 2280 9664
rect 1492 9172 1544 9178
rect 1492 9114 1544 9120
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 1688 5778 1716 9114
rect 3436 6769 3464 11494
rect 3792 11212 3844 11218
rect 3792 11154 3844 11160
rect 3804 11014 3832 11154
rect 3974 11112 4030 11121
rect 3974 11047 4030 11056
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3804 10810 3832 10950
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 3988 9897 4016 11047
rect 4080 11014 4108 11630
rect 6564 11558 6592 12242
rect 7012 12232 7064 12238
rect 7116 12186 7144 12854
rect 7064 12180 7144 12186
rect 7012 12174 7144 12180
rect 7024 12158 7144 12174
rect 7116 11694 7144 12158
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6564 11286 6592 11494
rect 6552 11280 6604 11286
rect 6552 11222 6604 11228
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 4080 10606 4108 10950
rect 4289 10908 4585 10928
rect 4345 10906 4369 10908
rect 4425 10906 4449 10908
rect 4505 10906 4529 10908
rect 4367 10854 4369 10906
rect 4431 10854 4443 10906
rect 4505 10854 4507 10906
rect 4345 10852 4369 10854
rect 4425 10852 4449 10854
rect 4505 10852 4529 10854
rect 4289 10832 4585 10852
rect 6932 10810 6960 11494
rect 7116 11082 7144 11630
rect 7484 11121 7512 12922
rect 7576 12918 7604 13110
rect 7852 12986 7880 13262
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7564 12912 7616 12918
rect 7564 12854 7616 12860
rect 8312 12753 8340 13903
rect 8298 12744 8354 12753
rect 8298 12679 8354 12688
rect 7622 12540 7918 12560
rect 7678 12538 7702 12540
rect 7758 12538 7782 12540
rect 7838 12538 7862 12540
rect 7700 12486 7702 12538
rect 7764 12486 7776 12538
rect 7838 12486 7840 12538
rect 7678 12484 7702 12486
rect 7758 12484 7782 12486
rect 7838 12484 7862 12486
rect 7622 12464 7918 12484
rect 8496 11898 8524 19479
rect 9232 12374 9260 27814
rect 9324 27112 9352 32302
rect 9416 31736 9444 34462
rect 9586 34439 9642 34448
rect 9600 34066 9628 34439
rect 9692 34066 9720 35040
rect 10060 35034 10088 39782
rect 10152 37874 10180 46650
rect 10244 45830 10272 49558
rect 10324 49088 10376 49094
rect 10324 49030 10376 49036
rect 10336 48686 10364 49030
rect 10324 48680 10376 48686
rect 10324 48622 10376 48628
rect 10324 48340 10376 48346
rect 10324 48282 10376 48288
rect 10232 45824 10284 45830
rect 10232 45766 10284 45772
rect 10232 45416 10284 45422
rect 10230 45384 10232 45393
rect 10284 45384 10286 45393
rect 10230 45319 10286 45328
rect 10232 44328 10284 44334
rect 10232 44270 10284 44276
rect 10244 42906 10272 44270
rect 10336 43994 10364 48282
rect 10428 48210 10456 56170
rect 10520 55876 10548 63514
rect 10612 62257 10640 65010
rect 10692 65000 10744 65006
rect 10692 64942 10744 64948
rect 10704 64841 10732 64942
rect 10690 64832 10746 64841
rect 10690 64767 10746 64776
rect 10796 64530 10824 65062
rect 10784 64524 10836 64530
rect 10784 64466 10836 64472
rect 10692 63436 10744 63442
rect 10692 63378 10744 63384
rect 10704 62966 10732 63378
rect 10692 62960 10744 62966
rect 10692 62902 10744 62908
rect 10796 62914 10824 64466
rect 10888 63016 10916 66150
rect 11348 65958 11376 66982
rect 11244 65952 11296 65958
rect 11244 65894 11296 65900
rect 11336 65952 11388 65958
rect 11336 65894 11388 65900
rect 11256 65793 11284 65894
rect 11242 65784 11298 65793
rect 11242 65719 11298 65728
rect 11336 65680 11388 65686
rect 11336 65622 11388 65628
rect 10956 65308 11252 65328
rect 11012 65306 11036 65308
rect 11092 65306 11116 65308
rect 11172 65306 11196 65308
rect 11034 65254 11036 65306
rect 11098 65254 11110 65306
rect 11172 65254 11174 65306
rect 11012 65252 11036 65254
rect 11092 65252 11116 65254
rect 11172 65252 11196 65254
rect 10956 65232 11252 65252
rect 11348 64462 11376 65622
rect 11336 64456 11388 64462
rect 11336 64398 11388 64404
rect 10956 64220 11252 64240
rect 11012 64218 11036 64220
rect 11092 64218 11116 64220
rect 11172 64218 11196 64220
rect 11034 64166 11036 64218
rect 11098 64166 11110 64218
rect 11172 64166 11174 64218
rect 11012 64164 11036 64166
rect 11092 64164 11116 64166
rect 11172 64164 11196 64166
rect 10956 64144 11252 64164
rect 11336 64048 11388 64054
rect 11336 63990 11388 63996
rect 11060 63844 11112 63850
rect 11060 63786 11112 63792
rect 11072 63730 11100 63786
rect 10980 63702 11100 63730
rect 11152 63776 11204 63782
rect 11152 63718 11204 63724
rect 10980 63374 11008 63702
rect 11164 63617 11192 63718
rect 11150 63608 11206 63617
rect 11150 63543 11206 63552
rect 10968 63368 11020 63374
rect 10968 63310 11020 63316
rect 10956 63132 11252 63152
rect 11012 63130 11036 63132
rect 11092 63130 11116 63132
rect 11172 63130 11196 63132
rect 11034 63078 11036 63130
rect 11098 63078 11110 63130
rect 11172 63078 11174 63130
rect 11012 63076 11036 63078
rect 11092 63076 11116 63078
rect 11172 63076 11196 63078
rect 10956 63056 11252 63076
rect 10888 62988 11008 63016
rect 10796 62886 10916 62914
rect 10692 62824 10744 62830
rect 10692 62766 10744 62772
rect 10598 62248 10654 62257
rect 10598 62183 10654 62192
rect 10704 62150 10732 62766
rect 10782 62656 10838 62665
rect 10782 62591 10838 62600
rect 10692 62144 10744 62150
rect 10692 62086 10744 62092
rect 10600 60648 10652 60654
rect 10600 60590 10652 60596
rect 10612 59974 10640 60590
rect 10600 59968 10652 59974
rect 10600 59910 10652 59916
rect 10612 59770 10640 59910
rect 10600 59764 10652 59770
rect 10600 59706 10652 59712
rect 10704 59650 10732 62086
rect 10796 59809 10824 62591
rect 10888 60761 10916 62886
rect 10980 62830 11008 62988
rect 10968 62824 11020 62830
rect 10968 62766 11020 62772
rect 11348 62354 11376 63990
rect 11440 63374 11468 67646
rect 11532 65550 11560 70071
rect 11612 68672 11664 68678
rect 11612 68614 11664 68620
rect 11624 68338 11652 68614
rect 11612 68332 11664 68338
rect 11612 68274 11664 68280
rect 11624 68241 11652 68274
rect 11610 68232 11666 68241
rect 11610 68167 11666 68176
rect 11612 67856 11664 67862
rect 11612 67798 11664 67804
rect 11624 67046 11652 67798
rect 11612 67040 11664 67046
rect 11612 66982 11664 66988
rect 11624 66230 11652 66982
rect 11612 66224 11664 66230
rect 11612 66166 11664 66172
rect 11612 65952 11664 65958
rect 11612 65894 11664 65900
rect 11520 65544 11572 65550
rect 11520 65486 11572 65492
rect 11624 65362 11652 65894
rect 11532 65334 11652 65362
rect 11428 63368 11480 63374
rect 11428 63310 11480 63316
rect 11532 62665 11560 65334
rect 11612 63572 11664 63578
rect 11612 63514 11664 63520
rect 11518 62656 11574 62665
rect 11518 62591 11574 62600
rect 11336 62348 11388 62354
rect 11336 62290 11388 62296
rect 10956 62044 11252 62064
rect 11012 62042 11036 62044
rect 11092 62042 11116 62044
rect 11172 62042 11196 62044
rect 11034 61990 11036 62042
rect 11098 61990 11110 62042
rect 11172 61990 11174 62042
rect 11012 61988 11036 61990
rect 11092 61988 11116 61990
rect 11172 61988 11196 61990
rect 10956 61968 11252 61988
rect 11348 61946 11376 62290
rect 11520 62280 11572 62286
rect 11520 62222 11572 62228
rect 11532 61946 11560 62222
rect 11336 61940 11388 61946
rect 11336 61882 11388 61888
rect 11520 61940 11572 61946
rect 11520 61882 11572 61888
rect 11058 61296 11114 61305
rect 11058 61231 11060 61240
rect 11112 61231 11114 61240
rect 11060 61202 11112 61208
rect 11348 61198 11376 61882
rect 11520 61600 11572 61606
rect 11520 61542 11572 61548
rect 11428 61260 11480 61266
rect 11428 61202 11480 61208
rect 11336 61192 11388 61198
rect 11336 61134 11388 61140
rect 10956 60956 11252 60976
rect 11012 60954 11036 60956
rect 11092 60954 11116 60956
rect 11172 60954 11196 60956
rect 11034 60902 11036 60954
rect 11098 60902 11110 60954
rect 11172 60902 11174 60954
rect 11012 60900 11036 60902
rect 11092 60900 11116 60902
rect 11172 60900 11196 60902
rect 10956 60880 11252 60900
rect 11440 60858 11468 61202
rect 11428 60852 11480 60858
rect 11348 60812 11428 60840
rect 10874 60752 10930 60761
rect 10874 60687 10930 60696
rect 10876 60172 10928 60178
rect 10876 60114 10928 60120
rect 10782 59800 10838 59809
rect 10782 59735 10838 59744
rect 10612 59622 10732 59650
rect 10784 59628 10836 59634
rect 10612 59226 10640 59622
rect 10784 59570 10836 59576
rect 10692 59560 10744 59566
rect 10690 59528 10692 59537
rect 10744 59528 10746 59537
rect 10690 59463 10746 59472
rect 10692 59424 10744 59430
rect 10692 59366 10744 59372
rect 10600 59220 10652 59226
rect 10600 59162 10652 59168
rect 10612 58478 10640 59162
rect 10704 59129 10732 59366
rect 10690 59120 10746 59129
rect 10690 59055 10746 59064
rect 10600 58472 10652 58478
rect 10600 58414 10652 58420
rect 10612 56914 10640 58414
rect 10704 57934 10732 59055
rect 10692 57928 10744 57934
rect 10692 57870 10744 57876
rect 10692 57792 10744 57798
rect 10692 57734 10744 57740
rect 10600 56908 10652 56914
rect 10600 56850 10652 56856
rect 10704 56137 10732 57734
rect 10690 56128 10746 56137
rect 10690 56063 10746 56072
rect 10520 55848 10732 55876
rect 10508 55752 10560 55758
rect 10508 55694 10560 55700
rect 10600 55752 10652 55758
rect 10600 55694 10652 55700
rect 10520 55418 10548 55694
rect 10508 55412 10560 55418
rect 10508 55354 10560 55360
rect 10612 54670 10640 55694
rect 10600 54664 10652 54670
rect 10600 54606 10652 54612
rect 10506 54088 10562 54097
rect 10506 54023 10562 54032
rect 10520 52426 10548 54023
rect 10612 53990 10640 54606
rect 10600 53984 10652 53990
rect 10600 53926 10652 53932
rect 10598 53680 10654 53689
rect 10598 53615 10600 53624
rect 10652 53615 10654 53624
rect 10600 53586 10652 53592
rect 10612 53242 10640 53586
rect 10600 53236 10652 53242
rect 10600 53178 10652 53184
rect 10600 52896 10652 52902
rect 10600 52838 10652 52844
rect 10612 52601 10640 52838
rect 10598 52592 10654 52601
rect 10598 52527 10654 52536
rect 10508 52420 10560 52426
rect 10508 52362 10560 52368
rect 10600 51876 10652 51882
rect 10600 51818 10652 51824
rect 10508 51536 10560 51542
rect 10508 51478 10560 51484
rect 10520 50862 10548 51478
rect 10508 50856 10560 50862
rect 10508 50798 10560 50804
rect 10520 49745 10548 50798
rect 10612 49774 10640 51818
rect 10704 50969 10732 55848
rect 10796 54738 10824 59570
rect 10888 59226 10916 60114
rect 10956 59868 11252 59888
rect 11012 59866 11036 59868
rect 11092 59866 11116 59868
rect 11172 59866 11196 59868
rect 11034 59814 11036 59866
rect 11098 59814 11110 59866
rect 11172 59814 11174 59866
rect 11012 59812 11036 59814
rect 11092 59812 11116 59814
rect 11172 59812 11196 59814
rect 10956 59792 11252 59812
rect 10876 59220 10928 59226
rect 10876 59162 10928 59168
rect 10956 58780 11252 58800
rect 11012 58778 11036 58780
rect 11092 58778 11116 58780
rect 11172 58778 11196 58780
rect 11034 58726 11036 58778
rect 11098 58726 11110 58778
rect 11172 58726 11174 58778
rect 11012 58724 11036 58726
rect 11092 58724 11116 58726
rect 11172 58724 11196 58726
rect 10956 58704 11252 58724
rect 11244 58608 11296 58614
rect 11244 58550 11296 58556
rect 11152 58132 11204 58138
rect 11152 58074 11204 58080
rect 10876 57928 10928 57934
rect 11164 57905 11192 58074
rect 10876 57870 10928 57876
rect 11150 57896 11206 57905
rect 10888 57458 10916 57870
rect 11256 57866 11284 58550
rect 11150 57831 11206 57840
rect 11244 57860 11296 57866
rect 11244 57802 11296 57808
rect 10956 57692 11252 57712
rect 11012 57690 11036 57692
rect 11092 57690 11116 57692
rect 11172 57690 11196 57692
rect 11034 57638 11036 57690
rect 11098 57638 11110 57690
rect 11172 57638 11174 57690
rect 11012 57636 11036 57638
rect 11092 57636 11116 57638
rect 11172 57636 11196 57638
rect 10956 57616 11252 57636
rect 10966 57488 11022 57497
rect 10876 57452 10928 57458
rect 10966 57423 11022 57432
rect 10876 57394 10928 57400
rect 10980 57390 11008 57423
rect 10968 57384 11020 57390
rect 10968 57326 11020 57332
rect 10956 56604 11252 56624
rect 11012 56602 11036 56604
rect 11092 56602 11116 56604
rect 11172 56602 11196 56604
rect 11034 56550 11036 56602
rect 11098 56550 11110 56602
rect 11172 56550 11174 56602
rect 11012 56548 11036 56550
rect 11092 56548 11116 56550
rect 11172 56548 11196 56550
rect 10956 56528 11252 56548
rect 11152 56296 11204 56302
rect 11152 56238 11204 56244
rect 10966 56128 11022 56137
rect 10966 56063 11022 56072
rect 10980 55962 11008 56063
rect 11164 55962 11192 56238
rect 10968 55956 11020 55962
rect 10968 55898 11020 55904
rect 11152 55956 11204 55962
rect 11152 55898 11204 55904
rect 11164 55729 11192 55898
rect 11150 55720 11206 55729
rect 10876 55684 10928 55690
rect 11150 55655 11206 55664
rect 10876 55626 10928 55632
rect 10888 55214 10916 55626
rect 10956 55516 11252 55536
rect 11012 55514 11036 55516
rect 11092 55514 11116 55516
rect 11172 55514 11196 55516
rect 11034 55462 11036 55514
rect 11098 55462 11110 55514
rect 11172 55462 11174 55514
rect 11012 55460 11036 55462
rect 11092 55460 11116 55462
rect 11172 55460 11196 55462
rect 10956 55440 11252 55460
rect 10876 55208 10928 55214
rect 10876 55150 10928 55156
rect 10784 54732 10836 54738
rect 10784 54674 10836 54680
rect 10796 54330 10824 54674
rect 10876 54528 10928 54534
rect 10876 54470 10928 54476
rect 10784 54324 10836 54330
rect 10784 54266 10836 54272
rect 10888 53718 10916 54470
rect 10956 54428 11252 54448
rect 11012 54426 11036 54428
rect 11092 54426 11116 54428
rect 11172 54426 11196 54428
rect 11034 54374 11036 54426
rect 11098 54374 11110 54426
rect 11172 54374 11174 54426
rect 11012 54372 11036 54374
rect 11092 54372 11116 54374
rect 11172 54372 11196 54374
rect 10956 54352 11252 54372
rect 10966 54224 11022 54233
rect 10966 54159 11022 54168
rect 10876 53712 10928 53718
rect 10876 53654 10928 53660
rect 10784 53644 10836 53650
rect 10784 53586 10836 53592
rect 10796 52698 10824 53586
rect 10980 53428 11008 54159
rect 11152 53984 11204 53990
rect 11152 53926 11204 53932
rect 11164 53786 11192 53926
rect 11152 53780 11204 53786
rect 11152 53722 11204 53728
rect 10888 53400 11008 53428
rect 10784 52692 10836 52698
rect 10784 52634 10836 52640
rect 10888 52562 10916 53400
rect 10956 53340 11252 53360
rect 11012 53338 11036 53340
rect 11092 53338 11116 53340
rect 11172 53338 11196 53340
rect 11034 53286 11036 53338
rect 11098 53286 11110 53338
rect 11172 53286 11174 53338
rect 11012 53284 11036 53286
rect 11092 53284 11116 53286
rect 11172 53284 11196 53286
rect 10956 53264 11252 53284
rect 11244 53168 11296 53174
rect 11244 53110 11296 53116
rect 11256 52630 11284 53110
rect 11348 52970 11376 60812
rect 11428 60794 11480 60800
rect 11428 60716 11480 60722
rect 11428 60658 11480 60664
rect 11440 58614 11468 60658
rect 11532 60081 11560 61542
rect 11518 60072 11574 60081
rect 11518 60007 11574 60016
rect 11520 59968 11572 59974
rect 11520 59910 11572 59916
rect 11428 58608 11480 58614
rect 11428 58550 11480 58556
rect 11428 58336 11480 58342
rect 11428 58278 11480 58284
rect 11440 55078 11468 58278
rect 11532 55418 11560 59910
rect 11624 59537 11652 63514
rect 11716 61606 11744 70382
rect 11796 70304 11848 70310
rect 11796 70246 11848 70252
rect 11808 69290 11836 70246
rect 11900 69426 11928 71130
rect 11980 70848 12032 70854
rect 11980 70790 12032 70796
rect 11992 70446 12020 70790
rect 11980 70440 12032 70446
rect 11980 70382 12032 70388
rect 12072 70440 12124 70446
rect 12072 70382 12124 70388
rect 11978 70000 12034 70009
rect 11978 69935 12034 69944
rect 11992 69834 12020 69935
rect 11980 69828 12032 69834
rect 11980 69770 12032 69776
rect 11888 69420 11940 69426
rect 11888 69362 11940 69368
rect 11796 69284 11848 69290
rect 11796 69226 11848 69232
rect 11796 66020 11848 66026
rect 11796 65962 11848 65968
rect 11704 61600 11756 61606
rect 11704 61542 11756 61548
rect 11808 60790 11836 65962
rect 11796 60784 11848 60790
rect 11796 60726 11848 60732
rect 11796 60648 11848 60654
rect 11796 60590 11848 60596
rect 11704 60104 11756 60110
rect 11704 60046 11756 60052
rect 11610 59528 11666 59537
rect 11610 59463 11666 59472
rect 11624 59226 11652 59463
rect 11612 59220 11664 59226
rect 11612 59162 11664 59168
rect 11612 59084 11664 59090
rect 11612 59026 11664 59032
rect 11624 58342 11652 59026
rect 11612 58336 11664 58342
rect 11612 58278 11664 58284
rect 11716 57934 11744 60046
rect 11704 57928 11756 57934
rect 11704 57870 11756 57876
rect 11612 57860 11664 57866
rect 11612 57802 11664 57808
rect 11624 57769 11652 57802
rect 11610 57760 11666 57769
rect 11610 57695 11666 57704
rect 11808 57610 11836 60590
rect 11624 57582 11836 57610
rect 11520 55412 11572 55418
rect 11520 55354 11572 55360
rect 11518 55312 11574 55321
rect 11518 55247 11520 55256
rect 11572 55247 11574 55256
rect 11520 55218 11572 55224
rect 11624 55162 11652 57582
rect 11796 57452 11848 57458
rect 11796 57394 11848 57400
rect 11704 56908 11756 56914
rect 11704 56850 11756 56856
rect 11716 56273 11744 56850
rect 11702 56264 11758 56273
rect 11702 56199 11758 56208
rect 11532 55134 11652 55162
rect 11428 55072 11480 55078
rect 11428 55014 11480 55020
rect 11428 54664 11480 54670
rect 11428 54606 11480 54612
rect 11440 53961 11468 54606
rect 11426 53952 11482 53961
rect 11426 53887 11482 53896
rect 11428 53780 11480 53786
rect 11428 53722 11480 53728
rect 11440 53242 11468 53722
rect 11428 53236 11480 53242
rect 11428 53178 11480 53184
rect 11532 53122 11560 55134
rect 11612 55072 11664 55078
rect 11612 55014 11664 55020
rect 11624 53972 11652 55014
rect 11716 54126 11744 56199
rect 11808 54874 11836 57394
rect 11900 56506 11928 69362
rect 11992 69358 12020 69770
rect 12084 69766 12112 70382
rect 12072 69760 12124 69766
rect 12072 69702 12124 69708
rect 12084 69494 12112 69702
rect 12072 69488 12124 69494
rect 12072 69430 12124 69436
rect 11980 69352 12032 69358
rect 11980 69294 12032 69300
rect 11992 69057 12020 69294
rect 11978 69048 12034 69057
rect 11978 68983 12034 68992
rect 12084 68678 12112 69430
rect 12348 69284 12400 69290
rect 12400 69244 12480 69272
rect 12348 69226 12400 69232
rect 12452 68882 12480 69244
rect 12440 68876 12492 68882
rect 12440 68818 12492 68824
rect 12072 68672 12124 68678
rect 12072 68614 12124 68620
rect 11980 67244 12032 67250
rect 11980 67186 12032 67192
rect 11992 67046 12020 67186
rect 11980 67040 12032 67046
rect 11980 66982 12032 66988
rect 11992 66774 12020 66982
rect 11980 66768 12032 66774
rect 11980 66710 12032 66716
rect 11992 66094 12020 66710
rect 11980 66088 12032 66094
rect 11980 66030 12032 66036
rect 11980 65544 12032 65550
rect 11980 65486 12032 65492
rect 11992 60722 12020 65486
rect 12084 63918 12112 68614
rect 12452 68134 12480 68818
rect 12440 68128 12492 68134
rect 12440 68070 12492 68076
rect 12164 67176 12216 67182
rect 12164 67118 12216 67124
rect 12176 66638 12204 67118
rect 12452 67114 12480 68070
rect 12256 67108 12308 67114
rect 12256 67050 12308 67056
rect 12440 67108 12492 67114
rect 12440 67050 12492 67056
rect 12164 66632 12216 66638
rect 12164 66574 12216 66580
rect 12176 64818 12204 66574
rect 12268 66502 12296 67050
rect 12440 66700 12492 66706
rect 12440 66642 12492 66648
rect 12256 66496 12308 66502
rect 12256 66438 12308 66444
rect 12268 65618 12296 66438
rect 12452 66230 12480 66642
rect 12544 66638 12572 72422
rect 12624 68672 12676 68678
rect 12624 68614 12676 68620
rect 12636 68270 12664 68614
rect 12624 68264 12676 68270
rect 12624 68206 12676 68212
rect 12532 66632 12584 66638
rect 12532 66574 12584 66580
rect 12532 66496 12584 66502
rect 12532 66438 12584 66444
rect 12440 66224 12492 66230
rect 12440 66166 12492 66172
rect 12256 65612 12308 65618
rect 12256 65554 12308 65560
rect 12452 65521 12480 66166
rect 12544 66094 12572 66438
rect 12532 66088 12584 66094
rect 12532 66030 12584 66036
rect 12544 65754 12572 66030
rect 12622 65920 12678 65929
rect 12622 65855 12678 65864
rect 12532 65748 12584 65754
rect 12532 65690 12584 65696
rect 12438 65512 12494 65521
rect 12438 65447 12494 65456
rect 12256 65408 12308 65414
rect 12256 65350 12308 65356
rect 12268 64954 12296 65350
rect 12348 65000 12400 65006
rect 12268 64948 12348 64954
rect 12268 64942 12400 64948
rect 12268 64926 12388 64942
rect 12176 64790 12296 64818
rect 12072 63912 12124 63918
rect 12072 63854 12124 63860
rect 12084 63578 12112 63854
rect 12072 63572 12124 63578
rect 12072 63514 12124 63520
rect 12164 62688 12216 62694
rect 12164 62630 12216 62636
rect 12070 62112 12126 62121
rect 12070 62047 12126 62056
rect 11980 60716 12032 60722
rect 11980 60658 12032 60664
rect 12084 60602 12112 62047
rect 11992 60574 12112 60602
rect 11992 60518 12020 60574
rect 11980 60512 12032 60518
rect 11980 60454 12032 60460
rect 11888 56500 11940 56506
rect 11888 56442 11940 56448
rect 11900 56234 11928 56442
rect 11888 56228 11940 56234
rect 11888 56170 11940 56176
rect 11888 55616 11940 55622
rect 11888 55558 11940 55564
rect 11900 55185 11928 55558
rect 11992 55214 12020 60454
rect 12176 59090 12204 62630
rect 12164 59084 12216 59090
rect 12164 59026 12216 59032
rect 12164 58540 12216 58546
rect 12164 58482 12216 58488
rect 12072 58336 12124 58342
rect 12072 58278 12124 58284
rect 12084 57050 12112 58278
rect 12072 57044 12124 57050
rect 12072 56986 12124 56992
rect 12070 56536 12126 56545
rect 12070 56471 12126 56480
rect 12084 56438 12112 56471
rect 12072 56432 12124 56438
rect 12072 56374 12124 56380
rect 12176 55962 12204 58482
rect 12268 58426 12296 64790
rect 12360 62370 12388 64926
rect 12530 64832 12586 64841
rect 12530 64767 12586 64776
rect 12544 63850 12572 64767
rect 12532 63844 12584 63850
rect 12532 63786 12584 63792
rect 12544 63442 12572 63786
rect 12532 63436 12584 63442
rect 12532 63378 12584 63384
rect 12544 62694 12572 63378
rect 12636 63034 12664 65855
rect 12728 65532 12756 72576
rect 14289 72380 14585 72400
rect 14345 72378 14369 72380
rect 14425 72378 14449 72380
rect 14505 72378 14529 72380
rect 14367 72326 14369 72378
rect 14431 72326 14443 72378
rect 14505 72326 14507 72378
rect 14345 72324 14369 72326
rect 14425 72324 14449 72326
rect 14505 72324 14529 72326
rect 14289 72304 14585 72324
rect 12808 71528 12860 71534
rect 12808 71470 12860 71476
rect 16120 71528 16172 71534
rect 16120 71470 16172 71476
rect 12820 68678 12848 71470
rect 16028 71392 16080 71398
rect 16028 71334 16080 71340
rect 14289 71292 14585 71312
rect 14345 71290 14369 71292
rect 14425 71290 14449 71292
rect 14505 71290 14529 71292
rect 14367 71238 14369 71290
rect 14431 71238 14443 71290
rect 14505 71238 14507 71290
rect 14345 71236 14369 71238
rect 14425 71236 14449 71238
rect 14505 71236 14529 71238
rect 14289 71216 14585 71236
rect 14289 70204 14585 70224
rect 14345 70202 14369 70204
rect 14425 70202 14449 70204
rect 14505 70202 14529 70204
rect 14367 70150 14369 70202
rect 14431 70150 14443 70202
rect 14505 70150 14507 70202
rect 14345 70148 14369 70150
rect 14425 70148 14449 70150
rect 14505 70148 14529 70150
rect 14289 70128 14585 70148
rect 14289 69116 14585 69136
rect 14345 69114 14369 69116
rect 14425 69114 14449 69116
rect 14505 69114 14529 69116
rect 14367 69062 14369 69114
rect 14431 69062 14443 69114
rect 14505 69062 14507 69114
rect 14345 69060 14369 69062
rect 14425 69060 14449 69062
rect 14505 69060 14529 69062
rect 14289 69040 14585 69060
rect 14096 68944 14148 68950
rect 14096 68886 14148 68892
rect 13912 68876 13964 68882
rect 13912 68818 13964 68824
rect 12808 68672 12860 68678
rect 12808 68614 12860 68620
rect 13360 68672 13412 68678
rect 13360 68614 13412 68620
rect 12820 68270 12848 68614
rect 13372 68270 13400 68614
rect 12808 68264 12860 68270
rect 12808 68206 12860 68212
rect 13176 68264 13228 68270
rect 13176 68206 13228 68212
rect 13360 68264 13412 68270
rect 13360 68206 13412 68212
rect 13450 68232 13506 68241
rect 12820 66026 12848 68206
rect 13188 67794 13216 68206
rect 13176 67788 13228 67794
rect 13176 67730 13228 67736
rect 13084 67584 13136 67590
rect 13084 67526 13136 67532
rect 12992 67176 13044 67182
rect 12912 67136 12992 67164
rect 12912 66706 12940 67136
rect 12992 67118 13044 67124
rect 12900 66700 12952 66706
rect 12900 66642 12952 66648
rect 12808 66020 12860 66026
rect 12808 65962 12860 65968
rect 12912 65958 12940 66642
rect 12992 66632 13044 66638
rect 12992 66574 13044 66580
rect 12900 65952 12952 65958
rect 12900 65894 12952 65900
rect 12728 65504 12848 65532
rect 12716 64932 12768 64938
rect 12716 64874 12768 64880
rect 12624 63028 12676 63034
rect 12624 62970 12676 62976
rect 12532 62688 12584 62694
rect 12532 62630 12584 62636
rect 12728 62490 12756 64874
rect 12716 62484 12768 62490
rect 12716 62426 12768 62432
rect 12360 62354 12480 62370
rect 12360 62348 12492 62354
rect 12360 62342 12440 62348
rect 12440 62290 12492 62296
rect 12452 62257 12480 62290
rect 12438 62248 12494 62257
rect 12438 62183 12494 62192
rect 12716 61736 12768 61742
rect 12716 61678 12768 61684
rect 12624 61668 12676 61674
rect 12624 61610 12676 61616
rect 12348 61056 12400 61062
rect 12348 60998 12400 61004
rect 12360 60738 12388 60998
rect 12438 60888 12494 60897
rect 12438 60823 12494 60832
rect 12452 60738 12480 60823
rect 12360 60710 12480 60738
rect 12452 60654 12480 60710
rect 12532 60716 12584 60722
rect 12532 60658 12584 60664
rect 12440 60648 12492 60654
rect 12440 60590 12492 60596
rect 12440 60172 12492 60178
rect 12440 60114 12492 60120
rect 12348 59492 12400 59498
rect 12348 59434 12400 59440
rect 12360 59226 12388 59434
rect 12348 59220 12400 59226
rect 12348 59162 12400 59168
rect 12452 59072 12480 60114
rect 12544 59566 12572 60658
rect 12532 59560 12584 59566
rect 12532 59502 12584 59508
rect 12452 59044 12572 59072
rect 12440 58948 12492 58954
rect 12440 58890 12492 58896
rect 12452 58478 12480 58890
rect 12440 58472 12492 58478
rect 12268 58398 12388 58426
rect 12440 58414 12492 58420
rect 12256 58336 12308 58342
rect 12256 58278 12308 58284
rect 12268 58138 12296 58278
rect 12256 58132 12308 58138
rect 12256 58074 12308 58080
rect 12256 57928 12308 57934
rect 12256 57870 12308 57876
rect 12268 57458 12296 57870
rect 12256 57452 12308 57458
rect 12256 57394 12308 57400
rect 12256 57248 12308 57254
rect 12256 57190 12308 57196
rect 12268 56710 12296 57190
rect 12256 56704 12308 56710
rect 12256 56646 12308 56652
rect 12164 55956 12216 55962
rect 12164 55898 12216 55904
rect 12176 55758 12204 55898
rect 12072 55752 12124 55758
rect 12072 55694 12124 55700
rect 12164 55752 12216 55758
rect 12164 55694 12216 55700
rect 12084 55622 12112 55694
rect 12072 55616 12124 55622
rect 12072 55558 12124 55564
rect 12084 55282 12112 55558
rect 12164 55412 12216 55418
rect 12164 55354 12216 55360
rect 12072 55276 12124 55282
rect 12072 55218 12124 55224
rect 11980 55208 12032 55214
rect 11886 55176 11942 55185
rect 11980 55150 12032 55156
rect 11886 55111 11942 55120
rect 11900 55078 11928 55111
rect 11888 55072 11940 55078
rect 11888 55014 11940 55020
rect 11796 54868 11848 54874
rect 11796 54810 11848 54816
rect 11704 54120 11756 54126
rect 11808 54108 11836 54810
rect 11980 54324 12032 54330
rect 11980 54266 12032 54272
rect 11888 54120 11940 54126
rect 11808 54080 11888 54108
rect 11704 54062 11756 54068
rect 11888 54062 11940 54068
rect 11624 53944 11744 53972
rect 11612 53644 11664 53650
rect 11612 53586 11664 53592
rect 11624 53417 11652 53586
rect 11610 53408 11666 53417
rect 11610 53343 11666 53352
rect 11440 53094 11560 53122
rect 11336 52964 11388 52970
rect 11336 52906 11388 52912
rect 11244 52624 11296 52630
rect 11244 52566 11296 52572
rect 11440 52562 11468 53094
rect 11624 53038 11652 53343
rect 11612 53032 11664 53038
rect 11612 52974 11664 52980
rect 11520 52964 11572 52970
rect 11520 52906 11572 52912
rect 10784 52556 10836 52562
rect 10784 52498 10836 52504
rect 10876 52556 10928 52562
rect 10876 52498 10928 52504
rect 11428 52556 11480 52562
rect 11428 52498 11480 52504
rect 10796 51814 10824 52498
rect 10888 52154 10916 52498
rect 11426 52456 11482 52465
rect 11426 52391 11482 52400
rect 10956 52252 11252 52272
rect 11012 52250 11036 52252
rect 11092 52250 11116 52252
rect 11172 52250 11196 52252
rect 11034 52198 11036 52250
rect 11098 52198 11110 52250
rect 11172 52198 11174 52250
rect 11012 52196 11036 52198
rect 11092 52196 11116 52198
rect 11172 52196 11196 52198
rect 10956 52176 11252 52196
rect 10876 52148 10928 52154
rect 11336 52148 11388 52154
rect 10928 52108 11100 52136
rect 10876 52090 10928 52096
rect 10876 51944 10928 51950
rect 10876 51886 10928 51892
rect 10784 51808 10836 51814
rect 10784 51750 10836 51756
rect 10888 51626 10916 51886
rect 10968 51876 11020 51882
rect 10968 51818 11020 51824
rect 10796 51598 10916 51626
rect 10980 51610 11008 51818
rect 10968 51604 11020 51610
rect 10796 51252 10824 51598
rect 10968 51546 11020 51552
rect 11072 51513 11100 52108
rect 11336 52090 11388 52096
rect 11244 52080 11296 52086
rect 11244 52022 11296 52028
rect 11058 51504 11114 51513
rect 10968 51468 11020 51474
rect 11058 51439 11114 51448
rect 10968 51410 11020 51416
rect 10980 51377 11008 51410
rect 10966 51368 11022 51377
rect 11256 51354 11284 52022
rect 11348 51610 11376 52090
rect 11440 51950 11468 52391
rect 11428 51944 11480 51950
rect 11428 51886 11480 51892
rect 11428 51808 11480 51814
rect 11428 51750 11480 51756
rect 11336 51604 11388 51610
rect 11336 51546 11388 51552
rect 11334 51504 11390 51513
rect 11334 51439 11336 51448
rect 11388 51439 11390 51448
rect 11336 51410 11388 51416
rect 11256 51326 11376 51354
rect 10966 51303 11022 51312
rect 10796 51224 10916 51252
rect 10782 51096 10838 51105
rect 10782 51031 10838 51040
rect 10690 50960 10746 50969
rect 10690 50895 10746 50904
rect 10692 50788 10744 50794
rect 10692 50730 10744 50736
rect 10600 49768 10652 49774
rect 10506 49736 10562 49745
rect 10600 49710 10652 49716
rect 10506 49671 10562 49680
rect 10508 49632 10560 49638
rect 10508 49574 10560 49580
rect 10520 48890 10548 49574
rect 10704 49366 10732 50730
rect 10796 50522 10824 51031
rect 10784 50516 10836 50522
rect 10784 50458 10836 50464
rect 10784 50176 10836 50182
rect 10784 50118 10836 50124
rect 10796 49774 10824 50118
rect 10784 49768 10836 49774
rect 10784 49710 10836 49716
rect 10600 49360 10652 49366
rect 10598 49328 10600 49337
rect 10692 49360 10744 49366
rect 10652 49328 10654 49337
rect 10692 49302 10744 49308
rect 10598 49263 10654 49272
rect 10612 48890 10640 49263
rect 10692 49156 10744 49162
rect 10692 49098 10744 49104
rect 10508 48884 10560 48890
rect 10508 48826 10560 48832
rect 10600 48884 10652 48890
rect 10600 48826 10652 48832
rect 10600 48748 10652 48754
rect 10520 48708 10600 48736
rect 10520 48210 10548 48708
rect 10600 48690 10652 48696
rect 10704 48346 10732 49098
rect 10692 48340 10744 48346
rect 10692 48282 10744 48288
rect 10416 48204 10468 48210
rect 10416 48146 10468 48152
rect 10508 48204 10560 48210
rect 10508 48146 10560 48152
rect 10692 48204 10744 48210
rect 10692 48146 10744 48152
rect 10428 47802 10456 48146
rect 10416 47796 10468 47802
rect 10416 47738 10468 47744
rect 10520 47462 10548 48146
rect 10600 48068 10652 48074
rect 10600 48010 10652 48016
rect 10612 47598 10640 48010
rect 10600 47592 10652 47598
rect 10600 47534 10652 47540
rect 10508 47456 10560 47462
rect 10508 47398 10560 47404
rect 10416 46028 10468 46034
rect 10416 45970 10468 45976
rect 10428 45558 10456 45970
rect 10416 45552 10468 45558
rect 10416 45494 10468 45500
rect 10324 43988 10376 43994
rect 10324 43930 10376 43936
rect 10322 43888 10378 43897
rect 10322 43823 10324 43832
rect 10376 43823 10378 43832
rect 10324 43794 10376 43800
rect 10416 43784 10468 43790
rect 10416 43726 10468 43732
rect 10324 43240 10376 43246
rect 10324 43182 10376 43188
rect 10232 42900 10284 42906
rect 10232 42842 10284 42848
rect 10230 42800 10286 42809
rect 10230 42735 10232 42744
rect 10284 42735 10286 42744
rect 10232 42706 10284 42712
rect 10230 42664 10286 42673
rect 10230 42599 10286 42608
rect 10244 42362 10272 42599
rect 10232 42356 10284 42362
rect 10232 42298 10284 42304
rect 10244 42158 10272 42298
rect 10232 42152 10284 42158
rect 10232 42094 10284 42100
rect 10244 41138 10272 42094
rect 10336 41818 10364 43182
rect 10428 42945 10456 43726
rect 10414 42936 10470 42945
rect 10414 42871 10470 42880
rect 10520 42786 10548 47398
rect 10600 47116 10652 47122
rect 10600 47058 10652 47064
rect 10612 46714 10640 47058
rect 10704 46986 10732 48146
rect 10796 48006 10824 49710
rect 10784 48000 10836 48006
rect 10784 47942 10836 47948
rect 10692 46980 10744 46986
rect 10692 46922 10744 46928
rect 10600 46708 10652 46714
rect 10600 46650 10652 46656
rect 10704 46594 10732 46922
rect 10428 42758 10548 42786
rect 10612 46566 10732 46594
rect 10324 41812 10376 41818
rect 10324 41754 10376 41760
rect 10232 41132 10284 41138
rect 10232 41074 10284 41080
rect 10336 41070 10364 41754
rect 10324 41064 10376 41070
rect 10324 41006 10376 41012
rect 10324 40928 10376 40934
rect 10324 40870 10376 40876
rect 10336 40633 10364 40870
rect 10322 40624 10378 40633
rect 10322 40559 10324 40568
rect 10376 40559 10378 40568
rect 10324 40530 10376 40536
rect 10232 40112 10284 40118
rect 10232 40054 10284 40060
rect 10244 39030 10272 40054
rect 10322 39128 10378 39137
rect 10322 39063 10324 39072
rect 10376 39063 10378 39072
rect 10324 39034 10376 39040
rect 10232 39024 10284 39030
rect 10428 38978 10456 42758
rect 10508 42628 10560 42634
rect 10508 42570 10560 42576
rect 10232 38966 10284 38972
rect 10336 38950 10456 38978
rect 10232 38888 10284 38894
rect 10232 38830 10284 38836
rect 10140 37868 10192 37874
rect 10140 37810 10192 37816
rect 10152 36854 10180 37810
rect 10244 36922 10272 38830
rect 10232 36916 10284 36922
rect 10232 36858 10284 36864
rect 10140 36848 10192 36854
rect 10140 36790 10192 36796
rect 10232 36780 10284 36786
rect 10232 36722 10284 36728
rect 10140 36712 10192 36718
rect 10140 36654 10192 36660
rect 9968 35006 10088 35034
rect 9772 34944 9824 34950
rect 9772 34886 9824 34892
rect 9784 34542 9812 34886
rect 9772 34536 9824 34542
rect 9772 34478 9824 34484
rect 9588 34060 9640 34066
rect 9588 34002 9640 34008
rect 9680 34060 9732 34066
rect 9680 34002 9732 34008
rect 9600 33386 9628 34002
rect 9680 33924 9732 33930
rect 9680 33866 9732 33872
rect 9588 33380 9640 33386
rect 9588 33322 9640 33328
rect 9692 32994 9720 33866
rect 9600 32978 9720 32994
rect 9588 32972 9720 32978
rect 9640 32966 9720 32972
rect 9588 32914 9640 32920
rect 9600 32026 9628 32914
rect 9784 32858 9812 34478
rect 9968 33318 9996 35006
rect 10048 34060 10100 34066
rect 10048 34002 10100 34008
rect 10060 33658 10088 34002
rect 10048 33652 10100 33658
rect 10048 33594 10100 33600
rect 9956 33312 10008 33318
rect 9956 33254 10008 33260
rect 9864 33040 9916 33046
rect 9862 33008 9864 33017
rect 9916 33008 9918 33017
rect 9862 32943 9918 32952
rect 9692 32830 9812 32858
rect 9864 32904 9916 32910
rect 9864 32846 9916 32852
rect 9588 32020 9640 32026
rect 9588 31962 9640 31968
rect 9416 31708 9628 31736
rect 9496 31272 9548 31278
rect 9494 31240 9496 31249
rect 9548 31240 9550 31249
rect 9494 31175 9550 31184
rect 9496 29708 9548 29714
rect 9496 29650 9548 29656
rect 9404 29504 9456 29510
rect 9404 29446 9456 29452
rect 9416 28218 9444 29446
rect 9508 29306 9536 29650
rect 9496 29300 9548 29306
rect 9496 29242 9548 29248
rect 9508 29102 9536 29242
rect 9496 29096 9548 29102
rect 9496 29038 9548 29044
rect 9404 28212 9456 28218
rect 9404 28154 9456 28160
rect 9324 27084 9444 27112
rect 9310 26480 9366 26489
rect 9310 26415 9312 26424
rect 9364 26415 9366 26424
rect 9312 26386 9364 26392
rect 9324 26042 9352 26386
rect 9312 26036 9364 26042
rect 9312 25978 9364 25984
rect 9416 25362 9444 27084
rect 9494 25664 9550 25673
rect 9494 25599 9550 25608
rect 9508 25498 9536 25599
rect 9496 25492 9548 25498
rect 9496 25434 9548 25440
rect 9404 25356 9456 25362
rect 9324 25316 9404 25344
rect 9324 17814 9352 25316
rect 9404 25298 9456 25304
rect 9496 22976 9548 22982
rect 9496 22918 9548 22924
rect 9508 22642 9536 22918
rect 9496 22636 9548 22642
rect 9496 22578 9548 22584
rect 9404 20528 9456 20534
rect 9402 20496 9404 20505
rect 9456 20496 9458 20505
rect 9402 20431 9458 20440
rect 9312 17808 9364 17814
rect 9312 17750 9364 17756
rect 9402 17776 9458 17785
rect 9402 17711 9458 17720
rect 9416 17338 9444 17711
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9494 13424 9550 13433
rect 9494 13359 9496 13368
rect 9548 13359 9550 13368
rect 9496 13330 9548 13336
rect 9494 13016 9550 13025
rect 9494 12951 9550 12960
rect 9220 12368 9272 12374
rect 9220 12310 9272 12316
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 7622 11452 7918 11472
rect 7678 11450 7702 11452
rect 7758 11450 7782 11452
rect 7838 11450 7862 11452
rect 7700 11398 7702 11450
rect 7764 11398 7776 11450
rect 7838 11398 7840 11450
rect 7678 11396 7702 11398
rect 7758 11396 7782 11398
rect 7838 11396 7862 11398
rect 7622 11376 7918 11396
rect 8114 11384 8170 11393
rect 8114 11319 8116 11328
rect 8168 11319 8170 11328
rect 8116 11290 8168 11296
rect 7470 11112 7526 11121
rect 7104 11076 7156 11082
rect 7470 11047 7526 11056
rect 7104 11018 7156 11024
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4264 10266 4292 10610
rect 8128 10606 8156 11290
rect 8758 10704 8814 10713
rect 8758 10639 8760 10648
rect 8812 10639 8814 10648
rect 8760 10610 8812 10616
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 8024 10600 8076 10606
rect 8024 10542 8076 10548
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4448 10198 4476 10542
rect 8036 10470 8064 10542
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 7622 10364 7918 10384
rect 7678 10362 7702 10364
rect 7758 10362 7782 10364
rect 7838 10362 7862 10364
rect 7700 10310 7702 10362
rect 7764 10310 7776 10362
rect 7838 10310 7840 10362
rect 7678 10308 7702 10310
rect 7758 10308 7782 10310
rect 7838 10308 7862 10310
rect 7622 10288 7918 10308
rect 4436 10192 4488 10198
rect 4436 10134 4488 10140
rect 7840 9920 7892 9926
rect 3974 9888 4030 9897
rect 8036 9908 8064 10406
rect 8114 10296 8170 10305
rect 8114 10231 8170 10240
rect 8128 10198 8156 10231
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 7892 9880 8064 9908
rect 7840 9862 7892 9868
rect 3974 9823 4030 9832
rect 4289 9820 4585 9840
rect 4345 9818 4369 9820
rect 4425 9818 4449 9820
rect 4505 9818 4529 9820
rect 4367 9766 4369 9818
rect 4431 9766 4443 9818
rect 4505 9766 4507 9818
rect 4345 9764 4369 9766
rect 4425 9764 4449 9766
rect 4505 9764 4529 9766
rect 4289 9744 4585 9764
rect 7852 9518 7880 9862
rect 8128 9722 8156 10134
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 7840 9512 7892 9518
rect 7838 9480 7840 9489
rect 7892 9480 7894 9489
rect 7838 9415 7894 9424
rect 8220 9382 8248 10066
rect 8404 9722 8432 10542
rect 8482 10432 8538 10441
rect 8482 10367 8538 10376
rect 8496 10198 8524 10367
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8208 9376 8260 9382
rect 8576 9376 8628 9382
rect 8208 9318 8260 9324
rect 8574 9344 8576 9353
rect 8628 9344 8630 9353
rect 7622 9276 7918 9296
rect 8574 9279 8630 9288
rect 7678 9274 7702 9276
rect 7758 9274 7782 9276
rect 7838 9274 7862 9276
rect 7700 9222 7702 9274
rect 7764 9222 7776 9274
rect 7838 9222 7840 9274
rect 7678 9220 7702 9222
rect 7758 9220 7782 9222
rect 7838 9220 7862 9222
rect 7622 9200 7918 9220
rect 4289 8732 4585 8752
rect 4345 8730 4369 8732
rect 4425 8730 4449 8732
rect 4505 8730 4529 8732
rect 4367 8678 4369 8730
rect 4431 8678 4443 8730
rect 4505 8678 4507 8730
rect 4345 8676 4369 8678
rect 4425 8676 4449 8678
rect 4505 8676 4529 8678
rect 4289 8656 4585 8676
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 7622 8188 7918 8208
rect 7678 8186 7702 8188
rect 7758 8186 7782 8188
rect 7838 8186 7862 8188
rect 7700 8134 7702 8186
rect 7764 8134 7776 8186
rect 7838 8134 7840 8186
rect 7678 8132 7702 8134
rect 7758 8132 7782 8134
rect 7838 8132 7862 8134
rect 7622 8112 7918 8132
rect 8772 7970 8800 8434
rect 8680 7954 8800 7970
rect 8680 7948 8812 7954
rect 8680 7942 8760 7948
rect 4289 7644 4585 7664
rect 4345 7642 4369 7644
rect 4425 7642 4449 7644
rect 4505 7642 4529 7644
rect 4367 7590 4369 7642
rect 4431 7590 4443 7642
rect 4505 7590 4507 7642
rect 4345 7588 4369 7590
rect 4425 7588 4449 7590
rect 4505 7588 4529 7590
rect 4289 7568 4585 7588
rect 8680 7546 8708 7942
rect 8760 7890 8812 7896
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8864 7834 8892 7890
rect 8772 7806 8892 7834
rect 8942 7848 8998 7857
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8772 7478 8800 7806
rect 8942 7783 8998 7792
rect 8760 7472 8812 7478
rect 8758 7440 8760 7449
rect 8812 7440 8814 7449
rect 8758 7375 8814 7384
rect 5632 7336 5684 7342
rect 5722 7304 5778 7313
rect 5684 7284 5722 7290
rect 5632 7278 5722 7284
rect 5644 7262 5722 7278
rect 5722 7239 5778 7248
rect 7288 7268 7340 7274
rect 5540 7200 5592 7206
rect 4066 7168 4122 7177
rect 4066 7103 4122 7112
rect 5538 7168 5540 7177
rect 5592 7168 5594 7177
rect 5538 7103 5594 7112
rect 3422 6760 3478 6769
rect 3422 6695 3478 6704
rect 4080 5953 4108 7103
rect 5736 7002 5764 7239
rect 7288 7210 7340 7216
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 7300 6769 7328 7210
rect 7622 7100 7918 7120
rect 7678 7098 7702 7100
rect 7758 7098 7782 7100
rect 7838 7098 7862 7100
rect 7700 7046 7702 7098
rect 7764 7046 7776 7098
rect 7838 7046 7840 7098
rect 7678 7044 7702 7046
rect 7758 7044 7782 7046
rect 7838 7044 7862 7046
rect 7622 7024 7918 7044
rect 7286 6760 7342 6769
rect 7286 6695 7342 6704
rect 4289 6556 4585 6576
rect 4345 6554 4369 6556
rect 4425 6554 4449 6556
rect 4505 6554 4529 6556
rect 4367 6502 4369 6554
rect 4431 6502 4443 6554
rect 4505 6502 4507 6554
rect 4345 6500 4369 6502
rect 4425 6500 4449 6502
rect 4505 6500 4529 6502
rect 4289 6480 4585 6500
rect 7622 6012 7918 6032
rect 7678 6010 7702 6012
rect 7758 6010 7782 6012
rect 7838 6010 7862 6012
rect 7700 5958 7702 6010
rect 7764 5958 7776 6010
rect 7838 5958 7840 6010
rect 7678 5956 7702 5958
rect 7758 5956 7782 5958
rect 7838 5956 7862 5958
rect 4066 5944 4122 5953
rect 7622 5936 7918 5956
rect 4066 5879 4122 5888
rect 8956 5846 8984 7783
rect 8944 5840 8996 5846
rect 3790 5808 3846 5817
rect 1676 5772 1728 5778
rect 1676 5714 1728 5720
rect 2228 5772 2280 5778
rect 8944 5782 8996 5788
rect 7380 5772 7432 5778
rect 3790 5743 3792 5752
rect 2228 5714 2280 5720
rect 3844 5743 3846 5752
rect 3792 5714 3844 5720
rect 7300 5732 7380 5760
rect 1688 5370 1716 5714
rect 2240 5658 2268 5714
rect 2148 5630 2268 5658
rect 1676 5364 1728 5370
rect 1676 5306 1728 5312
rect 1688 4826 1716 5306
rect 2148 5166 2176 5630
rect 4289 5468 4585 5488
rect 4345 5466 4369 5468
rect 4425 5466 4449 5468
rect 4505 5466 4529 5468
rect 4367 5414 4369 5466
rect 4431 5414 4443 5466
rect 4505 5414 4507 5466
rect 4345 5412 4369 5414
rect 4425 5412 4449 5414
rect 4505 5412 4529 5414
rect 4289 5392 4585 5412
rect 2136 5160 2188 5166
rect 2134 5128 2136 5137
rect 2188 5128 2190 5137
rect 2134 5063 2190 5072
rect 7300 5030 7328 5732
rect 7380 5714 7432 5720
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7760 5370 7788 5646
rect 7748 5364 7800 5370
rect 7748 5306 7800 5312
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 1400 4820 1452 4826
rect 1400 4762 1452 4768
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1412 4146 1440 4762
rect 4066 4720 4122 4729
rect 4066 4655 4122 4664
rect 3054 4584 3110 4593
rect 3054 4519 3110 4528
rect 1674 4312 1730 4321
rect 1674 4247 1730 4256
rect 1688 4146 1716 4247
rect 3068 4146 3096 4519
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 1688 3738 1716 4082
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 4080 3505 4108 4655
rect 4289 4380 4585 4400
rect 4345 4378 4369 4380
rect 4425 4378 4449 4380
rect 4505 4378 4529 4380
rect 4367 4326 4369 4378
rect 4431 4326 4443 4378
rect 4505 4326 4507 4378
rect 4345 4324 4369 4326
rect 4425 4324 4449 4326
rect 4505 4324 4529 4326
rect 4289 4304 4585 4324
rect 4066 3496 4122 3505
rect 4066 3431 4122 3440
rect 4289 3292 4585 3312
rect 4345 3290 4369 3292
rect 4425 3290 4449 3292
rect 4505 3290 4529 3292
rect 4367 3238 4369 3290
rect 4431 3238 4443 3290
rect 4505 3238 4507 3290
rect 4345 3236 4369 3238
rect 4425 3236 4449 3238
rect 4505 3236 4529 3238
rect 4289 3216 4585 3236
rect 7300 2689 7328 4966
rect 7622 4924 7918 4944
rect 7678 4922 7702 4924
rect 7758 4922 7782 4924
rect 7838 4922 7862 4924
rect 7700 4870 7702 4922
rect 7764 4870 7776 4922
rect 7838 4870 7840 4922
rect 7678 4868 7702 4870
rect 7758 4868 7782 4870
rect 7838 4868 7862 4870
rect 7622 4848 7918 4868
rect 7622 3836 7918 3856
rect 7678 3834 7702 3836
rect 7758 3834 7782 3836
rect 7838 3834 7862 3836
rect 7700 3782 7702 3834
rect 7764 3782 7776 3834
rect 7838 3782 7840 3834
rect 7678 3780 7702 3782
rect 7758 3780 7782 3782
rect 7838 3780 7862 3782
rect 7622 3760 7918 3780
rect 7622 2748 7918 2768
rect 7678 2746 7702 2748
rect 7758 2746 7782 2748
rect 7838 2746 7862 2748
rect 7700 2694 7702 2746
rect 7764 2694 7776 2746
rect 7838 2694 7840 2746
rect 7678 2692 7702 2694
rect 7758 2692 7782 2694
rect 7838 2692 7862 2694
rect 7286 2680 7342 2689
rect 7622 2672 7918 2692
rect 7286 2615 7342 2624
rect 3422 2544 3478 2553
rect 3422 2479 3478 2488
rect 3436 1873 3464 2479
rect 4289 2204 4585 2224
rect 4345 2202 4369 2204
rect 4425 2202 4449 2204
rect 4505 2202 4529 2204
rect 4367 2150 4369 2202
rect 4431 2150 4443 2202
rect 4505 2150 4507 2202
rect 4345 2148 4369 2150
rect 4425 2148 4449 2150
rect 4505 2148 4529 2150
rect 4289 2128 4585 2148
rect 3422 1864 3478 1873
rect 3422 1799 3478 1808
rect 9324 377 9352 11698
rect 9402 10568 9458 10577
rect 9402 10503 9404 10512
rect 9456 10503 9458 10512
rect 9404 10474 9456 10480
rect 9508 10062 9536 12951
rect 9600 11762 9628 31708
rect 9692 22250 9720 32830
rect 9772 32768 9824 32774
rect 9772 32710 9824 32716
rect 9784 25838 9812 32710
rect 9876 32026 9904 32846
rect 9968 32774 9996 33254
rect 10046 32872 10102 32881
rect 10046 32807 10102 32816
rect 9956 32768 10008 32774
rect 9956 32710 10008 32716
rect 9864 32020 9916 32026
rect 9916 31980 9996 32008
rect 9864 31962 9916 31968
rect 9864 31748 9916 31754
rect 9864 31690 9916 31696
rect 9876 31278 9904 31690
rect 9968 31278 9996 31980
rect 9864 31272 9916 31278
rect 9864 31214 9916 31220
rect 9956 31272 10008 31278
rect 9956 31214 10008 31220
rect 9876 30938 9904 31214
rect 9956 31136 10008 31142
rect 9956 31078 10008 31084
rect 9864 30932 9916 30938
rect 9864 30874 9916 30880
rect 9864 25900 9916 25906
rect 9864 25842 9916 25848
rect 9772 25832 9824 25838
rect 9772 25774 9824 25780
rect 9876 25294 9904 25842
rect 9864 25288 9916 25294
rect 9864 25230 9916 25236
rect 9876 24886 9904 25230
rect 9864 24880 9916 24886
rect 9864 24822 9916 24828
rect 9864 24132 9916 24138
rect 9864 24074 9916 24080
rect 9770 24032 9826 24041
rect 9770 23967 9826 23976
rect 9784 22438 9812 23967
rect 9876 22506 9904 24074
rect 9968 23186 9996 31078
rect 10060 25430 10088 32807
rect 10152 29714 10180 36654
rect 10244 34066 10272 36722
rect 10232 34060 10284 34066
rect 10232 34002 10284 34008
rect 10336 33046 10364 38950
rect 10416 38888 10468 38894
rect 10416 38830 10468 38836
rect 10428 38350 10456 38830
rect 10520 38729 10548 42570
rect 10612 38962 10640 46566
rect 10784 46164 10836 46170
rect 10784 46106 10836 46112
rect 10692 46096 10744 46102
rect 10690 46064 10692 46073
rect 10744 46064 10746 46073
rect 10690 45999 10746 46008
rect 10796 45626 10824 46106
rect 10888 46102 10916 51224
rect 10956 51164 11252 51184
rect 11012 51162 11036 51164
rect 11092 51162 11116 51164
rect 11172 51162 11196 51164
rect 11034 51110 11036 51162
rect 11098 51110 11110 51162
rect 11172 51110 11174 51162
rect 11012 51108 11036 51110
rect 11092 51108 11116 51110
rect 11172 51108 11196 51110
rect 10956 51088 11252 51108
rect 10966 50960 11022 50969
rect 10966 50895 11022 50904
rect 10980 50425 11008 50895
rect 11244 50856 11296 50862
rect 11244 50798 11296 50804
rect 11256 50522 11284 50798
rect 11244 50516 11296 50522
rect 11244 50458 11296 50464
rect 10966 50416 11022 50425
rect 10966 50351 10968 50360
rect 11020 50351 11022 50360
rect 10968 50322 11020 50328
rect 10980 50291 11008 50322
rect 10956 50076 11252 50096
rect 11012 50074 11036 50076
rect 11092 50074 11116 50076
rect 11172 50074 11196 50076
rect 11034 50022 11036 50074
rect 11098 50022 11110 50074
rect 11172 50022 11174 50074
rect 11012 50020 11036 50022
rect 11092 50020 11116 50022
rect 11172 50020 11196 50022
rect 10956 50000 11252 50020
rect 10966 49872 11022 49881
rect 10966 49807 11022 49816
rect 11060 49836 11112 49842
rect 10980 49162 11008 49807
rect 11060 49778 11112 49784
rect 11072 49434 11100 49778
rect 11060 49428 11112 49434
rect 11060 49370 11112 49376
rect 10968 49156 11020 49162
rect 10968 49098 11020 49104
rect 10956 48988 11252 49008
rect 11012 48986 11036 48988
rect 11092 48986 11116 48988
rect 11172 48986 11196 48988
rect 11034 48934 11036 48986
rect 11098 48934 11110 48986
rect 11172 48934 11174 48986
rect 11012 48932 11036 48934
rect 11092 48932 11116 48934
rect 11172 48932 11196 48934
rect 10956 48912 11252 48932
rect 11060 48816 11112 48822
rect 10966 48784 11022 48793
rect 11060 48758 11112 48764
rect 10966 48719 11022 48728
rect 10980 48686 11008 48719
rect 10968 48680 11020 48686
rect 10968 48622 11020 48628
rect 11072 48142 11100 48758
rect 11244 48680 11296 48686
rect 11242 48648 11244 48657
rect 11296 48648 11298 48657
rect 11242 48583 11298 48592
rect 11256 48346 11284 48583
rect 11244 48340 11296 48346
rect 11244 48282 11296 48288
rect 11060 48136 11112 48142
rect 11060 48078 11112 48084
rect 10956 47900 11252 47920
rect 11012 47898 11036 47900
rect 11092 47898 11116 47900
rect 11172 47898 11196 47900
rect 11034 47846 11036 47898
rect 11098 47846 11110 47898
rect 11172 47846 11174 47898
rect 11012 47844 11036 47846
rect 11092 47844 11116 47846
rect 11172 47844 11196 47846
rect 10956 47824 11252 47844
rect 10966 47696 11022 47705
rect 10966 47631 11022 47640
rect 10980 47122 11008 47631
rect 10968 47116 11020 47122
rect 10968 47058 11020 47064
rect 10956 46812 11252 46832
rect 11012 46810 11036 46812
rect 11092 46810 11116 46812
rect 11172 46810 11196 46812
rect 11034 46758 11036 46810
rect 11098 46758 11110 46810
rect 11172 46758 11174 46810
rect 11012 46756 11036 46758
rect 11092 46756 11116 46758
rect 11172 46756 11196 46758
rect 10956 46736 11252 46756
rect 10968 46640 11020 46646
rect 10968 46582 11020 46588
rect 10876 46096 10928 46102
rect 10876 46038 10928 46044
rect 10980 45812 11008 46582
rect 10888 45784 11008 45812
rect 10784 45620 10836 45626
rect 10888 45608 10916 45784
rect 10956 45724 11252 45744
rect 11012 45722 11036 45724
rect 11092 45722 11116 45724
rect 11172 45722 11196 45724
rect 11034 45670 11036 45722
rect 11098 45670 11110 45722
rect 11172 45670 11174 45722
rect 11012 45668 11036 45670
rect 11092 45668 11116 45670
rect 11172 45668 11196 45670
rect 10956 45648 11252 45668
rect 10888 45580 11008 45608
rect 10784 45562 10836 45568
rect 10692 45552 10744 45558
rect 10692 45494 10744 45500
rect 10704 43330 10732 45494
rect 10796 43450 10824 45562
rect 10874 45520 10930 45529
rect 10874 45455 10930 45464
rect 10888 44946 10916 45455
rect 10876 44940 10928 44946
rect 10876 44882 10928 44888
rect 10888 44441 10916 44882
rect 10980 44810 11008 45580
rect 10968 44804 11020 44810
rect 10968 44746 11020 44752
rect 10956 44636 11252 44656
rect 11012 44634 11036 44636
rect 11092 44634 11116 44636
rect 11172 44634 11196 44636
rect 11034 44582 11036 44634
rect 11098 44582 11110 44634
rect 11172 44582 11174 44634
rect 11012 44580 11036 44582
rect 11092 44580 11116 44582
rect 11172 44580 11196 44582
rect 10956 44560 11252 44580
rect 10874 44432 10930 44441
rect 10874 44367 10930 44376
rect 10876 44328 10928 44334
rect 10876 44270 10928 44276
rect 10784 43444 10836 43450
rect 10888 43432 10916 44270
rect 10956 43548 11252 43568
rect 11012 43546 11036 43548
rect 11092 43546 11116 43548
rect 11172 43546 11196 43548
rect 11034 43494 11036 43546
rect 11098 43494 11110 43546
rect 11172 43494 11174 43546
rect 11012 43492 11036 43494
rect 11092 43492 11116 43494
rect 11172 43492 11196 43494
rect 10956 43472 11252 43492
rect 10888 43404 11008 43432
rect 10784 43386 10836 43392
rect 10704 43302 10916 43330
rect 10784 43172 10836 43178
rect 10784 43114 10836 43120
rect 10796 42838 10824 43114
rect 10784 42832 10836 42838
rect 10784 42774 10836 42780
rect 10692 42764 10744 42770
rect 10692 42706 10744 42712
rect 10704 42566 10732 42706
rect 10782 42664 10838 42673
rect 10782 42599 10784 42608
rect 10836 42599 10838 42608
rect 10784 42570 10836 42576
rect 10692 42560 10744 42566
rect 10692 42502 10744 42508
rect 10704 42362 10732 42502
rect 10692 42356 10744 42362
rect 10692 42298 10744 42304
rect 10692 42152 10744 42158
rect 10692 42094 10744 42100
rect 10704 41664 10732 42094
rect 10796 41818 10824 42570
rect 10784 41812 10836 41818
rect 10784 41754 10836 41760
rect 10704 41636 10824 41664
rect 10796 41018 10824 41636
rect 10704 40990 10824 41018
rect 10888 41002 10916 43302
rect 10980 42809 11008 43404
rect 10966 42800 11022 42809
rect 10966 42735 11022 42744
rect 10956 42460 11252 42480
rect 11012 42458 11036 42460
rect 11092 42458 11116 42460
rect 11172 42458 11196 42460
rect 11034 42406 11036 42458
rect 11098 42406 11110 42458
rect 11172 42406 11174 42458
rect 11012 42404 11036 42406
rect 11092 42404 11116 42406
rect 11172 42404 11196 42406
rect 10956 42384 11252 42404
rect 10956 41372 11252 41392
rect 11012 41370 11036 41372
rect 11092 41370 11116 41372
rect 11172 41370 11196 41372
rect 11034 41318 11036 41370
rect 11098 41318 11110 41370
rect 11172 41318 11174 41370
rect 11012 41316 11036 41318
rect 11092 41316 11116 41318
rect 11172 41316 11196 41318
rect 10956 41296 11252 41316
rect 10876 40996 10928 41002
rect 10600 38956 10652 38962
rect 10600 38898 10652 38904
rect 10600 38820 10652 38826
rect 10600 38762 10652 38768
rect 10506 38720 10562 38729
rect 10506 38655 10562 38664
rect 10508 38548 10560 38554
rect 10508 38490 10560 38496
rect 10520 38457 10548 38490
rect 10506 38448 10562 38457
rect 10506 38383 10562 38392
rect 10416 38344 10468 38350
rect 10416 38286 10468 38292
rect 10416 38208 10468 38214
rect 10416 38150 10468 38156
rect 10428 37942 10456 38150
rect 10416 37936 10468 37942
rect 10416 37878 10468 37884
rect 10416 37664 10468 37670
rect 10416 37606 10468 37612
rect 10324 33040 10376 33046
rect 10230 33008 10286 33017
rect 10324 32982 10376 32988
rect 10230 32943 10232 32952
rect 10284 32943 10286 32952
rect 10232 32914 10284 32920
rect 10232 32768 10284 32774
rect 10232 32710 10284 32716
rect 10244 32366 10272 32710
rect 10336 32570 10364 32982
rect 10324 32564 10376 32570
rect 10324 32506 10376 32512
rect 10232 32360 10284 32366
rect 10230 32328 10232 32337
rect 10284 32328 10286 32337
rect 10230 32263 10286 32272
rect 10324 32292 10376 32298
rect 10324 32234 10376 32240
rect 10230 32192 10286 32201
rect 10230 32127 10286 32136
rect 10244 30841 10272 32127
rect 10230 30832 10286 30841
rect 10230 30767 10286 30776
rect 10140 29708 10192 29714
rect 10140 29650 10192 29656
rect 10232 29708 10284 29714
rect 10232 29650 10284 29656
rect 10244 29306 10272 29650
rect 10232 29300 10284 29306
rect 10232 29242 10284 29248
rect 10140 29096 10192 29102
rect 10140 29038 10192 29044
rect 10152 28626 10180 29038
rect 10140 28620 10192 28626
rect 10140 28562 10192 28568
rect 10152 27878 10180 28562
rect 10140 27872 10192 27878
rect 10140 27814 10192 27820
rect 10336 27690 10364 32234
rect 10428 28762 10456 37606
rect 10520 36922 10548 38383
rect 10508 36916 10560 36922
rect 10508 36858 10560 36864
rect 10506 36816 10562 36825
rect 10506 36751 10562 36760
rect 10520 36718 10548 36751
rect 10508 36712 10560 36718
rect 10508 36654 10560 36660
rect 10520 36378 10548 36654
rect 10508 36372 10560 36378
rect 10508 36314 10560 36320
rect 10612 35170 10640 38762
rect 10520 35142 10640 35170
rect 10520 33658 10548 35142
rect 10704 35034 10732 40990
rect 10876 40938 10928 40944
rect 10874 40624 10930 40633
rect 10784 40588 10836 40594
rect 10874 40559 10876 40568
rect 10784 40530 10836 40536
rect 10928 40559 10930 40568
rect 10876 40530 10928 40536
rect 10796 40066 10824 40530
rect 10956 40284 11252 40304
rect 11012 40282 11036 40284
rect 11092 40282 11116 40284
rect 11172 40282 11196 40284
rect 11034 40230 11036 40282
rect 11098 40230 11110 40282
rect 11172 40230 11174 40282
rect 11012 40228 11036 40230
rect 11092 40228 11116 40230
rect 11172 40228 11196 40230
rect 10956 40208 11252 40228
rect 10968 40112 11020 40118
rect 10796 40038 10916 40066
rect 10968 40054 11020 40060
rect 10888 39846 10916 40038
rect 10876 39840 10928 39846
rect 10874 39808 10876 39817
rect 10928 39808 10930 39817
rect 10874 39743 10930 39752
rect 10980 39658 11008 40054
rect 11244 39840 11296 39846
rect 11244 39782 11296 39788
rect 10796 39630 11008 39658
rect 10796 38554 10824 39630
rect 11256 39506 11284 39782
rect 10876 39500 10928 39506
rect 10876 39442 10928 39448
rect 11244 39500 11296 39506
rect 11244 39442 11296 39448
rect 10888 38554 10916 39442
rect 11256 39370 11284 39442
rect 11244 39364 11296 39370
rect 11244 39306 11296 39312
rect 10956 39196 11252 39216
rect 11012 39194 11036 39196
rect 11092 39194 11116 39196
rect 11172 39194 11196 39196
rect 11034 39142 11036 39194
rect 11098 39142 11110 39194
rect 11172 39142 11174 39194
rect 11012 39140 11036 39142
rect 11092 39140 11116 39142
rect 11172 39140 11196 39142
rect 10956 39120 11252 39140
rect 10968 38956 11020 38962
rect 10968 38898 11020 38904
rect 10784 38548 10836 38554
rect 10784 38490 10836 38496
rect 10876 38548 10928 38554
rect 10876 38490 10928 38496
rect 10980 38486 11008 38898
rect 11060 38888 11112 38894
rect 11060 38830 11112 38836
rect 11072 38729 11100 38830
rect 11058 38720 11114 38729
rect 11058 38655 11114 38664
rect 11242 38720 11298 38729
rect 11242 38655 11298 38664
rect 10968 38480 11020 38486
rect 10968 38422 11020 38428
rect 10784 38412 10836 38418
rect 10784 38354 10836 38360
rect 10876 38412 10928 38418
rect 10876 38354 10928 38360
rect 10796 37670 10824 38354
rect 10888 37670 10916 38354
rect 11256 38282 11284 38655
rect 11244 38276 11296 38282
rect 11244 38218 11296 38224
rect 10956 38108 11252 38128
rect 11012 38106 11036 38108
rect 11092 38106 11116 38108
rect 11172 38106 11196 38108
rect 11034 38054 11036 38106
rect 11098 38054 11110 38106
rect 11172 38054 11174 38106
rect 11012 38052 11036 38054
rect 11092 38052 11116 38054
rect 11172 38052 11196 38054
rect 10956 38032 11252 38052
rect 11242 37904 11298 37913
rect 11242 37839 11298 37848
rect 10968 37732 11020 37738
rect 10968 37674 11020 37680
rect 10784 37664 10836 37670
rect 10784 37606 10836 37612
rect 10876 37664 10928 37670
rect 10876 37606 10928 37612
rect 10784 37120 10836 37126
rect 10784 37062 10836 37068
rect 10612 35006 10732 35034
rect 10508 33652 10560 33658
rect 10508 33594 10560 33600
rect 10520 33289 10548 33594
rect 10506 33280 10562 33289
rect 10506 33215 10562 33224
rect 10612 31890 10640 35006
rect 10796 34932 10824 37062
rect 10888 36922 10916 37606
rect 10980 37194 11008 37674
rect 11256 37466 11284 37839
rect 11348 37482 11376 51326
rect 11440 50402 11468 51750
rect 11532 50810 11560 52906
rect 11716 52884 11744 53944
rect 11888 53576 11940 53582
rect 11888 53518 11940 53524
rect 11796 53168 11848 53174
rect 11794 53136 11796 53145
rect 11848 53136 11850 53145
rect 11794 53071 11850 53080
rect 11796 53032 11848 53038
rect 11796 52974 11848 52980
rect 11624 52856 11744 52884
rect 11624 52086 11652 52856
rect 11704 52624 11756 52630
rect 11704 52566 11756 52572
rect 11612 52080 11664 52086
rect 11612 52022 11664 52028
rect 11612 51808 11664 51814
rect 11612 51750 11664 51756
rect 11624 51649 11652 51750
rect 11610 51640 11666 51649
rect 11610 51575 11666 51584
rect 11612 51400 11664 51406
rect 11612 51342 11664 51348
rect 11624 50930 11652 51342
rect 11612 50924 11664 50930
rect 11612 50866 11664 50872
rect 11532 50782 11652 50810
rect 11624 50436 11652 50782
rect 11716 50561 11744 52566
rect 11808 52426 11836 52974
rect 11900 52737 11928 53518
rect 11886 52728 11942 52737
rect 11886 52663 11942 52672
rect 11888 52488 11940 52494
rect 11888 52430 11940 52436
rect 11796 52420 11848 52426
rect 11796 52362 11848 52368
rect 11808 51105 11836 52362
rect 11794 51096 11850 51105
rect 11794 51031 11850 51040
rect 11794 50960 11850 50969
rect 11794 50895 11850 50904
rect 11702 50552 11758 50561
rect 11702 50487 11758 50496
rect 11624 50408 11744 50436
rect 11440 50386 11560 50402
rect 11440 50380 11572 50386
rect 11440 50374 11520 50380
rect 11520 50322 11572 50328
rect 11532 49774 11560 50322
rect 11610 50280 11666 50289
rect 11610 50215 11666 50224
rect 11520 49768 11572 49774
rect 11520 49710 11572 49716
rect 11428 49224 11480 49230
rect 11428 49166 11480 49172
rect 11440 48890 11468 49166
rect 11428 48884 11480 48890
rect 11428 48826 11480 48832
rect 11426 48376 11482 48385
rect 11426 48311 11482 48320
rect 11440 46714 11468 48311
rect 11532 47530 11560 49710
rect 11624 49094 11652 50215
rect 11612 49088 11664 49094
rect 11612 49030 11664 49036
rect 11624 47705 11652 49030
rect 11610 47696 11666 47705
rect 11610 47631 11666 47640
rect 11520 47524 11572 47530
rect 11520 47466 11572 47472
rect 11716 47274 11744 50408
rect 11808 48278 11836 50895
rect 11900 50425 11928 52430
rect 11992 51241 12020 54266
rect 12084 53666 12112 55218
rect 12176 54126 12204 55354
rect 12164 54120 12216 54126
rect 12164 54062 12216 54068
rect 12268 53786 12296 56646
rect 12360 54233 12388 58398
rect 12544 58120 12572 59044
rect 12452 58092 12572 58120
rect 12452 57066 12480 58092
rect 12532 57996 12584 58002
rect 12532 57938 12584 57944
rect 12544 57390 12572 57938
rect 12532 57384 12584 57390
rect 12532 57326 12584 57332
rect 12452 57050 12572 57066
rect 12452 57044 12584 57050
rect 12452 57038 12532 57044
rect 12532 56986 12584 56992
rect 12440 56976 12492 56982
rect 12438 56944 12440 56953
rect 12492 56944 12494 56953
rect 12438 56879 12494 56888
rect 12544 56302 12572 56986
rect 12636 56914 12664 61610
rect 12728 60654 12756 61678
rect 12716 60648 12768 60654
rect 12716 60590 12768 60596
rect 12728 60314 12756 60590
rect 12716 60308 12768 60314
rect 12716 60250 12768 60256
rect 12728 60042 12756 60250
rect 12716 60036 12768 60042
rect 12716 59978 12768 59984
rect 12716 59560 12768 59566
rect 12716 59502 12768 59508
rect 12728 59158 12756 59502
rect 12716 59152 12768 59158
rect 12716 59094 12768 59100
rect 12820 58970 12848 65504
rect 12912 64938 12940 65894
rect 12900 64932 12952 64938
rect 12900 64874 12952 64880
rect 13004 64546 13032 66574
rect 13096 64682 13124 67526
rect 13188 67386 13216 67730
rect 13176 67380 13228 67386
rect 13176 67322 13228 67328
rect 13268 67108 13320 67114
rect 13268 67050 13320 67056
rect 13280 66094 13308 67050
rect 13372 66162 13400 68206
rect 13450 68167 13506 68176
rect 13360 66156 13412 66162
rect 13360 66098 13412 66104
rect 13268 66088 13320 66094
rect 13268 66030 13320 66036
rect 13280 65686 13308 66030
rect 13268 65680 13320 65686
rect 13268 65622 13320 65628
rect 13176 65612 13228 65618
rect 13176 65554 13228 65560
rect 13188 65210 13216 65554
rect 13176 65204 13228 65210
rect 13176 65146 13228 65152
rect 13096 64654 13216 64682
rect 12912 64518 13032 64546
rect 13084 64524 13136 64530
rect 12912 63209 12940 64518
rect 13084 64466 13136 64472
rect 12992 64456 13044 64462
rect 12992 64398 13044 64404
rect 13004 63238 13032 64398
rect 13096 63918 13124 64466
rect 13084 63912 13136 63918
rect 13082 63880 13084 63889
rect 13136 63880 13138 63889
rect 13082 63815 13138 63824
rect 13082 63744 13138 63753
rect 13082 63679 13138 63688
rect 12992 63232 13044 63238
rect 12898 63200 12954 63209
rect 12992 63174 13044 63180
rect 12898 63135 12954 63144
rect 12912 61169 12940 63135
rect 13096 62914 13124 63679
rect 13004 62886 13124 62914
rect 12898 61160 12954 61169
rect 12898 61095 12954 61104
rect 13004 61044 13032 62886
rect 13084 62824 13136 62830
rect 13084 62766 13136 62772
rect 12728 58942 12848 58970
rect 12912 61016 13032 61044
rect 12728 57322 12756 58942
rect 12808 58880 12860 58886
rect 12808 58822 12860 58828
rect 12820 58478 12848 58822
rect 12808 58472 12860 58478
rect 12808 58414 12860 58420
rect 12808 57996 12860 58002
rect 12808 57938 12860 57944
rect 12820 57594 12848 57938
rect 12808 57588 12860 57594
rect 12808 57530 12860 57536
rect 12716 57316 12768 57322
rect 12716 57258 12768 57264
rect 12624 56908 12676 56914
rect 12624 56850 12676 56856
rect 12728 56545 12756 57258
rect 12820 57254 12848 57530
rect 12808 57248 12860 57254
rect 12808 57190 12860 57196
rect 12808 56704 12860 56710
rect 12808 56646 12860 56652
rect 12714 56536 12770 56545
rect 12714 56471 12770 56480
rect 12820 56386 12848 56646
rect 12728 56358 12848 56386
rect 12532 56296 12584 56302
rect 12584 56244 12664 56250
rect 12532 56238 12664 56244
rect 12544 56222 12664 56238
rect 12532 56160 12584 56166
rect 12532 56102 12584 56108
rect 12544 56001 12572 56102
rect 12530 55992 12586 56001
rect 12530 55927 12586 55936
rect 12532 55888 12584 55894
rect 12532 55830 12584 55836
rect 12544 55162 12572 55830
rect 12452 55134 12572 55162
rect 12346 54224 12402 54233
rect 12346 54159 12402 54168
rect 12348 54120 12400 54126
rect 12348 54062 12400 54068
rect 12256 53780 12308 53786
rect 12256 53722 12308 53728
rect 12084 53638 12296 53666
rect 12072 53576 12124 53582
rect 12072 53518 12124 53524
rect 12084 52902 12112 53518
rect 12072 52896 12124 52902
rect 12072 52838 12124 52844
rect 12084 51388 12112 52838
rect 12164 52692 12216 52698
rect 12164 52634 12216 52640
rect 12176 51542 12204 52634
rect 12268 52494 12296 53638
rect 12256 52488 12308 52494
rect 12256 52430 12308 52436
rect 12256 52352 12308 52358
rect 12256 52294 12308 52300
rect 12268 52018 12296 52294
rect 12256 52012 12308 52018
rect 12256 51954 12308 51960
rect 12164 51536 12216 51542
rect 12164 51478 12216 51484
rect 12256 51468 12308 51474
rect 12256 51410 12308 51416
rect 12084 51360 12204 51388
rect 12072 51264 12124 51270
rect 11978 51232 12034 51241
rect 12072 51206 12124 51212
rect 11978 51167 12034 51176
rect 11980 51060 12032 51066
rect 11980 51002 12032 51008
rect 11886 50416 11942 50425
rect 11886 50351 11942 50360
rect 11888 50244 11940 50250
rect 11888 50186 11940 50192
rect 11900 49978 11928 50186
rect 11888 49972 11940 49978
rect 11888 49914 11940 49920
rect 11900 48793 11928 49914
rect 11992 49910 12020 51002
rect 11980 49904 12032 49910
rect 11980 49846 12032 49852
rect 12084 49774 12112 51206
rect 12072 49768 12124 49774
rect 12072 49710 12124 49716
rect 12084 49434 12112 49710
rect 12072 49428 12124 49434
rect 12072 49370 12124 49376
rect 11980 49292 12032 49298
rect 11980 49234 12032 49240
rect 11886 48784 11942 48793
rect 11886 48719 11942 48728
rect 11992 48618 12020 49234
rect 12084 48890 12112 49370
rect 12072 48884 12124 48890
rect 12072 48826 12124 48832
rect 11980 48612 12032 48618
rect 11980 48554 12032 48560
rect 11796 48272 11848 48278
rect 11796 48214 11848 48220
rect 11808 47598 11836 48214
rect 11796 47592 11848 47598
rect 11796 47534 11848 47540
rect 11888 47592 11940 47598
rect 11888 47534 11940 47540
rect 11716 47246 11836 47274
rect 11702 47152 11758 47161
rect 11702 47087 11758 47096
rect 11610 47016 11666 47025
rect 11520 46980 11572 46986
rect 11610 46951 11666 46960
rect 11520 46922 11572 46928
rect 11428 46708 11480 46714
rect 11428 46650 11480 46656
rect 11428 46504 11480 46510
rect 11428 46446 11480 46452
rect 11440 45830 11468 46446
rect 11428 45824 11480 45830
rect 11428 45766 11480 45772
rect 11440 45422 11468 45766
rect 11532 45529 11560 46922
rect 11624 46170 11652 46951
rect 11612 46164 11664 46170
rect 11612 46106 11664 46112
rect 11518 45520 11574 45529
rect 11518 45455 11574 45464
rect 11624 45422 11652 46106
rect 11428 45416 11480 45422
rect 11428 45358 11480 45364
rect 11612 45416 11664 45422
rect 11612 45358 11664 45364
rect 11428 45076 11480 45082
rect 11428 45018 11480 45024
rect 11440 42362 11468 45018
rect 11612 44940 11664 44946
rect 11612 44882 11664 44888
rect 11520 44804 11572 44810
rect 11520 44746 11572 44752
rect 11532 44470 11560 44746
rect 11624 44538 11652 44882
rect 11612 44532 11664 44538
rect 11612 44474 11664 44480
rect 11520 44464 11572 44470
rect 11520 44406 11572 44412
rect 11520 43852 11572 43858
rect 11520 43794 11572 43800
rect 11532 43450 11560 43794
rect 11520 43444 11572 43450
rect 11520 43386 11572 43392
rect 11532 42838 11560 43386
rect 11520 42832 11572 42838
rect 11520 42774 11572 42780
rect 11428 42356 11480 42362
rect 11428 42298 11480 42304
rect 11624 42265 11652 44474
rect 11610 42256 11666 42265
rect 11610 42191 11666 42200
rect 11612 42152 11664 42158
rect 11612 42094 11664 42100
rect 11520 41676 11572 41682
rect 11520 41618 11572 41624
rect 11532 41449 11560 41618
rect 11518 41440 11574 41449
rect 11518 41375 11574 41384
rect 11624 41256 11652 42094
rect 11532 41228 11652 41256
rect 11428 41132 11480 41138
rect 11428 41074 11480 41080
rect 11440 40050 11468 41074
rect 11428 40044 11480 40050
rect 11428 39986 11480 39992
rect 11532 39930 11560 41228
rect 11612 41132 11664 41138
rect 11612 41074 11664 41080
rect 11440 39902 11560 39930
rect 11440 37874 11468 39902
rect 11624 39522 11652 41074
rect 11716 40730 11744 47087
rect 11808 45529 11836 47246
rect 11794 45520 11850 45529
rect 11794 45455 11850 45464
rect 11900 45422 11928 47534
rect 11888 45416 11940 45422
rect 11808 45364 11888 45370
rect 11808 45358 11940 45364
rect 11808 45342 11928 45358
rect 11808 44742 11836 45342
rect 11796 44736 11848 44742
rect 11796 44678 11848 44684
rect 11704 40724 11756 40730
rect 11704 40666 11756 40672
rect 11704 39976 11756 39982
rect 11702 39944 11704 39953
rect 11756 39944 11758 39953
rect 11702 39879 11758 39888
rect 11716 39681 11744 39879
rect 11702 39672 11758 39681
rect 11702 39607 11758 39616
rect 11624 39494 11744 39522
rect 11612 39432 11664 39438
rect 11518 39400 11574 39409
rect 11612 39374 11664 39380
rect 11518 39335 11574 39344
rect 11428 37868 11480 37874
rect 11428 37810 11480 37816
rect 11244 37460 11296 37466
rect 11348 37454 11468 37482
rect 11244 37402 11296 37408
rect 11336 37324 11388 37330
rect 11336 37266 11388 37272
rect 10968 37188 11020 37194
rect 10968 37130 11020 37136
rect 10956 37020 11252 37040
rect 11012 37018 11036 37020
rect 11092 37018 11116 37020
rect 11172 37018 11196 37020
rect 11034 36966 11036 37018
rect 11098 36966 11110 37018
rect 11172 36966 11174 37018
rect 11012 36964 11036 36966
rect 11092 36964 11116 36966
rect 11172 36964 11196 36966
rect 10956 36944 11252 36964
rect 10876 36916 10928 36922
rect 10876 36858 10928 36864
rect 11348 36582 11376 37266
rect 11336 36576 11388 36582
rect 11336 36518 11388 36524
rect 10876 36372 10928 36378
rect 10876 36314 10928 36320
rect 10704 34904 10824 34932
rect 10704 31929 10732 34904
rect 10782 34504 10838 34513
rect 10782 34439 10838 34448
rect 10690 31920 10746 31929
rect 10600 31884 10652 31890
rect 10690 31855 10746 31864
rect 10600 31826 10652 31832
rect 10612 30938 10640 31826
rect 10692 31748 10744 31754
rect 10692 31690 10744 31696
rect 10600 30932 10652 30938
rect 10600 30874 10652 30880
rect 10704 30870 10732 31690
rect 10796 31498 10824 34439
rect 10888 31686 10916 36314
rect 11348 36242 11376 36518
rect 11336 36236 11388 36242
rect 11336 36178 11388 36184
rect 10956 35932 11252 35952
rect 11012 35930 11036 35932
rect 11092 35930 11116 35932
rect 11172 35930 11196 35932
rect 11034 35878 11036 35930
rect 11098 35878 11110 35930
rect 11172 35878 11174 35930
rect 11012 35876 11036 35878
rect 11092 35876 11116 35878
rect 11172 35876 11196 35878
rect 10956 35856 11252 35876
rect 11348 35834 11376 36178
rect 11336 35828 11388 35834
rect 11336 35770 11388 35776
rect 11440 35630 11468 37454
rect 11532 36650 11560 39335
rect 11520 36644 11572 36650
rect 11520 36586 11572 36592
rect 11428 35624 11480 35630
rect 11428 35566 11480 35572
rect 10956 34844 11252 34864
rect 11012 34842 11036 34844
rect 11092 34842 11116 34844
rect 11172 34842 11196 34844
rect 11034 34790 11036 34842
rect 11098 34790 11110 34842
rect 11172 34790 11174 34842
rect 11012 34788 11036 34790
rect 11092 34788 11116 34790
rect 11172 34788 11196 34790
rect 10956 34768 11252 34788
rect 11426 34096 11482 34105
rect 11426 34031 11482 34040
rect 10956 33756 11252 33776
rect 11012 33754 11036 33756
rect 11092 33754 11116 33756
rect 11172 33754 11196 33756
rect 11034 33702 11036 33754
rect 11098 33702 11110 33754
rect 11172 33702 11174 33754
rect 11012 33700 11036 33702
rect 11092 33700 11116 33702
rect 11172 33700 11196 33702
rect 10956 33680 11252 33700
rect 11336 32768 11388 32774
rect 11336 32710 11388 32716
rect 10956 32668 11252 32688
rect 11012 32666 11036 32668
rect 11092 32666 11116 32668
rect 11172 32666 11196 32668
rect 11034 32614 11036 32666
rect 11098 32614 11110 32666
rect 11172 32614 11174 32666
rect 11012 32612 11036 32614
rect 11092 32612 11116 32614
rect 11172 32612 11196 32614
rect 10956 32592 11252 32612
rect 11060 32428 11112 32434
rect 11060 32370 11112 32376
rect 11072 31890 11100 32370
rect 11348 32230 11376 32710
rect 11336 32224 11388 32230
rect 11336 32166 11388 32172
rect 11060 31884 11112 31890
rect 11060 31826 11112 31832
rect 11348 31793 11376 32166
rect 11334 31784 11390 31793
rect 11334 31719 11390 31728
rect 10876 31680 10928 31686
rect 10876 31622 10928 31628
rect 11336 31680 11388 31686
rect 11336 31622 11388 31628
rect 10956 31580 11252 31600
rect 11012 31578 11036 31580
rect 11092 31578 11116 31580
rect 11172 31578 11196 31580
rect 11034 31526 11036 31578
rect 11098 31526 11110 31578
rect 11172 31526 11174 31578
rect 11012 31524 11036 31526
rect 11092 31524 11116 31526
rect 11172 31524 11196 31526
rect 10956 31504 11252 31524
rect 10796 31470 10916 31498
rect 10782 31376 10838 31385
rect 10782 31311 10784 31320
rect 10836 31311 10838 31320
rect 10784 31282 10836 31288
rect 10888 31192 10916 31470
rect 11348 31278 11376 31622
rect 11336 31272 11388 31278
rect 11336 31214 11388 31220
rect 10796 31164 10916 31192
rect 10692 30864 10744 30870
rect 10598 30832 10654 30841
rect 10692 30806 10744 30812
rect 10598 30767 10654 30776
rect 10506 30288 10562 30297
rect 10506 30223 10562 30232
rect 10520 30190 10548 30223
rect 10508 30184 10560 30190
rect 10508 30126 10560 30132
rect 10416 28756 10468 28762
rect 10416 28698 10468 28704
rect 10336 27662 10456 27690
rect 10324 27532 10376 27538
rect 10324 27474 10376 27480
rect 10336 27130 10364 27474
rect 10324 27124 10376 27130
rect 10324 27066 10376 27072
rect 10140 26240 10192 26246
rect 10140 26182 10192 26188
rect 10152 25838 10180 26182
rect 10428 25838 10456 27662
rect 10508 27328 10560 27334
rect 10508 27270 10560 27276
rect 10520 27033 10548 27270
rect 10506 27024 10562 27033
rect 10506 26959 10562 26968
rect 10140 25832 10192 25838
rect 10140 25774 10192 25780
rect 10416 25832 10468 25838
rect 10416 25774 10468 25780
rect 10048 25424 10100 25430
rect 10048 25366 10100 25372
rect 10060 24410 10088 25366
rect 10048 24404 10100 24410
rect 10048 24346 10100 24352
rect 10046 24304 10102 24313
rect 10046 24239 10048 24248
rect 10100 24239 10102 24248
rect 10048 24210 10100 24216
rect 10060 23730 10088 24210
rect 10048 23724 10100 23730
rect 10048 23666 10100 23672
rect 10152 23594 10180 25774
rect 10428 25498 10456 25774
rect 10416 25492 10468 25498
rect 10416 25434 10468 25440
rect 10416 25220 10468 25226
rect 10416 25162 10468 25168
rect 10232 24744 10284 24750
rect 10232 24686 10284 24692
rect 10244 24342 10272 24686
rect 10232 24336 10284 24342
rect 10232 24278 10284 24284
rect 10140 23588 10192 23594
rect 10140 23530 10192 23536
rect 9956 23180 10008 23186
rect 9956 23122 10008 23128
rect 9968 22710 9996 23122
rect 10244 22953 10272 24278
rect 10428 23186 10456 25162
rect 10612 23304 10640 30767
rect 10690 30560 10746 30569
rect 10690 30495 10746 30504
rect 10704 29510 10732 30495
rect 10692 29504 10744 29510
rect 10692 29446 10744 29452
rect 10704 26246 10732 29446
rect 10692 26240 10744 26246
rect 10692 26182 10744 26188
rect 10796 24750 10824 31164
rect 11060 31136 11112 31142
rect 10888 31084 11060 31090
rect 10888 31078 11112 31084
rect 10888 31062 11100 31078
rect 10888 29306 10916 31062
rect 11348 30870 11376 31214
rect 11336 30864 11388 30870
rect 11334 30832 11336 30841
rect 11388 30832 11390 30841
rect 11334 30767 11390 30776
rect 11348 30741 11376 30767
rect 11336 30660 11388 30666
rect 11336 30602 11388 30608
rect 10956 30492 11252 30512
rect 11012 30490 11036 30492
rect 11092 30490 11116 30492
rect 11172 30490 11196 30492
rect 11034 30438 11036 30490
rect 11098 30438 11110 30490
rect 11172 30438 11174 30490
rect 11012 30436 11036 30438
rect 11092 30436 11116 30438
rect 11172 30436 11196 30438
rect 10956 30416 11252 30436
rect 10966 29744 11022 29753
rect 10966 29679 10968 29688
rect 11020 29679 11022 29688
rect 10968 29650 11020 29656
rect 10956 29404 11252 29424
rect 11012 29402 11036 29404
rect 11092 29402 11116 29404
rect 11172 29402 11196 29404
rect 11034 29350 11036 29402
rect 11098 29350 11110 29402
rect 11172 29350 11174 29402
rect 11012 29348 11036 29350
rect 11092 29348 11116 29350
rect 11172 29348 11196 29350
rect 10956 29328 11252 29348
rect 10876 29300 10928 29306
rect 10876 29242 10928 29248
rect 10956 28316 11252 28336
rect 11012 28314 11036 28316
rect 11092 28314 11116 28316
rect 11172 28314 11196 28316
rect 11034 28262 11036 28314
rect 11098 28262 11110 28314
rect 11172 28262 11174 28314
rect 11012 28260 11036 28262
rect 11092 28260 11116 28262
rect 11172 28260 11196 28262
rect 10956 28240 11252 28260
rect 11348 27674 11376 30602
rect 11336 27668 11388 27674
rect 11336 27610 11388 27616
rect 11336 27532 11388 27538
rect 11336 27474 11388 27480
rect 10956 27228 11252 27248
rect 11012 27226 11036 27228
rect 11092 27226 11116 27228
rect 11172 27226 11196 27228
rect 11034 27174 11036 27226
rect 11098 27174 11110 27226
rect 11172 27174 11174 27226
rect 11012 27172 11036 27174
rect 11092 27172 11116 27174
rect 11172 27172 11196 27174
rect 10956 27152 11252 27172
rect 11348 27112 11376 27474
rect 11164 27084 11376 27112
rect 11164 26926 11192 27084
rect 11152 26920 11204 26926
rect 11152 26862 11204 26868
rect 10876 26784 10928 26790
rect 10876 26726 10928 26732
rect 10888 25770 10916 26726
rect 11164 26353 11192 26862
rect 11440 26568 11468 34031
rect 11518 33144 11574 33153
rect 11518 33079 11574 33088
rect 11532 31890 11560 33079
rect 11520 31884 11572 31890
rect 11520 31826 11572 31832
rect 11532 31249 11560 31826
rect 11518 31240 11574 31249
rect 11518 31175 11574 31184
rect 11624 30666 11652 39374
rect 11716 32366 11744 39494
rect 11808 36310 11836 44678
rect 11888 43988 11940 43994
rect 11888 43930 11940 43936
rect 11900 41274 11928 43930
rect 11992 42158 12020 48554
rect 12070 48104 12126 48113
rect 12070 48039 12126 48048
rect 12084 45082 12112 48039
rect 12072 45076 12124 45082
rect 12072 45018 12124 45024
rect 12084 44713 12112 45018
rect 12176 44946 12204 51360
rect 12268 50250 12296 51410
rect 12256 50244 12308 50250
rect 12256 50186 12308 50192
rect 12254 50144 12310 50153
rect 12254 50079 12310 50088
rect 12268 49298 12296 50079
rect 12256 49292 12308 49298
rect 12256 49234 12308 49240
rect 12256 48680 12308 48686
rect 12256 48622 12308 48628
rect 12268 47598 12296 48622
rect 12256 47592 12308 47598
rect 12256 47534 12308 47540
rect 12268 46986 12296 47534
rect 12360 47433 12388 54062
rect 12452 53990 12480 55134
rect 12636 54618 12664 56222
rect 12728 55894 12756 56358
rect 12716 55888 12768 55894
rect 12716 55830 12768 55836
rect 12808 55820 12860 55826
rect 12808 55762 12860 55768
rect 12820 55078 12848 55762
rect 12808 55072 12860 55078
rect 12808 55014 12860 55020
rect 12716 54868 12768 54874
rect 12716 54810 12768 54816
rect 12544 54590 12664 54618
rect 12544 54330 12572 54590
rect 12624 54528 12676 54534
rect 12624 54470 12676 54476
rect 12532 54324 12584 54330
rect 12532 54266 12584 54272
rect 12532 54188 12584 54194
rect 12532 54130 12584 54136
rect 12440 53984 12492 53990
rect 12440 53926 12492 53932
rect 12544 53938 12572 54130
rect 12636 54126 12664 54470
rect 12624 54120 12676 54126
rect 12622 54088 12624 54097
rect 12676 54088 12678 54097
rect 12622 54023 12678 54032
rect 12452 53514 12480 53926
rect 12544 53910 12664 53938
rect 12532 53780 12584 53786
rect 12532 53722 12584 53728
rect 12440 53508 12492 53514
rect 12440 53450 12492 53456
rect 12544 52902 12572 53722
rect 12532 52896 12584 52902
rect 12532 52838 12584 52844
rect 12440 51536 12492 51542
rect 12440 51478 12492 51484
rect 12452 51066 12480 51478
rect 12544 51474 12572 52838
rect 12532 51468 12584 51474
rect 12532 51410 12584 51416
rect 12636 51354 12664 53910
rect 12544 51326 12664 51354
rect 12440 51060 12492 51066
rect 12440 51002 12492 51008
rect 12440 50312 12492 50318
rect 12440 50254 12492 50260
rect 12452 49978 12480 50254
rect 12440 49972 12492 49978
rect 12440 49914 12492 49920
rect 12440 49836 12492 49842
rect 12440 49778 12492 49784
rect 12452 48890 12480 49778
rect 12544 49230 12572 51326
rect 12624 51264 12676 51270
rect 12624 51206 12676 51212
rect 12636 49314 12664 51206
rect 12728 49722 12756 54810
rect 12820 53650 12848 55014
rect 12912 54874 12940 61016
rect 12992 60104 13044 60110
rect 12992 60046 13044 60052
rect 13004 59566 13032 60046
rect 12992 59560 13044 59566
rect 12992 59502 13044 59508
rect 13096 58290 13124 62766
rect 13188 61266 13216 64654
rect 13464 64433 13492 68167
rect 13924 68134 13952 68818
rect 14108 68134 14136 68886
rect 15016 68808 15068 68814
rect 15016 68750 15068 68756
rect 15936 68808 15988 68814
rect 15936 68750 15988 68756
rect 13912 68128 13964 68134
rect 13910 68096 13912 68105
rect 14096 68128 14148 68134
rect 13964 68096 13966 68105
rect 14096 68070 14148 68076
rect 13910 68031 13966 68040
rect 14289 68028 14585 68048
rect 14345 68026 14369 68028
rect 14425 68026 14449 68028
rect 14505 68026 14529 68028
rect 14367 67974 14369 68026
rect 14431 67974 14443 68026
rect 14505 67974 14507 68026
rect 14345 67972 14369 67974
rect 14425 67972 14449 67974
rect 14505 67972 14529 67974
rect 14289 67952 14585 67972
rect 14094 67824 14150 67833
rect 14094 67759 14150 67768
rect 13728 67720 13780 67726
rect 13728 67662 13780 67668
rect 13740 67028 13768 67662
rect 13820 67040 13872 67046
rect 13740 67000 13820 67028
rect 13636 65544 13688 65550
rect 13636 65486 13688 65492
rect 13648 64938 13676 65486
rect 13636 64932 13688 64938
rect 13636 64874 13688 64880
rect 13740 64818 13768 67000
rect 13820 66982 13872 66988
rect 14004 66292 14056 66298
rect 14004 66234 14056 66240
rect 13910 65920 13966 65929
rect 13910 65855 13966 65864
rect 13924 65754 13952 65855
rect 13912 65748 13964 65754
rect 13912 65690 13964 65696
rect 14016 65618 14044 66234
rect 14004 65612 14056 65618
rect 14004 65554 14056 65560
rect 14004 65000 14056 65006
rect 14004 64942 14056 64948
rect 13648 64790 13768 64818
rect 13450 64424 13506 64433
rect 13450 64359 13506 64368
rect 13268 63776 13320 63782
rect 13464 63753 13492 64359
rect 13268 63718 13320 63724
rect 13450 63744 13506 63753
rect 13280 61878 13308 63718
rect 13450 63679 13506 63688
rect 13360 63232 13412 63238
rect 13360 63174 13412 63180
rect 13372 62694 13400 63174
rect 13360 62688 13412 62694
rect 13360 62630 13412 62636
rect 13372 62354 13400 62630
rect 13360 62348 13412 62354
rect 13360 62290 13412 62296
rect 13268 61872 13320 61878
rect 13268 61814 13320 61820
rect 13280 61742 13308 61814
rect 13648 61810 13676 64790
rect 14016 63918 14044 64942
rect 14004 63912 14056 63918
rect 14004 63854 14056 63860
rect 13728 63368 13780 63374
rect 13728 63310 13780 63316
rect 13740 62150 13768 63310
rect 13820 62688 13872 62694
rect 13820 62630 13872 62636
rect 13728 62144 13780 62150
rect 13728 62086 13780 62092
rect 13832 61826 13860 62630
rect 14004 62280 14056 62286
rect 14004 62222 14056 62228
rect 13636 61804 13688 61810
rect 13636 61746 13688 61752
rect 13740 61798 13860 61826
rect 13268 61736 13320 61742
rect 13268 61678 13320 61684
rect 13280 61282 13308 61678
rect 13740 61674 13768 61798
rect 13728 61668 13780 61674
rect 13728 61610 13780 61616
rect 14016 61606 14044 62222
rect 14004 61600 14056 61606
rect 14004 61542 14056 61548
rect 13452 61328 13504 61334
rect 13176 61260 13228 61266
rect 13280 61254 13400 61282
rect 13452 61270 13504 61276
rect 13176 61202 13228 61208
rect 13188 60858 13216 61202
rect 13266 60888 13322 60897
rect 13176 60852 13228 60858
rect 13266 60823 13322 60832
rect 13176 60794 13228 60800
rect 13176 60172 13228 60178
rect 13176 60114 13228 60120
rect 13188 59770 13216 60114
rect 13176 59764 13228 59770
rect 13176 59706 13228 59712
rect 13004 58262 13124 58290
rect 13004 57361 13032 58262
rect 13188 58120 13216 59706
rect 13280 59430 13308 60823
rect 13268 59424 13320 59430
rect 13268 59366 13320 59372
rect 13268 59152 13320 59158
rect 13268 59094 13320 59100
rect 13096 58092 13216 58120
rect 12990 57352 13046 57361
rect 12990 57287 13046 57296
rect 12992 56908 13044 56914
rect 12992 56850 13044 56856
rect 13004 56166 13032 56850
rect 12992 56160 13044 56166
rect 12992 56102 13044 56108
rect 12900 54868 12952 54874
rect 12900 54810 12952 54816
rect 12900 54596 12952 54602
rect 12900 54538 12952 54544
rect 12912 54126 12940 54538
rect 12900 54120 12952 54126
rect 12900 54062 12952 54068
rect 12808 53644 12860 53650
rect 12808 53586 12860 53592
rect 12912 53582 12940 54062
rect 12900 53576 12952 53582
rect 12900 53518 12952 53524
rect 12808 53508 12860 53514
rect 12808 53450 12860 53456
rect 12820 51066 12848 53450
rect 12900 53440 12952 53446
rect 12900 53382 12952 53388
rect 12912 53009 12940 53382
rect 12898 53000 12954 53009
rect 12898 52935 12954 52944
rect 12912 52737 12940 52935
rect 12898 52728 12954 52737
rect 12898 52663 12954 52672
rect 12900 52488 12952 52494
rect 12900 52430 12952 52436
rect 12912 52018 12940 52430
rect 12900 52012 12952 52018
rect 12900 51954 12952 51960
rect 12900 51536 12952 51542
rect 12898 51504 12900 51513
rect 12952 51504 12954 51513
rect 12898 51439 12954 51448
rect 12900 51400 12952 51406
rect 12900 51342 12952 51348
rect 12808 51060 12860 51066
rect 12808 51002 12860 51008
rect 12912 50912 12940 51342
rect 13004 50969 13032 56102
rect 13096 55894 13124 58092
rect 13176 57996 13228 58002
rect 13176 57938 13228 57944
rect 13188 57322 13216 57938
rect 13176 57316 13228 57322
rect 13176 57258 13228 57264
rect 13084 55888 13136 55894
rect 13084 55830 13136 55836
rect 13084 55752 13136 55758
rect 13084 55694 13136 55700
rect 13096 54738 13124 55694
rect 13280 55298 13308 59094
rect 13188 55270 13308 55298
rect 13084 54732 13136 54738
rect 13084 54674 13136 54680
rect 13084 53644 13136 53650
rect 13084 53586 13136 53592
rect 13096 52902 13124 53586
rect 13188 53106 13216 55270
rect 13268 55140 13320 55146
rect 13268 55082 13320 55088
rect 13280 54602 13308 55082
rect 13268 54596 13320 54602
rect 13268 54538 13320 54544
rect 13176 53100 13228 53106
rect 13176 53042 13228 53048
rect 13176 52964 13228 52970
rect 13176 52906 13228 52912
rect 13084 52896 13136 52902
rect 13084 52838 13136 52844
rect 12820 50884 12940 50912
rect 12990 50960 13046 50969
rect 12990 50895 13046 50904
rect 12820 50726 12848 50884
rect 12808 50720 12860 50726
rect 12808 50662 12860 50668
rect 12900 50720 12952 50726
rect 12900 50662 12952 50668
rect 12820 50318 12848 50662
rect 12808 50312 12860 50318
rect 12808 50254 12860 50260
rect 12820 49842 12848 50254
rect 12912 49842 12940 50662
rect 12808 49836 12860 49842
rect 12808 49778 12860 49784
rect 12900 49836 12952 49842
rect 12900 49778 12952 49784
rect 12728 49694 13032 49722
rect 12898 49600 12954 49609
rect 12898 49535 12954 49544
rect 12636 49298 12756 49314
rect 12636 49292 12768 49298
rect 12636 49286 12716 49292
rect 12716 49234 12768 49240
rect 12532 49224 12584 49230
rect 12532 49166 12584 49172
rect 12440 48884 12492 48890
rect 12440 48826 12492 48832
rect 12622 48784 12678 48793
rect 12440 48748 12492 48754
rect 12622 48719 12678 48728
rect 12440 48690 12492 48696
rect 12346 47424 12402 47433
rect 12346 47359 12402 47368
rect 12346 47288 12402 47297
rect 12346 47223 12402 47232
rect 12256 46980 12308 46986
rect 12256 46922 12308 46928
rect 12256 46368 12308 46374
rect 12256 46310 12308 46316
rect 12268 46170 12296 46310
rect 12256 46164 12308 46170
rect 12256 46106 12308 46112
rect 12360 45898 12388 47223
rect 12452 46322 12480 48690
rect 12636 48521 12664 48719
rect 12622 48512 12678 48521
rect 12622 48447 12678 48456
rect 12636 48278 12664 48447
rect 12728 48346 12756 49234
rect 12808 49224 12860 49230
rect 12808 49166 12860 49172
rect 12716 48340 12768 48346
rect 12716 48282 12768 48288
rect 12624 48272 12676 48278
rect 12624 48214 12676 48220
rect 12728 47841 12756 48282
rect 12714 47832 12770 47841
rect 12714 47767 12770 47776
rect 12820 47682 12848 49166
rect 12912 49094 12940 49535
rect 12900 49088 12952 49094
rect 12900 49030 12952 49036
rect 12900 48884 12952 48890
rect 12900 48826 12952 48832
rect 12912 48142 12940 48826
rect 12900 48136 12952 48142
rect 12900 48078 12952 48084
rect 12636 47654 12848 47682
rect 12452 46294 12572 46322
rect 12348 45892 12400 45898
rect 12348 45834 12400 45840
rect 12256 45620 12308 45626
rect 12256 45562 12308 45568
rect 12164 44940 12216 44946
rect 12164 44882 12216 44888
rect 12070 44704 12126 44713
rect 12126 44662 12204 44690
rect 12070 44639 12126 44648
rect 12070 44432 12126 44441
rect 12070 44367 12126 44376
rect 12084 43110 12112 44367
rect 12072 43104 12124 43110
rect 12072 43046 12124 43052
rect 11980 42152 12032 42158
rect 11980 42094 12032 42100
rect 11980 41676 12032 41682
rect 11980 41618 12032 41624
rect 11888 41268 11940 41274
rect 11888 41210 11940 41216
rect 11992 41138 12020 41618
rect 11980 41132 12032 41138
rect 11900 41092 11980 41120
rect 11900 39982 11928 41092
rect 11980 41074 12032 41080
rect 11980 40996 12032 41002
rect 11980 40938 12032 40944
rect 11992 40186 12020 40938
rect 11980 40180 12032 40186
rect 11980 40122 12032 40128
rect 11888 39976 11940 39982
rect 11888 39918 11940 39924
rect 11900 39642 11928 39918
rect 11888 39636 11940 39642
rect 11888 39578 11940 39584
rect 11980 39500 12032 39506
rect 11980 39442 12032 39448
rect 11992 38894 12020 39442
rect 11980 38888 12032 38894
rect 11978 38856 11980 38865
rect 12032 38856 12034 38865
rect 11978 38791 12034 38800
rect 11978 38176 12034 38185
rect 11978 38111 12034 38120
rect 11888 37868 11940 37874
rect 11888 37810 11940 37816
rect 11900 37670 11928 37810
rect 11992 37806 12020 38111
rect 12084 37806 12112 43046
rect 12176 42226 12204 44662
rect 12164 42220 12216 42226
rect 12164 42162 12216 42168
rect 12164 41608 12216 41614
rect 12164 41550 12216 41556
rect 12176 41070 12204 41550
rect 12268 41274 12296 45562
rect 12360 44334 12388 45834
rect 12440 45824 12492 45830
rect 12440 45766 12492 45772
rect 12452 45268 12480 45766
rect 12544 45626 12572 46294
rect 12532 45620 12584 45626
rect 12532 45562 12584 45568
rect 12532 45280 12584 45286
rect 12452 45240 12532 45268
rect 12532 45222 12584 45228
rect 12544 44878 12572 45222
rect 12440 44872 12492 44878
rect 12440 44814 12492 44820
rect 12532 44872 12584 44878
rect 12532 44814 12584 44820
rect 12452 44470 12480 44814
rect 12440 44464 12492 44470
rect 12440 44406 12492 44412
rect 12348 44328 12400 44334
rect 12348 44270 12400 44276
rect 12256 41268 12308 41274
rect 12256 41210 12308 41216
rect 12254 41168 12310 41177
rect 12254 41103 12310 41112
rect 12164 41064 12216 41070
rect 12164 41006 12216 41012
rect 12164 40588 12216 40594
rect 12164 40530 12216 40536
rect 12176 40186 12204 40530
rect 12164 40180 12216 40186
rect 12164 40122 12216 40128
rect 12164 39840 12216 39846
rect 12164 39782 12216 39788
rect 12176 38894 12204 39782
rect 12164 38888 12216 38894
rect 12164 38830 12216 38836
rect 11980 37800 12032 37806
rect 11980 37742 12032 37748
rect 12072 37800 12124 37806
rect 12072 37742 12124 37748
rect 11888 37664 11940 37670
rect 11888 37606 11940 37612
rect 11796 36304 11848 36310
rect 11796 36246 11848 36252
rect 11796 35624 11848 35630
rect 11796 35566 11848 35572
rect 11704 32360 11756 32366
rect 11704 32302 11756 32308
rect 11808 32212 11836 35566
rect 11900 32434 11928 37606
rect 11992 37398 12020 37742
rect 11980 37392 12032 37398
rect 11980 37334 12032 37340
rect 12084 37330 12112 37742
rect 12072 37324 12124 37330
rect 12072 37266 12124 37272
rect 11980 36644 12032 36650
rect 11980 36586 12032 36592
rect 11992 35630 12020 36586
rect 11980 35624 12032 35630
rect 11980 35566 12032 35572
rect 11888 32428 11940 32434
rect 11888 32370 11940 32376
rect 11716 32184 11836 32212
rect 11612 30660 11664 30666
rect 11612 30602 11664 30608
rect 11716 28948 11744 32184
rect 11978 31920 12034 31929
rect 11978 31855 12034 31864
rect 11886 31784 11942 31793
rect 11886 31719 11942 31728
rect 11900 30297 11928 31719
rect 11886 30288 11942 30297
rect 11886 30223 11942 30232
rect 11796 29028 11848 29034
rect 11796 28970 11848 28976
rect 11518 28928 11574 28937
rect 11624 28920 11744 28948
rect 11624 28914 11652 28920
rect 11574 28886 11652 28914
rect 11518 28863 11574 28872
rect 11518 27976 11574 27985
rect 11518 27911 11574 27920
rect 11532 26586 11560 27911
rect 11808 27062 11836 28970
rect 11992 28121 12020 31855
rect 12084 31142 12112 37266
rect 12176 37262 12204 38830
rect 12164 37256 12216 37262
rect 12164 37198 12216 37204
rect 12176 36378 12204 37198
rect 12268 36650 12296 41103
rect 12360 40497 12388 44270
rect 12452 43994 12480 44406
rect 12532 44328 12584 44334
rect 12532 44270 12584 44276
rect 12440 43988 12492 43994
rect 12440 43930 12492 43936
rect 12544 43790 12572 44270
rect 12532 43784 12584 43790
rect 12532 43726 12584 43732
rect 12544 43353 12572 43726
rect 12636 43450 12664 47654
rect 12806 47560 12862 47569
rect 12716 47524 12768 47530
rect 12806 47495 12862 47504
rect 12716 47466 12768 47472
rect 12728 46186 12756 47466
rect 12820 47258 12848 47495
rect 12912 47462 12940 48078
rect 12900 47456 12952 47462
rect 12900 47398 12952 47404
rect 12808 47252 12860 47258
rect 12808 47194 12860 47200
rect 12820 46510 12848 47194
rect 12912 47054 12940 47398
rect 12900 47048 12952 47054
rect 12900 46990 12952 46996
rect 12912 46578 12940 46990
rect 12900 46572 12952 46578
rect 12900 46514 12952 46520
rect 12808 46504 12860 46510
rect 12808 46446 12860 46452
rect 12728 46170 12848 46186
rect 12716 46164 12848 46170
rect 12768 46158 12848 46164
rect 12716 46106 12768 46112
rect 12716 46028 12768 46034
rect 12716 45970 12768 45976
rect 12728 45082 12756 45970
rect 12820 45558 12848 46158
rect 13004 46050 13032 49694
rect 13096 46170 13124 52838
rect 13188 51950 13216 52906
rect 13280 52630 13308 54538
rect 13268 52624 13320 52630
rect 13268 52566 13320 52572
rect 13268 52420 13320 52426
rect 13268 52362 13320 52368
rect 13176 51944 13228 51950
rect 13176 51886 13228 51892
rect 13176 51400 13228 51406
rect 13176 51342 13228 51348
rect 13188 51066 13216 51342
rect 13280 51270 13308 52362
rect 13268 51264 13320 51270
rect 13268 51206 13320 51212
rect 13372 51105 13400 61254
rect 13464 60518 13492 61270
rect 13820 61260 13872 61266
rect 13820 61202 13872 61208
rect 13636 61192 13688 61198
rect 13636 61134 13688 61140
rect 13452 60512 13504 60518
rect 13452 60454 13504 60460
rect 13464 59770 13492 60454
rect 13452 59764 13504 59770
rect 13452 59706 13504 59712
rect 13544 59696 13596 59702
rect 13544 59638 13596 59644
rect 13556 59566 13584 59638
rect 13544 59560 13596 59566
rect 13544 59502 13596 59508
rect 13452 59424 13504 59430
rect 13452 59366 13504 59372
rect 13464 57338 13492 59366
rect 13556 57934 13584 59502
rect 13648 58562 13676 61134
rect 13832 59226 13860 61202
rect 14108 60761 14136 67759
rect 14372 67312 14424 67318
rect 14370 67280 14372 67289
rect 14424 67280 14426 67289
rect 14370 67215 14426 67224
rect 14289 66940 14585 66960
rect 14345 66938 14369 66940
rect 14425 66938 14449 66940
rect 14505 66938 14529 66940
rect 14367 66886 14369 66938
rect 14431 66886 14443 66938
rect 14505 66886 14507 66938
rect 14345 66884 14369 66886
rect 14425 66884 14449 66886
rect 14505 66884 14529 66886
rect 14289 66864 14585 66884
rect 14372 66700 14424 66706
rect 14372 66642 14424 66648
rect 14384 66298 14412 66642
rect 14372 66292 14424 66298
rect 14372 66234 14424 66240
rect 14740 65952 14792 65958
rect 14738 65920 14740 65929
rect 14792 65920 14794 65929
rect 14289 65852 14585 65872
rect 14738 65855 14794 65864
rect 14345 65850 14369 65852
rect 14425 65850 14449 65852
rect 14505 65850 14529 65852
rect 14367 65798 14369 65850
rect 14431 65798 14443 65850
rect 14505 65798 14507 65850
rect 14345 65796 14369 65798
rect 14425 65796 14449 65798
rect 14505 65796 14529 65798
rect 14289 65776 14585 65796
rect 14289 64764 14585 64784
rect 14345 64762 14369 64764
rect 14425 64762 14449 64764
rect 14505 64762 14529 64764
rect 14367 64710 14369 64762
rect 14431 64710 14443 64762
rect 14505 64710 14507 64762
rect 14345 64708 14369 64710
rect 14425 64708 14449 64710
rect 14505 64708 14529 64710
rect 14289 64688 14585 64708
rect 14370 64560 14426 64569
rect 14370 64495 14426 64504
rect 14384 64462 14412 64495
rect 14372 64456 14424 64462
rect 14372 64398 14424 64404
rect 14289 63676 14585 63696
rect 14345 63674 14369 63676
rect 14425 63674 14449 63676
rect 14505 63674 14529 63676
rect 14367 63622 14369 63674
rect 14431 63622 14443 63674
rect 14505 63622 14507 63674
rect 14345 63620 14369 63622
rect 14425 63620 14449 63622
rect 14505 63620 14529 63622
rect 14289 63600 14585 63620
rect 14740 63436 14792 63442
rect 14740 63378 14792 63384
rect 14752 63034 14780 63378
rect 14832 63232 14884 63238
rect 14832 63174 14884 63180
rect 14740 63028 14792 63034
rect 14740 62970 14792 62976
rect 14289 62588 14585 62608
rect 14345 62586 14369 62588
rect 14425 62586 14449 62588
rect 14505 62586 14529 62588
rect 14367 62534 14369 62586
rect 14431 62534 14443 62586
rect 14505 62534 14507 62586
rect 14345 62532 14369 62534
rect 14425 62532 14449 62534
rect 14505 62532 14529 62534
rect 14289 62512 14585 62532
rect 14280 62348 14332 62354
rect 14280 62290 14332 62296
rect 14292 61878 14320 62290
rect 14752 61946 14780 62970
rect 14740 61940 14792 61946
rect 14740 61882 14792 61888
rect 14280 61872 14332 61878
rect 14280 61814 14332 61820
rect 14648 61872 14700 61878
rect 14648 61814 14700 61820
rect 14289 61500 14585 61520
rect 14345 61498 14369 61500
rect 14425 61498 14449 61500
rect 14505 61498 14529 61500
rect 14367 61446 14369 61498
rect 14431 61446 14443 61498
rect 14505 61446 14507 61498
rect 14345 61444 14369 61446
rect 14425 61444 14449 61446
rect 14505 61444 14529 61446
rect 14289 61424 14585 61444
rect 14660 61266 14688 61814
rect 14752 61742 14780 61882
rect 14740 61736 14792 61742
rect 14740 61678 14792 61684
rect 14648 61260 14700 61266
rect 14648 61202 14700 61208
rect 14660 60790 14688 61202
rect 14738 61024 14794 61033
rect 14738 60959 14794 60968
rect 14648 60784 14700 60790
rect 14094 60752 14150 60761
rect 14752 60761 14780 60959
rect 14648 60726 14700 60732
rect 14738 60752 14794 60761
rect 14094 60687 14150 60696
rect 14738 60687 14794 60696
rect 14289 60412 14585 60432
rect 14345 60410 14369 60412
rect 14425 60410 14449 60412
rect 14505 60410 14529 60412
rect 14367 60358 14369 60410
rect 14431 60358 14443 60410
rect 14505 60358 14507 60410
rect 14345 60356 14369 60358
rect 14425 60356 14449 60358
rect 14505 60356 14529 60358
rect 14289 60336 14585 60356
rect 14738 60344 14794 60353
rect 14738 60279 14740 60288
rect 14792 60279 14794 60288
rect 14740 60250 14792 60256
rect 14186 60208 14242 60217
rect 14186 60143 14242 60152
rect 14094 60072 14150 60081
rect 14004 60036 14056 60042
rect 14094 60007 14150 60016
rect 14004 59978 14056 59984
rect 14016 59770 14044 59978
rect 14108 59770 14136 60007
rect 14004 59764 14056 59770
rect 14004 59706 14056 59712
rect 14096 59764 14148 59770
rect 14096 59706 14148 59712
rect 14002 59528 14058 59537
rect 14002 59463 14058 59472
rect 13820 59220 13872 59226
rect 13820 59162 13872 59168
rect 13648 58534 13768 58562
rect 13636 58472 13688 58478
rect 13636 58414 13688 58420
rect 13544 57928 13596 57934
rect 13544 57870 13596 57876
rect 13464 57310 13584 57338
rect 13452 57248 13504 57254
rect 13452 57190 13504 57196
rect 13464 54534 13492 57190
rect 13452 54528 13504 54534
rect 13452 54470 13504 54476
rect 13464 52562 13492 54470
rect 13452 52556 13504 52562
rect 13452 52498 13504 52504
rect 13452 52420 13504 52426
rect 13452 52362 13504 52368
rect 13358 51096 13414 51105
rect 13176 51060 13228 51066
rect 13464 51066 13492 52362
rect 13358 51031 13414 51040
rect 13452 51060 13504 51066
rect 13176 51002 13228 51008
rect 13452 51002 13504 51008
rect 13450 50960 13506 50969
rect 13176 50924 13228 50930
rect 13450 50895 13506 50904
rect 13176 50866 13228 50872
rect 13188 50522 13216 50866
rect 13358 50824 13414 50833
rect 13268 50788 13320 50794
rect 13358 50759 13414 50768
rect 13268 50730 13320 50736
rect 13176 50516 13228 50522
rect 13176 50458 13228 50464
rect 13176 50380 13228 50386
rect 13176 50322 13228 50328
rect 13188 50289 13216 50322
rect 13174 50280 13230 50289
rect 13174 50215 13230 50224
rect 13176 49836 13228 49842
rect 13176 49778 13228 49784
rect 13188 46889 13216 49778
rect 13280 48226 13308 50730
rect 13372 50386 13400 50759
rect 13360 50380 13412 50386
rect 13360 50322 13412 50328
rect 13372 49978 13400 50322
rect 13360 49972 13412 49978
rect 13360 49914 13412 49920
rect 13358 49872 13414 49881
rect 13358 49807 13414 49816
rect 13372 48754 13400 49807
rect 13360 48748 13412 48754
rect 13360 48690 13412 48696
rect 13280 48198 13400 48226
rect 13268 48136 13320 48142
rect 13266 48104 13268 48113
rect 13320 48104 13322 48113
rect 13266 48039 13322 48048
rect 13280 47802 13308 48039
rect 13268 47796 13320 47802
rect 13268 47738 13320 47744
rect 13268 47048 13320 47054
rect 13268 46990 13320 46996
rect 13174 46880 13230 46889
rect 13174 46815 13230 46824
rect 13280 46730 13308 46990
rect 13188 46714 13308 46730
rect 13176 46708 13308 46714
rect 13228 46702 13308 46708
rect 13176 46650 13228 46656
rect 13280 46617 13308 46702
rect 13266 46608 13322 46617
rect 13176 46572 13228 46578
rect 13266 46543 13322 46552
rect 13176 46514 13228 46520
rect 13084 46164 13136 46170
rect 13084 46106 13136 46112
rect 13188 46102 13216 46514
rect 13268 46504 13320 46510
rect 13268 46446 13320 46452
rect 13176 46096 13228 46102
rect 13004 46022 13124 46050
rect 13280 46073 13308 46446
rect 13176 46038 13228 46044
rect 13266 46064 13322 46073
rect 12900 45960 12952 45966
rect 12900 45902 12952 45908
rect 12992 45960 13044 45966
rect 12992 45902 13044 45908
rect 12912 45626 12940 45902
rect 12900 45620 12952 45626
rect 12900 45562 12952 45568
rect 12808 45552 12860 45558
rect 12808 45494 12860 45500
rect 12808 45416 12860 45422
rect 12808 45358 12860 45364
rect 12716 45076 12768 45082
rect 12716 45018 12768 45024
rect 12728 44402 12756 45018
rect 12716 44396 12768 44402
rect 12716 44338 12768 44344
rect 12716 44260 12768 44266
rect 12716 44202 12768 44208
rect 12728 43994 12756 44202
rect 12716 43988 12768 43994
rect 12716 43930 12768 43936
rect 12716 43648 12768 43654
rect 12716 43590 12768 43596
rect 12624 43444 12676 43450
rect 12624 43386 12676 43392
rect 12530 43344 12586 43353
rect 12530 43279 12586 43288
rect 12624 43172 12676 43178
rect 12624 43114 12676 43120
rect 12440 42900 12492 42906
rect 12440 42842 12492 42848
rect 12452 41188 12480 42842
rect 12532 42016 12584 42022
rect 12532 41958 12584 41964
rect 12544 41614 12572 41958
rect 12532 41608 12584 41614
rect 12532 41550 12584 41556
rect 12452 41160 12572 41188
rect 12440 40588 12492 40594
rect 12440 40530 12492 40536
rect 12346 40488 12402 40497
rect 12346 40423 12402 40432
rect 12348 40180 12400 40186
rect 12348 40122 12400 40128
rect 12360 39642 12388 40122
rect 12348 39636 12400 39642
rect 12348 39578 12400 39584
rect 12452 39574 12480 40530
rect 12544 39982 12572 41160
rect 12636 41138 12664 43114
rect 12728 42906 12756 43590
rect 12716 42900 12768 42906
rect 12716 42842 12768 42848
rect 12716 41472 12768 41478
rect 12716 41414 12768 41420
rect 12624 41132 12676 41138
rect 12624 41074 12676 41080
rect 12728 41070 12756 41414
rect 12716 41064 12768 41070
rect 12716 41006 12768 41012
rect 12624 40996 12676 41002
rect 12624 40938 12676 40944
rect 12636 40390 12664 40938
rect 12624 40384 12676 40390
rect 12624 40326 12676 40332
rect 12532 39976 12584 39982
rect 12532 39918 12584 39924
rect 12440 39568 12492 39574
rect 12440 39510 12492 39516
rect 12544 39420 12572 39918
rect 12452 39392 12572 39420
rect 12348 39024 12400 39030
rect 12348 38966 12400 38972
rect 12360 38486 12388 38966
rect 12452 38758 12480 39392
rect 12532 39092 12584 39098
rect 12532 39034 12584 39040
rect 12440 38752 12492 38758
rect 12440 38694 12492 38700
rect 12440 38548 12492 38554
rect 12440 38490 12492 38496
rect 12348 38480 12400 38486
rect 12348 38422 12400 38428
rect 12346 38312 12402 38321
rect 12346 38247 12402 38256
rect 12360 37466 12388 38247
rect 12452 37738 12480 38490
rect 12440 37732 12492 37738
rect 12440 37674 12492 37680
rect 12348 37460 12400 37466
rect 12348 37402 12400 37408
rect 12360 36922 12388 37402
rect 12452 37398 12480 37674
rect 12440 37392 12492 37398
rect 12440 37334 12492 37340
rect 12348 36916 12400 36922
rect 12348 36858 12400 36864
rect 12256 36644 12308 36650
rect 12256 36586 12308 36592
rect 12164 36372 12216 36378
rect 12164 36314 12216 36320
rect 12164 35760 12216 35766
rect 12164 35702 12216 35708
rect 12072 31136 12124 31142
rect 12072 31078 12124 31084
rect 12072 30048 12124 30054
rect 12072 29990 12124 29996
rect 12084 28966 12112 29990
rect 12072 28960 12124 28966
rect 12072 28902 12124 28908
rect 12084 28558 12112 28902
rect 12072 28552 12124 28558
rect 12176 28529 12204 35702
rect 12360 35698 12388 36858
rect 12452 36718 12480 37334
rect 12440 36712 12492 36718
rect 12440 36654 12492 36660
rect 12544 35834 12572 39034
rect 12636 37874 12664 40326
rect 12716 39432 12768 39438
rect 12716 39374 12768 39380
rect 12728 39098 12756 39374
rect 12716 39092 12768 39098
rect 12716 39034 12768 39040
rect 12820 38554 12848 45358
rect 12912 45014 12940 45562
rect 13004 45354 13032 45902
rect 12992 45348 13044 45354
rect 12992 45290 13044 45296
rect 13004 45082 13032 45290
rect 12992 45076 13044 45082
rect 12992 45018 13044 45024
rect 12900 45008 12952 45014
rect 12900 44950 12952 44956
rect 12900 44872 12952 44878
rect 12900 44814 12952 44820
rect 12912 43790 12940 44814
rect 13096 43858 13124 46022
rect 13266 45999 13322 46008
rect 13176 45960 13228 45966
rect 13176 45902 13228 45908
rect 13084 43852 13136 43858
rect 13084 43794 13136 43800
rect 12900 43784 12952 43790
rect 12900 43726 12952 43732
rect 12912 39438 12940 43726
rect 13096 43110 13124 43794
rect 13084 43104 13136 43110
rect 13084 43046 13136 43052
rect 13084 42696 13136 42702
rect 13188 42673 13216 45902
rect 13280 44146 13308 45999
rect 13372 44266 13400 48198
rect 13360 44260 13412 44266
rect 13360 44202 13412 44208
rect 13280 44118 13400 44146
rect 13268 43988 13320 43994
rect 13268 43930 13320 43936
rect 13280 42838 13308 43930
rect 13268 42832 13320 42838
rect 13268 42774 13320 42780
rect 13084 42638 13136 42644
rect 13174 42664 13230 42673
rect 13096 42362 13124 42638
rect 13174 42599 13230 42608
rect 13176 42560 13228 42566
rect 13176 42502 13228 42508
rect 13084 42356 13136 42362
rect 13084 42298 13136 42304
rect 12990 42256 13046 42265
rect 12990 42191 12992 42200
rect 13044 42191 13046 42200
rect 12992 42162 13044 42168
rect 13004 41682 13032 42162
rect 12992 41676 13044 41682
rect 12992 41618 13044 41624
rect 13188 41614 13216 42502
rect 13268 42220 13320 42226
rect 13268 42162 13320 42168
rect 13176 41608 13228 41614
rect 13174 41576 13176 41585
rect 13228 41576 13230 41585
rect 13174 41511 13230 41520
rect 12992 41064 13044 41070
rect 12992 41006 13044 41012
rect 12900 39432 12952 39438
rect 12900 39374 12952 39380
rect 13004 38962 13032 41006
rect 13084 40588 13136 40594
rect 13084 40530 13136 40536
rect 13096 39846 13124 40530
rect 13280 39930 13308 42162
rect 13188 39902 13308 39930
rect 13084 39840 13136 39846
rect 13082 39808 13084 39817
rect 13136 39808 13138 39817
rect 13082 39743 13138 39752
rect 13188 39624 13216 39902
rect 13268 39840 13320 39846
rect 13268 39782 13320 39788
rect 13096 39596 13216 39624
rect 12992 38956 13044 38962
rect 12992 38898 13044 38904
rect 12808 38548 12860 38554
rect 12808 38490 12860 38496
rect 12808 38276 12860 38282
rect 12808 38218 12860 38224
rect 12714 38176 12770 38185
rect 12714 38111 12770 38120
rect 12624 37868 12676 37874
rect 12624 37810 12676 37816
rect 12728 36378 12756 38111
rect 12820 36922 12848 38218
rect 12898 37360 12954 37369
rect 13096 37330 13124 39596
rect 13176 39500 13228 39506
rect 13176 39442 13228 39448
rect 12898 37295 12954 37304
rect 13084 37324 13136 37330
rect 12808 36916 12860 36922
rect 12808 36858 12860 36864
rect 12716 36372 12768 36378
rect 12716 36314 12768 36320
rect 12820 36310 12848 36858
rect 12912 36854 12940 37295
rect 13084 37266 13136 37272
rect 12900 36848 12952 36854
rect 12900 36790 12952 36796
rect 12808 36304 12860 36310
rect 12808 36246 12860 36252
rect 13082 36272 13138 36281
rect 13082 36207 13084 36216
rect 13136 36207 13138 36216
rect 13084 36178 13136 36184
rect 13096 35834 13124 36178
rect 12532 35828 12584 35834
rect 12532 35770 12584 35776
rect 13084 35828 13136 35834
rect 13084 35770 13136 35776
rect 12348 35692 12400 35698
rect 12348 35634 12400 35640
rect 13096 35222 13124 35770
rect 13084 35216 13136 35222
rect 13084 35158 13136 35164
rect 12806 33552 12862 33561
rect 12806 33487 12862 33496
rect 12622 33280 12678 33289
rect 12622 33215 12678 33224
rect 12636 32026 12664 33215
rect 12624 32020 12676 32026
rect 12624 31962 12676 31968
rect 12440 31884 12492 31890
rect 12440 31826 12492 31832
rect 12452 31210 12480 31826
rect 12440 31204 12492 31210
rect 12440 31146 12492 31152
rect 12716 30592 12768 30598
rect 12716 30534 12768 30540
rect 12728 30190 12756 30534
rect 12716 30184 12768 30190
rect 12716 30126 12768 30132
rect 12532 30048 12584 30054
rect 12532 29990 12584 29996
rect 12360 29668 12480 29696
rect 12256 29504 12308 29510
rect 12256 29446 12308 29452
rect 12268 29170 12296 29446
rect 12256 29164 12308 29170
rect 12256 29106 12308 29112
rect 12072 28494 12124 28500
rect 12162 28520 12218 28529
rect 12084 28422 12112 28494
rect 12162 28455 12218 28464
rect 12072 28416 12124 28422
rect 12072 28358 12124 28364
rect 11978 28112 12034 28121
rect 11978 28047 12034 28056
rect 11888 28008 11940 28014
rect 12084 27996 12112 28358
rect 11888 27950 11940 27956
rect 11992 27968 12112 27996
rect 11900 27334 11928 27950
rect 11888 27328 11940 27334
rect 11888 27270 11940 27276
rect 11796 27056 11848 27062
rect 11796 26998 11848 27004
rect 11808 26790 11836 26998
rect 11900 26858 11928 27270
rect 11888 26852 11940 26858
rect 11888 26794 11940 26800
rect 11796 26784 11848 26790
rect 11796 26726 11848 26732
rect 11348 26540 11468 26568
rect 11520 26580 11572 26586
rect 11150 26344 11206 26353
rect 11150 26279 11152 26288
rect 11204 26279 11206 26288
rect 11152 26250 11204 26256
rect 10956 26140 11252 26160
rect 11012 26138 11036 26140
rect 11092 26138 11116 26140
rect 11172 26138 11196 26140
rect 11034 26086 11036 26138
rect 11098 26086 11110 26138
rect 11172 26086 11174 26138
rect 11012 26084 11036 26086
rect 11092 26084 11116 26086
rect 11172 26084 11196 26086
rect 10956 26064 11252 26084
rect 10876 25764 10928 25770
rect 10876 25706 10928 25712
rect 10956 25052 11252 25072
rect 11012 25050 11036 25052
rect 11092 25050 11116 25052
rect 11172 25050 11196 25052
rect 11034 24998 11036 25050
rect 11098 24998 11110 25050
rect 11172 24998 11174 25050
rect 11012 24996 11036 24998
rect 11092 24996 11116 24998
rect 11172 24996 11196 24998
rect 10956 24976 11252 24996
rect 10784 24744 10836 24750
rect 10784 24686 10836 24692
rect 11348 24274 11376 26540
rect 11520 26522 11572 26528
rect 11428 26444 11480 26450
rect 11428 26386 11480 26392
rect 11440 25702 11468 26386
rect 11900 26314 11928 26794
rect 11888 26308 11940 26314
rect 11888 26250 11940 26256
rect 11428 25696 11480 25702
rect 11428 25638 11480 25644
rect 11440 24993 11468 25638
rect 11426 24984 11482 24993
rect 11426 24919 11482 24928
rect 11520 24608 11572 24614
rect 11520 24550 11572 24556
rect 10876 24268 10928 24274
rect 10876 24210 10928 24216
rect 11336 24268 11388 24274
rect 11336 24210 11388 24216
rect 10888 23798 10916 24210
rect 10956 23964 11252 23984
rect 11012 23962 11036 23964
rect 11092 23962 11116 23964
rect 11172 23962 11196 23964
rect 11034 23910 11036 23962
rect 11098 23910 11110 23962
rect 11172 23910 11174 23962
rect 11012 23908 11036 23910
rect 11092 23908 11116 23910
rect 11172 23908 11196 23910
rect 10956 23888 11252 23908
rect 11348 23866 11376 24210
rect 11336 23860 11388 23866
rect 11336 23802 11388 23808
rect 10876 23792 10928 23798
rect 10928 23740 11100 23746
rect 10876 23734 11100 23740
rect 10888 23718 11100 23734
rect 10888 23669 10916 23718
rect 11072 23322 11100 23718
rect 10520 23276 10640 23304
rect 11060 23316 11112 23322
rect 10416 23180 10468 23186
rect 10416 23122 10468 23128
rect 10230 22944 10286 22953
rect 10230 22879 10286 22888
rect 10428 22778 10456 23122
rect 10416 22772 10468 22778
rect 10416 22714 10468 22720
rect 9956 22704 10008 22710
rect 10520 22658 10548 23276
rect 11060 23258 11112 23264
rect 10600 23180 10652 23186
rect 10600 23122 10652 23128
rect 10612 22778 10640 23122
rect 11428 23112 11480 23118
rect 11428 23054 11480 23060
rect 10956 22876 11252 22896
rect 11012 22874 11036 22876
rect 11092 22874 11116 22876
rect 11172 22874 11196 22876
rect 11034 22822 11036 22874
rect 11098 22822 11110 22874
rect 11172 22822 11174 22874
rect 11012 22820 11036 22822
rect 11092 22820 11116 22822
rect 11172 22820 11196 22822
rect 10956 22800 11252 22820
rect 11440 22778 11468 23054
rect 10600 22772 10652 22778
rect 10600 22714 10652 22720
rect 11428 22772 11480 22778
rect 11428 22714 11480 22720
rect 9956 22646 10008 22652
rect 10428 22630 10548 22658
rect 10968 22704 11020 22710
rect 10968 22646 11020 22652
rect 11426 22672 11482 22681
rect 9864 22500 9916 22506
rect 9864 22442 9916 22448
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9862 22264 9918 22273
rect 9692 22222 9812 22250
rect 9680 22160 9732 22166
rect 9678 22128 9680 22137
rect 9732 22128 9734 22137
rect 9678 22063 9734 22072
rect 9784 19553 9812 22222
rect 9862 22199 9918 22208
rect 9876 22098 9904 22199
rect 9864 22092 9916 22098
rect 9864 22034 9916 22040
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 10060 21690 10088 22034
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 10244 21690 10272 21966
rect 10048 21684 10100 21690
rect 10048 21626 10100 21632
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 9864 20392 9916 20398
rect 9864 20334 9916 20340
rect 9876 19718 9904 20334
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 9770 19544 9826 19553
rect 9770 19479 9826 19488
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9692 16697 9720 17070
rect 9770 16960 9826 16969
rect 9876 16946 9904 19654
rect 10428 19360 10456 22630
rect 10508 22568 10560 22574
rect 10508 22510 10560 22516
rect 10520 22137 10548 22510
rect 10506 22128 10562 22137
rect 10980 22098 11008 22646
rect 11426 22607 11482 22616
rect 11336 22432 11388 22438
rect 11336 22374 11388 22380
rect 10506 22063 10562 22072
rect 10968 22092 11020 22098
rect 10968 22034 11020 22040
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 10704 21622 10732 21966
rect 10956 21788 11252 21808
rect 11012 21786 11036 21788
rect 11092 21786 11116 21788
rect 11172 21786 11196 21788
rect 11034 21734 11036 21786
rect 11098 21734 11110 21786
rect 11172 21734 11174 21786
rect 11012 21732 11036 21734
rect 11092 21732 11116 21734
rect 11172 21732 11196 21734
rect 10956 21712 11252 21732
rect 10692 21616 10744 21622
rect 10692 21558 10744 21564
rect 10956 20700 11252 20720
rect 11012 20698 11036 20700
rect 11092 20698 11116 20700
rect 11172 20698 11196 20700
rect 11034 20646 11036 20698
rect 11098 20646 11110 20698
rect 11172 20646 11174 20698
rect 11012 20644 11036 20646
rect 11092 20644 11116 20646
rect 11172 20644 11196 20646
rect 10956 20624 11252 20644
rect 10956 19612 11252 19632
rect 11012 19610 11036 19612
rect 11092 19610 11116 19612
rect 11172 19610 11196 19612
rect 11034 19558 11036 19610
rect 11098 19558 11110 19610
rect 11172 19558 11174 19610
rect 11012 19556 11036 19558
rect 11092 19556 11116 19558
rect 11172 19556 11196 19558
rect 10956 19536 11252 19556
rect 11348 19394 11376 22374
rect 9826 16918 9904 16946
rect 10152 19332 10456 19360
rect 11256 19366 11376 19394
rect 9770 16895 9826 16904
rect 9678 16688 9734 16697
rect 9678 16623 9680 16632
rect 9732 16623 9734 16632
rect 9680 16594 9732 16600
rect 9784 15502 9812 16895
rect 10152 15706 10180 19332
rect 11256 18873 11284 19366
rect 10782 18864 10838 18873
rect 11242 18864 11298 18873
rect 10782 18799 10784 18808
rect 10836 18799 10838 18808
rect 10876 18828 10928 18834
rect 10784 18770 10836 18776
rect 11242 18799 11298 18808
rect 11336 18828 11388 18834
rect 10876 18770 10928 18776
rect 11336 18770 11388 18776
rect 10796 17882 10824 18770
rect 10888 18426 10916 18770
rect 10956 18524 11252 18544
rect 11012 18522 11036 18524
rect 11092 18522 11116 18524
rect 11172 18522 11196 18524
rect 11034 18470 11036 18522
rect 11098 18470 11110 18522
rect 11172 18470 11174 18522
rect 11012 18468 11036 18470
rect 11092 18468 11116 18470
rect 11172 18468 11196 18470
rect 10956 18448 11252 18468
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10784 17876 10836 17882
rect 10784 17818 10836 17824
rect 11348 17746 11376 18770
rect 11336 17740 11388 17746
rect 11336 17682 11388 17688
rect 10956 17436 11252 17456
rect 11012 17434 11036 17436
rect 11092 17434 11116 17436
rect 11172 17434 11196 17436
rect 11034 17382 11036 17434
rect 11098 17382 11110 17434
rect 11172 17382 11174 17434
rect 11012 17380 11036 17382
rect 11092 17380 11116 17382
rect 11172 17380 11196 17382
rect 10956 17360 11252 17380
rect 11348 17338 11376 17682
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 11072 16538 11100 16934
rect 11334 16688 11390 16697
rect 11334 16623 11390 16632
rect 10888 16510 11100 16538
rect 10888 16250 10916 16510
rect 10956 16348 11252 16368
rect 11012 16346 11036 16348
rect 11092 16346 11116 16348
rect 11172 16346 11196 16348
rect 11034 16294 11036 16346
rect 11098 16294 11110 16346
rect 11172 16294 11174 16346
rect 11012 16292 11036 16294
rect 11092 16292 11116 16294
rect 11172 16292 11196 16294
rect 10956 16272 11252 16292
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 11348 16114 11376 16623
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 10876 15972 10928 15978
rect 10876 15914 10928 15920
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 9864 15564 9916 15570
rect 9864 15506 9916 15512
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9876 14822 9904 15506
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10244 14822 10272 15438
rect 10888 15162 10916 15914
rect 11440 15638 11468 22607
rect 11532 22030 11560 24550
rect 11900 23186 11928 26250
rect 11992 25265 12020 27968
rect 12084 25838 12112 25869
rect 12072 25832 12124 25838
rect 12070 25800 12072 25809
rect 12124 25800 12126 25809
rect 12070 25735 12126 25744
rect 12084 25498 12112 25735
rect 12164 25696 12216 25702
rect 12162 25664 12164 25673
rect 12216 25664 12218 25673
rect 12162 25599 12218 25608
rect 12072 25492 12124 25498
rect 12072 25434 12124 25440
rect 11978 25256 12034 25265
rect 11978 25191 12034 25200
rect 11992 23882 12020 25191
rect 11992 23866 12112 23882
rect 11980 23860 12112 23866
rect 12032 23854 12112 23860
rect 11980 23802 12032 23808
rect 11978 23760 12034 23769
rect 11978 23695 12034 23704
rect 11888 23180 11940 23186
rect 11888 23122 11940 23128
rect 11520 22024 11572 22030
rect 11520 21966 11572 21972
rect 11888 20324 11940 20330
rect 11888 20266 11940 20272
rect 11612 19236 11664 19242
rect 11612 19178 11664 19184
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11428 15632 11480 15638
rect 11428 15574 11480 15580
rect 10956 15260 11252 15280
rect 11012 15258 11036 15260
rect 11092 15258 11116 15260
rect 11172 15258 11196 15260
rect 11034 15206 11036 15258
rect 11098 15206 11110 15258
rect 11172 15206 11174 15258
rect 11012 15204 11036 15206
rect 11092 15204 11116 15206
rect 11172 15204 11196 15206
rect 10956 15184 11252 15204
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10888 14958 10916 15098
rect 10876 14952 10928 14958
rect 10796 14900 10876 14906
rect 10796 14894 10928 14900
rect 10796 14878 10916 14894
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 9876 14521 9904 14758
rect 9862 14512 9918 14521
rect 9862 14447 9918 14456
rect 9772 13184 9824 13190
rect 9770 13152 9772 13161
rect 9824 13152 9826 13161
rect 9770 13087 9826 13096
rect 9784 12782 9812 13087
rect 10244 13025 10272 14758
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10704 13870 10732 14418
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 10336 13394 10364 13670
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10336 13297 10364 13330
rect 10322 13288 10378 13297
rect 10322 13223 10378 13232
rect 10230 13016 10286 13025
rect 10230 12951 10286 12960
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10520 12374 10548 12582
rect 10508 12368 10560 12374
rect 10508 12310 10560 12316
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 10152 11694 10180 12242
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10520 11898 10548 12106
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10140 11688 10192 11694
rect 9586 11656 9642 11665
rect 10140 11630 10192 11636
rect 9586 11591 9642 11600
rect 9600 10130 9628 11591
rect 10152 11218 10180 11630
rect 10704 11558 10732 13806
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9692 10810 9720 11086
rect 10060 11082 10088 11154
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9784 10690 9812 10950
rect 9692 10662 9812 10690
rect 9692 10606 9720 10662
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9508 9586 9536 9998
rect 9600 9654 9628 10066
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9508 9042 9536 9522
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9508 8498 9536 8978
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9600 5760 9628 7482
rect 9692 7313 9720 10542
rect 10060 9382 10088 11018
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10152 10305 10180 10950
rect 10796 10554 10824 14878
rect 10956 14172 11252 14192
rect 11012 14170 11036 14172
rect 11092 14170 11116 14172
rect 11172 14170 11196 14172
rect 11034 14118 11036 14170
rect 11098 14118 11110 14170
rect 11172 14118 11174 14170
rect 11012 14116 11036 14118
rect 11092 14116 11116 14118
rect 11172 14116 11196 14118
rect 10956 14096 11252 14116
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10888 13394 10916 13670
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10888 12782 10916 13330
rect 10956 13084 11252 13104
rect 11012 13082 11036 13084
rect 11092 13082 11116 13084
rect 11172 13082 11196 13084
rect 11034 13030 11036 13082
rect 11098 13030 11110 13082
rect 11172 13030 11174 13082
rect 11012 13028 11036 13030
rect 11092 13028 11116 13030
rect 11172 13028 11196 13030
rect 10956 13008 11252 13028
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 11348 12594 11376 13466
rect 11532 13410 11560 18702
rect 11624 18086 11652 19178
rect 11796 19168 11848 19174
rect 11794 19136 11796 19145
rect 11848 19136 11850 19145
rect 11794 19071 11850 19080
rect 11900 18834 11928 20266
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 11888 18692 11940 18698
rect 11888 18634 11940 18640
rect 11900 18222 11928 18634
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11888 18216 11940 18222
rect 11888 18158 11940 18164
rect 11612 18080 11664 18086
rect 11612 18022 11664 18028
rect 11808 17882 11836 18158
rect 11796 17876 11848 17882
rect 11716 17836 11796 17864
rect 11612 16448 11664 16454
rect 11612 16390 11664 16396
rect 11624 16046 11652 16390
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11440 13394 11560 13410
rect 11428 13388 11560 13394
rect 11480 13382 11560 13388
rect 11428 13330 11480 13336
rect 11532 12850 11560 13382
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11520 12708 11572 12714
rect 11520 12650 11572 12656
rect 11256 12566 11376 12594
rect 11256 12238 11284 12566
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 10956 11996 11252 12016
rect 11012 11994 11036 11996
rect 11092 11994 11116 11996
rect 11172 11994 11196 11996
rect 11034 11942 11036 11994
rect 11098 11942 11110 11994
rect 11172 11942 11174 11994
rect 11012 11940 11036 11942
rect 11092 11940 11116 11942
rect 11172 11940 11196 11942
rect 10956 11920 11252 11940
rect 11348 11778 11376 12378
rect 11532 12186 11560 12650
rect 11624 12322 11652 15982
rect 11716 15094 11744 17836
rect 11796 17818 11848 17824
rect 11794 17640 11850 17649
rect 11794 17575 11850 17584
rect 11808 16590 11836 17575
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11900 16998 11928 17478
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 11704 15088 11756 15094
rect 11704 15030 11756 15036
rect 11716 14550 11744 15030
rect 11808 14958 11836 15302
rect 11796 14952 11848 14958
rect 11796 14894 11848 14900
rect 11704 14544 11756 14550
rect 11704 14486 11756 14492
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11716 12442 11744 14214
rect 11808 12850 11836 14894
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11624 12294 11744 12322
rect 11532 12158 11652 12186
rect 11624 12102 11652 12158
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 11256 11750 11376 11778
rect 11072 11393 11100 11698
rect 11058 11384 11114 11393
rect 11058 11319 11114 11328
rect 11256 11150 11284 11750
rect 11440 11694 11468 12038
rect 11428 11688 11480 11694
rect 11348 11636 11428 11642
rect 11716 11642 11744 12294
rect 11808 11694 11836 12378
rect 11900 12306 11928 16934
rect 11992 12442 12020 23695
rect 12084 23662 12112 23854
rect 12072 23656 12124 23662
rect 12072 23598 12124 23604
rect 12072 21344 12124 21350
rect 12072 21286 12124 21292
rect 12084 18465 12112 21286
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 12176 20058 12204 20198
rect 12164 20052 12216 20058
rect 12164 19994 12216 20000
rect 12164 19508 12216 19514
rect 12164 19450 12216 19456
rect 12176 19417 12204 19450
rect 12162 19408 12218 19417
rect 12162 19343 12218 19352
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 12070 18456 12126 18465
rect 12070 18391 12126 18400
rect 12176 18358 12204 19110
rect 12164 18352 12216 18358
rect 12164 18294 12216 18300
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 12084 13002 12112 18022
rect 12164 17264 12216 17270
rect 12164 17206 12216 17212
rect 12176 14074 12204 17206
rect 12268 16998 12296 29106
rect 12360 28762 12388 29668
rect 12452 29578 12480 29668
rect 12440 29572 12492 29578
rect 12440 29514 12492 29520
rect 12348 28756 12400 28762
rect 12348 28698 12400 28704
rect 12360 28082 12388 28698
rect 12440 28620 12492 28626
rect 12440 28562 12492 28568
rect 12348 28076 12400 28082
rect 12348 28018 12400 28024
rect 12452 28014 12480 28562
rect 12544 28490 12572 29990
rect 12624 29640 12676 29646
rect 12624 29582 12676 29588
rect 12636 29102 12664 29582
rect 12624 29096 12676 29102
rect 12624 29038 12676 29044
rect 12636 28966 12664 29038
rect 12624 28960 12676 28966
rect 12624 28902 12676 28908
rect 12636 28694 12664 28902
rect 12728 28762 12756 30126
rect 12716 28756 12768 28762
rect 12716 28698 12768 28704
rect 12624 28688 12676 28694
rect 12624 28630 12676 28636
rect 12532 28484 12584 28490
rect 12532 28426 12584 28432
rect 12440 28008 12492 28014
rect 12440 27950 12492 27956
rect 12544 27690 12572 28426
rect 12636 27878 12664 28630
rect 12624 27872 12676 27878
rect 12676 27820 12756 27826
rect 12624 27814 12756 27820
rect 12636 27798 12756 27814
rect 12544 27662 12664 27690
rect 12532 25764 12584 25770
rect 12532 25706 12584 25712
rect 12348 23248 12400 23254
rect 12348 23190 12400 23196
rect 12360 21690 12388 23190
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12452 22438 12480 23122
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 12544 22250 12572 25706
rect 12636 25430 12664 27662
rect 12728 27538 12756 27798
rect 12716 27532 12768 27538
rect 12716 27474 12768 27480
rect 12728 27402 12756 27474
rect 12716 27396 12768 27402
rect 12716 27338 12768 27344
rect 12728 27130 12756 27338
rect 12716 27124 12768 27130
rect 12716 27066 12768 27072
rect 12716 26376 12768 26382
rect 12716 26318 12768 26324
rect 12728 25702 12756 26318
rect 12820 26042 12848 33487
rect 12900 32224 12952 32230
rect 12900 32166 12952 32172
rect 12912 30326 12940 32166
rect 13188 31793 13216 39442
rect 13280 35494 13308 39782
rect 13372 38185 13400 44118
rect 13464 39506 13492 50895
rect 13556 50153 13584 57310
rect 13542 50144 13598 50153
rect 13542 50079 13598 50088
rect 13648 49960 13676 58414
rect 13740 56817 13768 58534
rect 13832 57934 13860 59162
rect 13912 59016 13964 59022
rect 13912 58958 13964 58964
rect 13820 57928 13872 57934
rect 13820 57870 13872 57876
rect 13924 57798 13952 58958
rect 13912 57792 13964 57798
rect 13912 57734 13964 57740
rect 13726 56808 13782 56817
rect 13726 56743 13782 56752
rect 13726 56264 13782 56273
rect 13726 56199 13728 56208
rect 13780 56199 13782 56208
rect 13728 56170 13780 56176
rect 13728 55888 13780 55894
rect 13728 55830 13780 55836
rect 13740 55457 13768 55830
rect 13912 55752 13964 55758
rect 13912 55694 13964 55700
rect 13726 55448 13782 55457
rect 13924 55418 13952 55694
rect 13726 55383 13782 55392
rect 13912 55412 13964 55418
rect 13740 54754 13768 55383
rect 13912 55354 13964 55360
rect 13820 55276 13872 55282
rect 13820 55218 13872 55224
rect 13832 54874 13860 55218
rect 13820 54868 13872 54874
rect 13820 54810 13872 54816
rect 13740 54726 13860 54754
rect 13728 54664 13780 54670
rect 13728 54606 13780 54612
rect 13740 53990 13768 54606
rect 13728 53984 13780 53990
rect 13728 53926 13780 53932
rect 13740 52057 13768 53926
rect 13832 52086 13860 54726
rect 14016 54108 14044 59463
rect 14096 58336 14148 58342
rect 14096 58278 14148 58284
rect 14108 58041 14136 58278
rect 14094 58032 14150 58041
rect 14094 57967 14150 57976
rect 14200 56794 14228 60143
rect 14844 59974 14872 63174
rect 15028 63034 15056 68750
rect 15108 68128 15160 68134
rect 15108 68070 15160 68076
rect 15120 66586 15148 68070
rect 15292 67788 15344 67794
rect 15292 67730 15344 67736
rect 15304 67046 15332 67730
rect 15948 67726 15976 68750
rect 15936 67720 15988 67726
rect 15936 67662 15988 67668
rect 15948 67182 15976 67662
rect 15384 67176 15436 67182
rect 15384 67118 15436 67124
rect 15936 67176 15988 67182
rect 15936 67118 15988 67124
rect 15292 67040 15344 67046
rect 15292 66982 15344 66988
rect 15200 66632 15252 66638
rect 15120 66580 15200 66586
rect 15120 66574 15252 66580
rect 15120 66558 15240 66574
rect 15120 65958 15148 66558
rect 15108 65952 15160 65958
rect 15108 65894 15160 65900
rect 15120 64938 15240 64954
rect 15108 64932 15240 64938
rect 15160 64926 15240 64932
rect 15108 64874 15160 64880
rect 15108 64524 15160 64530
rect 15108 64466 15160 64472
rect 15120 64122 15148 64466
rect 15108 64116 15160 64122
rect 15108 64058 15160 64064
rect 15120 63442 15148 64058
rect 15108 63436 15160 63442
rect 15108 63378 15160 63384
rect 15212 63345 15240 64926
rect 15198 63336 15254 63345
rect 15198 63271 15254 63280
rect 15016 63028 15068 63034
rect 15016 62970 15068 62976
rect 15016 62824 15068 62830
rect 15016 62766 15068 62772
rect 15028 61878 15056 62766
rect 15198 62384 15254 62393
rect 15198 62319 15254 62328
rect 15212 62286 15240 62319
rect 15200 62280 15252 62286
rect 15200 62222 15252 62228
rect 15304 62098 15332 66982
rect 15396 66094 15424 67118
rect 15948 66842 15976 67118
rect 15936 66836 15988 66842
rect 15936 66778 15988 66784
rect 15476 66156 15528 66162
rect 15476 66098 15528 66104
rect 15384 66088 15436 66094
rect 15384 66030 15436 66036
rect 15396 65754 15424 66030
rect 15384 65748 15436 65754
rect 15384 65690 15436 65696
rect 15396 63986 15424 65690
rect 15384 63980 15436 63986
rect 15384 63922 15436 63928
rect 15382 63880 15438 63889
rect 15382 63815 15438 63824
rect 15396 62529 15424 63815
rect 15382 62520 15438 62529
rect 15382 62455 15438 62464
rect 15212 62070 15332 62098
rect 15384 62144 15436 62150
rect 15384 62086 15436 62092
rect 15016 61872 15068 61878
rect 15016 61814 15068 61820
rect 14924 61600 14976 61606
rect 14924 61542 14976 61548
rect 14936 61033 14964 61542
rect 15016 61192 15068 61198
rect 15016 61134 15068 61140
rect 14922 61024 14978 61033
rect 14922 60959 14978 60968
rect 15028 60518 15056 61134
rect 15016 60512 15068 60518
rect 15016 60454 15068 60460
rect 14832 59968 14884 59974
rect 14832 59910 14884 59916
rect 14289 59324 14585 59344
rect 14345 59322 14369 59324
rect 14425 59322 14449 59324
rect 14505 59322 14529 59324
rect 14367 59270 14369 59322
rect 14431 59270 14443 59322
rect 14505 59270 14507 59322
rect 14345 59268 14369 59270
rect 14425 59268 14449 59270
rect 14505 59268 14529 59270
rect 14289 59248 14585 59268
rect 14830 59120 14886 59129
rect 14830 59055 14886 59064
rect 14844 59022 14872 59055
rect 14832 59016 14884 59022
rect 14832 58958 14884 58964
rect 14648 58880 14700 58886
rect 14648 58822 14700 58828
rect 14660 58682 14688 58822
rect 14648 58676 14700 58682
rect 14648 58618 14700 58624
rect 14289 58236 14585 58256
rect 14345 58234 14369 58236
rect 14425 58234 14449 58236
rect 14505 58234 14529 58236
rect 14367 58182 14369 58234
rect 14431 58182 14443 58234
rect 14505 58182 14507 58234
rect 14345 58180 14369 58182
rect 14425 58180 14449 58182
rect 14505 58180 14529 58182
rect 14289 58160 14585 58180
rect 14830 58032 14886 58041
rect 14830 57967 14886 57976
rect 14648 57520 14700 57526
rect 14648 57462 14700 57468
rect 14289 57148 14585 57168
rect 14345 57146 14369 57148
rect 14425 57146 14449 57148
rect 14505 57146 14529 57148
rect 14367 57094 14369 57146
rect 14431 57094 14443 57146
rect 14505 57094 14507 57146
rect 14345 57092 14369 57094
rect 14425 57092 14449 57094
rect 14505 57092 14529 57094
rect 14289 57072 14585 57092
rect 14108 56766 14228 56794
rect 14108 54210 14136 56766
rect 14188 56704 14240 56710
rect 14188 56646 14240 56652
rect 14200 56166 14228 56646
rect 14188 56160 14240 56166
rect 14188 56102 14240 56108
rect 14200 55826 14228 56102
rect 14289 56060 14585 56080
rect 14345 56058 14369 56060
rect 14425 56058 14449 56060
rect 14505 56058 14529 56060
rect 14367 56006 14369 56058
rect 14431 56006 14443 56058
rect 14505 56006 14507 56058
rect 14345 56004 14369 56006
rect 14425 56004 14449 56006
rect 14505 56004 14529 56006
rect 14289 55984 14585 56004
rect 14188 55820 14240 55826
rect 14188 55762 14240 55768
rect 14370 55448 14426 55457
rect 14370 55383 14426 55392
rect 14188 55344 14240 55350
rect 14186 55312 14188 55321
rect 14240 55312 14242 55321
rect 14186 55247 14242 55256
rect 14384 55214 14412 55383
rect 14372 55208 14424 55214
rect 14372 55150 14424 55156
rect 14289 54972 14585 54992
rect 14345 54970 14369 54972
rect 14425 54970 14449 54972
rect 14505 54970 14529 54972
rect 14367 54918 14369 54970
rect 14431 54918 14443 54970
rect 14505 54918 14507 54970
rect 14345 54916 14369 54918
rect 14425 54916 14449 54918
rect 14505 54916 14529 54918
rect 14289 54896 14585 54916
rect 14660 54777 14688 57462
rect 14740 55072 14792 55078
rect 14740 55014 14792 55020
rect 14646 54768 14702 54777
rect 14646 54703 14702 54712
rect 14108 54182 14228 54210
rect 14096 54120 14148 54126
rect 14016 54080 14096 54108
rect 14096 54062 14148 54068
rect 14004 53984 14056 53990
rect 14004 53926 14056 53932
rect 13912 52624 13964 52630
rect 13912 52566 13964 52572
rect 13924 52465 13952 52566
rect 13910 52456 13966 52465
rect 13910 52391 13966 52400
rect 14016 52306 14044 53926
rect 14200 53786 14228 54182
rect 14289 53884 14585 53904
rect 14345 53882 14369 53884
rect 14425 53882 14449 53884
rect 14505 53882 14529 53884
rect 14367 53830 14369 53882
rect 14431 53830 14443 53882
rect 14505 53830 14507 53882
rect 14345 53828 14369 53830
rect 14425 53828 14449 53830
rect 14505 53828 14529 53830
rect 14289 53808 14585 53828
rect 14188 53780 14240 53786
rect 14660 53768 14688 54703
rect 14188 53722 14240 53728
rect 14568 53740 14688 53768
rect 14096 53508 14148 53514
rect 14096 53450 14148 53456
rect 14108 52426 14136 53450
rect 14200 53106 14228 53722
rect 14188 53100 14240 53106
rect 14188 53042 14240 53048
rect 14568 53038 14596 53740
rect 14752 53689 14780 55014
rect 14738 53680 14794 53689
rect 14648 53644 14700 53650
rect 14738 53615 14794 53624
rect 14648 53586 14700 53592
rect 14660 53446 14688 53586
rect 14648 53440 14700 53446
rect 14648 53382 14700 53388
rect 14660 53174 14688 53382
rect 14648 53168 14700 53174
rect 14648 53110 14700 53116
rect 14556 53032 14608 53038
rect 14556 52974 14608 52980
rect 14188 52896 14240 52902
rect 14188 52838 14240 52844
rect 14096 52420 14148 52426
rect 14096 52362 14148 52368
rect 13924 52278 14044 52306
rect 13924 52154 13952 52278
rect 13912 52148 13964 52154
rect 13912 52090 13964 52096
rect 14004 52148 14056 52154
rect 14004 52090 14056 52096
rect 13820 52080 13872 52086
rect 13726 52048 13782 52057
rect 13820 52022 13872 52028
rect 13726 51983 13782 51992
rect 13726 51912 13782 51921
rect 13726 51847 13728 51856
rect 13780 51847 13782 51856
rect 13728 51818 13780 51824
rect 13728 51060 13780 51066
rect 13728 51002 13780 51008
rect 13740 50969 13768 51002
rect 13726 50960 13782 50969
rect 13726 50895 13782 50904
rect 13728 50856 13780 50862
rect 13728 50798 13780 50804
rect 13556 49932 13676 49960
rect 13556 48793 13584 49932
rect 13636 49632 13688 49638
rect 13636 49574 13688 49580
rect 13648 49094 13676 49574
rect 13740 49366 13768 50798
rect 13728 49360 13780 49366
rect 13728 49302 13780 49308
rect 13726 49192 13782 49201
rect 13726 49127 13782 49136
rect 13636 49088 13688 49094
rect 13636 49030 13688 49036
rect 13542 48784 13598 48793
rect 13542 48719 13598 48728
rect 13544 48544 13596 48550
rect 13544 48486 13596 48492
rect 13556 47002 13584 48486
rect 13648 47161 13676 49030
rect 13634 47152 13690 47161
rect 13634 47087 13690 47096
rect 13556 46974 13676 47002
rect 13542 46880 13598 46889
rect 13542 46815 13598 46824
rect 13556 46481 13584 46815
rect 13542 46472 13598 46481
rect 13542 46407 13598 46416
rect 13648 46322 13676 46974
rect 13556 46294 13676 46322
rect 13556 45490 13584 46294
rect 13636 46164 13688 46170
rect 13636 46106 13688 46112
rect 13544 45484 13596 45490
rect 13544 45426 13596 45432
rect 13542 45384 13598 45393
rect 13542 45319 13598 45328
rect 13556 44946 13584 45319
rect 13544 44940 13596 44946
rect 13544 44882 13596 44888
rect 13556 44538 13584 44882
rect 13544 44532 13596 44538
rect 13544 44474 13596 44480
rect 13542 44432 13598 44441
rect 13542 44367 13598 44376
rect 13556 43858 13584 44367
rect 13544 43852 13596 43858
rect 13544 43794 13596 43800
rect 13556 43450 13584 43794
rect 13544 43444 13596 43450
rect 13544 43386 13596 43392
rect 13544 43104 13596 43110
rect 13544 43046 13596 43052
rect 13556 42770 13584 43046
rect 13544 42764 13596 42770
rect 13544 42706 13596 42712
rect 13556 42294 13584 42706
rect 13544 42288 13596 42294
rect 13544 42230 13596 42236
rect 13544 42152 13596 42158
rect 13544 42094 13596 42100
rect 13556 41478 13584 42094
rect 13544 41472 13596 41478
rect 13544 41414 13596 41420
rect 13648 40610 13676 46106
rect 13740 44334 13768 49127
rect 13832 46186 13860 52022
rect 13912 51944 13964 51950
rect 13912 51886 13964 51892
rect 13924 51610 13952 51886
rect 13912 51604 13964 51610
rect 13912 51546 13964 51552
rect 13924 50862 13952 51546
rect 13912 50856 13964 50862
rect 13912 50798 13964 50804
rect 14016 50289 14044 52090
rect 14002 50280 14058 50289
rect 14002 50215 14058 50224
rect 14004 50176 14056 50182
rect 14004 50118 14056 50124
rect 13912 49972 13964 49978
rect 13912 49914 13964 49920
rect 13924 49094 13952 49914
rect 13912 49088 13964 49094
rect 13912 49030 13964 49036
rect 13912 48000 13964 48006
rect 13912 47942 13964 47948
rect 13924 46374 13952 47942
rect 13912 46368 13964 46374
rect 13912 46310 13964 46316
rect 13832 46158 13952 46186
rect 13728 44328 13780 44334
rect 13728 44270 13780 44276
rect 13820 44260 13872 44266
rect 13820 44202 13872 44208
rect 13832 44146 13860 44202
rect 13740 44118 13860 44146
rect 13740 43314 13768 44118
rect 13818 44024 13874 44033
rect 13818 43959 13874 43968
rect 13832 43450 13860 43959
rect 13820 43444 13872 43450
rect 13820 43386 13872 43392
rect 13818 43344 13874 43353
rect 13728 43308 13780 43314
rect 13818 43279 13874 43288
rect 13728 43250 13780 43256
rect 13832 43246 13860 43279
rect 13820 43240 13872 43246
rect 13820 43182 13872 43188
rect 13832 42922 13860 43182
rect 13740 42894 13860 42922
rect 13740 41682 13768 42894
rect 13820 42764 13872 42770
rect 13820 42706 13872 42712
rect 13832 42158 13860 42706
rect 13820 42152 13872 42158
rect 13820 42094 13872 42100
rect 13832 41818 13860 42094
rect 13820 41812 13872 41818
rect 13820 41754 13872 41760
rect 13728 41676 13780 41682
rect 13728 41618 13780 41624
rect 13556 40582 13676 40610
rect 13740 41154 13768 41618
rect 13740 41138 13860 41154
rect 13740 41132 13872 41138
rect 13740 41126 13820 41132
rect 13556 39982 13584 40582
rect 13636 40520 13688 40526
rect 13636 40462 13688 40468
rect 13544 39976 13596 39982
rect 13544 39918 13596 39924
rect 13452 39500 13504 39506
rect 13452 39442 13504 39448
rect 13452 39296 13504 39302
rect 13452 39238 13504 39244
rect 13464 38758 13492 39238
rect 13556 38894 13584 39918
rect 13648 39098 13676 40462
rect 13636 39092 13688 39098
rect 13636 39034 13688 39040
rect 13636 38956 13688 38962
rect 13636 38898 13688 38904
rect 13544 38888 13596 38894
rect 13544 38830 13596 38836
rect 13452 38752 13504 38758
rect 13452 38694 13504 38700
rect 13358 38176 13414 38185
rect 13358 38111 13414 38120
rect 13464 36378 13492 38694
rect 13648 38418 13676 38898
rect 13740 38826 13768 41126
rect 13820 41074 13872 41080
rect 13818 40624 13874 40633
rect 13818 40559 13820 40568
rect 13872 40559 13874 40568
rect 13820 40530 13872 40536
rect 13820 40452 13872 40458
rect 13820 40394 13872 40400
rect 13728 38820 13780 38826
rect 13728 38762 13780 38768
rect 13726 38584 13782 38593
rect 13726 38519 13728 38528
rect 13780 38519 13782 38528
rect 13728 38490 13780 38496
rect 13636 38412 13688 38418
rect 13636 38354 13688 38360
rect 13544 38276 13596 38282
rect 13544 38218 13596 38224
rect 13452 36372 13504 36378
rect 13452 36314 13504 36320
rect 13556 35766 13584 38218
rect 13648 38010 13676 38354
rect 13728 38344 13780 38350
rect 13728 38286 13780 38292
rect 13636 38004 13688 38010
rect 13636 37946 13688 37952
rect 13648 36922 13676 37946
rect 13740 37670 13768 38286
rect 13728 37664 13780 37670
rect 13728 37606 13780 37612
rect 13636 36916 13688 36922
rect 13636 36858 13688 36864
rect 13544 35760 13596 35766
rect 13544 35702 13596 35708
rect 13740 35494 13768 37606
rect 13268 35488 13320 35494
rect 13268 35430 13320 35436
rect 13544 35488 13596 35494
rect 13544 35430 13596 35436
rect 13728 35488 13780 35494
rect 13728 35430 13780 35436
rect 13268 32292 13320 32298
rect 13268 32234 13320 32240
rect 13174 31784 13230 31793
rect 13174 31719 13230 31728
rect 12900 30320 12952 30326
rect 12900 30262 12952 30268
rect 13176 30184 13228 30190
rect 13176 30126 13228 30132
rect 13188 29646 13216 30126
rect 13280 29850 13308 32234
rect 13268 29844 13320 29850
rect 13268 29786 13320 29792
rect 13176 29640 13228 29646
rect 13176 29582 13228 29588
rect 13084 28756 13136 28762
rect 13084 28698 13136 28704
rect 12900 28008 12952 28014
rect 12900 27950 12952 27956
rect 12912 27674 12940 27950
rect 12992 27872 13044 27878
rect 12992 27814 13044 27820
rect 12900 27668 12952 27674
rect 12900 27610 12952 27616
rect 13004 26382 13032 27814
rect 12992 26376 13044 26382
rect 12992 26318 13044 26324
rect 12808 26036 12860 26042
rect 12808 25978 12860 25984
rect 12992 25832 13044 25838
rect 12992 25774 13044 25780
rect 12716 25696 12768 25702
rect 12716 25638 12768 25644
rect 12624 25424 12676 25430
rect 12624 25366 12676 25372
rect 12728 25362 12756 25638
rect 12716 25356 12768 25362
rect 12716 25298 12768 25304
rect 12900 25356 12952 25362
rect 12900 25298 12952 25304
rect 12624 24676 12676 24682
rect 12624 24618 12676 24624
rect 12636 23594 12664 24618
rect 12728 24614 12756 25298
rect 12912 24698 12940 25298
rect 13004 24886 13032 25774
rect 12992 24880 13044 24886
rect 12992 24822 13044 24828
rect 12912 24670 13032 24698
rect 13004 24614 13032 24670
rect 12716 24608 12768 24614
rect 12716 24550 12768 24556
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 12624 23588 12676 23594
rect 12624 23530 12676 23536
rect 12452 22222 12572 22250
rect 12348 21684 12400 21690
rect 12348 21626 12400 21632
rect 12452 21146 12480 22222
rect 12532 21684 12584 21690
rect 12532 21626 12584 21632
rect 12544 21593 12572 21626
rect 12530 21584 12586 21593
rect 12530 21519 12586 21528
rect 12532 21412 12584 21418
rect 12532 21354 12584 21360
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12440 20800 12492 20806
rect 12440 20742 12492 20748
rect 12452 20482 12480 20742
rect 12360 20466 12480 20482
rect 12348 20460 12480 20466
rect 12400 20454 12480 20460
rect 12348 20402 12400 20408
rect 12348 19440 12400 19446
rect 12348 19382 12400 19388
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12360 16114 12388 19382
rect 12452 18970 12480 20454
rect 12544 20398 12572 21354
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12636 20244 12664 23530
rect 12728 22982 12756 24550
rect 12900 24268 12952 24274
rect 12900 24210 12952 24216
rect 12808 24200 12860 24206
rect 12808 24142 12860 24148
rect 12716 22976 12768 22982
rect 12716 22918 12768 22924
rect 12728 22098 12756 22918
rect 12820 22522 12848 24142
rect 12912 23662 12940 24210
rect 12900 23656 12952 23662
rect 12898 23624 12900 23633
rect 12952 23624 12954 23633
rect 12898 23559 12954 23568
rect 12898 23216 12954 23225
rect 12898 23151 12900 23160
rect 12952 23151 12954 23160
rect 12900 23122 12952 23128
rect 12912 22642 12940 23122
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 12820 22494 12940 22522
rect 12716 22092 12768 22098
rect 12716 22034 12768 22040
rect 12728 21418 12756 22034
rect 12716 21412 12768 21418
rect 12716 21354 12768 21360
rect 12808 21344 12860 21350
rect 12808 21286 12860 21292
rect 12716 21140 12768 21146
rect 12716 21082 12768 21088
rect 12544 20216 12664 20244
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12452 17882 12480 18906
rect 12544 18834 12572 20216
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12636 19417 12664 19790
rect 12622 19408 12678 19417
rect 12622 19343 12678 19352
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12544 18358 12572 18770
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12532 18352 12584 18358
rect 12532 18294 12584 18300
rect 12544 18154 12572 18294
rect 12532 18148 12584 18154
rect 12532 18090 12584 18096
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12452 17270 12480 17818
rect 12440 17264 12492 17270
rect 12440 17206 12492 17212
rect 12440 17128 12492 17134
rect 12492 17076 12572 17082
rect 12440 17070 12572 17076
rect 12452 17054 12572 17070
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12452 16794 12480 16934
rect 12544 16794 12572 17054
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12348 16108 12400 16114
rect 12348 16050 12400 16056
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12164 14068 12216 14074
rect 12216 14028 12296 14056
rect 12164 14010 12216 14016
rect 12084 12974 12204 13002
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11348 11630 11480 11636
rect 11348 11614 11468 11630
rect 11624 11614 11744 11642
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11348 11082 11376 11614
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 10956 10908 11252 10928
rect 11012 10906 11036 10908
rect 11092 10906 11116 10908
rect 11172 10906 11196 10908
rect 11034 10854 11036 10906
rect 11098 10854 11110 10906
rect 11172 10854 11174 10906
rect 11012 10852 11036 10854
rect 11092 10852 11116 10854
rect 11172 10852 11196 10854
rect 10956 10832 11252 10852
rect 10704 10526 10824 10554
rect 10138 10296 10194 10305
rect 10138 10231 10194 10240
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 9770 9072 9826 9081
rect 9770 9007 9772 9016
rect 9824 9007 9826 9016
rect 9772 8978 9824 8984
rect 9784 8634 9812 8978
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9678 7304 9734 7313
rect 9678 7239 9734 7248
rect 9692 6798 9720 7239
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9680 5772 9732 5778
rect 9600 5732 9680 5760
rect 9680 5714 9732 5720
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 9692 5370 9720 5714
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9876 5030 9904 5714
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9876 4729 9904 4966
rect 10060 4729 10088 9318
rect 10598 8936 10654 8945
rect 10598 8871 10654 8880
rect 10506 8528 10562 8537
rect 10612 8498 10640 8871
rect 10506 8463 10562 8472
rect 10600 8492 10652 8498
rect 10520 8430 10548 8463
rect 10600 8434 10652 8440
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10138 7984 10194 7993
rect 10138 7919 10194 7928
rect 10152 6866 10180 7919
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10336 7410 10364 7686
rect 10704 7546 10732 10526
rect 10782 10432 10838 10441
rect 10782 10367 10838 10376
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10152 6458 10180 6802
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10244 6458 10272 6734
rect 10796 6458 10824 10367
rect 11348 10266 11376 11018
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10888 8401 10916 9862
rect 10956 9820 11252 9840
rect 11012 9818 11036 9820
rect 11092 9818 11116 9820
rect 11172 9818 11196 9820
rect 11034 9766 11036 9818
rect 11098 9766 11110 9818
rect 11172 9766 11174 9818
rect 11012 9764 11036 9766
rect 11092 9764 11116 9766
rect 11172 9764 11196 9766
rect 10956 9744 11252 9764
rect 11440 9722 11468 11086
rect 11624 10713 11652 11614
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11610 10704 11666 10713
rect 11610 10639 11666 10648
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11336 9648 11388 9654
rect 11150 9616 11206 9625
rect 11336 9590 11388 9596
rect 11150 9551 11206 9560
rect 11164 9110 11192 9551
rect 11348 9382 11376 9590
rect 11532 9518 11560 10202
rect 11428 9512 11480 9518
rect 11428 9454 11480 9460
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 10956 8732 11252 8752
rect 11012 8730 11036 8732
rect 11092 8730 11116 8732
rect 11172 8730 11196 8732
rect 11034 8678 11036 8730
rect 11098 8678 11110 8730
rect 11172 8678 11174 8730
rect 11012 8676 11036 8678
rect 11092 8676 11116 8678
rect 11172 8676 11196 8678
rect 10956 8656 11252 8676
rect 11348 8634 11376 9318
rect 11440 9178 11468 9454
rect 11518 9344 11574 9353
rect 11518 9279 11574 9288
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 10874 8392 10930 8401
rect 10874 8327 10930 8336
rect 11336 8016 11388 8022
rect 11336 7958 11388 7964
rect 10956 7644 11252 7664
rect 11012 7642 11036 7644
rect 11092 7642 11116 7644
rect 11172 7642 11196 7644
rect 11034 7590 11036 7642
rect 11098 7590 11110 7642
rect 11172 7590 11174 7642
rect 11012 7588 11036 7590
rect 11092 7588 11116 7590
rect 11172 7588 11196 7590
rect 10956 7568 11252 7588
rect 11348 7342 11376 7958
rect 11440 7342 11468 9114
rect 11532 8634 11560 9279
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11624 8498 11652 10542
rect 11716 9353 11744 11494
rect 11808 11286 11836 11630
rect 11900 11626 11928 12242
rect 11888 11620 11940 11626
rect 11888 11562 11940 11568
rect 11900 11286 11928 11562
rect 11796 11280 11848 11286
rect 11796 11222 11848 11228
rect 11888 11280 11940 11286
rect 11888 11222 11940 11228
rect 11900 10810 11928 11222
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11794 10704 11850 10713
rect 11794 10639 11850 10648
rect 11702 9344 11758 9353
rect 11702 9279 11758 9288
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11624 8106 11652 8434
rect 11624 8078 11744 8106
rect 11610 7984 11666 7993
rect 11610 7919 11666 7928
rect 11520 7472 11572 7478
rect 11520 7414 11572 7420
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 10956 6556 11252 6576
rect 11012 6554 11036 6556
rect 11092 6554 11116 6556
rect 11172 6554 11196 6556
rect 11034 6502 11036 6554
rect 11098 6502 11110 6554
rect 11172 6502 11174 6554
rect 11012 6500 11036 6502
rect 11092 6500 11116 6502
rect 11172 6500 11196 6502
rect 10956 6480 11252 6500
rect 11532 6458 11560 7414
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11624 6322 11652 7919
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11716 6254 11744 8078
rect 11808 8022 11836 10639
rect 11888 9920 11940 9926
rect 11992 9908 12020 11154
rect 12084 11150 12112 12854
rect 12072 11144 12124 11150
rect 12072 11086 12124 11092
rect 11940 9880 12020 9908
rect 11888 9862 11940 9868
rect 11796 8016 11848 8022
rect 11796 7958 11848 7964
rect 11900 7857 11928 9862
rect 11980 9716 12032 9722
rect 11980 9658 12032 9664
rect 11992 8537 12020 9658
rect 11978 8528 12034 8537
rect 11978 8463 12034 8472
rect 11992 7954 12020 8463
rect 12084 8430 12112 11086
rect 12176 10130 12204 12974
rect 12268 12918 12296 14028
rect 12360 13841 12388 14962
rect 12452 14618 12480 16730
rect 12544 16153 12572 16730
rect 12530 16144 12586 16153
rect 12530 16079 12586 16088
rect 12544 15706 12572 16079
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12636 15586 12664 18566
rect 12544 15558 12664 15586
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 12346 13832 12402 13841
rect 12346 13767 12402 13776
rect 12452 13682 12480 13942
rect 12360 13654 12480 13682
rect 12256 12912 12308 12918
rect 12256 12854 12308 12860
rect 12256 12368 12308 12374
rect 12254 12336 12256 12345
rect 12308 12336 12310 12345
rect 12254 12271 12310 12280
rect 12254 11656 12310 11665
rect 12254 11591 12310 11600
rect 12268 11354 12296 11591
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12254 10568 12310 10577
rect 12254 10503 12310 10512
rect 12268 10266 12296 10503
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12360 9518 12388 13654
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12452 9654 12480 10746
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12360 9110 12388 9454
rect 12438 9344 12494 9353
rect 12438 9279 12494 9288
rect 12348 9104 12400 9110
rect 12348 9046 12400 9052
rect 12360 8430 12388 9046
rect 12452 8634 12480 9279
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12084 8090 12112 8366
rect 12452 8242 12480 8570
rect 12268 8214 12480 8242
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11886 7848 11942 7857
rect 11886 7783 11942 7792
rect 11796 7268 11848 7274
rect 11796 7210 11848 7216
rect 11704 6248 11756 6254
rect 11808 6225 11836 7210
rect 11992 6730 12020 7890
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 11980 6724 12032 6730
rect 11980 6666 12032 6672
rect 11704 6190 11756 6196
rect 11794 6216 11850 6225
rect 11716 5914 11744 6190
rect 11794 6151 11850 6160
rect 12176 5914 12204 6802
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 12164 5908 12216 5914
rect 12164 5850 12216 5856
rect 11428 5704 11480 5710
rect 11426 5672 11428 5681
rect 11480 5672 11482 5681
rect 11426 5607 11482 5616
rect 10956 5468 11252 5488
rect 11012 5466 11036 5468
rect 11092 5466 11116 5468
rect 11172 5466 11196 5468
rect 11034 5414 11036 5466
rect 11098 5414 11110 5466
rect 11172 5414 11174 5466
rect 11012 5412 11036 5414
rect 11092 5412 11116 5414
rect 11172 5412 11196 5414
rect 10956 5392 11252 5412
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 9862 4720 9918 4729
rect 9862 4655 9918 4664
rect 10046 4720 10102 4729
rect 10046 4655 10102 4664
rect 10244 4146 10272 5306
rect 10956 4380 11252 4400
rect 11012 4378 11036 4380
rect 11092 4378 11116 4380
rect 11172 4378 11196 4380
rect 11034 4326 11036 4378
rect 11098 4326 11110 4378
rect 11172 4326 11174 4378
rect 11012 4324 11036 4326
rect 11092 4324 11116 4326
rect 11172 4324 11196 4326
rect 10956 4304 11252 4324
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9508 2310 9536 2450
rect 9784 2446 9812 2586
rect 10060 2553 10088 3878
rect 10244 3738 10272 4082
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10244 2666 10272 3674
rect 10956 3292 11252 3312
rect 11012 3290 11036 3292
rect 11092 3290 11116 3292
rect 11172 3290 11196 3292
rect 11034 3238 11036 3290
rect 11098 3238 11110 3290
rect 11172 3238 11174 3290
rect 11012 3236 11036 3238
rect 11092 3236 11116 3238
rect 11172 3236 11196 3238
rect 10956 3216 11252 3236
rect 10152 2650 10272 2666
rect 10140 2644 10272 2650
rect 10192 2638 10272 2644
rect 10140 2586 10192 2592
rect 10046 2544 10102 2553
rect 10046 2479 10102 2488
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 12268 2310 12296 8214
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12452 5302 12480 7822
rect 12544 5778 12572 15558
rect 12728 14550 12756 21082
rect 12820 19854 12848 21286
rect 12808 19848 12860 19854
rect 12808 19790 12860 19796
rect 12820 19446 12848 19790
rect 12808 19440 12860 19446
rect 12808 19382 12860 19388
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12820 16250 12848 17138
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12820 16046 12848 16186
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 12912 15570 12940 22494
rect 13004 20398 13032 24550
rect 13096 22778 13124 28698
rect 13188 28694 13216 29582
rect 13176 28688 13228 28694
rect 13176 28630 13228 28636
rect 13280 28098 13308 29786
rect 13188 28070 13308 28098
rect 13360 28076 13412 28082
rect 13188 24274 13216 28070
rect 13360 28018 13412 28024
rect 13268 28008 13320 28014
rect 13268 27950 13320 27956
rect 13280 27606 13308 27950
rect 13268 27600 13320 27606
rect 13268 27542 13320 27548
rect 13280 26994 13308 27542
rect 13372 27334 13400 28018
rect 13360 27328 13412 27334
rect 13556 27282 13584 35430
rect 13636 35148 13688 35154
rect 13636 35090 13688 35096
rect 13648 34542 13676 35090
rect 13636 34536 13688 34542
rect 13636 34478 13688 34484
rect 13648 33969 13676 34478
rect 13634 33960 13690 33969
rect 13634 33895 13690 33904
rect 13636 32972 13688 32978
rect 13636 32914 13688 32920
rect 13648 32230 13676 32914
rect 13636 32224 13688 32230
rect 13636 32166 13688 32172
rect 13740 31890 13768 35430
rect 13728 31884 13780 31890
rect 13728 31826 13780 31832
rect 13832 31249 13860 40394
rect 13924 32842 13952 46158
rect 14016 45370 14044 50118
rect 14108 50017 14136 52362
rect 14094 50008 14150 50017
rect 14094 49943 14150 49952
rect 14096 49836 14148 49842
rect 14096 49778 14148 49784
rect 14108 49434 14136 49778
rect 14096 49428 14148 49434
rect 14096 49370 14148 49376
rect 14096 49292 14148 49298
rect 14096 49234 14148 49240
rect 14108 48550 14136 49234
rect 14200 48929 14228 52838
rect 14289 52796 14585 52816
rect 14345 52794 14369 52796
rect 14425 52794 14449 52796
rect 14505 52794 14529 52796
rect 14367 52742 14369 52794
rect 14431 52742 14443 52794
rect 14505 52742 14507 52794
rect 14345 52740 14369 52742
rect 14425 52740 14449 52742
rect 14505 52740 14529 52742
rect 14289 52720 14585 52740
rect 14660 52562 14688 53110
rect 14752 53106 14780 53615
rect 14740 53100 14792 53106
rect 14740 53042 14792 53048
rect 14648 52556 14700 52562
rect 14648 52498 14700 52504
rect 14280 52352 14332 52358
rect 14280 52294 14332 52300
rect 14740 52352 14792 52358
rect 14740 52294 14792 52300
rect 14292 51950 14320 52294
rect 14648 52012 14700 52018
rect 14648 51954 14700 51960
rect 14280 51944 14332 51950
rect 14280 51886 14332 51892
rect 14289 51708 14585 51728
rect 14345 51706 14369 51708
rect 14425 51706 14449 51708
rect 14505 51706 14529 51708
rect 14367 51654 14369 51706
rect 14431 51654 14443 51706
rect 14505 51654 14507 51706
rect 14345 51652 14369 51654
rect 14425 51652 14449 51654
rect 14505 51652 14529 51654
rect 14289 51632 14585 51652
rect 14289 50620 14585 50640
rect 14345 50618 14369 50620
rect 14425 50618 14449 50620
rect 14505 50618 14529 50620
rect 14367 50566 14369 50618
rect 14431 50566 14443 50618
rect 14505 50566 14507 50618
rect 14345 50564 14369 50566
rect 14425 50564 14449 50566
rect 14505 50564 14529 50566
rect 14289 50544 14585 50564
rect 14289 49532 14585 49552
rect 14345 49530 14369 49532
rect 14425 49530 14449 49532
rect 14505 49530 14529 49532
rect 14367 49478 14369 49530
rect 14431 49478 14443 49530
rect 14505 49478 14507 49530
rect 14345 49476 14369 49478
rect 14425 49476 14449 49478
rect 14505 49476 14529 49478
rect 14289 49456 14585 49476
rect 14280 49224 14332 49230
rect 14280 49166 14332 49172
rect 14186 48920 14242 48929
rect 14186 48855 14242 48864
rect 14292 48804 14320 49166
rect 14556 49088 14608 49094
rect 14556 49030 14608 49036
rect 14200 48776 14320 48804
rect 14096 48544 14148 48550
rect 14096 48486 14148 48492
rect 14108 48346 14136 48486
rect 14096 48340 14148 48346
rect 14096 48282 14148 48288
rect 14094 47288 14150 47297
rect 14094 47223 14096 47232
rect 14148 47223 14150 47232
rect 14096 47194 14148 47200
rect 14016 45342 14136 45370
rect 14004 45280 14056 45286
rect 14004 45222 14056 45228
rect 14016 42362 14044 45222
rect 14108 44470 14136 45342
rect 14096 44464 14148 44470
rect 14096 44406 14148 44412
rect 14096 44328 14148 44334
rect 14096 44270 14148 44276
rect 14004 42356 14056 42362
rect 14004 42298 14056 42304
rect 14004 41472 14056 41478
rect 14002 41440 14004 41449
rect 14056 41440 14058 41449
rect 14002 41375 14058 41384
rect 14004 41200 14056 41206
rect 14004 41142 14056 41148
rect 14016 36904 14044 41142
rect 14108 39420 14136 44270
rect 14200 43926 14228 48776
rect 14568 48618 14596 49030
rect 14556 48612 14608 48618
rect 14556 48554 14608 48560
rect 14289 48444 14585 48464
rect 14345 48442 14369 48444
rect 14425 48442 14449 48444
rect 14505 48442 14529 48444
rect 14367 48390 14369 48442
rect 14431 48390 14443 48442
rect 14505 48390 14507 48442
rect 14345 48388 14369 48390
rect 14425 48388 14449 48390
rect 14505 48388 14529 48390
rect 14289 48368 14585 48388
rect 14289 47356 14585 47376
rect 14345 47354 14369 47356
rect 14425 47354 14449 47356
rect 14505 47354 14529 47356
rect 14367 47302 14369 47354
rect 14431 47302 14443 47354
rect 14505 47302 14507 47354
rect 14345 47300 14369 47302
rect 14425 47300 14449 47302
rect 14505 47300 14529 47302
rect 14289 47280 14585 47300
rect 14289 46268 14585 46288
rect 14345 46266 14369 46268
rect 14425 46266 14449 46268
rect 14505 46266 14529 46268
rect 14367 46214 14369 46266
rect 14431 46214 14443 46266
rect 14505 46214 14507 46266
rect 14345 46212 14369 46214
rect 14425 46212 14449 46214
rect 14505 46212 14529 46214
rect 14289 46192 14585 46212
rect 14556 46096 14608 46102
rect 14556 46038 14608 46044
rect 14568 45268 14596 46038
rect 14660 46034 14688 51954
rect 14752 49366 14780 52294
rect 14844 50969 14872 57967
rect 14922 56808 14978 56817
rect 14922 56743 14978 56752
rect 14830 50960 14886 50969
rect 14830 50895 14886 50904
rect 14832 50720 14884 50726
rect 14832 50662 14884 50668
rect 14844 50454 14872 50662
rect 14832 50448 14884 50454
rect 14832 50390 14884 50396
rect 14844 49978 14872 50390
rect 14832 49972 14884 49978
rect 14832 49914 14884 49920
rect 14832 49700 14884 49706
rect 14832 49642 14884 49648
rect 14740 49360 14792 49366
rect 14740 49302 14792 49308
rect 14752 48890 14780 49302
rect 14844 49201 14872 49642
rect 14830 49192 14886 49201
rect 14830 49127 14886 49136
rect 14844 48890 14872 49127
rect 14740 48884 14792 48890
rect 14740 48826 14792 48832
rect 14832 48884 14884 48890
rect 14832 48826 14884 48832
rect 14832 48748 14884 48754
rect 14832 48690 14884 48696
rect 14740 48544 14792 48550
rect 14740 48486 14792 48492
rect 14752 46986 14780 48486
rect 14740 46980 14792 46986
rect 14740 46922 14792 46928
rect 14648 46028 14700 46034
rect 14648 45970 14700 45976
rect 14660 45422 14688 45970
rect 14648 45416 14700 45422
rect 14648 45358 14700 45364
rect 14568 45240 14688 45268
rect 14289 45180 14585 45200
rect 14345 45178 14369 45180
rect 14425 45178 14449 45180
rect 14505 45178 14529 45180
rect 14367 45126 14369 45178
rect 14431 45126 14443 45178
rect 14505 45126 14507 45178
rect 14345 45124 14369 45126
rect 14425 45124 14449 45126
rect 14505 45124 14529 45126
rect 14289 45104 14585 45124
rect 14556 44736 14608 44742
rect 14554 44704 14556 44713
rect 14608 44704 14610 44713
rect 14554 44639 14610 44648
rect 14289 44092 14585 44112
rect 14345 44090 14369 44092
rect 14425 44090 14449 44092
rect 14505 44090 14529 44092
rect 14367 44038 14369 44090
rect 14431 44038 14443 44090
rect 14505 44038 14507 44090
rect 14345 44036 14369 44038
rect 14425 44036 14449 44038
rect 14505 44036 14529 44038
rect 14289 44016 14585 44036
rect 14188 43920 14240 43926
rect 14188 43862 14240 43868
rect 14372 43920 14424 43926
rect 14372 43862 14424 43868
rect 14280 43852 14332 43858
rect 14280 43794 14332 43800
rect 14292 43382 14320 43794
rect 14280 43376 14332 43382
rect 14280 43318 14332 43324
rect 14188 43308 14240 43314
rect 14188 43250 14240 43256
rect 14200 42702 14228 43250
rect 14384 43178 14412 43862
rect 14372 43172 14424 43178
rect 14372 43114 14424 43120
rect 14289 43004 14585 43024
rect 14345 43002 14369 43004
rect 14425 43002 14449 43004
rect 14505 43002 14529 43004
rect 14367 42950 14369 43002
rect 14431 42950 14443 43002
rect 14505 42950 14507 43002
rect 14345 42948 14369 42950
rect 14425 42948 14449 42950
rect 14505 42948 14529 42950
rect 14289 42928 14585 42948
rect 14188 42696 14240 42702
rect 14188 42638 14240 42644
rect 14188 42356 14240 42362
rect 14188 42298 14240 42304
rect 14200 39574 14228 42298
rect 14289 41916 14585 41936
rect 14345 41914 14369 41916
rect 14425 41914 14449 41916
rect 14505 41914 14529 41916
rect 14367 41862 14369 41914
rect 14431 41862 14443 41914
rect 14505 41862 14507 41914
rect 14345 41860 14369 41862
rect 14425 41860 14449 41862
rect 14505 41860 14529 41862
rect 14289 41840 14585 41860
rect 14556 41132 14608 41138
rect 14556 41074 14608 41080
rect 14568 41041 14596 41074
rect 14554 41032 14610 41041
rect 14554 40967 14610 40976
rect 14289 40828 14585 40848
rect 14345 40826 14369 40828
rect 14425 40826 14449 40828
rect 14505 40826 14529 40828
rect 14367 40774 14369 40826
rect 14431 40774 14443 40826
rect 14505 40774 14507 40826
rect 14345 40772 14369 40774
rect 14425 40772 14449 40774
rect 14505 40772 14529 40774
rect 14289 40752 14585 40772
rect 14660 40594 14688 45240
rect 14752 44826 14780 46922
rect 14844 45665 14872 48690
rect 14830 45656 14886 45665
rect 14830 45591 14886 45600
rect 14832 45280 14884 45286
rect 14832 45222 14884 45228
rect 14844 45014 14872 45222
rect 14832 45008 14884 45014
rect 14832 44950 14884 44956
rect 14752 44798 14872 44826
rect 14740 44192 14792 44198
rect 14740 44134 14792 44140
rect 14752 41750 14780 44134
rect 14844 43654 14872 44798
rect 14936 44538 14964 56743
rect 15028 55049 15056 60454
rect 15014 55040 15070 55049
rect 15014 54975 15070 54984
rect 15108 53984 15160 53990
rect 15108 53926 15160 53932
rect 15120 53514 15148 53926
rect 15108 53508 15160 53514
rect 15108 53450 15160 53456
rect 15016 52964 15068 52970
rect 15016 52906 15068 52912
rect 15028 52562 15056 52906
rect 15016 52556 15068 52562
rect 15016 52498 15068 52504
rect 15108 52556 15160 52562
rect 15108 52498 15160 52504
rect 15028 51610 15056 52498
rect 15120 52154 15148 52498
rect 15108 52148 15160 52154
rect 15108 52090 15160 52096
rect 15016 51604 15068 51610
rect 15068 51564 15148 51592
rect 15016 51546 15068 51552
rect 15120 50930 15148 51564
rect 15016 50924 15068 50930
rect 15016 50866 15068 50872
rect 15108 50924 15160 50930
rect 15108 50866 15160 50872
rect 15028 49745 15056 50866
rect 15106 50280 15162 50289
rect 15106 50215 15162 50224
rect 15120 49774 15148 50215
rect 15108 49768 15160 49774
rect 15014 49736 15070 49745
rect 15108 49710 15160 49716
rect 15014 49671 15070 49680
rect 15016 49632 15068 49638
rect 15016 49574 15068 49580
rect 15028 49366 15056 49574
rect 15016 49360 15068 49366
rect 15016 49302 15068 49308
rect 15016 49224 15068 49230
rect 15016 49166 15068 49172
rect 14924 44532 14976 44538
rect 14924 44474 14976 44480
rect 14924 44396 14976 44402
rect 14924 44338 14976 44344
rect 14832 43648 14884 43654
rect 14832 43590 14884 43596
rect 14832 43172 14884 43178
rect 14832 43114 14884 43120
rect 14844 42566 14872 43114
rect 14936 43110 14964 44338
rect 15028 43897 15056 49166
rect 15120 46102 15148 49710
rect 15108 46096 15160 46102
rect 15108 46038 15160 46044
rect 15106 45928 15162 45937
rect 15106 45863 15162 45872
rect 15014 43888 15070 43897
rect 15014 43823 15070 43832
rect 15016 43648 15068 43654
rect 15016 43590 15068 43596
rect 14924 43104 14976 43110
rect 14924 43046 14976 43052
rect 14924 42628 14976 42634
rect 14924 42570 14976 42576
rect 14832 42560 14884 42566
rect 14832 42502 14884 42508
rect 14832 42356 14884 42362
rect 14832 42298 14884 42304
rect 14740 41744 14792 41750
rect 14740 41686 14792 41692
rect 14752 41070 14780 41686
rect 14740 41064 14792 41070
rect 14740 41006 14792 41012
rect 14648 40588 14700 40594
rect 14648 40530 14700 40536
rect 14648 40452 14700 40458
rect 14648 40394 14700 40400
rect 14289 39740 14585 39760
rect 14345 39738 14369 39740
rect 14425 39738 14449 39740
rect 14505 39738 14529 39740
rect 14367 39686 14369 39738
rect 14431 39686 14443 39738
rect 14505 39686 14507 39738
rect 14345 39684 14369 39686
rect 14425 39684 14449 39686
rect 14505 39684 14529 39686
rect 14289 39664 14585 39684
rect 14660 39642 14688 40394
rect 14648 39636 14700 39642
rect 14648 39578 14700 39584
rect 14188 39568 14240 39574
rect 14188 39510 14240 39516
rect 14372 39568 14424 39574
rect 14372 39510 14424 39516
rect 14646 39536 14702 39545
rect 14108 39392 14228 39420
rect 14096 37664 14148 37670
rect 14096 37606 14148 37612
rect 14108 37330 14136 37606
rect 14096 37324 14148 37330
rect 14096 37266 14148 37272
rect 14200 37126 14228 39392
rect 14384 39098 14412 39510
rect 14646 39471 14702 39480
rect 14372 39092 14424 39098
rect 14372 39034 14424 39040
rect 14289 38652 14585 38672
rect 14345 38650 14369 38652
rect 14425 38650 14449 38652
rect 14505 38650 14529 38652
rect 14367 38598 14369 38650
rect 14431 38598 14443 38650
rect 14505 38598 14507 38650
rect 14345 38596 14369 38598
rect 14425 38596 14449 38598
rect 14505 38596 14529 38598
rect 14289 38576 14585 38596
rect 14660 38321 14688 39471
rect 14752 38418 14780 41006
rect 14844 40934 14872 42298
rect 14936 41313 14964 42570
rect 14922 41304 14978 41313
rect 14922 41239 14978 41248
rect 15028 41154 15056 43590
rect 15120 43353 15148 45863
rect 15106 43344 15162 43353
rect 15106 43279 15162 43288
rect 15106 43208 15162 43217
rect 15106 43143 15162 43152
rect 15120 42906 15148 43143
rect 15108 42900 15160 42906
rect 15108 42842 15160 42848
rect 15108 42084 15160 42090
rect 15108 42026 15160 42032
rect 14936 41126 15056 41154
rect 14832 40928 14884 40934
rect 14832 40870 14884 40876
rect 14936 40746 14964 41126
rect 15016 40928 15068 40934
rect 15016 40870 15068 40876
rect 14844 40718 14964 40746
rect 14740 38412 14792 38418
rect 14740 38354 14792 38360
rect 14646 38312 14702 38321
rect 14646 38247 14702 38256
rect 14648 38208 14700 38214
rect 14648 38150 14700 38156
rect 14289 37564 14585 37584
rect 14345 37562 14369 37564
rect 14425 37562 14449 37564
rect 14505 37562 14529 37564
rect 14367 37510 14369 37562
rect 14431 37510 14443 37562
rect 14505 37510 14507 37562
rect 14345 37508 14369 37510
rect 14425 37508 14449 37510
rect 14505 37508 14529 37510
rect 14289 37488 14585 37508
rect 14556 37324 14608 37330
rect 14556 37266 14608 37272
rect 14188 37120 14240 37126
rect 14188 37062 14240 37068
rect 14568 36922 14596 37266
rect 14660 37262 14688 38150
rect 14752 37738 14780 38354
rect 14740 37732 14792 37738
rect 14740 37674 14792 37680
rect 14648 37256 14700 37262
rect 14648 37198 14700 37204
rect 14556 36916 14608 36922
rect 14016 36876 14228 36904
rect 14004 36780 14056 36786
rect 14004 36722 14056 36728
rect 13912 32836 13964 32842
rect 13912 32778 13964 32784
rect 13818 31240 13874 31249
rect 13818 31175 13874 31184
rect 13636 29504 13688 29510
rect 13636 29446 13688 29452
rect 13648 29102 13676 29446
rect 13636 29096 13688 29102
rect 13636 29038 13688 29044
rect 13912 28756 13964 28762
rect 13912 28698 13964 28704
rect 13924 28014 13952 28698
rect 13912 28008 13964 28014
rect 13912 27950 13964 27956
rect 13820 27872 13872 27878
rect 13820 27814 13872 27820
rect 13832 27538 13860 27814
rect 13820 27532 13872 27538
rect 13820 27474 13872 27480
rect 13360 27270 13412 27276
rect 13268 26988 13320 26994
rect 13268 26930 13320 26936
rect 13268 26784 13320 26790
rect 13268 26726 13320 26732
rect 13280 25362 13308 26726
rect 13372 26450 13400 27270
rect 13464 27254 13584 27282
rect 13360 26444 13412 26450
rect 13360 26386 13412 26392
rect 13372 25838 13400 26386
rect 13360 25832 13412 25838
rect 13360 25774 13412 25780
rect 13268 25356 13320 25362
rect 13268 25298 13320 25304
rect 13280 24682 13308 25298
rect 13372 25294 13400 25774
rect 13360 25288 13412 25294
rect 13464 25276 13492 27254
rect 13544 27124 13596 27130
rect 13544 27066 13596 27072
rect 13556 27033 13584 27066
rect 13542 27024 13598 27033
rect 13542 26959 13598 26968
rect 13832 26790 13860 27474
rect 13912 27328 13964 27334
rect 13912 27270 13964 27276
rect 13924 26926 13952 27270
rect 13912 26920 13964 26926
rect 13912 26862 13964 26868
rect 13820 26784 13872 26790
rect 13648 26732 13820 26738
rect 13648 26726 13872 26732
rect 13648 26710 13860 26726
rect 13648 25498 13676 26710
rect 13728 26308 13780 26314
rect 13728 26250 13780 26256
rect 13740 26194 13768 26250
rect 13740 26166 13860 26194
rect 13832 25838 13860 26166
rect 13820 25832 13872 25838
rect 13740 25780 13820 25786
rect 13740 25774 13872 25780
rect 13740 25758 13860 25774
rect 13636 25492 13688 25498
rect 13636 25434 13688 25440
rect 13464 25248 13676 25276
rect 13360 25230 13412 25236
rect 13268 24676 13320 24682
rect 13268 24618 13320 24624
rect 13176 24268 13228 24274
rect 13176 24210 13228 24216
rect 13268 23112 13320 23118
rect 13266 23080 13268 23089
rect 13320 23080 13322 23089
rect 13266 23015 13322 23024
rect 13372 22930 13400 25230
rect 13544 25152 13596 25158
rect 13544 25094 13596 25100
rect 13450 24984 13506 24993
rect 13450 24919 13506 24928
rect 13464 24342 13492 24919
rect 13452 24336 13504 24342
rect 13452 24278 13504 24284
rect 13280 22902 13400 22930
rect 13084 22772 13136 22778
rect 13084 22714 13136 22720
rect 13096 22574 13124 22714
rect 13084 22568 13136 22574
rect 13084 22510 13136 22516
rect 13176 21412 13228 21418
rect 13176 21354 13228 21360
rect 13188 21146 13216 21354
rect 13176 21140 13228 21146
rect 13176 21082 13228 21088
rect 13176 20800 13228 20806
rect 13176 20742 13228 20748
rect 12992 20392 13044 20398
rect 12992 20334 13044 20340
rect 13084 20324 13136 20330
rect 13084 20266 13136 20272
rect 12992 19780 13044 19786
rect 12992 19722 13044 19728
rect 13004 18630 13032 19722
rect 13096 19378 13124 20266
rect 13188 19446 13216 20742
rect 13176 19440 13228 19446
rect 13176 19382 13228 19388
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 13096 18970 13124 19314
rect 13176 19304 13228 19310
rect 13176 19246 13228 19252
rect 13084 18964 13136 18970
rect 13084 18906 13136 18912
rect 13188 18698 13216 19246
rect 13176 18692 13228 18698
rect 13176 18634 13228 18640
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12912 15162 12940 15506
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 12716 14544 12768 14550
rect 12716 14486 12768 14492
rect 12728 14006 12756 14486
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 12728 13870 12756 13942
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12624 13796 12676 13802
rect 12624 13738 12676 13744
rect 12636 13530 12664 13738
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12728 13326 12756 13670
rect 12912 13462 12940 14214
rect 12900 13456 12952 13462
rect 12900 13398 12952 13404
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 12636 12646 12664 13194
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12636 9042 12664 12582
rect 12728 12442 12756 13262
rect 12820 12850 12848 13330
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12728 11558 12756 12038
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12728 10266 12756 11086
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12636 8362 12664 8978
rect 12624 8356 12676 8362
rect 12624 8298 12676 8304
rect 12728 7886 12756 9862
rect 12820 8022 12848 12786
rect 12912 12782 12940 13398
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 13004 10441 13032 18566
rect 13280 13988 13308 22902
rect 13360 22568 13412 22574
rect 13360 22510 13412 22516
rect 13452 22568 13504 22574
rect 13452 22510 13504 22516
rect 13372 21010 13400 22510
rect 13464 21894 13492 22510
rect 13452 21888 13504 21894
rect 13452 21830 13504 21836
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13372 20602 13400 20946
rect 13360 20596 13412 20602
rect 13360 20538 13412 20544
rect 13360 19236 13412 19242
rect 13360 19178 13412 19184
rect 13372 17746 13400 19178
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 13372 17270 13400 17682
rect 13464 17542 13492 21830
rect 13556 19310 13584 25094
rect 13648 23662 13676 25248
rect 13636 23656 13688 23662
rect 13636 23598 13688 23604
rect 13648 23322 13676 23598
rect 13636 23316 13688 23322
rect 13636 23258 13688 23264
rect 13636 22704 13688 22710
rect 13636 22646 13688 22652
rect 13648 22545 13676 22646
rect 13634 22536 13690 22545
rect 13634 22471 13690 22480
rect 13740 22386 13768 25758
rect 13924 24818 13952 26862
rect 14016 24857 14044 36722
rect 14096 36712 14148 36718
rect 14096 36654 14148 36660
rect 14108 36378 14136 36654
rect 14096 36372 14148 36378
rect 14096 36314 14148 36320
rect 14200 35850 14228 36876
rect 14556 36858 14608 36864
rect 14289 36476 14585 36496
rect 14345 36474 14369 36476
rect 14425 36474 14449 36476
rect 14505 36474 14529 36476
rect 14367 36422 14369 36474
rect 14431 36422 14443 36474
rect 14505 36422 14507 36474
rect 14345 36420 14369 36422
rect 14425 36420 14449 36422
rect 14505 36420 14529 36422
rect 14289 36400 14585 36420
rect 14660 36378 14688 37198
rect 14648 36372 14700 36378
rect 14648 36314 14700 36320
rect 14556 36304 14608 36310
rect 14556 36246 14608 36252
rect 14280 36168 14332 36174
rect 14280 36110 14332 36116
rect 14108 35822 14228 35850
rect 14292 35834 14320 36110
rect 14280 35828 14332 35834
rect 14108 34513 14136 35822
rect 14280 35770 14332 35776
rect 14188 35624 14240 35630
rect 14188 35566 14240 35572
rect 14200 35290 14228 35566
rect 14568 35562 14596 36246
rect 14752 36242 14780 37674
rect 14740 36236 14792 36242
rect 14740 36178 14792 36184
rect 14556 35556 14608 35562
rect 14556 35498 14608 35504
rect 14752 35494 14780 36178
rect 14740 35488 14792 35494
rect 14740 35430 14792 35436
rect 14289 35388 14585 35408
rect 14345 35386 14369 35388
rect 14425 35386 14449 35388
rect 14505 35386 14529 35388
rect 14367 35334 14369 35386
rect 14431 35334 14443 35386
rect 14505 35334 14507 35386
rect 14345 35332 14369 35334
rect 14425 35332 14449 35334
rect 14505 35332 14529 35334
rect 14289 35312 14585 35332
rect 14188 35284 14240 35290
rect 14752 35272 14780 35430
rect 14188 35226 14240 35232
rect 14660 35244 14780 35272
rect 14660 35018 14688 35244
rect 14740 35148 14792 35154
rect 14740 35090 14792 35096
rect 14648 35012 14700 35018
rect 14648 34954 14700 34960
rect 14752 34746 14780 35090
rect 14740 34740 14792 34746
rect 14740 34682 14792 34688
rect 14648 34604 14700 34610
rect 14648 34546 14700 34552
rect 14094 34504 14150 34513
rect 14094 34439 14150 34448
rect 14289 34300 14585 34320
rect 14345 34298 14369 34300
rect 14425 34298 14449 34300
rect 14505 34298 14529 34300
rect 14367 34246 14369 34298
rect 14431 34246 14443 34298
rect 14505 34246 14507 34298
rect 14345 34244 14369 34246
rect 14425 34244 14449 34246
rect 14505 34244 14529 34246
rect 14289 34224 14585 34244
rect 14188 34060 14240 34066
rect 14188 34002 14240 34008
rect 14200 33318 14228 34002
rect 14096 33312 14148 33318
rect 14096 33254 14148 33260
rect 14188 33312 14240 33318
rect 14188 33254 14240 33260
rect 14108 33046 14136 33254
rect 14096 33040 14148 33046
rect 14096 32982 14148 32988
rect 14108 32298 14136 32982
rect 14200 32978 14228 33254
rect 14289 33212 14585 33232
rect 14345 33210 14369 33212
rect 14425 33210 14449 33212
rect 14505 33210 14529 33212
rect 14367 33158 14369 33210
rect 14431 33158 14443 33210
rect 14505 33158 14507 33210
rect 14345 33156 14369 33158
rect 14425 33156 14449 33158
rect 14505 33156 14529 33158
rect 14289 33136 14585 33156
rect 14660 32978 14688 34546
rect 14740 34536 14792 34542
rect 14740 34478 14792 34484
rect 14188 32972 14240 32978
rect 14188 32914 14240 32920
rect 14648 32972 14700 32978
rect 14648 32914 14700 32920
rect 14188 32836 14240 32842
rect 14188 32778 14240 32784
rect 14096 32292 14148 32298
rect 14096 32234 14148 32240
rect 14200 30297 14228 32778
rect 14660 32570 14688 32914
rect 14648 32564 14700 32570
rect 14648 32506 14700 32512
rect 14289 32124 14585 32144
rect 14345 32122 14369 32124
rect 14425 32122 14449 32124
rect 14505 32122 14529 32124
rect 14367 32070 14369 32122
rect 14431 32070 14443 32122
rect 14505 32070 14507 32122
rect 14345 32068 14369 32070
rect 14425 32068 14449 32070
rect 14505 32068 14529 32070
rect 14289 32048 14585 32068
rect 14660 31890 14688 32506
rect 14556 31884 14608 31890
rect 14556 31826 14608 31832
rect 14648 31884 14700 31890
rect 14648 31826 14700 31832
rect 14568 31124 14596 31826
rect 14660 31482 14688 31826
rect 14648 31476 14700 31482
rect 14648 31418 14700 31424
rect 14648 31136 14700 31142
rect 14568 31096 14648 31124
rect 14648 31078 14700 31084
rect 14289 31036 14585 31056
rect 14345 31034 14369 31036
rect 14425 31034 14449 31036
rect 14505 31034 14529 31036
rect 14367 30982 14369 31034
rect 14431 30982 14443 31034
rect 14505 30982 14507 31034
rect 14345 30980 14369 30982
rect 14425 30980 14449 30982
rect 14505 30980 14529 30982
rect 14289 30960 14585 30980
rect 14186 30288 14242 30297
rect 14186 30223 14242 30232
rect 14289 29948 14585 29968
rect 14345 29946 14369 29948
rect 14425 29946 14449 29948
rect 14505 29946 14529 29948
rect 14367 29894 14369 29946
rect 14431 29894 14443 29946
rect 14505 29894 14507 29946
rect 14345 29892 14369 29894
rect 14425 29892 14449 29894
rect 14505 29892 14529 29894
rect 14289 29872 14585 29892
rect 14372 29708 14424 29714
rect 14372 29650 14424 29656
rect 14384 29306 14412 29650
rect 14372 29300 14424 29306
rect 14372 29242 14424 29248
rect 14660 29170 14688 31078
rect 14648 29164 14700 29170
rect 14648 29106 14700 29112
rect 14289 28860 14585 28880
rect 14345 28858 14369 28860
rect 14425 28858 14449 28860
rect 14505 28858 14529 28860
rect 14367 28806 14369 28858
rect 14431 28806 14443 28858
rect 14505 28806 14507 28858
rect 14345 28804 14369 28806
rect 14425 28804 14449 28806
rect 14505 28804 14529 28806
rect 14289 28784 14585 28804
rect 14752 28762 14780 34478
rect 14844 34202 14872 40718
rect 14924 40588 14976 40594
rect 14924 40530 14976 40536
rect 14936 40186 14964 40530
rect 14924 40180 14976 40186
rect 14924 40122 14976 40128
rect 14936 37890 14964 40122
rect 15028 38010 15056 40870
rect 15120 39409 15148 42026
rect 15212 40769 15240 62070
rect 15396 61169 15424 62086
rect 15382 61160 15438 61169
rect 15382 61095 15438 61104
rect 15382 61024 15438 61033
rect 15382 60959 15438 60968
rect 15396 60081 15424 60959
rect 15382 60072 15438 60081
rect 15382 60007 15438 60016
rect 15488 57089 15516 66098
rect 15660 64456 15712 64462
rect 15660 64398 15712 64404
rect 15568 63912 15620 63918
rect 15568 63854 15620 63860
rect 15580 63578 15608 63854
rect 15672 63782 15700 64398
rect 15660 63776 15712 63782
rect 15660 63718 15712 63724
rect 15568 63572 15620 63578
rect 15568 63514 15620 63520
rect 15568 63436 15620 63442
rect 15568 63378 15620 63384
rect 15580 62286 15608 63378
rect 15568 62280 15620 62286
rect 15566 62248 15568 62257
rect 15620 62248 15622 62257
rect 15566 62183 15622 62192
rect 15568 61736 15620 61742
rect 15568 61678 15620 61684
rect 15580 57882 15608 61678
rect 15672 59242 15700 63718
rect 15752 63572 15804 63578
rect 15752 63514 15804 63520
rect 15764 62830 15792 63514
rect 15752 62824 15804 62830
rect 15752 62766 15804 62772
rect 15936 61600 15988 61606
rect 15936 61542 15988 61548
rect 15948 59566 15976 61542
rect 16040 60489 16068 71334
rect 16132 70854 16160 71470
rect 16120 70848 16172 70854
rect 16120 70790 16172 70796
rect 16132 68814 16160 70790
rect 16120 68808 16172 68814
rect 16120 68750 16172 68756
rect 16120 68672 16172 68678
rect 16120 68614 16172 68620
rect 16132 68270 16160 68614
rect 16120 68264 16172 68270
rect 16120 68206 16172 68212
rect 16132 66706 16160 68206
rect 16120 66700 16172 66706
rect 16120 66642 16172 66648
rect 16132 65754 16160 66642
rect 16120 65748 16172 65754
rect 16120 65690 16172 65696
rect 16132 65006 16160 65690
rect 16120 65000 16172 65006
rect 16120 64942 16172 64948
rect 16132 64530 16160 64942
rect 16120 64524 16172 64530
rect 16120 64466 16172 64472
rect 16212 63232 16264 63238
rect 16210 63200 16212 63209
rect 16264 63200 16266 63209
rect 16210 63135 16266 63144
rect 16120 61056 16172 61062
rect 16120 60998 16172 61004
rect 16132 60897 16160 60998
rect 16118 60888 16174 60897
rect 16118 60823 16174 60832
rect 16120 60648 16172 60654
rect 16120 60590 16172 60596
rect 16026 60480 16082 60489
rect 16026 60415 16082 60424
rect 16132 60314 16160 60590
rect 16120 60308 16172 60314
rect 16120 60250 16172 60256
rect 15936 59560 15988 59566
rect 15936 59502 15988 59508
rect 15672 59214 15884 59242
rect 15856 57905 15884 59214
rect 15948 58886 15976 59502
rect 15936 58880 15988 58886
rect 15936 58822 15988 58828
rect 15948 58138 15976 58822
rect 15936 58132 15988 58138
rect 15936 58074 15988 58080
rect 15842 57896 15898 57905
rect 15580 57854 15792 57882
rect 15568 57792 15620 57798
rect 15568 57734 15620 57740
rect 15474 57080 15530 57089
rect 15474 57015 15530 57024
rect 15384 55820 15436 55826
rect 15384 55762 15436 55768
rect 15292 55616 15344 55622
rect 15292 55558 15344 55564
rect 15304 55185 15332 55558
rect 15396 55214 15424 55762
rect 15476 55752 15528 55758
rect 15476 55694 15528 55700
rect 15384 55208 15436 55214
rect 15290 55176 15346 55185
rect 15384 55150 15436 55156
rect 15290 55111 15346 55120
rect 15382 55040 15438 55049
rect 15382 54975 15438 54984
rect 15292 54120 15344 54126
rect 15292 54062 15344 54068
rect 15304 53650 15332 54062
rect 15292 53644 15344 53650
rect 15292 53586 15344 53592
rect 15292 53100 15344 53106
rect 15292 53042 15344 53048
rect 15304 52329 15332 53042
rect 15396 52465 15424 54975
rect 15488 53417 15516 55694
rect 15580 54641 15608 57734
rect 15660 56840 15712 56846
rect 15660 56782 15712 56788
rect 15672 56166 15700 56782
rect 15660 56160 15712 56166
rect 15660 56102 15712 56108
rect 15566 54632 15622 54641
rect 15566 54567 15622 54576
rect 15474 53408 15530 53417
rect 15474 53343 15530 53352
rect 15568 53032 15620 53038
rect 15568 52974 15620 52980
rect 15476 52488 15528 52494
rect 15382 52456 15438 52465
rect 15476 52430 15528 52436
rect 15382 52391 15438 52400
rect 15290 52320 15346 52329
rect 15290 52255 15346 52264
rect 15384 51944 15436 51950
rect 15384 51886 15436 51892
rect 15396 51406 15424 51886
rect 15488 51456 15516 52430
rect 15580 51950 15608 52974
rect 15568 51944 15620 51950
rect 15568 51886 15620 51892
rect 15568 51468 15620 51474
rect 15488 51428 15568 51456
rect 15568 51410 15620 51416
rect 15384 51400 15436 51406
rect 15436 51360 15516 51388
rect 15384 51342 15436 51348
rect 15384 51264 15436 51270
rect 15384 51206 15436 51212
rect 15292 51060 15344 51066
rect 15292 51002 15344 51008
rect 15304 50969 15332 51002
rect 15290 50960 15346 50969
rect 15290 50895 15346 50904
rect 15292 50720 15344 50726
rect 15292 50662 15344 50668
rect 15304 49366 15332 50662
rect 15396 49842 15424 51206
rect 15488 50726 15516 51360
rect 15476 50720 15528 50726
rect 15476 50662 15528 50668
rect 15384 49836 15436 49842
rect 15384 49778 15436 49784
rect 15292 49360 15344 49366
rect 15292 49302 15344 49308
rect 15384 49360 15436 49366
rect 15384 49302 15436 49308
rect 15292 48680 15344 48686
rect 15292 48622 15344 48628
rect 15304 45626 15332 48622
rect 15292 45620 15344 45626
rect 15292 45562 15344 45568
rect 15396 45472 15424 49302
rect 15488 48142 15516 50662
rect 15580 50386 15608 51410
rect 15568 50380 15620 50386
rect 15568 50322 15620 50328
rect 15580 49434 15608 50322
rect 15672 49473 15700 56102
rect 15764 52873 15792 57854
rect 15842 57831 15898 57840
rect 15948 57390 15976 58074
rect 16316 58041 16344 72655
rect 17498 72584 17554 72593
rect 17498 72519 17554 72528
rect 17512 71738 17540 72519
rect 17622 71836 17918 71856
rect 17678 71834 17702 71836
rect 17758 71834 17782 71836
rect 17838 71834 17862 71836
rect 17700 71782 17702 71834
rect 17764 71782 17776 71834
rect 17838 71782 17840 71834
rect 17678 71780 17702 71782
rect 17758 71780 17782 71782
rect 17838 71780 17862 71782
rect 17622 71760 17918 71780
rect 17500 71732 17552 71738
rect 17500 71674 17552 71680
rect 17622 70748 17918 70768
rect 17678 70746 17702 70748
rect 17758 70746 17782 70748
rect 17838 70746 17862 70748
rect 17700 70694 17702 70746
rect 17764 70694 17776 70746
rect 17838 70694 17840 70746
rect 17678 70692 17702 70694
rect 17758 70692 17782 70694
rect 17838 70692 17862 70694
rect 17622 70672 17918 70692
rect 17622 69660 17918 69680
rect 17678 69658 17702 69660
rect 17758 69658 17782 69660
rect 17838 69658 17862 69660
rect 17700 69606 17702 69658
rect 17764 69606 17776 69658
rect 17838 69606 17840 69658
rect 17678 69604 17702 69606
rect 17758 69604 17782 69606
rect 17838 69604 17862 69606
rect 17622 69584 17918 69604
rect 17498 68776 17554 68785
rect 17498 68711 17554 68720
rect 17512 68474 17540 68711
rect 17622 68572 17918 68592
rect 17678 68570 17702 68572
rect 17758 68570 17782 68572
rect 17838 68570 17862 68572
rect 17700 68518 17702 68570
rect 17764 68518 17776 68570
rect 17838 68518 17840 68570
rect 17678 68516 17702 68518
rect 17758 68516 17782 68518
rect 17838 68516 17862 68518
rect 17622 68496 17918 68516
rect 17500 68468 17552 68474
rect 17500 68410 17552 68416
rect 16396 68264 16448 68270
rect 16396 68206 16448 68212
rect 16408 65521 16436 68206
rect 17132 67720 17184 67726
rect 17132 67662 17184 67668
rect 17144 67289 17172 67662
rect 17622 67484 17918 67504
rect 17678 67482 17702 67484
rect 17758 67482 17782 67484
rect 17838 67482 17862 67484
rect 17700 67430 17702 67482
rect 17764 67430 17776 67482
rect 17838 67430 17840 67482
rect 17678 67428 17702 67430
rect 17758 67428 17782 67430
rect 17838 67428 17862 67430
rect 17622 67408 17918 67428
rect 17130 67280 17186 67289
rect 17130 67215 17186 67224
rect 16488 67176 16540 67182
rect 16488 67118 16540 67124
rect 17498 67144 17554 67153
rect 16394 65512 16450 65521
rect 16394 65447 16450 65456
rect 16396 65000 16448 65006
rect 16396 64942 16448 64948
rect 16408 63889 16436 64942
rect 16500 64569 16528 67118
rect 17498 67079 17554 67088
rect 17512 67046 17540 67079
rect 17500 67040 17552 67046
rect 17500 66982 17552 66988
rect 16672 66632 16724 66638
rect 16670 66600 16672 66609
rect 16724 66600 16726 66609
rect 16670 66535 16726 66544
rect 17622 66396 17918 66416
rect 17678 66394 17702 66396
rect 17758 66394 17782 66396
rect 17838 66394 17862 66396
rect 17700 66342 17702 66394
rect 17764 66342 17776 66394
rect 17838 66342 17840 66394
rect 17678 66340 17702 66342
rect 17758 66340 17782 66342
rect 17838 66340 17862 66342
rect 17622 66320 17918 66340
rect 16580 65952 16632 65958
rect 16580 65894 16632 65900
rect 16946 65920 17002 65929
rect 16486 64560 16542 64569
rect 16486 64495 16542 64504
rect 16488 63912 16540 63918
rect 16394 63880 16450 63889
rect 16488 63854 16540 63860
rect 16394 63815 16450 63824
rect 16500 61849 16528 63854
rect 16486 61840 16542 61849
rect 16486 61775 16542 61784
rect 16488 60648 16540 60654
rect 16488 60590 16540 60596
rect 16396 59560 16448 59566
rect 16396 59502 16448 59508
rect 16408 58449 16436 59502
rect 16500 59129 16528 60590
rect 16592 60217 16620 65894
rect 16946 65855 17002 65864
rect 16856 64456 16908 64462
rect 16854 64424 16856 64433
rect 16908 64424 16910 64433
rect 16854 64359 16910 64368
rect 16960 63034 16988 65855
rect 17498 65648 17554 65657
rect 17498 65583 17554 65592
rect 17512 65210 17540 65583
rect 17622 65308 17918 65328
rect 17678 65306 17702 65308
rect 17758 65306 17782 65308
rect 17838 65306 17862 65308
rect 17700 65254 17702 65306
rect 17764 65254 17776 65306
rect 17838 65254 17840 65306
rect 17678 65252 17702 65254
rect 17758 65252 17782 65254
rect 17838 65252 17862 65254
rect 17622 65232 17918 65252
rect 17500 65204 17552 65210
rect 17500 65146 17552 65152
rect 17622 64220 17918 64240
rect 17678 64218 17702 64220
rect 17758 64218 17782 64220
rect 17838 64218 17862 64220
rect 17700 64166 17702 64218
rect 17764 64166 17776 64218
rect 17838 64166 17840 64218
rect 17678 64164 17702 64166
rect 17758 64164 17782 64166
rect 17838 64164 17862 64166
rect 17622 64144 17918 64164
rect 17500 63776 17552 63782
rect 17500 63718 17552 63724
rect 16948 63028 17000 63034
rect 16948 62970 17000 62976
rect 17512 62801 17540 63718
rect 17622 63132 17918 63152
rect 17678 63130 17702 63132
rect 17758 63130 17782 63132
rect 17838 63130 17862 63132
rect 17700 63078 17702 63130
rect 17764 63078 17776 63130
rect 17838 63078 17840 63130
rect 17678 63076 17702 63078
rect 17758 63076 17782 63078
rect 17838 63076 17862 63078
rect 17622 63056 17918 63076
rect 17498 62792 17554 62801
rect 17498 62727 17554 62736
rect 17622 62044 17918 62064
rect 17678 62042 17702 62044
rect 17758 62042 17782 62044
rect 17838 62042 17862 62044
rect 17700 61990 17702 62042
rect 17764 61990 17776 62042
rect 17838 61990 17840 62042
rect 17678 61988 17702 61990
rect 17758 61988 17782 61990
rect 17838 61988 17862 61990
rect 17622 61968 17918 61988
rect 16672 61600 16724 61606
rect 16672 61542 16724 61548
rect 16684 60353 16712 61542
rect 17622 60956 17918 60976
rect 17678 60954 17702 60956
rect 17758 60954 17782 60956
rect 17838 60954 17862 60956
rect 17700 60902 17702 60954
rect 17764 60902 17776 60954
rect 17838 60902 17840 60954
rect 17678 60900 17702 60902
rect 17758 60900 17782 60902
rect 17838 60900 17862 60902
rect 17622 60880 17918 60900
rect 17498 60616 17554 60625
rect 17498 60551 17554 60560
rect 17512 60518 17540 60551
rect 17500 60512 17552 60518
rect 17500 60454 17552 60460
rect 16670 60344 16726 60353
rect 16670 60279 16726 60288
rect 16578 60208 16634 60217
rect 16578 60143 16634 60152
rect 17622 59868 17918 59888
rect 17678 59866 17702 59868
rect 17758 59866 17782 59868
rect 17838 59866 17862 59868
rect 17700 59814 17702 59866
rect 17764 59814 17776 59866
rect 17838 59814 17840 59866
rect 17678 59812 17702 59814
rect 17758 59812 17782 59814
rect 17838 59812 17862 59814
rect 17622 59792 17918 59812
rect 16486 59120 16542 59129
rect 16486 59055 16542 59064
rect 17622 58780 17918 58800
rect 17678 58778 17702 58780
rect 17758 58778 17782 58780
rect 17838 58778 17862 58780
rect 17700 58726 17702 58778
rect 17764 58726 17776 58778
rect 17838 58726 17840 58778
rect 17678 58724 17702 58726
rect 17758 58724 17782 58726
rect 17838 58724 17862 58726
rect 17622 58704 17918 58724
rect 16394 58440 16450 58449
rect 16394 58375 16450 58384
rect 16302 58032 16358 58041
rect 16302 57967 16358 57976
rect 17622 57692 17918 57712
rect 17678 57690 17702 57692
rect 17758 57690 17782 57692
rect 17838 57690 17862 57692
rect 17700 57638 17702 57690
rect 17764 57638 17776 57690
rect 17838 57638 17840 57690
rect 17678 57636 17702 57638
rect 17758 57636 17782 57638
rect 17838 57636 17862 57638
rect 17622 57616 17918 57636
rect 15936 57384 15988 57390
rect 16212 57384 16264 57390
rect 15936 57326 15988 57332
rect 16026 57352 16082 57361
rect 16212 57326 16264 57332
rect 16026 57287 16082 57296
rect 15936 54528 15988 54534
rect 15936 54470 15988 54476
rect 15844 54188 15896 54194
rect 15844 54130 15896 54136
rect 15750 52864 15806 52873
rect 15750 52799 15806 52808
rect 15856 51218 15884 54130
rect 15948 54126 15976 54470
rect 16040 54233 16068 57287
rect 16224 56409 16252 57326
rect 17316 57248 17368 57254
rect 17316 57190 17368 57196
rect 16672 56704 16724 56710
rect 16670 56672 16672 56681
rect 16724 56672 16726 56681
rect 16670 56607 16726 56616
rect 16210 56400 16266 56409
rect 16210 56335 16266 56344
rect 16396 56296 16448 56302
rect 16396 56238 16448 56244
rect 16304 55752 16356 55758
rect 16408 55729 16436 56238
rect 17328 55962 17356 57190
rect 17622 56604 17918 56624
rect 17678 56602 17702 56604
rect 17758 56602 17782 56604
rect 17838 56602 17862 56604
rect 17700 56550 17702 56602
rect 17764 56550 17776 56602
rect 17838 56550 17840 56602
rect 17678 56548 17702 56550
rect 17758 56548 17782 56550
rect 17838 56548 17862 56550
rect 17622 56528 17918 56548
rect 17500 56160 17552 56166
rect 17500 56102 17552 56108
rect 17316 55956 17368 55962
rect 17316 55898 17368 55904
rect 17512 55865 17540 56102
rect 17498 55856 17554 55865
rect 17408 55820 17460 55826
rect 17498 55791 17554 55800
rect 17408 55762 17460 55768
rect 17132 55752 17184 55758
rect 16304 55694 16356 55700
rect 16394 55720 16450 55729
rect 16316 55418 16344 55694
rect 17132 55694 17184 55700
rect 16394 55655 16450 55664
rect 17144 55457 17172 55694
rect 17130 55448 17186 55457
rect 16304 55412 16356 55418
rect 17130 55383 17132 55392
rect 16304 55354 16356 55360
rect 17184 55383 17186 55392
rect 17132 55354 17184 55360
rect 16120 54664 16172 54670
rect 16120 54606 16172 54612
rect 16026 54224 16082 54233
rect 16026 54159 16082 54168
rect 15936 54120 15988 54126
rect 15988 54080 16068 54108
rect 15936 54062 15988 54068
rect 15936 53644 15988 53650
rect 15936 53586 15988 53592
rect 15948 53038 15976 53586
rect 15936 53032 15988 53038
rect 15936 52974 15988 52980
rect 15948 52902 15976 52974
rect 15936 52896 15988 52902
rect 15936 52838 15988 52844
rect 15948 52358 15976 52838
rect 15936 52352 15988 52358
rect 15936 52294 15988 52300
rect 15948 52018 15976 52294
rect 15936 52012 15988 52018
rect 15936 51954 15988 51960
rect 16040 51474 16068 54080
rect 16132 53990 16160 54606
rect 16120 53984 16172 53990
rect 16120 53926 16172 53932
rect 16028 51468 16080 51474
rect 16028 51410 16080 51416
rect 15856 51190 15976 51218
rect 15752 50924 15804 50930
rect 15752 50866 15804 50872
rect 15764 50386 15792 50866
rect 15752 50380 15804 50386
rect 15752 50322 15804 50328
rect 15658 49464 15714 49473
rect 15568 49428 15620 49434
rect 15658 49399 15714 49408
rect 15568 49370 15620 49376
rect 15580 48890 15608 49370
rect 15764 49366 15792 50322
rect 15844 50312 15896 50318
rect 15844 50254 15896 50260
rect 15752 49360 15804 49366
rect 15658 49328 15714 49337
rect 15752 49302 15804 49308
rect 15658 49263 15714 49272
rect 15568 48884 15620 48890
rect 15568 48826 15620 48832
rect 15476 48136 15528 48142
rect 15476 48078 15528 48084
rect 15476 48000 15528 48006
rect 15476 47942 15528 47948
rect 15488 47462 15516 47942
rect 15568 47524 15620 47530
rect 15568 47466 15620 47472
rect 15476 47456 15528 47462
rect 15476 47398 15528 47404
rect 15488 46986 15516 47398
rect 15580 47190 15608 47466
rect 15568 47184 15620 47190
rect 15566 47152 15568 47161
rect 15620 47152 15622 47161
rect 15566 47087 15622 47096
rect 15580 47061 15608 47087
rect 15672 47002 15700 49263
rect 15752 48136 15804 48142
rect 15752 48078 15804 48084
rect 15476 46980 15528 46986
rect 15476 46922 15528 46928
rect 15580 46974 15700 47002
rect 15476 45960 15528 45966
rect 15476 45902 15528 45908
rect 15304 45444 15424 45472
rect 15304 42702 15332 45444
rect 15488 45422 15516 45902
rect 15476 45416 15528 45422
rect 15476 45358 15528 45364
rect 15384 45280 15436 45286
rect 15384 45222 15436 45228
rect 15396 44266 15424 45222
rect 15384 44260 15436 44266
rect 15384 44202 15436 44208
rect 15396 43110 15424 44202
rect 15384 43104 15436 43110
rect 15384 43046 15436 43052
rect 15292 42696 15344 42702
rect 15292 42638 15344 42644
rect 15304 42362 15332 42638
rect 15292 42356 15344 42362
rect 15292 42298 15344 42304
rect 15290 42256 15346 42265
rect 15290 42191 15346 42200
rect 15198 40760 15254 40769
rect 15198 40695 15254 40704
rect 15200 40656 15252 40662
rect 15200 40598 15252 40604
rect 15212 40186 15240 40598
rect 15200 40180 15252 40186
rect 15200 40122 15252 40128
rect 15200 39908 15252 39914
rect 15200 39850 15252 39856
rect 15106 39400 15162 39409
rect 15106 39335 15162 39344
rect 15212 39302 15240 39850
rect 15304 39574 15332 42191
rect 15396 41682 15424 43046
rect 15384 41676 15436 41682
rect 15384 41618 15436 41624
rect 15396 41274 15424 41618
rect 15488 41585 15516 45358
rect 15580 45354 15608 46974
rect 15660 45620 15712 45626
rect 15660 45562 15712 45568
rect 15568 45348 15620 45354
rect 15568 45290 15620 45296
rect 15568 45076 15620 45082
rect 15568 45018 15620 45024
rect 15580 43994 15608 45018
rect 15672 44198 15700 45562
rect 15764 45558 15792 48078
rect 15856 47598 15884 50254
rect 15948 48210 15976 51190
rect 16040 50522 16068 51410
rect 16132 51241 16160 53926
rect 16212 53644 16264 53650
rect 16212 53586 16264 53592
rect 16224 52698 16252 53586
rect 16212 52692 16264 52698
rect 16212 52634 16264 52640
rect 16224 51950 16252 52634
rect 16316 52086 16344 55354
rect 17144 55323 17172 55354
rect 17420 55282 17448 55762
rect 17622 55516 17918 55536
rect 17678 55514 17702 55516
rect 17758 55514 17782 55516
rect 17838 55514 17862 55516
rect 17700 55462 17702 55514
rect 17764 55462 17776 55514
rect 17838 55462 17840 55514
rect 17678 55460 17702 55462
rect 17758 55460 17782 55462
rect 17838 55460 17862 55462
rect 17622 55440 17918 55460
rect 17408 55276 17460 55282
rect 17408 55218 17460 55224
rect 16764 55072 16816 55078
rect 16764 55014 16816 55020
rect 16396 54596 16448 54602
rect 16396 54538 16448 54544
rect 16408 54126 16436 54538
rect 16396 54120 16448 54126
rect 16396 54062 16448 54068
rect 16672 54120 16724 54126
rect 16672 54062 16724 54068
rect 16304 52080 16356 52086
rect 16304 52022 16356 52028
rect 16212 51944 16264 51950
rect 16264 51904 16344 51932
rect 16212 51886 16264 51892
rect 16212 51468 16264 51474
rect 16212 51410 16264 51416
rect 16118 51232 16174 51241
rect 16118 51167 16174 51176
rect 16118 50960 16174 50969
rect 16118 50895 16174 50904
rect 16028 50516 16080 50522
rect 16028 50458 16080 50464
rect 16040 49978 16068 50458
rect 16028 49972 16080 49978
rect 16028 49914 16080 49920
rect 16026 49872 16082 49881
rect 16026 49807 16082 49816
rect 15936 48204 15988 48210
rect 15936 48146 15988 48152
rect 15844 47592 15896 47598
rect 15844 47534 15896 47540
rect 15844 47456 15896 47462
rect 15844 47398 15896 47404
rect 15752 45552 15804 45558
rect 15752 45494 15804 45500
rect 15764 44946 15792 45494
rect 15752 44940 15804 44946
rect 15752 44882 15804 44888
rect 15764 44334 15792 44882
rect 15856 44742 15884 47398
rect 15948 47258 15976 48146
rect 15936 47252 15988 47258
rect 15936 47194 15988 47200
rect 15936 45960 15988 45966
rect 15936 45902 15988 45908
rect 15948 45121 15976 45902
rect 15934 45112 15990 45121
rect 15934 45047 15990 45056
rect 15936 45008 15988 45014
rect 15936 44950 15988 44956
rect 15844 44736 15896 44742
rect 15844 44678 15896 44684
rect 15752 44328 15804 44334
rect 15752 44270 15804 44276
rect 15660 44192 15712 44198
rect 15660 44134 15712 44140
rect 15658 44024 15714 44033
rect 15568 43988 15620 43994
rect 15658 43959 15714 43968
rect 15568 43930 15620 43936
rect 15580 42838 15608 43930
rect 15568 42832 15620 42838
rect 15568 42774 15620 42780
rect 15568 42628 15620 42634
rect 15568 42570 15620 42576
rect 15580 42362 15608 42570
rect 15568 42356 15620 42362
rect 15568 42298 15620 42304
rect 15580 41818 15608 42298
rect 15568 41812 15620 41818
rect 15568 41754 15620 41760
rect 15566 41712 15622 41721
rect 15566 41647 15622 41656
rect 15474 41576 15530 41585
rect 15474 41511 15530 41520
rect 15580 41460 15608 41647
rect 15488 41432 15608 41460
rect 15384 41268 15436 41274
rect 15384 41210 15436 41216
rect 15292 39568 15344 39574
rect 15292 39510 15344 39516
rect 15292 39432 15344 39438
rect 15292 39374 15344 39380
rect 15200 39296 15252 39302
rect 15200 39238 15252 39244
rect 15016 38004 15068 38010
rect 15016 37946 15068 37952
rect 15106 37904 15162 37913
rect 14936 37862 15056 37890
rect 14924 37800 14976 37806
rect 14924 37742 14976 37748
rect 14936 37466 14964 37742
rect 14924 37460 14976 37466
rect 14924 37402 14976 37408
rect 14936 36582 14964 37402
rect 14924 36576 14976 36582
rect 14924 36518 14976 36524
rect 14936 36242 14964 36518
rect 14924 36236 14976 36242
rect 14924 36178 14976 36184
rect 14936 35834 14964 36178
rect 14924 35828 14976 35834
rect 14924 35770 14976 35776
rect 14924 35556 14976 35562
rect 14924 35498 14976 35504
rect 14936 35290 14964 35498
rect 14924 35284 14976 35290
rect 14924 35226 14976 35232
rect 14936 34610 14964 35226
rect 14924 34604 14976 34610
rect 14924 34546 14976 34552
rect 14832 34196 14884 34202
rect 14832 34138 14884 34144
rect 14830 34096 14886 34105
rect 14830 34031 14832 34040
rect 14884 34031 14886 34040
rect 14832 34002 14884 34008
rect 14844 33658 14872 34002
rect 14924 33992 14976 33998
rect 14924 33934 14976 33940
rect 14832 33652 14884 33658
rect 14832 33594 14884 33600
rect 14832 33312 14884 33318
rect 14832 33254 14884 33260
rect 14844 31890 14872 33254
rect 14936 33046 14964 33934
rect 14924 33040 14976 33046
rect 14924 32982 14976 32988
rect 14832 31884 14884 31890
rect 14832 31826 14884 31832
rect 14844 31414 14872 31826
rect 14832 31408 14884 31414
rect 14832 31350 14884 31356
rect 14830 30288 14886 30297
rect 14830 30223 14886 30232
rect 14740 28756 14792 28762
rect 14740 28698 14792 28704
rect 14648 28620 14700 28626
rect 14648 28562 14700 28568
rect 14660 27878 14688 28562
rect 14648 27872 14700 27878
rect 14648 27814 14700 27820
rect 14289 27772 14585 27792
rect 14345 27770 14369 27772
rect 14425 27770 14449 27772
rect 14505 27770 14529 27772
rect 14367 27718 14369 27770
rect 14431 27718 14443 27770
rect 14505 27718 14507 27770
rect 14345 27716 14369 27718
rect 14425 27716 14449 27718
rect 14505 27716 14529 27718
rect 14289 27696 14585 27716
rect 14188 27532 14240 27538
rect 14188 27474 14240 27480
rect 14200 27130 14228 27474
rect 14648 27464 14700 27470
rect 14648 27406 14700 27412
rect 14188 27124 14240 27130
rect 14188 27066 14240 27072
rect 14188 26920 14240 26926
rect 14188 26862 14240 26868
rect 14096 26444 14148 26450
rect 14096 26386 14148 26392
rect 14108 25770 14136 26386
rect 14200 26382 14228 26862
rect 14289 26684 14585 26704
rect 14345 26682 14369 26684
rect 14425 26682 14449 26684
rect 14505 26682 14529 26684
rect 14367 26630 14369 26682
rect 14431 26630 14443 26682
rect 14505 26630 14507 26682
rect 14345 26628 14369 26630
rect 14425 26628 14449 26630
rect 14505 26628 14529 26630
rect 14289 26608 14585 26628
rect 14188 26376 14240 26382
rect 14188 26318 14240 26324
rect 14096 25764 14148 25770
rect 14096 25706 14148 25712
rect 14289 25596 14585 25616
rect 14345 25594 14369 25596
rect 14425 25594 14449 25596
rect 14505 25594 14529 25596
rect 14367 25542 14369 25594
rect 14431 25542 14443 25594
rect 14505 25542 14507 25594
rect 14345 25540 14369 25542
rect 14425 25540 14449 25542
rect 14505 25540 14529 25542
rect 14289 25520 14585 25540
rect 14002 24848 14058 24857
rect 13912 24812 13964 24818
rect 14002 24783 14058 24792
rect 13912 24754 13964 24760
rect 14188 24744 14240 24750
rect 14188 24686 14240 24692
rect 14004 24676 14056 24682
rect 14004 24618 14056 24624
rect 13820 24608 13872 24614
rect 13820 24550 13872 24556
rect 13832 22817 13860 24550
rect 14016 24410 14044 24618
rect 14200 24410 14228 24686
rect 14289 24508 14585 24528
rect 14345 24506 14369 24508
rect 14425 24506 14449 24508
rect 14505 24506 14529 24508
rect 14367 24454 14369 24506
rect 14431 24454 14443 24506
rect 14505 24454 14507 24506
rect 14345 24452 14369 24454
rect 14425 24452 14449 24454
rect 14505 24452 14529 24454
rect 14289 24432 14585 24452
rect 14004 24404 14056 24410
rect 14004 24346 14056 24352
rect 14188 24404 14240 24410
rect 14188 24346 14240 24352
rect 14556 24268 14608 24274
rect 14556 24210 14608 24216
rect 14568 23866 14596 24210
rect 14556 23860 14608 23866
rect 14556 23802 14608 23808
rect 14660 23769 14688 27406
rect 14844 24750 14872 30223
rect 15028 27538 15056 37862
rect 15106 37839 15162 37848
rect 15120 37262 15148 37839
rect 15108 37256 15160 37262
rect 15108 37198 15160 37204
rect 15108 37120 15160 37126
rect 15108 37062 15160 37068
rect 15120 32881 15148 37062
rect 15212 36922 15240 39238
rect 15304 38894 15332 39374
rect 15396 39098 15424 41210
rect 15488 41138 15516 41432
rect 15566 41304 15622 41313
rect 15566 41239 15622 41248
rect 15476 41132 15528 41138
rect 15476 41074 15528 41080
rect 15476 40928 15528 40934
rect 15476 40870 15528 40876
rect 15488 40458 15516 40870
rect 15476 40452 15528 40458
rect 15476 40394 15528 40400
rect 15476 39296 15528 39302
rect 15476 39238 15528 39244
rect 15384 39092 15436 39098
rect 15384 39034 15436 39040
rect 15292 38888 15344 38894
rect 15292 38830 15344 38836
rect 15292 38548 15344 38554
rect 15292 38490 15344 38496
rect 15200 36916 15252 36922
rect 15200 36858 15252 36864
rect 15304 36854 15332 38490
rect 15382 37496 15438 37505
rect 15382 37431 15384 37440
rect 15436 37431 15438 37440
rect 15384 37402 15436 37408
rect 15382 37224 15438 37233
rect 15382 37159 15438 37168
rect 15292 36848 15344 36854
rect 15292 36790 15344 36796
rect 15200 36372 15252 36378
rect 15200 36314 15252 36320
rect 15212 33114 15240 36314
rect 15304 35766 15332 36790
rect 15292 35760 15344 35766
rect 15292 35702 15344 35708
rect 15304 34678 15332 35702
rect 15292 34672 15344 34678
rect 15292 34614 15344 34620
rect 15200 33108 15252 33114
rect 15200 33050 15252 33056
rect 15106 32872 15162 32881
rect 15106 32807 15162 32816
rect 15212 32366 15240 33050
rect 15396 32450 15424 37159
rect 15304 32422 15424 32450
rect 15200 32360 15252 32366
rect 15200 32302 15252 32308
rect 15304 32298 15332 32422
rect 15384 32360 15436 32366
rect 15384 32302 15436 32308
rect 15292 32292 15344 32298
rect 15292 32234 15344 32240
rect 15304 31346 15332 32234
rect 15396 31906 15424 32302
rect 15488 32026 15516 39238
rect 15580 38418 15608 41239
rect 15672 41206 15700 43959
rect 15764 43858 15792 44270
rect 15752 43852 15804 43858
rect 15752 43794 15804 43800
rect 15856 43489 15884 44678
rect 15948 43654 15976 44950
rect 16040 43858 16068 49807
rect 16132 47462 16160 50895
rect 16224 50454 16252 51410
rect 16212 50448 16264 50454
rect 16212 50390 16264 50396
rect 16212 50312 16264 50318
rect 16212 50254 16264 50260
rect 16224 49910 16252 50254
rect 16212 49904 16264 49910
rect 16316 49881 16344 51904
rect 16408 51474 16436 54062
rect 16684 53582 16712 54062
rect 16672 53576 16724 53582
rect 16672 53518 16724 53524
rect 16580 53440 16632 53446
rect 16578 53408 16580 53417
rect 16632 53408 16634 53417
rect 16578 53343 16634 53352
rect 16684 53038 16712 53518
rect 16672 53032 16724 53038
rect 16776 53009 16804 55014
rect 16856 54732 16908 54738
rect 16856 54674 16908 54680
rect 16868 54330 16896 54674
rect 17132 54664 17184 54670
rect 17132 54606 17184 54612
rect 16948 54596 17000 54602
rect 16948 54538 17000 54544
rect 16856 54324 16908 54330
rect 16856 54266 16908 54272
rect 16854 53136 16910 53145
rect 16854 53071 16910 53080
rect 16672 52974 16724 52980
rect 16762 53000 16818 53009
rect 16762 52935 16818 52944
rect 16868 52562 16896 53071
rect 16856 52556 16908 52562
rect 16856 52498 16908 52504
rect 16868 52154 16896 52498
rect 16856 52148 16908 52154
rect 16856 52090 16908 52096
rect 16672 52080 16724 52086
rect 16672 52022 16724 52028
rect 16396 51468 16448 51474
rect 16396 51410 16448 51416
rect 16684 50946 16712 52022
rect 16764 51944 16816 51950
rect 16764 51886 16816 51892
rect 16776 51474 16804 51886
rect 16764 51468 16816 51474
rect 16764 51410 16816 51416
rect 16500 50918 16712 50946
rect 16396 49972 16448 49978
rect 16396 49914 16448 49920
rect 16212 49846 16264 49852
rect 16302 49872 16358 49881
rect 16302 49807 16358 49816
rect 16304 49768 16356 49774
rect 16304 49710 16356 49716
rect 16212 49700 16264 49706
rect 16212 49642 16264 49648
rect 16120 47456 16172 47462
rect 16120 47398 16172 47404
rect 16224 46458 16252 49642
rect 16316 48686 16344 49710
rect 16304 48680 16356 48686
rect 16304 48622 16356 48628
rect 16304 48272 16356 48278
rect 16304 48214 16356 48220
rect 16316 47802 16344 48214
rect 16304 47796 16356 47802
rect 16304 47738 16356 47744
rect 16408 47666 16436 49914
rect 16500 48278 16528 50918
rect 16580 50856 16632 50862
rect 16632 50804 16712 50810
rect 16580 50798 16712 50804
rect 16592 50782 16712 50798
rect 16580 50720 16632 50726
rect 16580 50662 16632 50668
rect 16592 48550 16620 50662
rect 16684 49910 16712 50782
rect 16672 49904 16724 49910
rect 16672 49846 16724 49852
rect 16670 49736 16726 49745
rect 16670 49671 16726 49680
rect 16684 49366 16712 49671
rect 16764 49632 16816 49638
rect 16764 49574 16816 49580
rect 16672 49360 16724 49366
rect 16672 49302 16724 49308
rect 16776 49298 16804 49574
rect 16764 49292 16816 49298
rect 16764 49234 16816 49240
rect 16672 49224 16724 49230
rect 16670 49192 16672 49201
rect 16724 49192 16726 49201
rect 16670 49127 16726 49136
rect 16684 48754 16712 49127
rect 16672 48748 16724 48754
rect 16672 48690 16724 48696
rect 16672 48612 16724 48618
rect 16672 48554 16724 48560
rect 16580 48544 16632 48550
rect 16580 48486 16632 48492
rect 16684 48498 16712 48554
rect 16776 48498 16804 49234
rect 16488 48272 16540 48278
rect 16488 48214 16540 48220
rect 16396 47660 16448 47666
rect 16396 47602 16448 47608
rect 16488 47524 16540 47530
rect 16488 47466 16540 47472
rect 16394 47152 16450 47161
rect 16394 47087 16450 47096
rect 16302 47016 16358 47025
rect 16302 46951 16358 46960
rect 16132 46430 16252 46458
rect 16132 44962 16160 46430
rect 16212 46368 16264 46374
rect 16212 46310 16264 46316
rect 16224 45082 16252 46310
rect 16212 45076 16264 45082
rect 16212 45018 16264 45024
rect 16132 44934 16252 44962
rect 16028 43852 16080 43858
rect 16028 43794 16080 43800
rect 15936 43648 15988 43654
rect 15936 43590 15988 43596
rect 15842 43480 15898 43489
rect 15842 43415 15898 43424
rect 15948 43246 15976 43590
rect 16040 43450 16068 43794
rect 16120 43784 16172 43790
rect 16120 43726 16172 43732
rect 16028 43444 16080 43450
rect 16028 43386 16080 43392
rect 15936 43240 15988 43246
rect 15856 43188 15936 43194
rect 15856 43182 15988 43188
rect 15856 43166 15976 43182
rect 15856 42158 15884 43166
rect 16040 42809 16068 43386
rect 16026 42800 16082 42809
rect 15936 42764 15988 42770
rect 16026 42735 16082 42744
rect 15936 42706 15988 42712
rect 15948 42566 15976 42706
rect 15936 42560 15988 42566
rect 15936 42502 15988 42508
rect 16028 42560 16080 42566
rect 16028 42502 16080 42508
rect 15948 42401 15976 42502
rect 15934 42392 15990 42401
rect 15934 42327 15990 42336
rect 15936 42288 15988 42294
rect 15936 42230 15988 42236
rect 15844 42152 15896 42158
rect 15844 42094 15896 42100
rect 15752 42084 15804 42090
rect 15752 42026 15804 42032
rect 15764 41750 15792 42026
rect 15844 41812 15896 41818
rect 15844 41754 15896 41760
rect 15752 41744 15804 41750
rect 15750 41712 15752 41721
rect 15804 41712 15806 41721
rect 15750 41647 15806 41656
rect 15752 41608 15804 41614
rect 15752 41550 15804 41556
rect 15660 41200 15712 41206
rect 15660 41142 15712 41148
rect 15660 40928 15712 40934
rect 15660 40870 15712 40876
rect 15672 39506 15700 40870
rect 15660 39500 15712 39506
rect 15660 39442 15712 39448
rect 15658 39264 15714 39273
rect 15658 39199 15714 39208
rect 15568 38412 15620 38418
rect 15568 38354 15620 38360
rect 15580 38010 15608 38354
rect 15672 38282 15700 39199
rect 15660 38276 15712 38282
rect 15660 38218 15712 38224
rect 15764 38162 15792 41550
rect 15856 40594 15884 41754
rect 15948 41682 15976 42230
rect 15936 41676 15988 41682
rect 15936 41618 15988 41624
rect 15936 41540 15988 41546
rect 15936 41482 15988 41488
rect 15948 41070 15976 41482
rect 15936 41064 15988 41070
rect 15936 41006 15988 41012
rect 15844 40588 15896 40594
rect 15844 40530 15896 40536
rect 15856 39914 15884 40530
rect 15936 40180 15988 40186
rect 15936 40122 15988 40128
rect 15844 39908 15896 39914
rect 15844 39850 15896 39856
rect 15948 39794 15976 40122
rect 15856 39766 15976 39794
rect 15856 38554 15884 39766
rect 15934 39536 15990 39545
rect 15934 39471 15936 39480
rect 15988 39471 15990 39480
rect 15936 39442 15988 39448
rect 15948 38826 15976 39442
rect 15936 38820 15988 38826
rect 15936 38762 15988 38768
rect 15844 38548 15896 38554
rect 15844 38490 15896 38496
rect 15764 38134 15884 38162
rect 15568 38004 15620 38010
rect 15568 37946 15620 37952
rect 15856 37924 15884 38134
rect 15764 37896 15884 37924
rect 15568 37800 15620 37806
rect 15568 37742 15620 37748
rect 15580 37330 15608 37742
rect 15660 37732 15712 37738
rect 15660 37674 15712 37680
rect 15672 37330 15700 37674
rect 15568 37324 15620 37330
rect 15568 37266 15620 37272
rect 15660 37324 15712 37330
rect 15660 37266 15712 37272
rect 15580 34746 15608 37266
rect 15672 35834 15700 37266
rect 15660 35828 15712 35834
rect 15660 35770 15712 35776
rect 15658 35728 15714 35737
rect 15658 35663 15714 35672
rect 15568 34740 15620 34746
rect 15568 34682 15620 34688
rect 15566 34504 15622 34513
rect 15566 34439 15622 34448
rect 15580 33658 15608 34439
rect 15672 34202 15700 35663
rect 15660 34196 15712 34202
rect 15660 34138 15712 34144
rect 15568 33652 15620 33658
rect 15568 33594 15620 33600
rect 15580 33561 15608 33594
rect 15566 33552 15622 33561
rect 15566 33487 15622 33496
rect 15580 33454 15608 33487
rect 15568 33448 15620 33454
rect 15568 33390 15620 33396
rect 15764 32978 15792 37896
rect 15948 37806 15976 38762
rect 15936 37800 15988 37806
rect 15936 37742 15988 37748
rect 15936 37664 15988 37670
rect 15936 37606 15988 37612
rect 15948 37398 15976 37606
rect 15936 37392 15988 37398
rect 15936 37334 15988 37340
rect 15936 37256 15988 37262
rect 15936 37198 15988 37204
rect 15844 36712 15896 36718
rect 15844 36654 15896 36660
rect 15856 35834 15884 36654
rect 15844 35828 15896 35834
rect 15844 35770 15896 35776
rect 15856 35630 15884 35770
rect 15844 35624 15896 35630
rect 15844 35566 15896 35572
rect 15948 35562 15976 37198
rect 15936 35556 15988 35562
rect 15936 35498 15988 35504
rect 15936 34944 15988 34950
rect 15936 34886 15988 34892
rect 15844 34060 15896 34066
rect 15844 34002 15896 34008
rect 15856 33658 15884 34002
rect 15844 33652 15896 33658
rect 15844 33594 15896 33600
rect 15856 33114 15884 33594
rect 15948 33318 15976 34886
rect 15936 33312 15988 33318
rect 15936 33254 15988 33260
rect 15844 33108 15896 33114
rect 15844 33050 15896 33056
rect 15752 32972 15804 32978
rect 15752 32914 15804 32920
rect 15764 32570 15792 32914
rect 15936 32836 15988 32842
rect 15936 32778 15988 32784
rect 15752 32564 15804 32570
rect 15672 32524 15752 32552
rect 15568 32224 15620 32230
rect 15568 32166 15620 32172
rect 15476 32020 15528 32026
rect 15476 31962 15528 31968
rect 15396 31878 15516 31906
rect 15292 31340 15344 31346
rect 15292 31282 15344 31288
rect 15384 31272 15436 31278
rect 15290 31240 15346 31249
rect 15384 31214 15436 31220
rect 15290 31175 15346 31184
rect 15200 30592 15252 30598
rect 15120 30540 15200 30546
rect 15120 30534 15252 30540
rect 15120 30518 15240 30534
rect 15120 30326 15148 30518
rect 15108 30320 15160 30326
rect 15108 30262 15160 30268
rect 15200 30184 15252 30190
rect 15120 30132 15200 30138
rect 15120 30126 15252 30132
rect 15120 30110 15240 30126
rect 15120 28694 15148 30110
rect 15304 29850 15332 31175
rect 15396 30666 15424 31214
rect 15488 30818 15516 31878
rect 15580 30938 15608 32166
rect 15568 30932 15620 30938
rect 15568 30874 15620 30880
rect 15488 30790 15608 30818
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 15384 30660 15436 30666
rect 15384 30602 15436 30608
rect 15488 30394 15516 30670
rect 15476 30388 15528 30394
rect 15476 30330 15528 30336
rect 15292 29844 15344 29850
rect 15292 29786 15344 29792
rect 15304 29730 15332 29786
rect 15304 29702 15424 29730
rect 15396 29102 15424 29702
rect 15384 29096 15436 29102
rect 15384 29038 15436 29044
rect 15108 28688 15160 28694
rect 15108 28630 15160 28636
rect 15384 28008 15436 28014
rect 15384 27950 15436 27956
rect 15396 27674 15424 27950
rect 15384 27668 15436 27674
rect 15384 27610 15436 27616
rect 15016 27532 15068 27538
rect 15016 27474 15068 27480
rect 15016 26852 15068 26858
rect 15016 26794 15068 26800
rect 14832 24744 14884 24750
rect 14752 24692 14832 24698
rect 14752 24686 14884 24692
rect 14752 24670 14872 24686
rect 14646 23760 14702 23769
rect 14646 23695 14702 23704
rect 14096 23656 14148 23662
rect 14096 23598 14148 23604
rect 13912 23180 13964 23186
rect 13912 23122 13964 23128
rect 13818 22808 13874 22817
rect 13818 22743 13874 22752
rect 13648 22358 13768 22386
rect 13648 21962 13676 22358
rect 13636 21956 13688 21962
rect 13636 21898 13688 21904
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13556 19145 13584 19246
rect 13542 19136 13598 19145
rect 13542 19071 13598 19080
rect 13648 18850 13676 21898
rect 13832 21486 13860 22743
rect 13924 21894 13952 23122
rect 13912 21888 13964 21894
rect 13912 21830 13964 21836
rect 13820 21480 13872 21486
rect 13820 21422 13872 21428
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13740 20806 13768 21286
rect 13832 21146 13860 21422
rect 13820 21140 13872 21146
rect 13820 21082 13872 21088
rect 13728 20800 13780 20806
rect 13728 20742 13780 20748
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13832 19961 13860 20198
rect 13818 19952 13874 19961
rect 13818 19887 13874 19896
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 13740 19514 13768 19790
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 13832 19446 13860 19654
rect 13820 19440 13872 19446
rect 13820 19382 13872 19388
rect 13556 18822 13676 18850
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13360 17264 13412 17270
rect 13360 17206 13412 17212
rect 13372 16794 13400 17206
rect 13360 16788 13412 16794
rect 13360 16730 13412 16736
rect 13372 16658 13400 16730
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13372 16250 13400 16594
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13360 16244 13412 16250
rect 13360 16186 13412 16192
rect 13464 15366 13492 16390
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13188 13960 13308 13988
rect 13188 13530 13216 13960
rect 13372 13870 13400 14554
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 13096 12102 13124 12718
rect 13280 12306 13308 13806
rect 13464 13716 13492 15302
rect 13372 13688 13492 13716
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 13280 11898 13308 12242
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13280 10606 13308 11834
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 12990 10432 13046 10441
rect 12990 10367 13046 10376
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12912 9722 12940 10066
rect 12900 9716 12952 9722
rect 12900 9658 12952 9664
rect 13280 9518 13308 10542
rect 13372 10198 13400 13688
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13464 12782 13492 13262
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13556 12238 13584 18822
rect 13832 18358 13860 19382
rect 13636 18352 13688 18358
rect 13634 18320 13636 18329
rect 13820 18352 13872 18358
rect 13688 18320 13690 18329
rect 13820 18294 13872 18300
rect 13634 18255 13690 18264
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 13648 15042 13676 17478
rect 13740 16998 13768 17614
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13740 16114 13768 16934
rect 13820 16516 13872 16522
rect 13820 16458 13872 16464
rect 13728 16108 13780 16114
rect 13728 16050 13780 16056
rect 13832 15570 13860 16458
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13832 15450 13860 15506
rect 13740 15422 13860 15450
rect 13740 15162 13768 15422
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13648 15014 13860 15042
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13740 13376 13768 14894
rect 13832 14482 13860 15014
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13832 13977 13860 14214
rect 13818 13968 13874 13977
rect 13818 13903 13874 13912
rect 13820 13388 13872 13394
rect 13740 13348 13820 13376
rect 13820 13330 13872 13336
rect 13728 13184 13780 13190
rect 13924 13138 13952 21830
rect 14004 18828 14056 18834
rect 14004 18770 14056 18776
rect 14016 17542 14044 18770
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 13780 13132 13952 13138
rect 13728 13126 13952 13132
rect 13740 13110 13952 13126
rect 13726 12744 13782 12753
rect 13726 12679 13728 12688
rect 13780 12679 13782 12688
rect 13728 12650 13780 12656
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13556 11218 13584 12174
rect 13636 11824 13688 11830
rect 13634 11792 13636 11801
rect 13688 11792 13690 11801
rect 13740 11762 13768 12242
rect 13832 12238 13860 13110
rect 14016 13002 14044 17478
rect 14108 16640 14136 23598
rect 14289 23420 14585 23440
rect 14345 23418 14369 23420
rect 14425 23418 14449 23420
rect 14505 23418 14529 23420
rect 14367 23366 14369 23418
rect 14431 23366 14443 23418
rect 14505 23366 14507 23418
rect 14345 23364 14369 23366
rect 14425 23364 14449 23366
rect 14505 23364 14529 23366
rect 14289 23344 14585 23364
rect 14556 23180 14608 23186
rect 14556 23122 14608 23128
rect 14568 22642 14596 23122
rect 14556 22636 14608 22642
rect 14556 22578 14608 22584
rect 14568 22522 14596 22578
rect 14568 22494 14688 22522
rect 14289 22332 14585 22352
rect 14345 22330 14369 22332
rect 14425 22330 14449 22332
rect 14505 22330 14529 22332
rect 14367 22278 14369 22330
rect 14431 22278 14443 22330
rect 14505 22278 14507 22330
rect 14345 22276 14369 22278
rect 14425 22276 14449 22278
rect 14505 22276 14529 22278
rect 14289 22256 14585 22276
rect 14660 22234 14688 22494
rect 14648 22228 14700 22234
rect 14648 22170 14700 22176
rect 14370 22128 14426 22137
rect 14370 22063 14426 22072
rect 14188 21616 14240 21622
rect 14188 21558 14240 21564
rect 14200 21146 14228 21558
rect 14384 21554 14412 22063
rect 14660 21554 14688 22170
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 14752 21486 14780 24670
rect 15028 23633 15056 26794
rect 15108 26376 15160 26382
rect 15108 26318 15160 26324
rect 15120 24954 15148 26318
rect 15476 26036 15528 26042
rect 15476 25978 15528 25984
rect 15292 25492 15344 25498
rect 15292 25434 15344 25440
rect 15200 25356 15252 25362
rect 15200 25298 15252 25304
rect 15108 24948 15160 24954
rect 15108 24890 15160 24896
rect 15212 24886 15240 25298
rect 15200 24880 15252 24886
rect 15200 24822 15252 24828
rect 15108 24200 15160 24206
rect 15160 24148 15240 24154
rect 15108 24142 15240 24148
rect 15120 24126 15240 24142
rect 15108 23656 15160 23662
rect 15014 23624 15070 23633
rect 15212 23610 15240 24126
rect 15160 23604 15240 23610
rect 15108 23598 15240 23604
rect 15120 23582 15240 23598
rect 15014 23559 15070 23568
rect 15028 23254 15056 23559
rect 14924 23248 14976 23254
rect 14924 23190 14976 23196
rect 15016 23248 15068 23254
rect 15016 23190 15068 23196
rect 14832 22772 14884 22778
rect 14832 22714 14884 22720
rect 14740 21480 14792 21486
rect 14740 21422 14792 21428
rect 14289 21244 14585 21264
rect 14345 21242 14369 21244
rect 14425 21242 14449 21244
rect 14505 21242 14529 21244
rect 14367 21190 14369 21242
rect 14431 21190 14443 21242
rect 14505 21190 14507 21242
rect 14345 21188 14369 21190
rect 14425 21188 14449 21190
rect 14505 21188 14529 21190
rect 14289 21168 14585 21188
rect 14188 21140 14240 21146
rect 14188 21082 14240 21088
rect 14844 20602 14872 22714
rect 14936 22710 14964 23190
rect 14924 22704 14976 22710
rect 14924 22646 14976 22652
rect 15212 22642 15240 23582
rect 15200 22636 15252 22642
rect 15200 22578 15252 22584
rect 15198 22536 15254 22545
rect 15198 22471 15254 22480
rect 15016 22092 15068 22098
rect 15016 22034 15068 22040
rect 14924 22024 14976 22030
rect 14924 21966 14976 21972
rect 14936 21350 14964 21966
rect 15028 21690 15056 22034
rect 15016 21684 15068 21690
rect 15016 21626 15068 21632
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 14924 21344 14976 21350
rect 14924 21286 14976 21292
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 14936 20482 14964 21286
rect 14844 20454 14964 20482
rect 14289 20156 14585 20176
rect 14345 20154 14369 20156
rect 14425 20154 14449 20156
rect 14505 20154 14529 20156
rect 14367 20102 14369 20154
rect 14431 20102 14443 20154
rect 14505 20102 14507 20154
rect 14345 20100 14369 20102
rect 14425 20100 14449 20102
rect 14505 20100 14529 20102
rect 14289 20080 14585 20100
rect 14738 19816 14794 19825
rect 14738 19751 14740 19760
rect 14792 19751 14794 19760
rect 14740 19722 14792 19728
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 14200 19281 14228 19654
rect 14186 19272 14242 19281
rect 14186 19207 14242 19216
rect 14740 19236 14792 19242
rect 14200 18850 14228 19207
rect 14740 19178 14792 19184
rect 14289 19068 14585 19088
rect 14345 19066 14369 19068
rect 14425 19066 14449 19068
rect 14505 19066 14529 19068
rect 14367 19014 14369 19066
rect 14431 19014 14443 19066
rect 14505 19014 14507 19066
rect 14345 19012 14369 19014
rect 14425 19012 14449 19014
rect 14505 19012 14529 19014
rect 14289 18992 14585 19012
rect 14200 18834 14320 18850
rect 14200 18828 14332 18834
rect 14200 18822 14280 18828
rect 14280 18770 14332 18776
rect 14752 18766 14780 19178
rect 14740 18760 14792 18766
rect 14740 18702 14792 18708
rect 14646 18456 14702 18465
rect 14646 18391 14648 18400
rect 14700 18391 14702 18400
rect 14648 18362 14700 18368
rect 14752 18222 14780 18702
rect 14740 18216 14792 18222
rect 14568 18154 14688 18170
rect 14740 18158 14792 18164
rect 14556 18148 14688 18154
rect 14608 18142 14688 18148
rect 14556 18090 14608 18096
rect 14289 17980 14585 18000
rect 14345 17978 14369 17980
rect 14425 17978 14449 17980
rect 14505 17978 14529 17980
rect 14367 17926 14369 17978
rect 14431 17926 14443 17978
rect 14505 17926 14507 17978
rect 14345 17924 14369 17926
rect 14425 17924 14449 17926
rect 14505 17924 14529 17926
rect 14289 17904 14585 17924
rect 14372 17740 14424 17746
rect 14372 17682 14424 17688
rect 14384 17066 14412 17682
rect 14372 17060 14424 17066
rect 14372 17002 14424 17008
rect 14289 16892 14585 16912
rect 14345 16890 14369 16892
rect 14425 16890 14449 16892
rect 14505 16890 14529 16892
rect 14367 16838 14369 16890
rect 14431 16838 14443 16890
rect 14505 16838 14507 16890
rect 14345 16836 14369 16838
rect 14425 16836 14449 16838
rect 14505 16836 14529 16838
rect 14289 16816 14585 16836
rect 14188 16652 14240 16658
rect 14108 16612 14188 16640
rect 14188 16594 14240 16600
rect 14200 16250 14228 16594
rect 14188 16244 14240 16250
rect 13924 12974 14044 13002
rect 14108 16204 14188 16232
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13634 11727 13690 11736
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13556 10810 13584 11154
rect 13740 11014 13768 11698
rect 13832 11694 13860 12174
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 13740 10538 13768 10950
rect 13924 10674 13952 12974
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 14016 11558 14044 12174
rect 14004 11552 14056 11558
rect 14004 11494 14056 11500
rect 14016 11234 14044 11494
rect 14108 11354 14136 16204
rect 14188 16186 14240 16192
rect 14289 15804 14585 15824
rect 14345 15802 14369 15804
rect 14425 15802 14449 15804
rect 14505 15802 14529 15804
rect 14367 15750 14369 15802
rect 14431 15750 14443 15802
rect 14505 15750 14507 15802
rect 14345 15748 14369 15750
rect 14425 15748 14449 15750
rect 14505 15748 14529 15750
rect 14289 15728 14585 15748
rect 14280 15428 14332 15434
rect 14280 15370 14332 15376
rect 14292 15337 14320 15370
rect 14278 15328 14334 15337
rect 14278 15263 14334 15272
rect 14289 14716 14585 14736
rect 14345 14714 14369 14716
rect 14425 14714 14449 14716
rect 14505 14714 14529 14716
rect 14367 14662 14369 14714
rect 14431 14662 14443 14714
rect 14505 14662 14507 14714
rect 14345 14660 14369 14662
rect 14425 14660 14449 14662
rect 14505 14660 14529 14662
rect 14289 14640 14585 14660
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14476 14006 14504 14418
rect 14568 14074 14596 14418
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14464 14000 14516 14006
rect 14464 13942 14516 13948
rect 14289 13628 14585 13648
rect 14345 13626 14369 13628
rect 14425 13626 14449 13628
rect 14505 13626 14529 13628
rect 14367 13574 14369 13626
rect 14431 13574 14443 13626
rect 14505 13574 14507 13626
rect 14345 13572 14369 13574
rect 14425 13572 14449 13574
rect 14505 13572 14529 13574
rect 14289 13552 14585 13572
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14200 12345 14228 13194
rect 14384 12986 14412 13330
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14289 12540 14585 12560
rect 14345 12538 14369 12540
rect 14425 12538 14449 12540
rect 14505 12538 14529 12540
rect 14367 12486 14369 12538
rect 14431 12486 14443 12538
rect 14505 12486 14507 12538
rect 14345 12484 14369 12486
rect 14425 12484 14449 12486
rect 14505 12484 14529 12486
rect 14289 12464 14585 12484
rect 14186 12336 14242 12345
rect 14186 12271 14188 12280
rect 14240 12271 14242 12280
rect 14188 12242 14240 12248
rect 14200 12211 14228 12242
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 11937 14228 12038
rect 14186 11928 14242 11937
rect 14186 11863 14242 11872
rect 14200 11694 14228 11863
rect 14188 11688 14240 11694
rect 14280 11688 14332 11694
rect 14188 11630 14240 11636
rect 14278 11656 14280 11665
rect 14332 11656 14334 11665
rect 14278 11591 14334 11600
rect 14289 11452 14585 11472
rect 14345 11450 14369 11452
rect 14425 11450 14449 11452
rect 14505 11450 14529 11452
rect 14367 11398 14369 11450
rect 14431 11398 14443 11450
rect 14505 11398 14507 11450
rect 14345 11396 14369 11398
rect 14425 11396 14449 11398
rect 14505 11396 14529 11398
rect 14289 11376 14585 11396
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 14016 11206 14136 11234
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 13820 10600 13872 10606
rect 13818 10568 13820 10577
rect 13872 10568 13874 10577
rect 13728 10532 13780 10538
rect 13818 10503 13874 10512
rect 13728 10474 13780 10480
rect 13360 10192 13412 10198
rect 13360 10134 13412 10140
rect 13740 10146 13768 10474
rect 13832 10266 13860 10503
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13740 10118 13860 10146
rect 13832 9926 13860 10118
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13268 9512 13320 9518
rect 13174 9480 13230 9489
rect 13268 9454 13320 9460
rect 13832 9450 13860 9862
rect 13174 9415 13230 9424
rect 13820 9444 13872 9450
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 13004 8945 13032 8978
rect 12990 8936 13046 8945
rect 13188 8906 13216 9415
rect 13820 9386 13872 9392
rect 13832 9178 13860 9386
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13924 9042 13952 10610
rect 14108 10606 14136 11206
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 14016 9625 14044 10066
rect 14108 9994 14136 10542
rect 14096 9988 14148 9994
rect 14096 9930 14148 9936
rect 14002 9616 14058 9625
rect 14002 9551 14058 9560
rect 14096 9512 14148 9518
rect 14200 9489 14228 11086
rect 14289 10364 14585 10384
rect 14345 10362 14369 10364
rect 14425 10362 14449 10364
rect 14505 10362 14529 10364
rect 14367 10310 14369 10362
rect 14431 10310 14443 10362
rect 14505 10310 14507 10362
rect 14345 10308 14369 10310
rect 14425 10308 14449 10310
rect 14505 10308 14529 10310
rect 14289 10288 14585 10308
rect 14096 9454 14148 9460
rect 14186 9480 14242 9489
rect 14108 9178 14136 9454
rect 14186 9415 14242 9424
rect 14289 9276 14585 9296
rect 14345 9274 14369 9276
rect 14425 9274 14449 9276
rect 14505 9274 14529 9276
rect 14367 9222 14369 9274
rect 14431 9222 14443 9274
rect 14505 9222 14507 9274
rect 14345 9220 14369 9222
rect 14425 9220 14449 9222
rect 14505 9220 14529 9222
rect 14289 9200 14585 9220
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 12990 8871 13046 8880
rect 13176 8900 13228 8906
rect 13004 8566 13032 8871
rect 13176 8842 13228 8848
rect 13280 8634 13308 8978
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 12992 8560 13044 8566
rect 12992 8502 13044 8508
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 12808 8016 12860 8022
rect 12808 7958 12860 7964
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12728 7002 12756 7822
rect 12820 7546 12848 7958
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 13188 6882 13216 7346
rect 13372 7342 13400 8298
rect 13820 7812 13872 7818
rect 13820 7754 13872 7760
rect 13832 7342 13860 7754
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13372 7002 13400 7278
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13268 6928 13320 6934
rect 13188 6876 13268 6882
rect 13188 6870 13320 6876
rect 13188 6854 13308 6870
rect 13188 6458 13216 6854
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13188 5846 13216 6394
rect 13636 6384 13688 6390
rect 13634 6352 13636 6361
rect 13688 6352 13690 6361
rect 13634 6287 13690 6296
rect 13268 6180 13320 6186
rect 13268 6122 13320 6128
rect 13280 5914 13308 6122
rect 13832 5914 13860 6666
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13176 5840 13228 5846
rect 13176 5782 13228 5788
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12544 5370 12572 5714
rect 13280 5370 13308 5850
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 13268 5364 13320 5370
rect 13268 5306 13320 5312
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 12544 5114 12572 5306
rect 13924 5166 13952 6734
rect 14016 6254 14044 8570
rect 14186 8392 14242 8401
rect 14186 8327 14242 8336
rect 14200 7954 14228 8327
rect 14289 8188 14585 8208
rect 14345 8186 14369 8188
rect 14425 8186 14449 8188
rect 14505 8186 14529 8188
rect 14367 8134 14369 8186
rect 14431 8134 14443 8186
rect 14505 8134 14507 8186
rect 14345 8132 14369 8134
rect 14425 8132 14449 8134
rect 14505 8132 14529 8134
rect 14289 8112 14585 8132
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14200 6458 14228 7890
rect 14289 7100 14585 7120
rect 14345 7098 14369 7100
rect 14425 7098 14449 7100
rect 14505 7098 14529 7100
rect 14367 7046 14369 7098
rect 14431 7046 14443 7098
rect 14505 7046 14507 7098
rect 14345 7044 14369 7046
rect 14425 7044 14449 7046
rect 14505 7044 14529 7046
rect 14289 7024 14585 7044
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14660 6322 14688 18142
rect 14752 17610 14780 18158
rect 14740 17604 14792 17610
rect 14740 17546 14792 17552
rect 14752 17202 14780 17546
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 14740 17060 14792 17066
rect 14740 17002 14792 17008
rect 14752 14414 14780 17002
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14752 12102 14780 13262
rect 14844 12186 14872 20454
rect 15028 20346 15056 21490
rect 15212 21457 15240 22471
rect 15304 21622 15332 25434
rect 15488 23168 15516 25978
rect 15580 25945 15608 30790
rect 15566 25936 15622 25945
rect 15672 25922 15700 32524
rect 15752 32506 15804 32512
rect 15752 32020 15804 32026
rect 15752 31962 15804 31968
rect 15764 30870 15792 31962
rect 15844 31952 15896 31958
rect 15844 31894 15896 31900
rect 15856 31346 15884 31894
rect 15948 31822 15976 32778
rect 15936 31816 15988 31822
rect 15936 31758 15988 31764
rect 15948 31482 15976 31758
rect 15936 31476 15988 31482
rect 15936 31418 15988 31424
rect 15844 31340 15896 31346
rect 15844 31282 15896 31288
rect 15844 31204 15896 31210
rect 15844 31146 15896 31152
rect 15752 30864 15804 30870
rect 15752 30806 15804 30812
rect 15856 30410 15884 31146
rect 15948 30734 15976 31418
rect 15936 30728 15988 30734
rect 15936 30670 15988 30676
rect 15764 30382 15884 30410
rect 15764 26246 15792 30382
rect 15948 30326 15976 30670
rect 15844 30320 15896 30326
rect 15842 30288 15844 30297
rect 15936 30320 15988 30326
rect 15896 30288 15898 30297
rect 15936 30262 15988 30268
rect 15842 30223 15898 30232
rect 15948 29646 15976 30262
rect 16040 29850 16068 42502
rect 16132 37262 16160 43726
rect 16224 40633 16252 44934
rect 16316 41177 16344 46951
rect 16408 45948 16436 47087
rect 16500 46050 16528 47466
rect 16592 46170 16620 48486
rect 16684 48470 16804 48498
rect 16580 46164 16632 46170
rect 16580 46106 16632 46112
rect 16500 46034 16620 46050
rect 16500 46028 16632 46034
rect 16500 46022 16580 46028
rect 16580 45970 16632 45976
rect 16408 45920 16528 45948
rect 16396 44260 16448 44266
rect 16396 44202 16448 44208
rect 16408 43858 16436 44202
rect 16396 43852 16448 43858
rect 16396 43794 16448 43800
rect 16394 43752 16450 43761
rect 16394 43687 16450 43696
rect 16408 42809 16436 43687
rect 16394 42800 16450 42809
rect 16394 42735 16450 42744
rect 16396 42560 16448 42566
rect 16396 42502 16448 42508
rect 16408 42158 16436 42502
rect 16396 42152 16448 42158
rect 16396 42094 16448 42100
rect 16408 41682 16436 42094
rect 16396 41676 16448 41682
rect 16396 41618 16448 41624
rect 16394 41576 16450 41585
rect 16394 41511 16450 41520
rect 16408 41274 16436 41511
rect 16396 41268 16448 41274
rect 16396 41210 16448 41216
rect 16302 41168 16358 41177
rect 16302 41103 16358 41112
rect 16396 41132 16448 41138
rect 16396 41074 16448 41080
rect 16304 40996 16356 41002
rect 16304 40938 16356 40944
rect 16210 40624 16266 40633
rect 16210 40559 16266 40568
rect 16316 40390 16344 40938
rect 16304 40384 16356 40390
rect 16304 40326 16356 40332
rect 16316 39982 16344 40326
rect 16304 39976 16356 39982
rect 16304 39918 16356 39924
rect 16302 39536 16358 39545
rect 16302 39471 16304 39480
rect 16356 39471 16358 39480
rect 16304 39442 16356 39448
rect 16212 39024 16264 39030
rect 16212 38966 16264 38972
rect 16120 37256 16172 37262
rect 16120 37198 16172 37204
rect 16132 36582 16160 37198
rect 16120 36576 16172 36582
rect 16120 36518 16172 36524
rect 16132 31278 16160 36518
rect 16224 35154 16252 38966
rect 16304 38888 16356 38894
rect 16304 38830 16356 38836
rect 16316 38350 16344 38830
rect 16304 38344 16356 38350
rect 16304 38286 16356 38292
rect 16316 37738 16344 38286
rect 16304 37732 16356 37738
rect 16304 37674 16356 37680
rect 16408 36938 16436 41074
rect 16500 39953 16528 45920
rect 16592 45490 16620 45970
rect 16580 45484 16632 45490
rect 16580 45426 16632 45432
rect 16672 44940 16724 44946
rect 16672 44882 16724 44888
rect 16684 44470 16712 44882
rect 16672 44464 16724 44470
rect 16672 44406 16724 44412
rect 16580 44192 16632 44198
rect 16580 44134 16632 44140
rect 16486 39944 16542 39953
rect 16486 39879 16542 39888
rect 16488 39092 16540 39098
rect 16488 39034 16540 39040
rect 16500 38894 16528 39034
rect 16488 38888 16540 38894
rect 16488 38830 16540 38836
rect 16500 38010 16528 38830
rect 16488 38004 16540 38010
rect 16488 37946 16540 37952
rect 16500 37806 16528 37946
rect 16488 37800 16540 37806
rect 16488 37742 16540 37748
rect 16316 36910 16436 36938
rect 16212 35148 16264 35154
rect 16212 35090 16264 35096
rect 16224 34746 16252 35090
rect 16316 35086 16344 36910
rect 16488 36848 16540 36854
rect 16488 36790 16540 36796
rect 16396 36780 16448 36786
rect 16396 36722 16448 36728
rect 16408 36378 16436 36722
rect 16500 36530 16528 36790
rect 16592 36650 16620 44134
rect 16672 43240 16724 43246
rect 16672 43182 16724 43188
rect 16684 42906 16712 43182
rect 16672 42900 16724 42906
rect 16672 42842 16724 42848
rect 16684 42634 16712 42842
rect 16672 42628 16724 42634
rect 16672 42570 16724 42576
rect 16776 42514 16804 48470
rect 16868 47122 16896 52090
rect 16856 47116 16908 47122
rect 16856 47058 16908 47064
rect 16960 47025 16988 54538
rect 17144 53990 17172 54606
rect 17132 53984 17184 53990
rect 17132 53926 17184 53932
rect 17040 53440 17092 53446
rect 17040 53382 17092 53388
rect 17052 53242 17080 53382
rect 17040 53236 17092 53242
rect 17040 53178 17092 53184
rect 17052 51542 17080 53178
rect 17144 52426 17172 53926
rect 17420 53417 17448 55218
rect 18144 55208 18196 55214
rect 18144 55150 18196 55156
rect 17622 54428 17918 54448
rect 17678 54426 17702 54428
rect 17758 54426 17782 54428
rect 17838 54426 17862 54428
rect 17700 54374 17702 54426
rect 17764 54374 17776 54426
rect 17838 54374 17840 54426
rect 17678 54372 17702 54374
rect 17758 54372 17782 54374
rect 17838 54372 17862 54374
rect 17622 54352 17918 54372
rect 17406 53408 17462 53417
rect 17406 53343 17462 53352
rect 17622 53340 17918 53360
rect 17678 53338 17702 53340
rect 17758 53338 17782 53340
rect 17838 53338 17862 53340
rect 17700 53286 17702 53338
rect 17764 53286 17776 53338
rect 17838 53286 17840 53338
rect 17678 53284 17702 53286
rect 17758 53284 17782 53286
rect 17838 53284 17862 53286
rect 17622 53264 17918 53284
rect 17960 53032 18012 53038
rect 17958 53000 17960 53009
rect 18012 53000 18014 53009
rect 17958 52935 18014 52944
rect 17960 52896 18012 52902
rect 17960 52838 18012 52844
rect 17132 52420 17184 52426
rect 17132 52362 17184 52368
rect 17144 51610 17172 52362
rect 17622 52252 17918 52272
rect 17678 52250 17702 52252
rect 17758 52250 17782 52252
rect 17838 52250 17862 52252
rect 17700 52198 17702 52250
rect 17764 52198 17776 52250
rect 17838 52198 17840 52250
rect 17678 52196 17702 52198
rect 17758 52196 17782 52198
rect 17838 52196 17862 52198
rect 17622 52176 17918 52196
rect 17972 52154 18000 52838
rect 17960 52148 18012 52154
rect 17960 52090 18012 52096
rect 17498 51912 17554 51921
rect 17408 51876 17460 51882
rect 17498 51847 17554 51856
rect 17408 51818 17460 51824
rect 17132 51604 17184 51610
rect 17132 51546 17184 51552
rect 17040 51536 17092 51542
rect 17040 51478 17092 51484
rect 17040 50992 17092 50998
rect 17040 50934 17092 50940
rect 17052 47161 17080 50934
rect 17144 50862 17172 51546
rect 17316 51468 17368 51474
rect 17316 51410 17368 51416
rect 17328 50930 17356 51410
rect 17316 50924 17368 50930
rect 17316 50866 17368 50872
rect 17132 50856 17184 50862
rect 17132 50798 17184 50804
rect 17144 50522 17172 50798
rect 17132 50516 17184 50522
rect 17184 50476 17264 50504
rect 17132 50458 17184 50464
rect 17132 50380 17184 50386
rect 17132 50322 17184 50328
rect 17144 49586 17172 50322
rect 17236 49774 17264 50476
rect 17328 50386 17356 50866
rect 17316 50380 17368 50386
rect 17316 50322 17368 50328
rect 17224 49768 17276 49774
rect 17224 49710 17276 49716
rect 17144 49558 17264 49586
rect 17038 47152 17094 47161
rect 17038 47087 17094 47096
rect 17132 47116 17184 47122
rect 17132 47058 17184 47064
rect 16946 47016 17002 47025
rect 16856 46980 16908 46986
rect 16946 46951 17002 46960
rect 16856 46922 16908 46928
rect 16868 45472 16896 46922
rect 17040 46504 17092 46510
rect 17040 46446 17092 46452
rect 16868 45444 16988 45472
rect 16856 45348 16908 45354
rect 16856 45290 16908 45296
rect 16684 42486 16804 42514
rect 16684 41070 16712 42486
rect 16762 41712 16818 41721
rect 16762 41647 16764 41656
rect 16816 41647 16818 41656
rect 16764 41618 16816 41624
rect 16672 41064 16724 41070
rect 16672 41006 16724 41012
rect 16580 36644 16632 36650
rect 16580 36586 16632 36592
rect 16500 36502 16620 36530
rect 16592 36378 16620 36502
rect 16396 36372 16448 36378
rect 16396 36314 16448 36320
rect 16580 36372 16632 36378
rect 16580 36314 16632 36320
rect 16488 36304 16540 36310
rect 16488 36246 16540 36252
rect 16396 36168 16448 36174
rect 16396 36110 16448 36116
rect 16304 35080 16356 35086
rect 16304 35022 16356 35028
rect 16316 34746 16344 35022
rect 16408 35018 16436 36110
rect 16500 35834 16528 36246
rect 16580 36032 16632 36038
rect 16580 35974 16632 35980
rect 16488 35828 16540 35834
rect 16488 35770 16540 35776
rect 16592 35630 16620 35974
rect 16580 35624 16632 35630
rect 16580 35566 16632 35572
rect 16488 35148 16540 35154
rect 16488 35090 16540 35096
rect 16396 35012 16448 35018
rect 16396 34954 16448 34960
rect 16212 34740 16264 34746
rect 16212 34682 16264 34688
rect 16304 34740 16356 34746
rect 16304 34682 16356 34688
rect 16224 34626 16252 34682
rect 16224 34598 16436 34626
rect 16304 34128 16356 34134
rect 16304 34070 16356 34076
rect 16212 33992 16264 33998
rect 16212 33934 16264 33940
rect 16224 33318 16252 33934
rect 16212 33312 16264 33318
rect 16212 33254 16264 33260
rect 16120 31272 16172 31278
rect 16120 31214 16172 31220
rect 16120 31136 16172 31142
rect 16120 31078 16172 31084
rect 16132 30190 16160 31078
rect 16120 30184 16172 30190
rect 16120 30126 16172 30132
rect 16028 29844 16080 29850
rect 16028 29786 16080 29792
rect 15936 29640 15988 29646
rect 15936 29582 15988 29588
rect 15948 29306 15976 29582
rect 15936 29300 15988 29306
rect 15936 29242 15988 29248
rect 15844 29028 15896 29034
rect 15844 28970 15896 28976
rect 15856 28064 15884 28970
rect 15948 28218 15976 29242
rect 16040 28762 16068 29786
rect 16224 29594 16252 33254
rect 16316 32910 16344 34070
rect 16304 32904 16356 32910
rect 16304 32846 16356 32852
rect 16304 31884 16356 31890
rect 16304 31826 16356 31832
rect 16316 30938 16344 31826
rect 16304 30932 16356 30938
rect 16304 30874 16356 30880
rect 16316 30394 16344 30874
rect 16304 30388 16356 30394
rect 16304 30330 16356 30336
rect 16316 29714 16344 30330
rect 16304 29708 16356 29714
rect 16304 29650 16356 29656
rect 16132 29566 16252 29594
rect 16028 28756 16080 28762
rect 16028 28698 16080 28704
rect 15936 28212 15988 28218
rect 15936 28154 15988 28160
rect 15856 28036 15976 28064
rect 15844 27940 15896 27946
rect 15844 27882 15896 27888
rect 15752 26240 15804 26246
rect 15752 26182 15804 26188
rect 15764 26042 15792 26182
rect 15752 26036 15804 26042
rect 15752 25978 15804 25984
rect 15672 25894 15792 25922
rect 15566 25871 15622 25880
rect 15660 25832 15712 25838
rect 15660 25774 15712 25780
rect 15568 25356 15620 25362
rect 15568 25298 15620 25304
rect 15580 24954 15608 25298
rect 15672 24993 15700 25774
rect 15764 25362 15792 25894
rect 15752 25356 15804 25362
rect 15752 25298 15804 25304
rect 15658 24984 15714 24993
rect 15568 24948 15620 24954
rect 15658 24919 15714 24928
rect 15568 24890 15620 24896
rect 15658 24848 15714 24857
rect 15764 24818 15792 25298
rect 15658 24783 15714 24792
rect 15752 24812 15804 24818
rect 15672 24750 15700 24783
rect 15752 24754 15804 24760
rect 15660 24744 15712 24750
rect 15660 24686 15712 24692
rect 15856 23662 15884 27882
rect 15948 23798 15976 28036
rect 16028 27396 16080 27402
rect 16028 27338 16080 27344
rect 16040 26790 16068 27338
rect 16028 26784 16080 26790
rect 16028 26726 16080 26732
rect 16040 26042 16068 26726
rect 16028 26036 16080 26042
rect 16028 25978 16080 25984
rect 16132 24993 16160 29566
rect 16212 29504 16264 29510
rect 16212 29446 16264 29452
rect 16224 27606 16252 29446
rect 16316 28694 16344 29650
rect 16304 28688 16356 28694
rect 16304 28630 16356 28636
rect 16304 28552 16356 28558
rect 16304 28494 16356 28500
rect 16316 27985 16344 28494
rect 16302 27976 16358 27985
rect 16302 27911 16304 27920
rect 16356 27911 16358 27920
rect 16304 27882 16356 27888
rect 16316 27674 16344 27882
rect 16304 27668 16356 27674
rect 16304 27610 16356 27616
rect 16212 27600 16264 27606
rect 16212 27542 16264 27548
rect 16224 26586 16252 27542
rect 16212 26580 16264 26586
rect 16212 26522 16264 26528
rect 16408 25650 16436 34598
rect 16500 34066 16528 35090
rect 16488 34060 16540 34066
rect 16488 34002 16540 34008
rect 16592 33402 16620 35566
rect 16500 33374 16620 33402
rect 16500 30666 16528 33374
rect 16580 33312 16632 33318
rect 16580 33254 16632 33260
rect 16592 32230 16620 33254
rect 16580 32224 16632 32230
rect 16580 32166 16632 32172
rect 16592 31278 16620 32166
rect 16580 31272 16632 31278
rect 16580 31214 16632 31220
rect 16488 30660 16540 30666
rect 16488 30602 16540 30608
rect 16592 30598 16620 31214
rect 16580 30592 16632 30598
rect 16580 30534 16632 30540
rect 16592 30190 16620 30534
rect 16580 30184 16632 30190
rect 16580 30126 16632 30132
rect 16592 29510 16620 30126
rect 16580 29504 16632 29510
rect 16500 29464 16580 29492
rect 16500 27402 16528 29464
rect 16580 29446 16632 29452
rect 16580 28960 16632 28966
rect 16580 28902 16632 28908
rect 16592 28762 16620 28902
rect 16580 28756 16632 28762
rect 16580 28698 16632 28704
rect 16684 28694 16712 41006
rect 16776 40882 16804 41618
rect 16868 41206 16896 45290
rect 16960 44538 16988 45444
rect 16948 44532 17000 44538
rect 16948 44474 17000 44480
rect 16948 43852 17000 43858
rect 16948 43794 17000 43800
rect 16960 43314 16988 43794
rect 16948 43308 17000 43314
rect 16948 43250 17000 43256
rect 16960 42158 16988 43250
rect 16948 42152 17000 42158
rect 16948 42094 17000 42100
rect 16960 41818 16988 42094
rect 16948 41812 17000 41818
rect 16948 41754 17000 41760
rect 17052 41449 17080 46446
rect 17144 46374 17172 47058
rect 17236 46481 17264 49558
rect 17316 48748 17368 48754
rect 17316 48690 17368 48696
rect 17328 48346 17356 48690
rect 17316 48340 17368 48346
rect 17316 48282 17368 48288
rect 17316 48204 17368 48210
rect 17316 48146 17368 48152
rect 17328 46714 17356 48146
rect 17316 46708 17368 46714
rect 17316 46650 17368 46656
rect 17222 46472 17278 46481
rect 17222 46407 17278 46416
rect 17132 46368 17184 46374
rect 17184 46316 17264 46322
rect 17132 46310 17264 46316
rect 17144 46294 17264 46310
rect 17132 46164 17184 46170
rect 17132 46106 17184 46112
rect 17038 41440 17094 41449
rect 17038 41375 17094 41384
rect 17038 41304 17094 41313
rect 16948 41268 17000 41274
rect 17038 41239 17094 41248
rect 16948 41210 17000 41216
rect 16856 41200 16908 41206
rect 16856 41142 16908 41148
rect 16776 40854 16896 40882
rect 16764 40724 16816 40730
rect 16764 40666 16816 40672
rect 16776 40066 16804 40666
rect 16868 40458 16896 40854
rect 16856 40452 16908 40458
rect 16856 40394 16908 40400
rect 16776 40038 16896 40066
rect 16868 39982 16896 40038
rect 16764 39976 16816 39982
rect 16764 39918 16816 39924
rect 16856 39976 16908 39982
rect 16856 39918 16908 39924
rect 16776 39438 16804 39918
rect 16868 39506 16896 39918
rect 16960 39794 16988 41210
rect 17052 39930 17080 41239
rect 17144 40168 17172 46106
rect 17236 40361 17264 46294
rect 17328 46170 17356 46650
rect 17316 46164 17368 46170
rect 17316 46106 17368 46112
rect 17328 45354 17356 46106
rect 17316 45348 17368 45354
rect 17316 45290 17368 45296
rect 17316 44328 17368 44334
rect 17316 44270 17368 44276
rect 17328 43110 17356 44270
rect 17316 43104 17368 43110
rect 17316 43046 17368 43052
rect 17316 42220 17368 42226
rect 17316 42162 17368 42168
rect 17328 40934 17356 42162
rect 17420 41426 17448 51818
rect 17512 51610 17540 51847
rect 17500 51604 17552 51610
rect 17500 51546 17552 51552
rect 17512 50862 17540 51546
rect 17622 51164 17918 51184
rect 17678 51162 17702 51164
rect 17758 51162 17782 51164
rect 17838 51162 17862 51164
rect 17700 51110 17702 51162
rect 17764 51110 17776 51162
rect 17838 51110 17840 51162
rect 17678 51108 17702 51110
rect 17758 51108 17782 51110
rect 17838 51108 17862 51110
rect 17622 51088 17918 51108
rect 17500 50856 17552 50862
rect 17500 50798 17552 50804
rect 17512 49774 17540 50798
rect 18052 50720 18104 50726
rect 18052 50662 18104 50668
rect 18064 50250 18092 50662
rect 18052 50244 18104 50250
rect 18052 50186 18104 50192
rect 18156 50153 18184 55150
rect 18142 50144 18198 50153
rect 17622 50076 17918 50096
rect 18142 50079 18198 50088
rect 17678 50074 17702 50076
rect 17758 50074 17782 50076
rect 17838 50074 17862 50076
rect 17700 50022 17702 50074
rect 17764 50022 17776 50074
rect 17838 50022 17840 50074
rect 17678 50020 17702 50022
rect 17758 50020 17782 50022
rect 17838 50020 17862 50022
rect 17622 50000 17918 50020
rect 17500 49768 17552 49774
rect 17500 49710 17552 49716
rect 17512 49434 17540 49710
rect 17500 49428 17552 49434
rect 17500 49370 17552 49376
rect 17500 49292 17552 49298
rect 17500 49234 17552 49240
rect 17512 48770 17540 49234
rect 17622 48988 17918 49008
rect 17678 48986 17702 48988
rect 17758 48986 17782 48988
rect 17838 48986 17862 48988
rect 17700 48934 17702 48986
rect 17764 48934 17776 48986
rect 17838 48934 17840 48986
rect 17678 48932 17702 48934
rect 17758 48932 17782 48934
rect 17838 48932 17862 48934
rect 17622 48912 17918 48932
rect 17512 48754 17632 48770
rect 17500 48748 17632 48754
rect 17552 48742 17632 48748
rect 17500 48690 17552 48696
rect 17500 48612 17552 48618
rect 17500 48554 17552 48560
rect 17512 41546 17540 48554
rect 17604 48278 17632 48742
rect 17592 48272 17644 48278
rect 17592 48214 17644 48220
rect 17622 47900 17918 47920
rect 17678 47898 17702 47900
rect 17758 47898 17782 47900
rect 17838 47898 17862 47900
rect 17700 47846 17702 47898
rect 17764 47846 17776 47898
rect 17838 47846 17840 47898
rect 17678 47844 17702 47846
rect 17758 47844 17782 47846
rect 17838 47844 17862 47846
rect 17622 47824 17918 47844
rect 17960 47660 18012 47666
rect 17960 47602 18012 47608
rect 17622 46812 17918 46832
rect 17678 46810 17702 46812
rect 17758 46810 17782 46812
rect 17838 46810 17862 46812
rect 17700 46758 17702 46810
rect 17764 46758 17776 46810
rect 17838 46758 17840 46810
rect 17678 46756 17702 46758
rect 17758 46756 17782 46758
rect 17838 46756 17862 46758
rect 17622 46736 17918 46756
rect 17622 45724 17918 45744
rect 17678 45722 17702 45724
rect 17758 45722 17782 45724
rect 17838 45722 17862 45724
rect 17700 45670 17702 45722
rect 17764 45670 17776 45722
rect 17838 45670 17840 45722
rect 17678 45668 17702 45670
rect 17758 45668 17782 45670
rect 17838 45668 17862 45670
rect 17622 45648 17918 45668
rect 17592 45416 17644 45422
rect 17592 45358 17644 45364
rect 17604 45082 17632 45358
rect 17592 45076 17644 45082
rect 17592 45018 17644 45024
rect 17622 44636 17918 44656
rect 17678 44634 17702 44636
rect 17758 44634 17782 44636
rect 17838 44634 17862 44636
rect 17700 44582 17702 44634
rect 17764 44582 17776 44634
rect 17838 44582 17840 44634
rect 17678 44580 17702 44582
rect 17758 44580 17782 44582
rect 17838 44580 17862 44582
rect 17622 44560 17918 44580
rect 17592 44328 17644 44334
rect 17592 44270 17644 44276
rect 17604 43926 17632 44270
rect 17592 43920 17644 43926
rect 17592 43862 17644 43868
rect 17622 43548 17918 43568
rect 17678 43546 17702 43548
rect 17758 43546 17782 43548
rect 17838 43546 17862 43548
rect 17700 43494 17702 43546
rect 17764 43494 17776 43546
rect 17838 43494 17840 43546
rect 17678 43492 17702 43494
rect 17758 43492 17782 43494
rect 17838 43492 17862 43494
rect 17622 43472 17918 43492
rect 17622 42460 17918 42480
rect 17678 42458 17702 42460
rect 17758 42458 17782 42460
rect 17838 42458 17862 42460
rect 17700 42406 17702 42458
rect 17764 42406 17776 42458
rect 17838 42406 17840 42458
rect 17678 42404 17702 42406
rect 17758 42404 17782 42406
rect 17838 42404 17862 42406
rect 17622 42384 17918 42404
rect 17776 42288 17828 42294
rect 17776 42230 17828 42236
rect 17788 41857 17816 42230
rect 17972 42226 18000 47602
rect 18144 46436 18196 46442
rect 18144 46378 18196 46384
rect 18052 43104 18104 43110
rect 18052 43046 18104 43052
rect 17960 42220 18012 42226
rect 17960 42162 18012 42168
rect 17958 42120 18014 42129
rect 17958 42055 18014 42064
rect 17774 41848 17830 41857
rect 17774 41783 17830 41792
rect 17500 41540 17552 41546
rect 17500 41482 17552 41488
rect 17420 41398 17540 41426
rect 17408 41200 17460 41206
rect 17408 41142 17460 41148
rect 17316 40928 17368 40934
rect 17316 40870 17368 40876
rect 17316 40384 17368 40390
rect 17222 40352 17278 40361
rect 17316 40326 17368 40332
rect 17222 40287 17278 40296
rect 17224 40180 17276 40186
rect 17144 40140 17224 40168
rect 17224 40122 17276 40128
rect 17236 40089 17264 40122
rect 17222 40080 17278 40089
rect 17222 40015 17278 40024
rect 17052 39902 17264 39930
rect 17132 39840 17184 39846
rect 16960 39766 17080 39794
rect 17132 39782 17184 39788
rect 16856 39500 16908 39506
rect 16856 39442 16908 39448
rect 16764 39432 16816 39438
rect 16764 39374 16816 39380
rect 16776 38826 16804 39374
rect 16868 38876 16896 39442
rect 16948 38888 17000 38894
rect 16868 38848 16948 38876
rect 16764 38820 16816 38826
rect 16764 38762 16816 38768
rect 16776 36854 16804 38762
rect 16868 38554 16896 38848
rect 16948 38830 17000 38836
rect 17052 38706 17080 39766
rect 16960 38678 17080 38706
rect 16856 38548 16908 38554
rect 16856 38490 16908 38496
rect 16856 38412 16908 38418
rect 16856 38354 16908 38360
rect 16868 38010 16896 38354
rect 16856 38004 16908 38010
rect 16856 37946 16908 37952
rect 16856 37868 16908 37874
rect 16856 37810 16908 37816
rect 16764 36848 16816 36854
rect 16764 36790 16816 36796
rect 16868 34610 16896 37810
rect 16856 34604 16908 34610
rect 16856 34546 16908 34552
rect 16868 34202 16896 34546
rect 16856 34196 16908 34202
rect 16856 34138 16908 34144
rect 16868 32722 16896 34138
rect 16776 32694 16896 32722
rect 16672 28688 16724 28694
rect 16672 28630 16724 28636
rect 16580 28620 16632 28626
rect 16580 28562 16632 28568
rect 16592 27402 16620 28562
rect 16488 27396 16540 27402
rect 16488 27338 16540 27344
rect 16580 27396 16632 27402
rect 16580 27338 16632 27344
rect 16488 27056 16540 27062
rect 16488 26998 16540 27004
rect 16316 25622 16436 25650
rect 16118 24984 16174 24993
rect 16118 24919 16174 24928
rect 16212 24676 16264 24682
rect 16212 24618 16264 24624
rect 15936 23792 15988 23798
rect 15936 23734 15988 23740
rect 15844 23656 15896 23662
rect 15844 23598 15896 23604
rect 16224 23526 16252 24618
rect 15936 23520 15988 23526
rect 15936 23462 15988 23468
rect 16212 23520 16264 23526
rect 16212 23462 16264 23468
rect 15488 23140 15700 23168
rect 15476 23044 15528 23050
rect 15476 22986 15528 22992
rect 15384 21956 15436 21962
rect 15384 21898 15436 21904
rect 15292 21616 15344 21622
rect 15292 21558 15344 21564
rect 15198 21448 15254 21457
rect 15198 21383 15254 21392
rect 15106 21312 15162 21321
rect 15106 21247 15162 21256
rect 15120 21010 15148 21247
rect 15108 21004 15160 21010
rect 15108 20946 15160 20952
rect 15120 20602 15148 20946
rect 15108 20596 15160 20602
rect 15108 20538 15160 20544
rect 15200 20392 15252 20398
rect 15028 20340 15200 20346
rect 15028 20334 15252 20340
rect 15028 20318 15240 20334
rect 14924 20256 14976 20262
rect 14924 20198 14976 20204
rect 14936 18834 14964 20198
rect 15028 19310 15056 20318
rect 15396 20097 15424 21898
rect 15488 20913 15516 22986
rect 15672 22166 15700 23140
rect 15660 22160 15712 22166
rect 15660 22102 15712 22108
rect 15660 22024 15712 22030
rect 15660 21966 15712 21972
rect 15568 21888 15620 21894
rect 15568 21830 15620 21836
rect 15580 21418 15608 21830
rect 15672 21690 15700 21966
rect 15660 21684 15712 21690
rect 15660 21626 15712 21632
rect 15568 21412 15620 21418
rect 15568 21354 15620 21360
rect 15580 21078 15608 21354
rect 15568 21072 15620 21078
rect 15568 21014 15620 21020
rect 15672 21010 15700 21626
rect 15948 21321 15976 23462
rect 16120 23112 16172 23118
rect 16120 23054 16172 23060
rect 16028 22976 16080 22982
rect 16028 22918 16080 22924
rect 16040 22681 16068 22918
rect 16132 22817 16160 23054
rect 16118 22808 16174 22817
rect 16118 22743 16120 22752
rect 16172 22743 16174 22752
rect 16120 22714 16172 22720
rect 16026 22672 16082 22681
rect 16026 22607 16082 22616
rect 16224 22098 16252 23462
rect 16212 22092 16264 22098
rect 16212 22034 16264 22040
rect 15934 21312 15990 21321
rect 15934 21247 15990 21256
rect 16316 21010 16344 25622
rect 16394 25528 16450 25537
rect 16394 25463 16450 25472
rect 16408 24290 16436 25463
rect 16500 24834 16528 26998
rect 16592 26518 16620 27338
rect 16580 26512 16632 26518
rect 16580 26454 16632 26460
rect 16776 25276 16804 32694
rect 16856 32292 16908 32298
rect 16856 32234 16908 32240
rect 16868 30870 16896 32234
rect 16960 30938 16988 38678
rect 17144 37346 17172 39782
rect 17052 37318 17172 37346
rect 17052 33674 17080 37318
rect 17132 37256 17184 37262
rect 17132 37198 17184 37204
rect 17144 36553 17172 37198
rect 17130 36544 17186 36553
rect 17130 36479 17186 36488
rect 17132 35080 17184 35086
rect 17132 35022 17184 35028
rect 17144 34513 17172 35022
rect 17130 34504 17186 34513
rect 17130 34439 17186 34448
rect 17132 33992 17184 33998
rect 17130 33960 17132 33969
rect 17184 33960 17186 33969
rect 17130 33895 17186 33904
rect 17052 33646 17172 33674
rect 17038 33552 17094 33561
rect 17038 33487 17094 33496
rect 17052 33454 17080 33487
rect 17040 33448 17092 33454
rect 17040 33390 17092 33396
rect 17144 33266 17172 33646
rect 17052 33238 17172 33266
rect 16948 30932 17000 30938
rect 16948 30874 17000 30880
rect 16856 30864 16908 30870
rect 16856 30806 16908 30812
rect 16856 30660 16908 30666
rect 16856 30602 16908 30608
rect 16868 30002 16896 30602
rect 16960 30190 16988 30874
rect 16948 30184 17000 30190
rect 16948 30126 17000 30132
rect 16868 29974 16988 30002
rect 16856 27668 16908 27674
rect 16856 27610 16908 27616
rect 16868 26994 16896 27610
rect 16856 26988 16908 26994
rect 16856 26930 16908 26936
rect 16868 26586 16896 26930
rect 16856 26580 16908 26586
rect 16856 26522 16908 26528
rect 16868 26042 16896 26522
rect 16856 26036 16908 26042
rect 16856 25978 16908 25984
rect 16868 25906 16896 25978
rect 16856 25900 16908 25906
rect 16856 25842 16908 25848
rect 16960 25276 16988 29974
rect 17052 26926 17080 33238
rect 17130 33144 17186 33153
rect 17130 33079 17186 33088
rect 17144 33046 17172 33079
rect 17132 33040 17184 33046
rect 17132 32982 17184 32988
rect 17130 32872 17186 32881
rect 17130 32807 17186 32816
rect 17144 29850 17172 32807
rect 17236 29866 17264 39902
rect 17328 39642 17356 40326
rect 17316 39636 17368 39642
rect 17316 39578 17368 39584
rect 17316 38548 17368 38554
rect 17316 38490 17368 38496
rect 17328 37806 17356 38490
rect 17316 37800 17368 37806
rect 17316 37742 17368 37748
rect 17420 37466 17448 41142
rect 17408 37460 17460 37466
rect 17408 37402 17460 37408
rect 17512 37312 17540 41398
rect 17622 41372 17918 41392
rect 17678 41370 17702 41372
rect 17758 41370 17782 41372
rect 17838 41370 17862 41372
rect 17700 41318 17702 41370
rect 17764 41318 17776 41370
rect 17838 41318 17840 41370
rect 17678 41316 17702 41318
rect 17758 41316 17782 41318
rect 17838 41316 17862 41318
rect 17622 41296 17918 41316
rect 17972 41274 18000 42055
rect 17960 41268 18012 41274
rect 17960 41210 18012 41216
rect 17592 41064 17644 41070
rect 17592 41006 17644 41012
rect 17604 40730 17632 41006
rect 17592 40724 17644 40730
rect 17592 40666 17644 40672
rect 17622 40284 17918 40304
rect 17678 40282 17702 40284
rect 17758 40282 17782 40284
rect 17838 40282 17862 40284
rect 17700 40230 17702 40282
rect 17764 40230 17776 40282
rect 17838 40230 17840 40282
rect 17678 40228 17702 40230
rect 17758 40228 17782 40230
rect 17838 40228 17862 40230
rect 17622 40208 17918 40228
rect 17622 39196 17918 39216
rect 17678 39194 17702 39196
rect 17758 39194 17782 39196
rect 17838 39194 17862 39196
rect 17700 39142 17702 39194
rect 17764 39142 17776 39194
rect 17838 39142 17840 39194
rect 17678 39140 17702 39142
rect 17758 39140 17782 39142
rect 17838 39140 17862 39142
rect 17622 39120 17918 39140
rect 18064 38826 18092 43046
rect 18156 40594 18184 46378
rect 18420 45960 18472 45966
rect 18420 45902 18472 45908
rect 18236 45280 18288 45286
rect 18236 45222 18288 45228
rect 18248 42673 18276 45222
rect 18328 45076 18380 45082
rect 18328 45018 18380 45024
rect 18234 42664 18290 42673
rect 18234 42599 18290 42608
rect 18340 42294 18368 45018
rect 18432 43314 18460 45902
rect 18420 43308 18472 43314
rect 18420 43250 18472 43256
rect 18328 42288 18380 42294
rect 18328 42230 18380 42236
rect 18328 41540 18380 41546
rect 18328 41482 18380 41488
rect 18340 41206 18368 41482
rect 18328 41200 18380 41206
rect 18328 41142 18380 41148
rect 18144 40588 18196 40594
rect 18144 40530 18196 40536
rect 18156 40186 18184 40530
rect 18144 40180 18196 40186
rect 18144 40122 18196 40128
rect 18432 39846 18460 43250
rect 18420 39840 18472 39846
rect 18420 39782 18472 39788
rect 18234 39536 18290 39545
rect 18234 39471 18290 39480
rect 18248 39098 18276 39471
rect 18236 39092 18288 39098
rect 18236 39034 18288 39040
rect 18052 38820 18104 38826
rect 18052 38762 18104 38768
rect 17622 38108 17918 38128
rect 17678 38106 17702 38108
rect 17758 38106 17782 38108
rect 17838 38106 17862 38108
rect 17700 38054 17702 38106
rect 17764 38054 17776 38106
rect 17838 38054 17840 38106
rect 17678 38052 17702 38054
rect 17758 38052 17782 38054
rect 17838 38052 17862 38054
rect 17622 38032 17918 38052
rect 17960 38004 18012 38010
rect 17960 37946 18012 37952
rect 17328 37284 17540 37312
rect 17328 31822 17356 37284
rect 17498 37224 17554 37233
rect 17408 37188 17460 37194
rect 17498 37159 17554 37168
rect 17408 37130 17460 37136
rect 17420 36854 17448 37130
rect 17408 36848 17460 36854
rect 17408 36790 17460 36796
rect 17408 36712 17460 36718
rect 17408 36654 17460 36660
rect 17420 36378 17448 36654
rect 17408 36372 17460 36378
rect 17408 36314 17460 36320
rect 17420 35290 17448 36314
rect 17512 35766 17540 37159
rect 17622 37020 17918 37040
rect 17678 37018 17702 37020
rect 17758 37018 17782 37020
rect 17838 37018 17862 37020
rect 17700 36966 17702 37018
rect 17764 36966 17776 37018
rect 17838 36966 17840 37018
rect 17678 36964 17702 36966
rect 17758 36964 17782 36966
rect 17838 36964 17862 36966
rect 17622 36944 17918 36964
rect 17684 36644 17736 36650
rect 17684 36586 17736 36592
rect 17868 36644 17920 36650
rect 17868 36586 17920 36592
rect 17696 36020 17724 36586
rect 17880 36122 17908 36586
rect 17972 36242 18000 37946
rect 18052 37120 18104 37126
rect 18052 37062 18104 37068
rect 18064 36922 18092 37062
rect 18052 36916 18104 36922
rect 18104 36876 18184 36904
rect 18052 36858 18104 36864
rect 17960 36236 18012 36242
rect 17960 36178 18012 36184
rect 17880 36094 18092 36122
rect 17696 35992 18000 36020
rect 17622 35932 17918 35952
rect 17678 35930 17702 35932
rect 17758 35930 17782 35932
rect 17838 35930 17862 35932
rect 17700 35878 17702 35930
rect 17764 35878 17776 35930
rect 17838 35878 17840 35930
rect 17678 35876 17702 35878
rect 17758 35876 17782 35878
rect 17838 35876 17862 35878
rect 17622 35856 17918 35876
rect 17500 35760 17552 35766
rect 17500 35702 17552 35708
rect 17408 35284 17460 35290
rect 17408 35226 17460 35232
rect 17420 34542 17448 35226
rect 17498 35184 17554 35193
rect 17498 35119 17554 35128
rect 17512 34678 17540 35119
rect 17622 34844 17918 34864
rect 17678 34842 17702 34844
rect 17758 34842 17782 34844
rect 17838 34842 17862 34844
rect 17700 34790 17702 34842
rect 17764 34790 17776 34842
rect 17838 34790 17840 34842
rect 17678 34788 17702 34790
rect 17758 34788 17782 34790
rect 17838 34788 17862 34790
rect 17622 34768 17918 34788
rect 17500 34672 17552 34678
rect 17500 34614 17552 34620
rect 17408 34536 17460 34542
rect 17408 34478 17460 34484
rect 17622 33756 17918 33776
rect 17678 33754 17702 33756
rect 17758 33754 17782 33756
rect 17838 33754 17862 33756
rect 17700 33702 17702 33754
rect 17764 33702 17776 33754
rect 17838 33702 17840 33754
rect 17678 33700 17702 33702
rect 17758 33700 17782 33702
rect 17838 33700 17862 33702
rect 17622 33680 17918 33700
rect 17500 33584 17552 33590
rect 17500 33526 17552 33532
rect 17408 33040 17460 33046
rect 17406 33008 17408 33017
rect 17460 33008 17462 33017
rect 17406 32943 17462 32952
rect 17420 32366 17448 32943
rect 17512 32473 17540 33526
rect 17622 32668 17918 32688
rect 17678 32666 17702 32668
rect 17758 32666 17782 32668
rect 17838 32666 17862 32668
rect 17700 32614 17702 32666
rect 17764 32614 17776 32666
rect 17838 32614 17840 32666
rect 17678 32612 17702 32614
rect 17758 32612 17782 32614
rect 17838 32612 17862 32614
rect 17622 32592 17918 32612
rect 17498 32464 17554 32473
rect 17498 32399 17554 32408
rect 17408 32360 17460 32366
rect 17408 32302 17460 32308
rect 17776 32292 17828 32298
rect 17776 32234 17828 32240
rect 17408 32224 17460 32230
rect 17408 32166 17460 32172
rect 17316 31816 17368 31822
rect 17316 31758 17368 31764
rect 17328 31278 17356 31758
rect 17316 31272 17368 31278
rect 17316 31214 17368 31220
rect 17132 29844 17184 29850
rect 17236 29838 17356 29866
rect 17132 29786 17184 29792
rect 17144 29102 17172 29786
rect 17222 29744 17278 29753
rect 17222 29679 17278 29688
rect 17132 29096 17184 29102
rect 17132 29038 17184 29044
rect 17236 28694 17264 29679
rect 17224 28688 17276 28694
rect 17224 28630 17276 28636
rect 17328 28014 17356 29838
rect 17420 28506 17448 32166
rect 17500 31952 17552 31958
rect 17500 31894 17552 31900
rect 17512 31278 17540 31894
rect 17788 31793 17816 32234
rect 17972 32230 18000 35992
rect 18064 35873 18092 36094
rect 18050 35864 18106 35873
rect 18156 35834 18184 36876
rect 18050 35799 18106 35808
rect 18144 35828 18196 35834
rect 18144 35770 18196 35776
rect 18052 33312 18104 33318
rect 18052 33254 18104 33260
rect 18064 32366 18092 33254
rect 18420 32904 18472 32910
rect 18420 32846 18472 32852
rect 18432 32570 18460 32846
rect 18420 32564 18472 32570
rect 18420 32506 18472 32512
rect 18052 32360 18104 32366
rect 18052 32302 18104 32308
rect 17960 32224 18012 32230
rect 17960 32166 18012 32172
rect 17774 31784 17830 31793
rect 17774 31719 17830 31728
rect 17622 31580 17918 31600
rect 17678 31578 17702 31580
rect 17758 31578 17782 31580
rect 17838 31578 17862 31580
rect 17700 31526 17702 31578
rect 17764 31526 17776 31578
rect 17838 31526 17840 31578
rect 17678 31524 17702 31526
rect 17758 31524 17782 31526
rect 17838 31524 17862 31526
rect 17622 31504 17918 31524
rect 17500 31272 17552 31278
rect 17500 31214 17552 31220
rect 17512 30190 17540 31214
rect 17776 31204 17828 31210
rect 17776 31146 17828 31152
rect 17788 31113 17816 31146
rect 17774 31104 17830 31113
rect 17774 31039 17830 31048
rect 17622 30492 17918 30512
rect 17678 30490 17702 30492
rect 17758 30490 17782 30492
rect 17838 30490 17862 30492
rect 17700 30438 17702 30490
rect 17764 30438 17776 30490
rect 17838 30438 17840 30490
rect 17678 30436 17702 30438
rect 17758 30436 17782 30438
rect 17838 30436 17862 30438
rect 17622 30416 17918 30436
rect 17866 30288 17922 30297
rect 17866 30223 17868 30232
rect 17920 30223 17922 30232
rect 17868 30194 17920 30200
rect 17500 30184 17552 30190
rect 17500 30126 17552 30132
rect 17500 29504 17552 29510
rect 17500 29446 17552 29452
rect 17512 29102 17540 29446
rect 17622 29404 17918 29424
rect 17678 29402 17702 29404
rect 17758 29402 17782 29404
rect 17838 29402 17862 29404
rect 17700 29350 17702 29402
rect 17764 29350 17776 29402
rect 17838 29350 17840 29402
rect 17678 29348 17702 29350
rect 17758 29348 17782 29350
rect 17838 29348 17862 29350
rect 17622 29328 17918 29348
rect 17500 29096 17552 29102
rect 17776 29096 17828 29102
rect 17500 29038 17552 29044
rect 17774 29064 17776 29073
rect 17828 29064 17830 29073
rect 17512 28626 17540 29038
rect 17774 28999 17830 29008
rect 17500 28620 17552 28626
rect 17500 28562 17552 28568
rect 17420 28478 17540 28506
rect 17408 28416 17460 28422
rect 17408 28358 17460 28364
rect 17420 28014 17448 28358
rect 17316 28008 17368 28014
rect 17316 27950 17368 27956
rect 17408 28008 17460 28014
rect 17408 27950 17460 27956
rect 17132 27600 17184 27606
rect 17132 27542 17184 27548
rect 17144 27130 17172 27542
rect 17420 27538 17448 27950
rect 17512 27826 17540 28478
rect 17622 28316 17918 28336
rect 17678 28314 17702 28316
rect 17758 28314 17782 28316
rect 17838 28314 17862 28316
rect 17700 28262 17702 28314
rect 17764 28262 17776 28314
rect 17838 28262 17840 28314
rect 17678 28260 17702 28262
rect 17758 28260 17782 28262
rect 17838 28260 17862 28262
rect 17622 28240 17918 28260
rect 17774 28112 17830 28121
rect 17774 28047 17776 28056
rect 17828 28047 17830 28056
rect 17776 28018 17828 28024
rect 17512 27798 17632 27826
rect 17498 27704 17554 27713
rect 17498 27639 17554 27648
rect 17408 27532 17460 27538
rect 17408 27474 17460 27480
rect 17316 27464 17368 27470
rect 17316 27406 17368 27412
rect 17132 27124 17184 27130
rect 17132 27066 17184 27072
rect 17040 26920 17092 26926
rect 17040 26862 17092 26868
rect 17038 25936 17094 25945
rect 17038 25871 17094 25880
rect 17052 25838 17080 25871
rect 17040 25832 17092 25838
rect 17040 25774 17092 25780
rect 17040 25288 17092 25294
rect 16776 25248 16896 25276
rect 16960 25248 17040 25276
rect 16764 25152 16816 25158
rect 16764 25094 16816 25100
rect 16670 24984 16726 24993
rect 16670 24919 16726 24928
rect 16500 24818 16620 24834
rect 16500 24812 16632 24818
rect 16500 24806 16580 24812
rect 16580 24754 16632 24760
rect 16408 24262 16528 24290
rect 16394 24168 16450 24177
rect 16394 24103 16450 24112
rect 15660 21004 15712 21010
rect 15660 20946 15712 20952
rect 16028 21004 16080 21010
rect 16028 20946 16080 20952
rect 16304 21004 16356 21010
rect 16304 20946 16356 20952
rect 15474 20904 15530 20913
rect 15474 20839 15530 20848
rect 16040 20602 16068 20946
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 15844 20392 15896 20398
rect 15844 20334 15896 20340
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15382 20088 15438 20097
rect 15382 20023 15438 20032
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 15200 19780 15252 19786
rect 15200 19722 15252 19728
rect 15016 19304 15068 19310
rect 15016 19246 15068 19252
rect 14924 18828 14976 18834
rect 14924 18770 14976 18776
rect 15212 18737 15240 19722
rect 15304 19174 15332 19858
rect 15292 19168 15344 19174
rect 15344 19128 15424 19156
rect 15292 19110 15344 19116
rect 15198 18728 15254 18737
rect 15108 18692 15160 18698
rect 15198 18663 15254 18672
rect 15108 18634 15160 18640
rect 15014 18456 15070 18465
rect 15014 18391 15070 18400
rect 14924 18216 14976 18222
rect 14924 18158 14976 18164
rect 14936 17542 14964 18158
rect 14924 17536 14976 17542
rect 14924 17478 14976 17484
rect 14936 16454 14964 17478
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 14936 15502 14964 15846
rect 14924 15496 14976 15502
rect 14924 15438 14976 15444
rect 14936 14890 14964 15438
rect 14924 14884 14976 14890
rect 14924 14826 14976 14832
rect 15028 14498 15056 18391
rect 15120 18057 15148 18634
rect 15198 18320 15254 18329
rect 15198 18255 15254 18264
rect 15106 18048 15162 18057
rect 15106 17983 15162 17992
rect 15108 17740 15160 17746
rect 15108 17682 15160 17688
rect 15120 17270 15148 17682
rect 15212 17649 15240 18255
rect 15198 17640 15254 17649
rect 15198 17575 15254 17584
rect 15108 17264 15160 17270
rect 15108 17206 15160 17212
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15304 16522 15332 17070
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15396 16046 15424 19128
rect 15580 17354 15608 20198
rect 15856 19922 15884 20334
rect 16316 20058 16344 20946
rect 16408 20754 16436 24103
rect 16500 21962 16528 24262
rect 16592 24154 16620 24754
rect 16684 24410 16712 24919
rect 16672 24404 16724 24410
rect 16672 24346 16724 24352
rect 16592 24126 16712 24154
rect 16580 23180 16632 23186
rect 16580 23122 16632 23128
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 16592 21894 16620 23122
rect 16684 22574 16712 24126
rect 16776 23730 16804 25094
rect 16868 24410 16896 25248
rect 17040 25230 17092 25236
rect 17052 24750 17080 25230
rect 17040 24744 17092 24750
rect 17040 24686 17092 24692
rect 16856 24404 16908 24410
rect 16856 24346 16908 24352
rect 16764 23724 16816 23730
rect 16764 23666 16816 23672
rect 16868 23594 16896 24346
rect 17040 24268 17092 24274
rect 17040 24210 17092 24216
rect 16948 23792 17000 23798
rect 16948 23734 17000 23740
rect 16764 23588 16816 23594
rect 16764 23530 16816 23536
rect 16856 23588 16908 23594
rect 16856 23530 16908 23536
rect 16776 22642 16804 23530
rect 16764 22636 16816 22642
rect 16764 22578 16816 22584
rect 16672 22568 16724 22574
rect 16724 22516 16804 22522
rect 16672 22510 16804 22516
rect 16684 22494 16804 22510
rect 16672 22092 16724 22098
rect 16672 22034 16724 22040
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 16580 21344 16632 21350
rect 16578 21312 16580 21321
rect 16632 21312 16634 21321
rect 16578 21247 16634 21256
rect 16684 21146 16712 22034
rect 16776 22030 16804 22494
rect 16856 22500 16908 22506
rect 16856 22442 16908 22448
rect 16868 22098 16896 22442
rect 16856 22092 16908 22098
rect 16856 22034 16908 22040
rect 16764 22024 16816 22030
rect 16764 21966 16816 21972
rect 16764 21412 16816 21418
rect 16764 21354 16816 21360
rect 16672 21140 16724 21146
rect 16672 21082 16724 21088
rect 16776 21078 16804 21354
rect 16764 21072 16816 21078
rect 16764 21014 16816 21020
rect 16868 20890 16896 22034
rect 16776 20862 16896 20890
rect 16776 20806 16804 20862
rect 16764 20800 16816 20806
rect 16408 20726 16528 20754
rect 16764 20742 16816 20748
rect 16500 20618 16528 20726
rect 16500 20590 16620 20618
rect 16592 20534 16620 20590
rect 16580 20528 16632 20534
rect 16580 20470 16632 20476
rect 16304 20052 16356 20058
rect 16304 19994 16356 20000
rect 15934 19952 15990 19961
rect 15844 19916 15896 19922
rect 15934 19887 15990 19896
rect 15844 19858 15896 19864
rect 15844 19304 15896 19310
rect 15844 19246 15896 19252
rect 15752 18828 15804 18834
rect 15752 18770 15804 18776
rect 15764 18086 15792 18770
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 15488 17326 15608 17354
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 15396 15706 15424 15982
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15108 15564 15160 15570
rect 15108 15506 15160 15512
rect 15120 15162 15148 15506
rect 15396 15434 15424 15642
rect 15384 15428 15436 15434
rect 15384 15370 15436 15376
rect 15108 15156 15160 15162
rect 15108 15098 15160 15104
rect 15382 14920 15438 14929
rect 15108 14884 15160 14890
rect 15382 14855 15438 14864
rect 15108 14826 15160 14832
rect 14936 14470 15056 14498
rect 14936 13462 14964 14470
rect 15016 14340 15068 14346
rect 15016 14282 15068 14288
rect 14924 13456 14976 13462
rect 14924 13398 14976 13404
rect 14936 12442 14964 13398
rect 14924 12436 14976 12442
rect 14924 12378 14976 12384
rect 14844 12158 14964 12186
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14752 10810 14780 11834
rect 14844 11694 14872 12038
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14844 11354 14872 11630
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14936 11234 14964 12158
rect 14844 11206 14964 11234
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14752 9518 14780 9998
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14752 8090 14780 9454
rect 14844 8430 14872 11206
rect 15028 10577 15056 14282
rect 15120 11762 15148 14826
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15304 13870 15332 14758
rect 15396 14618 15424 14855
rect 15384 14612 15436 14618
rect 15384 14554 15436 14560
rect 15292 13864 15344 13870
rect 15198 13832 15254 13841
rect 15292 13806 15344 13812
rect 15198 13767 15254 13776
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15014 10568 15070 10577
rect 15014 10503 15070 10512
rect 14924 10464 14976 10470
rect 14924 10406 14976 10412
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 14752 6730 14780 7890
rect 14740 6724 14792 6730
rect 14740 6666 14792 6672
rect 14752 6390 14780 6666
rect 14740 6384 14792 6390
rect 14740 6326 14792 6332
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 14016 6118 14044 6190
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14289 6012 14585 6032
rect 14345 6010 14369 6012
rect 14425 6010 14449 6012
rect 14505 6010 14529 6012
rect 14367 5958 14369 6010
rect 14431 5958 14443 6010
rect 14505 5958 14507 6010
rect 14345 5956 14369 5958
rect 14425 5956 14449 5958
rect 14505 5956 14529 5958
rect 14289 5936 14585 5956
rect 14660 5914 14688 6258
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14016 5234 14044 5850
rect 14094 5808 14150 5817
rect 14094 5743 14150 5752
rect 14646 5808 14702 5817
rect 14646 5743 14648 5752
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 12452 5086 12572 5114
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 12452 4978 12480 5086
rect 12360 4950 12480 4978
rect 12360 4146 12388 4950
rect 13924 4826 13952 5102
rect 14108 4826 14136 5743
rect 14700 5743 14702 5752
rect 14648 5714 14700 5720
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 13912 4820 13964 4826
rect 13912 4762 13964 4768
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14200 4622 14228 5102
rect 14648 5024 14700 5030
rect 14648 4966 14700 4972
rect 14289 4924 14585 4944
rect 14345 4922 14369 4924
rect 14425 4922 14449 4924
rect 14505 4922 14529 4924
rect 14367 4870 14369 4922
rect 14431 4870 14443 4922
rect 14505 4870 14507 4922
rect 14345 4868 14369 4870
rect 14425 4868 14449 4870
rect 14505 4868 14529 4870
rect 14289 4848 14585 4868
rect 14556 4752 14608 4758
rect 14660 4729 14688 4966
rect 14556 4694 14608 4700
rect 14646 4720 14702 4729
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14200 4282 14228 4558
rect 14568 4282 14596 4694
rect 14646 4655 14702 4664
rect 14844 4554 14872 8366
rect 14936 7410 14964 10406
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 15028 9518 15056 10066
rect 15120 9874 15148 11494
rect 15212 11257 15240 13767
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15304 12102 15332 12922
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15396 11914 15424 12718
rect 15304 11886 15424 11914
rect 15198 11248 15254 11257
rect 15304 11218 15332 11886
rect 15382 11792 15438 11801
rect 15382 11727 15438 11736
rect 15198 11183 15254 11192
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 15200 9920 15252 9926
rect 15120 9868 15200 9874
rect 15120 9862 15252 9868
rect 15120 9846 15240 9862
rect 15120 9586 15148 9846
rect 15304 9722 15332 10066
rect 15396 10033 15424 11727
rect 15488 11234 15516 17326
rect 15568 17264 15620 17270
rect 15568 17206 15620 17212
rect 15580 16017 15608 17206
rect 15660 17060 15712 17066
rect 15660 17002 15712 17008
rect 15672 16590 15700 17002
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15566 16008 15622 16017
rect 15566 15943 15622 15952
rect 15672 15366 15700 16050
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15566 13968 15622 13977
rect 15566 13903 15622 13912
rect 15580 12918 15608 13903
rect 15672 13433 15700 15302
rect 15658 13424 15714 13433
rect 15658 13359 15714 13368
rect 15660 13252 15712 13258
rect 15660 13194 15712 13200
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15672 12850 15700 13194
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15672 12186 15700 12786
rect 15764 12306 15792 18022
rect 15856 14822 15884 19246
rect 15948 16640 15976 19887
rect 16316 19446 16344 19994
rect 16304 19440 16356 19446
rect 16304 19382 16356 19388
rect 16776 19242 16804 20742
rect 16960 19530 16988 23734
rect 17052 23526 17080 24210
rect 17144 23662 17172 27066
rect 17328 26790 17356 27406
rect 17420 26926 17448 27474
rect 17512 27062 17540 27639
rect 17604 27606 17632 27798
rect 17592 27600 17644 27606
rect 17592 27542 17644 27548
rect 17622 27228 17918 27248
rect 17678 27226 17702 27228
rect 17758 27226 17782 27228
rect 17838 27226 17862 27228
rect 17700 27174 17702 27226
rect 17764 27174 17776 27226
rect 17838 27174 17840 27226
rect 17678 27172 17702 27174
rect 17758 27172 17782 27174
rect 17838 27172 17862 27174
rect 17622 27152 17918 27172
rect 17500 27056 17552 27062
rect 17500 26998 17552 27004
rect 17590 27024 17646 27033
rect 17590 26959 17646 26968
rect 17408 26920 17460 26926
rect 17408 26862 17460 26868
rect 17316 26784 17368 26790
rect 17316 26726 17368 26732
rect 17328 26382 17356 26726
rect 17316 26376 17368 26382
rect 17604 26364 17632 26959
rect 17316 26318 17368 26324
rect 17512 26336 17632 26364
rect 17328 25702 17356 26318
rect 17512 25974 17540 26336
rect 17622 26140 17918 26160
rect 17678 26138 17702 26140
rect 17758 26138 17782 26140
rect 17838 26138 17862 26140
rect 17700 26086 17702 26138
rect 17764 26086 17776 26138
rect 17838 26086 17840 26138
rect 17678 26084 17702 26086
rect 17758 26084 17782 26086
rect 17838 26084 17862 26086
rect 17622 26064 17918 26084
rect 17500 25968 17552 25974
rect 17500 25910 17552 25916
rect 17590 25936 17646 25945
rect 17590 25871 17646 25880
rect 17408 25832 17460 25838
rect 17408 25774 17460 25780
rect 17316 25696 17368 25702
rect 17316 25638 17368 25644
rect 17328 24562 17356 25638
rect 17420 25158 17448 25774
rect 17604 25378 17632 25871
rect 17512 25350 17632 25378
rect 17408 25152 17460 25158
rect 17408 25094 17460 25100
rect 17420 24750 17448 25094
rect 17512 24886 17540 25350
rect 17622 25052 17918 25072
rect 17678 25050 17702 25052
rect 17758 25050 17782 25052
rect 17838 25050 17862 25052
rect 17700 24998 17702 25050
rect 17764 24998 17776 25050
rect 17838 24998 17840 25050
rect 17678 24996 17702 24998
rect 17758 24996 17782 24998
rect 17838 24996 17862 24998
rect 17622 24976 17918 24996
rect 17500 24880 17552 24886
rect 17500 24822 17552 24828
rect 17590 24848 17646 24857
rect 17590 24783 17646 24792
rect 17408 24744 17460 24750
rect 17408 24686 17460 24692
rect 17328 24534 17448 24562
rect 17224 24336 17276 24342
rect 17224 24278 17276 24284
rect 17132 23656 17184 23662
rect 17132 23598 17184 23604
rect 17040 23520 17092 23526
rect 17040 23462 17092 23468
rect 17130 23488 17186 23497
rect 17052 23186 17080 23462
rect 17130 23423 17186 23432
rect 17040 23180 17092 23186
rect 17040 23122 17092 23128
rect 17040 22976 17092 22982
rect 17040 22918 17092 22924
rect 17052 21622 17080 22918
rect 17040 21616 17092 21622
rect 17040 21558 17092 21564
rect 17052 21418 17080 21558
rect 17040 21412 17092 21418
rect 17040 21354 17092 21360
rect 17144 21078 17172 23423
rect 17236 21554 17264 24278
rect 17420 23730 17448 24534
rect 17604 24154 17632 24783
rect 17512 24126 17632 24154
rect 17408 23724 17460 23730
rect 17408 23666 17460 23672
rect 17316 23520 17368 23526
rect 17316 23462 17368 23468
rect 17328 22794 17356 23462
rect 17420 22982 17448 23666
rect 17408 22976 17460 22982
rect 17408 22918 17460 22924
rect 17328 22766 17448 22794
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 17224 21412 17276 21418
rect 17224 21354 17276 21360
rect 17132 21072 17184 21078
rect 17132 21014 17184 21020
rect 17236 20806 17264 21354
rect 17224 20800 17276 20806
rect 17224 20742 17276 20748
rect 17236 19718 17264 20742
rect 17420 20398 17448 22766
rect 17512 22710 17540 24126
rect 17622 23964 17918 23984
rect 17678 23962 17702 23964
rect 17758 23962 17782 23964
rect 17838 23962 17862 23964
rect 17700 23910 17702 23962
rect 17764 23910 17776 23962
rect 17838 23910 17840 23962
rect 17678 23908 17702 23910
rect 17758 23908 17782 23910
rect 17838 23908 17862 23910
rect 17622 23888 17918 23908
rect 17622 22876 17918 22896
rect 17678 22874 17702 22876
rect 17758 22874 17782 22876
rect 17838 22874 17862 22876
rect 17700 22822 17702 22874
rect 17764 22822 17776 22874
rect 17838 22822 17840 22874
rect 17678 22820 17702 22822
rect 17758 22820 17782 22822
rect 17838 22820 17862 22822
rect 17622 22800 17918 22820
rect 17500 22704 17552 22710
rect 17500 22646 17552 22652
rect 17622 21788 17918 21808
rect 17678 21786 17702 21788
rect 17758 21786 17782 21788
rect 17838 21786 17862 21788
rect 17700 21734 17702 21786
rect 17764 21734 17776 21786
rect 17838 21734 17840 21786
rect 17678 21732 17702 21734
rect 17758 21732 17782 21734
rect 17838 21732 17862 21734
rect 17622 21712 17918 21732
rect 17500 21004 17552 21010
rect 17500 20946 17552 20952
rect 17512 20398 17540 20946
rect 17622 20700 17918 20720
rect 17678 20698 17702 20700
rect 17758 20698 17782 20700
rect 17838 20698 17862 20700
rect 17700 20646 17702 20698
rect 17764 20646 17776 20698
rect 17838 20646 17840 20698
rect 17678 20644 17702 20646
rect 17758 20644 17782 20646
rect 17838 20644 17862 20646
rect 17622 20624 17918 20644
rect 17408 20392 17460 20398
rect 17408 20334 17460 20340
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17420 20058 17448 20334
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17512 19922 17540 20334
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17224 19712 17276 19718
rect 17224 19654 17276 19660
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 16960 19502 17356 19530
rect 17328 19310 17356 19502
rect 17512 19378 17540 19654
rect 17622 19612 17918 19632
rect 17678 19610 17702 19612
rect 17758 19610 17782 19612
rect 17838 19610 17862 19612
rect 17700 19558 17702 19610
rect 17764 19558 17776 19610
rect 17838 19558 17840 19610
rect 17678 19556 17702 19558
rect 17758 19556 17782 19558
rect 17838 19556 17862 19558
rect 17622 19536 17918 19556
rect 17500 19372 17552 19378
rect 17500 19314 17552 19320
rect 17316 19304 17368 19310
rect 17316 19246 17368 19252
rect 16764 19236 16816 19242
rect 16764 19178 16816 19184
rect 16488 18828 16540 18834
rect 16488 18770 16540 18776
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16132 18222 16160 18702
rect 16396 18284 16448 18290
rect 16396 18226 16448 18232
rect 16120 18216 16172 18222
rect 16120 18158 16172 18164
rect 16132 17542 16160 18158
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 16132 16794 16160 17478
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 16120 16652 16172 16658
rect 15948 16612 16120 16640
rect 16120 16594 16172 16600
rect 15936 16176 15988 16182
rect 15936 16118 15988 16124
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15672 12158 15792 12186
rect 15764 12102 15792 12158
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15488 11206 15608 11234
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15382 10024 15438 10033
rect 15382 9959 15438 9968
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15198 9616 15254 9625
rect 15108 9580 15160 9586
rect 15198 9551 15254 9560
rect 15108 9522 15160 9528
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 15028 8022 15056 9454
rect 15212 9450 15240 9551
rect 15200 9444 15252 9450
rect 15200 9386 15252 9392
rect 15212 9042 15240 9386
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15120 8634 15148 8910
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15016 8016 15068 8022
rect 15016 7958 15068 7964
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 14924 6928 14976 6934
rect 14924 6870 14976 6876
rect 14936 5846 14964 6870
rect 14924 5840 14976 5846
rect 14924 5782 14976 5788
rect 15028 4758 15056 7822
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 15016 4752 15068 4758
rect 15016 4694 15068 4700
rect 14832 4548 14884 4554
rect 14832 4490 14884 4496
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 12348 4140 12400 4146
rect 15120 4128 15148 7278
rect 15212 7177 15240 8842
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15304 7274 15332 7890
rect 15292 7268 15344 7274
rect 15292 7210 15344 7216
rect 15198 7168 15254 7177
rect 15198 7103 15254 7112
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 15212 4690 15240 6666
rect 15304 6662 15332 7210
rect 15396 6934 15424 8026
rect 15384 6928 15436 6934
rect 15384 6870 15436 6876
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15304 5846 15332 6598
rect 15292 5840 15344 5846
rect 15292 5782 15344 5788
rect 15488 5166 15516 11086
rect 15580 9654 15608 11206
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15566 9208 15622 9217
rect 15566 9143 15622 9152
rect 15580 8566 15608 9143
rect 15672 8974 15700 11698
rect 15764 11694 15792 12038
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15568 8560 15620 8566
rect 15568 8502 15620 8508
rect 15672 8498 15700 8910
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15658 8392 15714 8401
rect 15658 8327 15660 8336
rect 15712 8327 15714 8336
rect 15660 8298 15712 8304
rect 15660 7880 15712 7886
rect 15658 7848 15660 7857
rect 15712 7848 15714 7857
rect 15658 7783 15714 7792
rect 15568 5296 15620 5302
rect 15568 5238 15620 5244
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15488 4758 15516 5102
rect 15476 4752 15528 4758
rect 15476 4694 15528 4700
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 15120 4100 15240 4128
rect 12348 4082 12400 4088
rect 14289 3836 14585 3856
rect 14345 3834 14369 3836
rect 14425 3834 14449 3836
rect 14505 3834 14529 3836
rect 14367 3782 14369 3834
rect 14431 3782 14443 3834
rect 14505 3782 14507 3834
rect 14345 3780 14369 3782
rect 14425 3780 14449 3782
rect 14505 3780 14529 3782
rect 14289 3760 14585 3780
rect 14289 2748 14585 2768
rect 14345 2746 14369 2748
rect 14425 2746 14449 2748
rect 14505 2746 14529 2748
rect 14367 2694 14369 2746
rect 14431 2694 14443 2746
rect 14505 2694 14507 2746
rect 14345 2692 14369 2694
rect 14425 2692 14449 2694
rect 14505 2692 14529 2694
rect 14289 2672 14585 2692
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 11336 2304 11388 2310
rect 11336 2246 11388 2252
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 9508 1465 9536 2246
rect 10956 2204 11252 2224
rect 11012 2202 11036 2204
rect 11092 2202 11116 2204
rect 11172 2202 11196 2204
rect 11034 2150 11036 2202
rect 11098 2150 11110 2202
rect 11172 2150 11174 2202
rect 11012 2148 11036 2150
rect 11092 2148 11116 2150
rect 11172 2148 11196 2150
rect 10956 2128 11252 2148
rect 9494 1456 9550 1465
rect 9494 1391 9550 1400
rect 11348 377 11376 2246
rect 15212 1057 15240 4100
rect 15580 3097 15608 5238
rect 15764 4758 15792 11630
rect 15856 10130 15884 13330
rect 15948 12374 15976 16118
rect 16132 15910 16160 16594
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 16224 15570 16252 18022
rect 16408 17542 16436 18226
rect 16500 17882 16528 18770
rect 16580 18692 16632 18698
rect 16580 18634 16632 18640
rect 16488 17876 16540 17882
rect 16488 17818 16540 17824
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16304 17128 16356 17134
rect 16304 17070 16356 17076
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 16316 15366 16344 17070
rect 16408 16114 16436 17478
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16500 15570 16528 17818
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16394 15464 16450 15473
rect 16394 15399 16450 15408
rect 16304 15360 16356 15366
rect 16026 15328 16082 15337
rect 16304 15302 16356 15308
rect 16026 15263 16082 15272
rect 15936 12368 15988 12374
rect 16040 12356 16068 15263
rect 16408 15094 16436 15399
rect 16500 15162 16528 15506
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16396 15088 16448 15094
rect 16396 15030 16448 15036
rect 16210 14648 16266 14657
rect 16210 14583 16266 14592
rect 16224 14346 16252 14583
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16212 14340 16264 14346
rect 16212 14282 16264 14288
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16316 13530 16344 14010
rect 16500 13870 16528 14418
rect 16592 14074 16620 18634
rect 17622 18524 17918 18544
rect 17678 18522 17702 18524
rect 17758 18522 17782 18524
rect 17838 18522 17862 18524
rect 17700 18470 17702 18522
rect 17764 18470 17776 18522
rect 17838 18470 17840 18522
rect 17678 18468 17702 18470
rect 17758 18468 17782 18470
rect 17838 18468 17862 18470
rect 16854 18456 16910 18465
rect 17622 18448 17918 18468
rect 16854 18391 16910 18400
rect 16868 18222 16896 18391
rect 16856 18216 16908 18222
rect 16856 18158 16908 18164
rect 17622 17436 17918 17456
rect 17678 17434 17702 17436
rect 17758 17434 17782 17436
rect 17838 17434 17862 17436
rect 17700 17382 17702 17434
rect 17764 17382 17776 17434
rect 17838 17382 17840 17434
rect 17678 17380 17702 17382
rect 17758 17380 17782 17382
rect 17838 17380 17862 17382
rect 17622 17360 17918 17380
rect 17622 16348 17918 16368
rect 17678 16346 17702 16348
rect 17758 16346 17782 16348
rect 17838 16346 17862 16348
rect 17700 16294 17702 16346
rect 17764 16294 17776 16346
rect 17838 16294 17840 16346
rect 17678 16292 17702 16294
rect 17758 16292 17782 16294
rect 17838 16292 17862 16294
rect 17622 16272 17918 16292
rect 17040 15904 17092 15910
rect 16946 15872 17002 15881
rect 17040 15846 17092 15852
rect 16946 15807 17002 15816
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16672 14952 16724 14958
rect 16672 14894 16724 14900
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16592 13870 16620 14010
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16316 12986 16344 13466
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16118 12880 16174 12889
rect 16118 12815 16174 12824
rect 16132 12782 16160 12815
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16394 12608 16450 12617
rect 16394 12543 16450 12552
rect 16040 12328 16160 12356
rect 15936 12310 15988 12316
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 15948 11694 15976 12174
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 15948 10606 15976 11630
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 15856 8430 15884 8774
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 16040 7857 16068 12174
rect 16026 7848 16082 7857
rect 16026 7783 16082 7792
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 15856 6458 15884 6802
rect 15934 6760 15990 6769
rect 15934 6695 15990 6704
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 15752 4752 15804 4758
rect 15752 4694 15804 4700
rect 15948 4690 15976 6695
rect 16028 5908 16080 5914
rect 16028 5850 16080 5856
rect 16040 5681 16068 5850
rect 16026 5672 16082 5681
rect 16026 5607 16082 5616
rect 16132 5137 16160 12328
rect 16408 12170 16436 12543
rect 16396 12164 16448 12170
rect 16396 12106 16448 12112
rect 16304 11688 16356 11694
rect 16304 11630 16356 11636
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16224 10198 16252 10610
rect 16316 10606 16344 11630
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 16212 10192 16264 10198
rect 16212 10134 16264 10140
rect 16224 9110 16252 10134
rect 16316 9926 16344 10542
rect 16408 10266 16436 10950
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16316 9382 16344 9522
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16212 9104 16264 9110
rect 16212 9046 16264 9052
rect 16316 9042 16344 9318
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16316 7886 16344 8978
rect 16408 8634 16436 9386
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16500 7410 16528 13806
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 16592 11898 16620 12242
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 16592 10742 16620 11834
rect 16684 11830 16712 14894
rect 16868 14890 16896 15302
rect 16960 14958 16988 15807
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16856 14884 16908 14890
rect 16856 14826 16908 14832
rect 16868 14482 16896 14826
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16854 14376 16910 14385
rect 16854 14311 16910 14320
rect 16764 14000 16816 14006
rect 16764 13942 16816 13948
rect 16776 13297 16804 13942
rect 16868 13802 16896 14311
rect 16856 13796 16908 13802
rect 16856 13738 16908 13744
rect 16868 13530 16896 13738
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16762 13288 16818 13297
rect 16762 13223 16818 13232
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16776 12306 16804 12922
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16762 11928 16818 11937
rect 16960 11914 16988 12582
rect 16818 11886 16988 11914
rect 16762 11863 16818 11872
rect 16672 11824 16724 11830
rect 16672 11766 16724 11772
rect 16580 10736 16632 10742
rect 16580 10678 16632 10684
rect 16592 10266 16620 10678
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16592 9518 16620 10202
rect 16684 9602 16712 11766
rect 16776 11354 16804 11863
rect 17052 11812 17080 15846
rect 17622 15260 17918 15280
rect 17678 15258 17702 15260
rect 17758 15258 17782 15260
rect 17838 15258 17862 15260
rect 17700 15206 17702 15258
rect 17764 15206 17776 15258
rect 17838 15206 17840 15258
rect 17678 15204 17702 15206
rect 17758 15204 17782 15206
rect 17838 15204 17862 15206
rect 17622 15184 17918 15204
rect 17622 14172 17918 14192
rect 17678 14170 17702 14172
rect 17758 14170 17782 14172
rect 17838 14170 17862 14172
rect 17700 14118 17702 14170
rect 17764 14118 17776 14170
rect 17838 14118 17840 14170
rect 17678 14116 17702 14118
rect 17758 14116 17782 14118
rect 17838 14116 17862 14118
rect 17622 14096 17918 14116
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 17144 12986 17172 13806
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 16960 11784 17080 11812
rect 16764 11348 16816 11354
rect 16764 11290 16816 11296
rect 16684 9574 16804 9602
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16672 9444 16724 9450
rect 16672 9386 16724 9392
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16212 7336 16264 7342
rect 16212 7278 16264 7284
rect 16224 6730 16252 7278
rect 16500 6984 16528 7346
rect 16500 6956 16620 6984
rect 16212 6724 16264 6730
rect 16212 6666 16264 6672
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 16302 6080 16358 6089
rect 16302 6015 16358 6024
rect 16118 5128 16174 5137
rect 16118 5063 16174 5072
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 15948 4282 15976 4626
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 15566 3088 15622 3097
rect 15566 3023 15622 3032
rect 16316 1737 16344 6015
rect 16396 5636 16448 5642
rect 16396 5578 16448 5584
rect 16408 3777 16436 5578
rect 16394 3768 16450 3777
rect 16394 3703 16450 3712
rect 16500 2417 16528 6666
rect 16592 5778 16620 6956
rect 16684 6089 16712 9386
rect 16776 6254 16804 9574
rect 16960 6866 16988 11784
rect 17328 11558 17356 12242
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17328 10169 17356 11494
rect 17314 10160 17370 10169
rect 17314 10095 17370 10104
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 16948 6860 17000 6866
rect 16868 6820 16948 6848
rect 16764 6248 16816 6254
rect 16764 6190 16816 6196
rect 16670 6080 16726 6089
rect 16670 6015 16726 6024
rect 16868 5914 16896 6820
rect 16948 6802 17000 6808
rect 17052 6798 17080 9590
rect 17420 6866 17448 13874
rect 17622 13084 17918 13104
rect 17678 13082 17702 13084
rect 17758 13082 17782 13084
rect 17838 13082 17862 13084
rect 17700 13030 17702 13082
rect 17764 13030 17776 13082
rect 17838 13030 17840 13082
rect 17678 13028 17702 13030
rect 17758 13028 17782 13030
rect 17838 13028 17862 13030
rect 17622 13008 17918 13028
rect 17622 11996 17918 12016
rect 17678 11994 17702 11996
rect 17758 11994 17782 11996
rect 17838 11994 17862 11996
rect 17700 11942 17702 11994
rect 17764 11942 17776 11994
rect 17838 11942 17840 11994
rect 17678 11940 17702 11942
rect 17758 11940 17782 11942
rect 17838 11940 17862 11942
rect 17622 11920 17918 11940
rect 17622 10908 17918 10928
rect 17678 10906 17702 10908
rect 17758 10906 17782 10908
rect 17838 10906 17862 10908
rect 17700 10854 17702 10906
rect 17764 10854 17776 10906
rect 17838 10854 17840 10906
rect 17678 10852 17702 10854
rect 17758 10852 17782 10854
rect 17838 10852 17862 10854
rect 17622 10832 17918 10852
rect 17622 9820 17918 9840
rect 17678 9818 17702 9820
rect 17758 9818 17782 9820
rect 17838 9818 17862 9820
rect 17700 9766 17702 9818
rect 17764 9766 17776 9818
rect 17838 9766 17840 9818
rect 17678 9764 17702 9766
rect 17758 9764 17782 9766
rect 17838 9764 17862 9766
rect 17622 9744 17918 9764
rect 17622 8732 17918 8752
rect 17678 8730 17702 8732
rect 17758 8730 17782 8732
rect 17838 8730 17862 8732
rect 17700 8678 17702 8730
rect 17764 8678 17776 8730
rect 17838 8678 17840 8730
rect 17678 8676 17702 8678
rect 17758 8676 17782 8678
rect 17838 8676 17862 8678
rect 17622 8656 17918 8676
rect 17622 7644 17918 7664
rect 17678 7642 17702 7644
rect 17758 7642 17782 7644
rect 17838 7642 17862 7644
rect 17700 7590 17702 7642
rect 17764 7590 17776 7642
rect 17838 7590 17840 7642
rect 17678 7588 17702 7590
rect 17758 7588 17782 7590
rect 17838 7588 17862 7590
rect 17622 7568 17918 7588
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 17406 6760 17462 6769
rect 17052 6474 17080 6734
rect 17406 6695 17408 6704
rect 17460 6695 17462 6704
rect 17408 6666 17460 6672
rect 16960 6458 17080 6474
rect 16948 6452 17080 6458
rect 17000 6446 17080 6452
rect 16948 6394 17000 6400
rect 17040 6384 17092 6390
rect 17040 6326 17092 6332
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16580 5772 16632 5778
rect 16580 5714 16632 5720
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 16592 5370 16620 5714
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 16960 4826 16988 5714
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 17052 4593 17080 6326
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 17144 5778 17172 6258
rect 17316 6248 17368 6254
rect 17420 6236 17448 6666
rect 17622 6556 17918 6576
rect 17678 6554 17702 6556
rect 17758 6554 17782 6556
rect 17838 6554 17862 6556
rect 17700 6502 17702 6554
rect 17764 6502 17776 6554
rect 17838 6502 17840 6554
rect 17678 6500 17702 6502
rect 17758 6500 17782 6502
rect 17838 6500 17862 6502
rect 17622 6480 17918 6500
rect 17500 6248 17552 6254
rect 17420 6208 17500 6236
rect 17316 6190 17368 6196
rect 17500 6190 17552 6196
rect 17328 5914 17356 6190
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 17144 5302 17172 5714
rect 17622 5468 17918 5488
rect 17678 5466 17702 5468
rect 17758 5466 17782 5468
rect 17838 5466 17862 5468
rect 17700 5414 17702 5466
rect 17764 5414 17776 5466
rect 17838 5414 17840 5466
rect 17678 5412 17702 5414
rect 17758 5412 17782 5414
rect 17838 5412 17862 5414
rect 17622 5392 17918 5412
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 17038 4584 17094 4593
rect 17038 4519 17094 4528
rect 17622 4380 17918 4400
rect 17678 4378 17702 4380
rect 17758 4378 17782 4380
rect 17838 4378 17862 4380
rect 17700 4326 17702 4378
rect 17764 4326 17776 4378
rect 17838 4326 17840 4378
rect 17678 4324 17702 4326
rect 17758 4324 17782 4326
rect 17838 4324 17862 4326
rect 17622 4304 17918 4324
rect 17622 3292 17918 3312
rect 17678 3290 17702 3292
rect 17758 3290 17782 3292
rect 17838 3290 17862 3292
rect 17700 3238 17702 3290
rect 17764 3238 17776 3290
rect 17838 3238 17840 3290
rect 17678 3236 17702 3238
rect 17758 3236 17782 3238
rect 17838 3236 17862 3238
rect 17622 3216 17918 3236
rect 16486 2408 16542 2417
rect 16486 2343 16542 2352
rect 17622 2204 17918 2224
rect 17678 2202 17702 2204
rect 17758 2202 17782 2204
rect 17838 2202 17862 2204
rect 17700 2150 17702 2202
rect 17764 2150 17776 2202
rect 17838 2150 17840 2202
rect 17678 2148 17702 2150
rect 17758 2148 17782 2150
rect 17838 2148 17862 2150
rect 17622 2128 17918 2148
rect 16302 1728 16358 1737
rect 16302 1663 16358 1672
rect 15198 1048 15254 1057
rect 15198 983 15254 992
rect 9310 368 9366 377
rect 9310 303 9366 312
rect 11334 368 11390 377
rect 11334 303 11390 312
<< via2 >>
rect 3606 79464 3662 79520
rect 2870 77832 2926 77888
rect 2134 77016 2190 77072
rect 2870 72256 2926 72312
rect 2870 69400 2926 69456
rect 2042 68992 2098 69048
rect 1306 67360 1362 67416
rect 1674 66680 1730 66736
rect 1766 65048 1822 65104
rect 1490 62600 1546 62656
rect 1490 60968 1546 61024
rect 1582 60288 1638 60344
rect 1398 59472 1454 59528
rect 1306 47368 1362 47424
rect 1582 57024 1638 57080
rect 1950 61784 2006 61840
rect 2962 69264 3018 69320
rect 2134 63416 2190 63472
rect 1858 53760 1914 53816
rect 1674 52572 1676 52592
rect 1676 52572 1728 52592
rect 1728 52572 1730 52592
rect 1674 52536 1730 52572
rect 1858 52264 1914 52320
rect 1490 51448 1546 51504
rect 1582 46960 1638 47016
rect 1766 45872 1822 45928
rect 1490 44240 1546 44296
rect 1582 43424 1638 43480
rect 1490 41792 1546 41848
rect 1582 41420 1584 41440
rect 1584 41420 1636 41440
rect 1636 41420 1638 41440
rect 1582 41384 1638 41420
rect 1582 40332 1584 40352
rect 1584 40332 1636 40352
rect 1636 40332 1638 40352
rect 1582 40296 1638 40332
rect 1950 49000 2006 49056
rect 2502 63416 2558 63472
rect 2502 63280 2558 63336
rect 2870 64232 2926 64288
rect 2686 63860 2688 63880
rect 2688 63860 2740 63880
rect 2740 63860 2742 63880
rect 2686 63824 2742 63860
rect 3054 69164 3056 69184
rect 3056 69164 3108 69184
rect 3108 69164 3110 69184
rect 3054 69128 3110 69164
rect 2686 60424 2742 60480
rect 2318 58112 2374 58168
rect 2502 60152 2558 60208
rect 3422 75384 3478 75440
rect 2318 54576 2374 54632
rect 2226 49680 2282 49736
rect 2134 48592 2190 48648
rect 2594 59608 2650 59664
rect 2502 49952 2558 50008
rect 2502 45872 2558 45928
rect 1950 42644 1952 42664
rect 1952 42644 2004 42664
rect 2004 42644 2006 42664
rect 1950 42608 2006 42644
rect 2410 45056 2466 45112
rect 2134 39480 2190 39536
rect 1858 36216 1914 36272
rect 1490 35400 1546 35456
rect 1398 33496 1454 33552
rect 1582 33768 1638 33824
rect 1582 32000 1638 32056
rect 1858 32272 1914 32328
rect 1766 31728 1822 31784
rect 1950 31864 2006 31920
rect 1582 30640 1638 30696
rect 1674 29824 1730 29880
rect 1582 28212 1638 28248
rect 1582 28192 1584 28212
rect 1584 28192 1636 28212
rect 1636 28192 1638 28212
rect 1674 28076 1730 28112
rect 1674 28056 1676 28076
rect 1676 28056 1728 28076
rect 1728 28056 1730 28076
rect 1582 26696 1638 26752
rect 1766 24792 1822 24848
rect 2134 29996 2136 30016
rect 2136 29996 2188 30016
rect 2188 29996 2190 30016
rect 2134 29960 2190 29996
rect 2134 29008 2190 29064
rect 1950 28500 1952 28520
rect 1952 28500 2004 28520
rect 2004 28500 2006 28520
rect 1950 28464 2006 28500
rect 2134 24248 2190 24304
rect 1674 22616 1730 22672
rect 1490 21800 1546 21856
rect 1766 19488 1822 19544
rect 1398 18672 1454 18728
rect 1674 17196 1730 17232
rect 1674 17176 1676 17196
rect 1676 17176 1728 17196
rect 1728 17176 1730 17196
rect 1214 15408 1270 15464
rect 1582 13096 1638 13152
rect 2318 34620 2320 34640
rect 2320 34620 2372 34640
rect 2372 34620 2374 34640
rect 2318 34584 2374 34620
rect 2502 43968 2558 44024
rect 2870 53080 2926 53136
rect 2778 51756 2780 51776
rect 2780 51756 2832 51776
rect 2832 51756 2834 51776
rect 2778 51720 2834 51756
rect 2870 49680 2926 49736
rect 2778 48184 2834 48240
rect 2686 40568 2742 40624
rect 2686 39344 2742 39400
rect 2594 38392 2650 38448
rect 3146 61104 3202 61160
rect 3054 57332 3056 57352
rect 3056 57332 3108 57352
rect 3108 57332 3110 57352
rect 3054 57296 3110 57332
rect 3146 52672 3202 52728
rect 3054 49816 3110 49872
rect 2870 47232 2926 47288
rect 2870 42744 2926 42800
rect 2870 41520 2926 41576
rect 2870 33088 2926 33144
rect 2778 25880 2834 25936
rect 2962 19760 3018 19816
rect 2778 17040 2834 17096
rect 2594 16224 2650 16280
rect 16026 78784 16082 78840
rect 3790 78668 3846 78704
rect 3790 78648 3792 78668
rect 3792 78648 3844 78668
rect 3844 78648 3846 78668
rect 4289 77274 4345 77276
rect 4369 77274 4425 77276
rect 4449 77274 4505 77276
rect 4529 77274 4585 77276
rect 4289 77222 4315 77274
rect 4315 77222 4345 77274
rect 4369 77222 4379 77274
rect 4379 77222 4425 77274
rect 4449 77222 4495 77274
rect 4495 77222 4505 77274
rect 4529 77222 4559 77274
rect 4559 77222 4585 77274
rect 4289 77220 4345 77222
rect 4369 77220 4425 77222
rect 4449 77220 4505 77222
rect 4529 77220 4585 77222
rect 4066 76200 4122 76256
rect 4289 76186 4345 76188
rect 4369 76186 4425 76188
rect 4449 76186 4505 76188
rect 4529 76186 4585 76188
rect 4289 76134 4315 76186
rect 4315 76134 4345 76186
rect 4369 76134 4379 76186
rect 4379 76134 4425 76186
rect 4449 76134 4495 76186
rect 4495 76134 4505 76186
rect 4529 76134 4559 76186
rect 4559 76134 4585 76186
rect 4289 76132 4345 76134
rect 4369 76132 4425 76134
rect 4449 76132 4505 76134
rect 4529 76132 4585 76134
rect 4289 75098 4345 75100
rect 4369 75098 4425 75100
rect 4449 75098 4505 75100
rect 4529 75098 4585 75100
rect 4289 75046 4315 75098
rect 4315 75046 4345 75098
rect 4369 75046 4379 75098
rect 4379 75046 4425 75098
rect 4449 75046 4495 75098
rect 4495 75046 4505 75098
rect 4529 75046 4559 75098
rect 4559 75046 4585 75098
rect 4289 75044 4345 75046
rect 4369 75044 4425 75046
rect 4449 75044 4505 75046
rect 4529 75044 4585 75046
rect 15934 78104 15990 78160
rect 7622 77818 7678 77820
rect 7702 77818 7758 77820
rect 7782 77818 7838 77820
rect 7862 77818 7918 77820
rect 7622 77766 7648 77818
rect 7648 77766 7678 77818
rect 7702 77766 7712 77818
rect 7712 77766 7758 77818
rect 7782 77766 7828 77818
rect 7828 77766 7838 77818
rect 7862 77766 7892 77818
rect 7892 77766 7918 77818
rect 7622 77764 7678 77766
rect 7702 77764 7758 77766
rect 7782 77764 7838 77766
rect 7862 77764 7918 77766
rect 14289 77818 14345 77820
rect 14369 77818 14425 77820
rect 14449 77818 14505 77820
rect 14529 77818 14585 77820
rect 14289 77766 14315 77818
rect 14315 77766 14345 77818
rect 14369 77766 14379 77818
rect 14379 77766 14425 77818
rect 14449 77766 14495 77818
rect 14495 77766 14505 77818
rect 14529 77766 14559 77818
rect 14559 77766 14585 77818
rect 14289 77764 14345 77766
rect 14369 77764 14425 77766
rect 14449 77764 14505 77766
rect 14529 77764 14585 77766
rect 10956 77274 11012 77276
rect 11036 77274 11092 77276
rect 11116 77274 11172 77276
rect 11196 77274 11252 77276
rect 10956 77222 10982 77274
rect 10982 77222 11012 77274
rect 11036 77222 11046 77274
rect 11046 77222 11092 77274
rect 11116 77222 11162 77274
rect 11162 77222 11172 77274
rect 11196 77222 11226 77274
rect 11226 77222 11252 77274
rect 10956 77220 11012 77222
rect 11036 77220 11092 77222
rect 11116 77220 11172 77222
rect 11196 77220 11252 77222
rect 17622 77274 17678 77276
rect 17702 77274 17758 77276
rect 17782 77274 17838 77276
rect 17862 77274 17918 77276
rect 17622 77222 17648 77274
rect 17648 77222 17678 77274
rect 17702 77222 17712 77274
rect 17712 77222 17758 77274
rect 17782 77222 17828 77274
rect 17828 77222 17838 77274
rect 17862 77222 17892 77274
rect 17892 77222 17918 77274
rect 17622 77220 17678 77222
rect 17702 77220 17758 77222
rect 17782 77220 17838 77222
rect 17862 77220 17918 77222
rect 7622 76730 7678 76732
rect 7702 76730 7758 76732
rect 7782 76730 7838 76732
rect 7862 76730 7918 76732
rect 7622 76678 7648 76730
rect 7648 76678 7678 76730
rect 7702 76678 7712 76730
rect 7712 76678 7758 76730
rect 7782 76678 7828 76730
rect 7828 76678 7838 76730
rect 7862 76678 7892 76730
rect 7892 76678 7918 76730
rect 7622 76676 7678 76678
rect 7702 76676 7758 76678
rect 7782 76676 7838 76678
rect 7862 76676 7918 76678
rect 14289 76730 14345 76732
rect 14369 76730 14425 76732
rect 14449 76730 14505 76732
rect 14529 76730 14585 76732
rect 14289 76678 14315 76730
rect 14315 76678 14345 76730
rect 14369 76678 14379 76730
rect 14379 76678 14425 76730
rect 14449 76678 14495 76730
rect 14495 76678 14505 76730
rect 14529 76678 14559 76730
rect 14559 76678 14585 76730
rect 14289 76676 14345 76678
rect 14369 76676 14425 76678
rect 14449 76676 14505 76678
rect 14529 76676 14585 76678
rect 10956 76186 11012 76188
rect 11036 76186 11092 76188
rect 11116 76186 11172 76188
rect 11196 76186 11252 76188
rect 10956 76134 10982 76186
rect 10982 76134 11012 76186
rect 11036 76134 11046 76186
rect 11046 76134 11092 76186
rect 11116 76134 11162 76186
rect 11162 76134 11172 76186
rect 11196 76134 11226 76186
rect 11226 76134 11252 76186
rect 10956 76132 11012 76134
rect 11036 76132 11092 76134
rect 11116 76132 11172 76134
rect 11196 76132 11252 76134
rect 17622 76186 17678 76188
rect 17702 76186 17758 76188
rect 17782 76186 17838 76188
rect 17862 76186 17918 76188
rect 17622 76134 17648 76186
rect 17648 76134 17678 76186
rect 17702 76134 17712 76186
rect 17712 76134 17758 76186
rect 17782 76134 17828 76186
rect 17828 76134 17838 76186
rect 17862 76134 17892 76186
rect 17892 76134 17918 76186
rect 17622 76132 17678 76134
rect 17702 76132 17758 76134
rect 17782 76132 17838 76134
rect 17862 76132 17918 76134
rect 7622 75642 7678 75644
rect 7702 75642 7758 75644
rect 7782 75642 7838 75644
rect 7862 75642 7918 75644
rect 7622 75590 7648 75642
rect 7648 75590 7678 75642
rect 7702 75590 7712 75642
rect 7712 75590 7758 75642
rect 7782 75590 7828 75642
rect 7828 75590 7838 75642
rect 7862 75590 7892 75642
rect 7892 75590 7918 75642
rect 7622 75588 7678 75590
rect 7702 75588 7758 75590
rect 7782 75588 7838 75590
rect 7862 75588 7918 75590
rect 14289 75642 14345 75644
rect 14369 75642 14425 75644
rect 14449 75642 14505 75644
rect 14529 75642 14585 75644
rect 14289 75590 14315 75642
rect 14315 75590 14345 75642
rect 14369 75590 14379 75642
rect 14379 75590 14425 75642
rect 14449 75590 14495 75642
rect 14495 75590 14505 75642
rect 14529 75590 14559 75642
rect 14559 75590 14585 75642
rect 14289 75588 14345 75590
rect 14369 75588 14425 75590
rect 14449 75588 14505 75590
rect 14529 75588 14585 75590
rect 4894 75284 4896 75304
rect 4896 75284 4948 75304
rect 4948 75284 4950 75304
rect 4894 75248 4950 75284
rect 7010 75248 7066 75304
rect 3882 73344 3938 73400
rect 4618 74568 4674 74624
rect 4289 74010 4345 74012
rect 4369 74010 4425 74012
rect 4449 74010 4505 74012
rect 4529 74010 4585 74012
rect 4289 73958 4315 74010
rect 4315 73958 4345 74010
rect 4369 73958 4379 74010
rect 4379 73958 4425 74010
rect 4449 73958 4495 74010
rect 4495 73958 4505 74010
rect 4529 73958 4559 74010
rect 4559 73958 4585 74010
rect 4289 73956 4345 73958
rect 4369 73956 4425 73958
rect 4449 73956 4505 73958
rect 4529 73956 4585 73958
rect 4342 73228 4398 73264
rect 4342 73208 4344 73228
rect 4344 73208 4396 73228
rect 4396 73208 4398 73228
rect 4250 73072 4306 73128
rect 4289 72922 4345 72924
rect 4369 72922 4425 72924
rect 4449 72922 4505 72924
rect 4529 72922 4585 72924
rect 4289 72870 4315 72922
rect 4315 72870 4345 72922
rect 4369 72870 4379 72922
rect 4379 72870 4425 72922
rect 4449 72870 4495 72922
rect 4495 72870 4505 72922
rect 4529 72870 4559 72922
rect 4559 72870 4585 72922
rect 4289 72868 4345 72870
rect 4369 72868 4425 72870
rect 4449 72868 4505 72870
rect 4529 72868 4585 72870
rect 4802 73752 4858 73808
rect 3698 71340 3700 71360
rect 3700 71340 3752 71360
rect 3752 71340 3754 71360
rect 3698 71304 3754 71340
rect 4289 71834 4345 71836
rect 4369 71834 4425 71836
rect 4449 71834 4505 71836
rect 4529 71834 4585 71836
rect 4289 71782 4315 71834
rect 4315 71782 4345 71834
rect 4369 71782 4379 71834
rect 4379 71782 4425 71834
rect 4449 71782 4495 71834
rect 4495 71782 4505 71834
rect 4529 71782 4559 71834
rect 4559 71782 4585 71834
rect 4289 71780 4345 71782
rect 4369 71780 4425 71782
rect 4449 71780 4505 71782
rect 4529 71780 4585 71782
rect 4289 70746 4345 70748
rect 4369 70746 4425 70748
rect 4449 70746 4505 70748
rect 4529 70746 4585 70748
rect 4289 70694 4315 70746
rect 4315 70694 4345 70746
rect 4369 70694 4379 70746
rect 4379 70694 4425 70746
rect 4449 70694 4495 70746
rect 4495 70694 4505 70746
rect 4529 70694 4559 70746
rect 4559 70694 4585 70746
rect 4289 70692 4345 70694
rect 4369 70692 4425 70694
rect 4449 70692 4505 70694
rect 4529 70692 4585 70694
rect 4710 70352 4766 70408
rect 3974 69808 4030 69864
rect 3606 68992 3662 69048
rect 3514 65864 3570 65920
rect 3330 60560 3386 60616
rect 3238 49136 3294 49192
rect 3238 46688 3294 46744
rect 3238 45872 3294 45928
rect 3238 43288 3294 43344
rect 3422 59372 3424 59392
rect 3424 59372 3476 59392
rect 3476 59372 3478 59392
rect 3422 59336 3478 59372
rect 4289 69658 4345 69660
rect 4369 69658 4425 69660
rect 4449 69658 4505 69660
rect 4529 69658 4585 69660
rect 4289 69606 4315 69658
rect 4315 69606 4345 69658
rect 4369 69606 4379 69658
rect 4379 69606 4425 69658
rect 4449 69606 4495 69658
rect 4495 69606 4505 69658
rect 4529 69606 4559 69658
rect 4559 69606 4585 69658
rect 4289 69604 4345 69606
rect 4369 69604 4425 69606
rect 4449 69604 4505 69606
rect 4529 69604 4585 69606
rect 4710 69536 4766 69592
rect 4289 68570 4345 68572
rect 4369 68570 4425 68572
rect 4449 68570 4505 68572
rect 4529 68570 4585 68572
rect 4289 68518 4315 68570
rect 4315 68518 4345 68570
rect 4369 68518 4379 68570
rect 4379 68518 4425 68570
rect 4449 68518 4495 68570
rect 4495 68518 4505 68570
rect 4529 68518 4559 68570
rect 4559 68518 4585 68570
rect 4289 68516 4345 68518
rect 4369 68516 4425 68518
rect 4449 68516 4505 68518
rect 4529 68516 4585 68518
rect 4158 68176 4214 68232
rect 4066 63996 4068 64016
rect 4068 63996 4120 64016
rect 4120 63996 4122 64016
rect 4066 63960 4122 63996
rect 4289 67482 4345 67484
rect 4369 67482 4425 67484
rect 4449 67482 4505 67484
rect 4529 67482 4585 67484
rect 4289 67430 4315 67482
rect 4315 67430 4345 67482
rect 4369 67430 4379 67482
rect 4379 67430 4425 67482
rect 4449 67430 4495 67482
rect 4495 67430 4505 67482
rect 4529 67430 4559 67482
rect 4559 67430 4585 67482
rect 4289 67428 4345 67430
rect 4369 67428 4425 67430
rect 4449 67428 4505 67430
rect 4529 67428 4585 67430
rect 4289 66394 4345 66396
rect 4369 66394 4425 66396
rect 4449 66394 4505 66396
rect 4529 66394 4585 66396
rect 4289 66342 4315 66394
rect 4315 66342 4345 66394
rect 4369 66342 4379 66394
rect 4379 66342 4425 66394
rect 4449 66342 4495 66394
rect 4495 66342 4505 66394
rect 4529 66342 4559 66394
rect 4559 66342 4585 66394
rect 4289 66340 4345 66342
rect 4369 66340 4425 66342
rect 4449 66340 4505 66342
rect 4529 66340 4585 66342
rect 4710 68720 4766 68776
rect 4289 65306 4345 65308
rect 4369 65306 4425 65308
rect 4449 65306 4505 65308
rect 4529 65306 4585 65308
rect 4289 65254 4315 65306
rect 4315 65254 4345 65306
rect 4369 65254 4379 65306
rect 4379 65254 4425 65306
rect 4449 65254 4495 65306
rect 4495 65254 4505 65306
rect 4529 65254 4559 65306
rect 4559 65254 4585 65306
rect 4289 65252 4345 65254
rect 4369 65252 4425 65254
rect 4449 65252 4505 65254
rect 4529 65252 4585 65254
rect 5078 73652 5080 73672
rect 5080 73652 5132 73672
rect 5132 73652 5134 73672
rect 5078 73616 5134 73652
rect 5998 73344 6054 73400
rect 5078 68740 5134 68776
rect 5078 68720 5080 68740
rect 5080 68720 5132 68740
rect 5132 68720 5134 68740
rect 4289 64218 4345 64220
rect 4369 64218 4425 64220
rect 4449 64218 4505 64220
rect 4529 64218 4585 64220
rect 4289 64166 4315 64218
rect 4315 64166 4345 64218
rect 4369 64166 4379 64218
rect 4379 64166 4425 64218
rect 4449 64166 4495 64218
rect 4495 64166 4505 64218
rect 4529 64166 4559 64218
rect 4559 64166 4585 64218
rect 4289 64164 4345 64166
rect 4369 64164 4425 64166
rect 4449 64164 4505 64166
rect 4529 64164 4585 64166
rect 4158 63824 4214 63880
rect 4526 63316 4528 63336
rect 4528 63316 4580 63336
rect 4580 63316 4582 63336
rect 4526 63280 4582 63316
rect 4289 63130 4345 63132
rect 4369 63130 4425 63132
rect 4449 63130 4505 63132
rect 4529 63130 4585 63132
rect 4289 63078 4315 63130
rect 4315 63078 4345 63130
rect 4369 63078 4379 63130
rect 4379 63078 4425 63130
rect 4449 63078 4495 63130
rect 4495 63078 4505 63130
rect 4529 63078 4559 63130
rect 4559 63078 4585 63130
rect 4289 63076 4345 63078
rect 4369 63076 4425 63078
rect 4449 63076 4505 63078
rect 4529 63076 4585 63078
rect 3790 61104 3846 61160
rect 3790 60560 3846 60616
rect 3698 60052 3700 60072
rect 3700 60052 3752 60072
rect 3752 60052 3754 60072
rect 3698 60016 3754 60052
rect 3698 56208 3754 56264
rect 3514 51720 3570 51776
rect 3606 51312 3662 51368
rect 3422 48184 3478 48240
rect 3606 46008 3662 46064
rect 3790 42744 3846 42800
rect 3698 40180 3754 40216
rect 3698 40160 3700 40180
rect 3700 40160 3752 40180
rect 3752 40160 3754 40180
rect 3238 38256 3294 38312
rect 3514 37848 3570 37904
rect 3422 36760 3478 36816
rect 3790 37032 3846 37088
rect 3974 57840 4030 57896
rect 4289 62042 4345 62044
rect 4369 62042 4425 62044
rect 4449 62042 4505 62044
rect 4529 62042 4585 62044
rect 4289 61990 4315 62042
rect 4315 61990 4345 62042
rect 4369 61990 4379 62042
rect 4379 61990 4425 62042
rect 4449 61990 4495 62042
rect 4495 61990 4505 62042
rect 4529 61990 4559 62042
rect 4559 61990 4585 62042
rect 4289 61988 4345 61990
rect 4369 61988 4425 61990
rect 4449 61988 4505 61990
rect 4529 61988 4585 61990
rect 4289 60954 4345 60956
rect 4369 60954 4425 60956
rect 4449 60954 4505 60956
rect 4529 60954 4585 60956
rect 4289 60902 4315 60954
rect 4315 60902 4345 60954
rect 4369 60902 4379 60954
rect 4379 60902 4425 60954
rect 4449 60902 4495 60954
rect 4495 60902 4505 60954
rect 4529 60902 4559 60954
rect 4559 60902 4585 60954
rect 4289 60900 4345 60902
rect 4369 60900 4425 60902
rect 4449 60900 4505 60902
rect 4529 60900 4585 60902
rect 4342 60460 4344 60480
rect 4344 60460 4396 60480
rect 4396 60460 4398 60480
rect 4342 60424 4398 60460
rect 4289 59866 4345 59868
rect 4369 59866 4425 59868
rect 4449 59866 4505 59868
rect 4529 59866 4585 59868
rect 4289 59814 4315 59866
rect 4315 59814 4345 59866
rect 4369 59814 4379 59866
rect 4379 59814 4425 59866
rect 4449 59814 4495 59866
rect 4495 59814 4505 59866
rect 4529 59814 4559 59866
rect 4559 59814 4585 59866
rect 4289 59812 4345 59814
rect 4369 59812 4425 59814
rect 4449 59812 4505 59814
rect 4529 59812 4585 59814
rect 4618 59200 4674 59256
rect 4289 58778 4345 58780
rect 4369 58778 4425 58780
rect 4449 58778 4505 58780
rect 4529 58778 4585 58780
rect 4289 58726 4315 58778
rect 4315 58726 4345 58778
rect 4369 58726 4379 58778
rect 4379 58726 4425 58778
rect 4449 58726 4495 58778
rect 4495 58726 4505 58778
rect 4529 58726 4559 58778
rect 4559 58726 4585 58778
rect 4289 58724 4345 58726
rect 4369 58724 4425 58726
rect 4449 58724 4505 58726
rect 4529 58724 4585 58726
rect 4289 57690 4345 57692
rect 4369 57690 4425 57692
rect 4449 57690 4505 57692
rect 4529 57690 4585 57692
rect 4289 57638 4315 57690
rect 4315 57638 4345 57690
rect 4369 57638 4379 57690
rect 4379 57638 4425 57690
rect 4449 57638 4495 57690
rect 4495 57638 4505 57690
rect 4529 57638 4559 57690
rect 4559 57638 4585 57690
rect 4289 57636 4345 57638
rect 4369 57636 4425 57638
rect 4449 57636 4505 57638
rect 4529 57636 4585 57638
rect 4289 56602 4345 56604
rect 4369 56602 4425 56604
rect 4449 56602 4505 56604
rect 4529 56602 4585 56604
rect 4289 56550 4315 56602
rect 4315 56550 4345 56602
rect 4369 56550 4379 56602
rect 4379 56550 4425 56602
rect 4449 56550 4495 56602
rect 4495 56550 4505 56602
rect 4529 56550 4559 56602
rect 4559 56550 4585 56602
rect 4289 56548 4345 56550
rect 4369 56548 4425 56550
rect 4449 56548 4505 56550
rect 4529 56548 4585 56550
rect 4802 56208 4858 56264
rect 4289 55514 4345 55516
rect 4369 55514 4425 55516
rect 4449 55514 4505 55516
rect 4529 55514 4585 55516
rect 4289 55462 4315 55514
rect 4315 55462 4345 55514
rect 4369 55462 4379 55514
rect 4379 55462 4425 55514
rect 4449 55462 4495 55514
rect 4495 55462 4505 55514
rect 4529 55462 4559 55514
rect 4559 55462 4585 55514
rect 4289 55460 4345 55462
rect 4369 55460 4425 55462
rect 4449 55460 4505 55462
rect 4529 55460 4585 55462
rect 4434 55020 4436 55040
rect 4436 55020 4488 55040
rect 4488 55020 4490 55040
rect 4434 54984 4490 55020
rect 4289 54426 4345 54428
rect 4369 54426 4425 54428
rect 4449 54426 4505 54428
rect 4529 54426 4585 54428
rect 4289 54374 4315 54426
rect 4315 54374 4345 54426
rect 4369 54374 4379 54426
rect 4379 54374 4425 54426
rect 4449 54374 4495 54426
rect 4495 54374 4505 54426
rect 4529 54374 4559 54426
rect 4559 54374 4585 54426
rect 4289 54372 4345 54374
rect 4369 54372 4425 54374
rect 4449 54372 4505 54374
rect 4529 54372 4585 54374
rect 4342 53508 4398 53544
rect 4342 53488 4344 53508
rect 4344 53488 4396 53508
rect 4396 53488 4398 53508
rect 4289 53338 4345 53340
rect 4369 53338 4425 53340
rect 4449 53338 4505 53340
rect 4529 53338 4585 53340
rect 4289 53286 4315 53338
rect 4315 53286 4345 53338
rect 4369 53286 4379 53338
rect 4379 53286 4425 53338
rect 4449 53286 4495 53338
rect 4495 53286 4505 53338
rect 4529 53286 4559 53338
rect 4559 53286 4585 53338
rect 4289 53284 4345 53286
rect 4369 53284 4425 53286
rect 4449 53284 4505 53286
rect 4529 53284 4585 53286
rect 4526 53080 4582 53136
rect 4289 52250 4345 52252
rect 4369 52250 4425 52252
rect 4449 52250 4505 52252
rect 4529 52250 4585 52252
rect 4289 52198 4315 52250
rect 4315 52198 4345 52250
rect 4369 52198 4379 52250
rect 4379 52198 4425 52250
rect 4449 52198 4495 52250
rect 4495 52198 4505 52250
rect 4529 52198 4559 52250
rect 4559 52198 4585 52250
rect 4289 52196 4345 52198
rect 4369 52196 4425 52198
rect 4449 52196 4505 52198
rect 4529 52196 4585 52198
rect 4289 51162 4345 51164
rect 4369 51162 4425 51164
rect 4449 51162 4505 51164
rect 4529 51162 4585 51164
rect 4289 51110 4315 51162
rect 4315 51110 4345 51162
rect 4369 51110 4379 51162
rect 4379 51110 4425 51162
rect 4449 51110 4495 51162
rect 4495 51110 4505 51162
rect 4529 51110 4559 51162
rect 4559 51110 4585 51162
rect 4289 51108 4345 51110
rect 4369 51108 4425 51110
rect 4449 51108 4505 51110
rect 4529 51108 4585 51110
rect 5354 69128 5410 69184
rect 5262 67088 5318 67144
rect 4986 60560 5042 60616
rect 4986 58792 5042 58848
rect 5078 56072 5134 56128
rect 5446 66136 5502 66192
rect 5446 63960 5502 64016
rect 5630 63416 5686 63472
rect 5170 52128 5226 52184
rect 4710 51040 4766 51096
rect 4066 50224 4122 50280
rect 4289 50074 4345 50076
rect 4369 50074 4425 50076
rect 4449 50074 4505 50076
rect 4529 50074 4585 50076
rect 4289 50022 4315 50074
rect 4315 50022 4345 50074
rect 4369 50022 4379 50074
rect 4379 50022 4425 50074
rect 4449 50022 4495 50074
rect 4495 50022 4505 50074
rect 4529 50022 4559 50074
rect 4559 50022 4585 50074
rect 4289 50020 4345 50022
rect 4369 50020 4425 50022
rect 4449 50020 4505 50022
rect 4529 50020 4585 50022
rect 4289 48986 4345 48988
rect 4369 48986 4425 48988
rect 4449 48986 4505 48988
rect 4529 48986 4585 48988
rect 4289 48934 4315 48986
rect 4315 48934 4345 48986
rect 4369 48934 4379 48986
rect 4379 48934 4425 48986
rect 4449 48934 4495 48986
rect 4495 48934 4505 48986
rect 4529 48934 4559 48986
rect 4559 48934 4585 48986
rect 4289 48932 4345 48934
rect 4369 48932 4425 48934
rect 4449 48932 4505 48934
rect 4529 48932 4585 48934
rect 4289 47898 4345 47900
rect 4369 47898 4425 47900
rect 4449 47898 4505 47900
rect 4529 47898 4585 47900
rect 4289 47846 4315 47898
rect 4315 47846 4345 47898
rect 4369 47846 4379 47898
rect 4379 47846 4425 47898
rect 4449 47846 4495 47898
rect 4495 47846 4505 47898
rect 4529 47846 4559 47898
rect 4559 47846 4585 47898
rect 4289 47844 4345 47846
rect 4369 47844 4425 47846
rect 4449 47844 4505 47846
rect 4529 47844 4585 47846
rect 4158 47504 4214 47560
rect 3974 44376 4030 44432
rect 4289 46810 4345 46812
rect 4369 46810 4425 46812
rect 4449 46810 4505 46812
rect 4529 46810 4585 46812
rect 4289 46758 4315 46810
rect 4315 46758 4345 46810
rect 4369 46758 4379 46810
rect 4379 46758 4425 46810
rect 4449 46758 4495 46810
rect 4495 46758 4505 46810
rect 4529 46758 4559 46810
rect 4559 46758 4585 46810
rect 4289 46756 4345 46758
rect 4369 46756 4425 46758
rect 4449 46756 4505 46758
rect 4529 46756 4585 46758
rect 4526 46572 4582 46608
rect 4526 46552 4528 46572
rect 4528 46552 4580 46572
rect 4580 46552 4582 46572
rect 4289 45722 4345 45724
rect 4369 45722 4425 45724
rect 4449 45722 4505 45724
rect 4529 45722 4585 45724
rect 4289 45670 4315 45722
rect 4315 45670 4345 45722
rect 4369 45670 4379 45722
rect 4379 45670 4425 45722
rect 4449 45670 4495 45722
rect 4495 45670 4505 45722
rect 4529 45670 4559 45722
rect 4559 45670 4585 45722
rect 4289 45668 4345 45670
rect 4369 45668 4425 45670
rect 4449 45668 4505 45670
rect 4529 45668 4585 45670
rect 4250 45076 4306 45112
rect 4250 45056 4252 45076
rect 4252 45056 4304 45076
rect 4304 45056 4306 45076
rect 4289 44634 4345 44636
rect 4369 44634 4425 44636
rect 4449 44634 4505 44636
rect 4529 44634 4585 44636
rect 4289 44582 4315 44634
rect 4315 44582 4345 44634
rect 4369 44582 4379 44634
rect 4379 44582 4425 44634
rect 4449 44582 4495 44634
rect 4495 44582 4505 44634
rect 4529 44582 4559 44634
rect 4559 44582 4585 44634
rect 4289 44580 4345 44582
rect 4369 44580 4425 44582
rect 4449 44580 4505 44582
rect 4529 44580 4585 44582
rect 3974 43016 4030 43072
rect 3974 42880 4030 42936
rect 3974 35028 3976 35048
rect 3976 35028 4028 35048
rect 4028 35028 4030 35048
rect 3974 34992 4030 35028
rect 3790 32952 3846 33008
rect 3698 30640 3754 30696
rect 3422 26288 3478 26344
rect 3238 25744 3294 25800
rect 3146 25200 3202 25256
rect 3330 23432 3386 23488
rect 3146 23024 3202 23080
rect 3422 21528 3478 21584
rect 3422 20984 3478 21040
rect 3330 20440 3386 20496
rect 3514 20304 3570 20360
rect 3790 18808 3846 18864
rect 3790 17856 3846 17912
rect 3514 17720 3570 17776
rect 3146 17620 3148 17640
rect 3148 17620 3200 17640
rect 3200 17620 3202 17640
rect 3146 17584 3202 17620
rect 3146 15988 3148 16008
rect 3148 15988 3200 16008
rect 3200 15988 3202 16008
rect 3146 15952 3202 15988
rect 4289 43546 4345 43548
rect 4369 43546 4425 43548
rect 4449 43546 4505 43548
rect 4529 43546 4585 43548
rect 4289 43494 4315 43546
rect 4315 43494 4345 43546
rect 4369 43494 4379 43546
rect 4379 43494 4425 43546
rect 4449 43494 4495 43546
rect 4495 43494 4505 43546
rect 4529 43494 4559 43546
rect 4559 43494 4585 43546
rect 4289 43492 4345 43494
rect 4369 43492 4425 43494
rect 4449 43492 4505 43494
rect 4529 43492 4585 43494
rect 4289 42458 4345 42460
rect 4369 42458 4425 42460
rect 4449 42458 4505 42460
rect 4529 42458 4585 42460
rect 4289 42406 4315 42458
rect 4315 42406 4345 42458
rect 4369 42406 4379 42458
rect 4379 42406 4425 42458
rect 4449 42406 4495 42458
rect 4495 42406 4505 42458
rect 4529 42406 4559 42458
rect 4559 42406 4585 42458
rect 4289 42404 4345 42406
rect 4369 42404 4425 42406
rect 4449 42404 4505 42406
rect 4529 42404 4585 42406
rect 4289 41370 4345 41372
rect 4369 41370 4425 41372
rect 4449 41370 4505 41372
rect 4529 41370 4585 41372
rect 4289 41318 4315 41370
rect 4315 41318 4345 41370
rect 4369 41318 4379 41370
rect 4379 41318 4425 41370
rect 4449 41318 4495 41370
rect 4495 41318 4505 41370
rect 4529 41318 4559 41370
rect 4559 41318 4585 41370
rect 4289 41316 4345 41318
rect 4369 41316 4425 41318
rect 4449 41316 4505 41318
rect 4529 41316 4585 41318
rect 4250 41112 4306 41168
rect 4710 47232 4766 47288
rect 4289 40282 4345 40284
rect 4369 40282 4425 40284
rect 4449 40282 4505 40284
rect 4529 40282 4585 40284
rect 4289 40230 4315 40282
rect 4315 40230 4345 40282
rect 4369 40230 4379 40282
rect 4379 40230 4425 40282
rect 4449 40230 4495 40282
rect 4495 40230 4505 40282
rect 4529 40230 4559 40282
rect 4559 40230 4585 40282
rect 4289 40228 4345 40230
rect 4369 40228 4425 40230
rect 4449 40228 4505 40230
rect 4529 40228 4585 40230
rect 4342 39888 4398 39944
rect 4289 39194 4345 39196
rect 4369 39194 4425 39196
rect 4449 39194 4505 39196
rect 4529 39194 4585 39196
rect 4289 39142 4315 39194
rect 4315 39142 4345 39194
rect 4369 39142 4379 39194
rect 4379 39142 4425 39194
rect 4449 39142 4495 39194
rect 4495 39142 4505 39194
rect 4529 39142 4559 39194
rect 4559 39142 4585 39194
rect 4289 39140 4345 39142
rect 4369 39140 4425 39142
rect 4449 39140 4505 39142
rect 4529 39140 4585 39142
rect 4289 38106 4345 38108
rect 4369 38106 4425 38108
rect 4449 38106 4505 38108
rect 4529 38106 4585 38108
rect 4289 38054 4315 38106
rect 4315 38054 4345 38106
rect 4369 38054 4379 38106
rect 4379 38054 4425 38106
rect 4449 38054 4495 38106
rect 4495 38054 4505 38106
rect 4529 38054 4559 38106
rect 4559 38054 4585 38106
rect 4289 38052 4345 38054
rect 4369 38052 4425 38054
rect 4449 38052 4505 38054
rect 4529 38052 4585 38054
rect 4289 37018 4345 37020
rect 4369 37018 4425 37020
rect 4449 37018 4505 37020
rect 4529 37018 4585 37020
rect 4289 36966 4315 37018
rect 4315 36966 4345 37018
rect 4369 36966 4379 37018
rect 4379 36966 4425 37018
rect 4449 36966 4495 37018
rect 4495 36966 4505 37018
rect 4529 36966 4559 37018
rect 4559 36966 4585 37018
rect 4289 36964 4345 36966
rect 4369 36964 4425 36966
rect 4449 36964 4505 36966
rect 4529 36964 4585 36966
rect 4289 35930 4345 35932
rect 4369 35930 4425 35932
rect 4449 35930 4505 35932
rect 4529 35930 4585 35932
rect 4289 35878 4315 35930
rect 4315 35878 4345 35930
rect 4369 35878 4379 35930
rect 4379 35878 4425 35930
rect 4449 35878 4495 35930
rect 4495 35878 4505 35930
rect 4529 35878 4559 35930
rect 4559 35878 4585 35930
rect 4289 35876 4345 35878
rect 4369 35876 4425 35878
rect 4449 35876 4505 35878
rect 4529 35876 4585 35878
rect 4894 51040 4950 51096
rect 5354 60424 5410 60480
rect 5262 51584 5318 51640
rect 4986 47096 5042 47152
rect 5078 46824 5134 46880
rect 5814 69420 5870 69456
rect 5814 69400 5816 69420
rect 5816 69400 5868 69420
rect 5868 69400 5870 69420
rect 7010 73616 7066 73672
rect 6918 73208 6974 73264
rect 7102 72140 7158 72176
rect 7102 72120 7104 72140
rect 7104 72120 7156 72140
rect 7156 72120 7158 72140
rect 10956 75098 11012 75100
rect 11036 75098 11092 75100
rect 11116 75098 11172 75100
rect 11196 75098 11252 75100
rect 10956 75046 10982 75098
rect 10982 75046 11012 75098
rect 11036 75046 11046 75098
rect 11046 75046 11092 75098
rect 11116 75046 11162 75098
rect 11162 75046 11172 75098
rect 11196 75046 11226 75098
rect 11226 75046 11252 75098
rect 10956 75044 11012 75046
rect 11036 75044 11092 75046
rect 11116 75044 11172 75046
rect 11196 75044 11252 75046
rect 17622 75098 17678 75100
rect 17702 75098 17758 75100
rect 17782 75098 17838 75100
rect 17862 75098 17918 75100
rect 17622 75046 17648 75098
rect 17648 75046 17678 75098
rect 17702 75046 17712 75098
rect 17712 75046 17758 75098
rect 17782 75046 17828 75098
rect 17828 75046 17838 75098
rect 17862 75046 17892 75098
rect 17892 75046 17918 75098
rect 17622 75044 17678 75046
rect 17702 75044 17758 75046
rect 17782 75044 17838 75046
rect 17862 75044 17918 75046
rect 7622 74554 7678 74556
rect 7702 74554 7758 74556
rect 7782 74554 7838 74556
rect 7862 74554 7918 74556
rect 7622 74502 7648 74554
rect 7648 74502 7678 74554
rect 7702 74502 7712 74554
rect 7712 74502 7758 74554
rect 7782 74502 7828 74554
rect 7828 74502 7838 74554
rect 7862 74502 7892 74554
rect 7892 74502 7918 74554
rect 7622 74500 7678 74502
rect 7702 74500 7758 74502
rect 7782 74500 7838 74502
rect 7862 74500 7918 74502
rect 14289 74554 14345 74556
rect 14369 74554 14425 74556
rect 14449 74554 14505 74556
rect 14529 74554 14585 74556
rect 14289 74502 14315 74554
rect 14315 74502 14345 74554
rect 14369 74502 14379 74554
rect 14379 74502 14425 74554
rect 14449 74502 14495 74554
rect 14495 74502 14505 74554
rect 14529 74502 14559 74554
rect 14559 74502 14585 74554
rect 14289 74500 14345 74502
rect 14369 74500 14425 74502
rect 14449 74500 14505 74502
rect 14529 74500 14585 74502
rect 7622 73466 7678 73468
rect 7702 73466 7758 73468
rect 7782 73466 7838 73468
rect 7862 73466 7918 73468
rect 7622 73414 7648 73466
rect 7648 73414 7678 73466
rect 7702 73414 7712 73466
rect 7712 73414 7758 73466
rect 7782 73414 7828 73466
rect 7828 73414 7838 73466
rect 7862 73414 7892 73466
rect 7892 73414 7918 73466
rect 7622 73412 7678 73414
rect 7702 73412 7758 73414
rect 7782 73412 7838 73414
rect 7862 73412 7918 73414
rect 5446 59200 5502 59256
rect 5538 58112 5594 58168
rect 5630 57296 5686 57352
rect 5630 52944 5686 53000
rect 5538 51720 5594 51776
rect 5446 51176 5502 51232
rect 5354 49000 5410 49056
rect 5262 43832 5318 43888
rect 5170 42336 5226 42392
rect 5170 42200 5226 42256
rect 5078 41792 5134 41848
rect 4289 34842 4345 34844
rect 4369 34842 4425 34844
rect 4449 34842 4505 34844
rect 4529 34842 4585 34844
rect 4289 34790 4315 34842
rect 4315 34790 4345 34842
rect 4369 34790 4379 34842
rect 4379 34790 4425 34842
rect 4449 34790 4495 34842
rect 4495 34790 4505 34842
rect 4529 34790 4559 34842
rect 4559 34790 4585 34842
rect 4289 34788 4345 34790
rect 4369 34788 4425 34790
rect 4449 34788 4505 34790
rect 4529 34788 4585 34790
rect 4289 33754 4345 33756
rect 4369 33754 4425 33756
rect 4449 33754 4505 33756
rect 4529 33754 4585 33756
rect 4289 33702 4315 33754
rect 4315 33702 4345 33754
rect 4369 33702 4379 33754
rect 4379 33702 4425 33754
rect 4449 33702 4495 33754
rect 4495 33702 4505 33754
rect 4529 33702 4559 33754
rect 4559 33702 4585 33754
rect 4289 33700 4345 33702
rect 4369 33700 4425 33702
rect 4449 33700 4505 33702
rect 4529 33700 4585 33702
rect 4894 33940 4896 33960
rect 4896 33940 4948 33960
rect 4948 33940 4950 33960
rect 4894 33904 4950 33940
rect 4289 32666 4345 32668
rect 4369 32666 4425 32668
rect 4449 32666 4505 32668
rect 4529 32666 4585 32668
rect 4289 32614 4315 32666
rect 4315 32614 4345 32666
rect 4369 32614 4379 32666
rect 4379 32614 4425 32666
rect 4449 32614 4495 32666
rect 4495 32614 4505 32666
rect 4529 32614 4559 32666
rect 4559 32614 4585 32666
rect 4289 32612 4345 32614
rect 4369 32612 4425 32614
rect 4449 32612 4505 32614
rect 4529 32612 4585 32614
rect 4289 31578 4345 31580
rect 4369 31578 4425 31580
rect 4449 31578 4505 31580
rect 4529 31578 4585 31580
rect 4289 31526 4315 31578
rect 4315 31526 4345 31578
rect 4369 31526 4379 31578
rect 4379 31526 4425 31578
rect 4449 31526 4495 31578
rect 4495 31526 4505 31578
rect 4529 31526 4559 31578
rect 4559 31526 4585 31578
rect 4289 31524 4345 31526
rect 4369 31524 4425 31526
rect 4449 31524 4505 31526
rect 4529 31524 4585 31526
rect 4066 30776 4122 30832
rect 4986 30504 5042 30560
rect 4289 30490 4345 30492
rect 4369 30490 4425 30492
rect 4449 30490 4505 30492
rect 4529 30490 4585 30492
rect 4289 30438 4315 30490
rect 4315 30438 4345 30490
rect 4369 30438 4379 30490
rect 4379 30438 4425 30490
rect 4449 30438 4495 30490
rect 4495 30438 4505 30490
rect 4529 30438 4559 30490
rect 4559 30438 4585 30490
rect 4289 30436 4345 30438
rect 4369 30436 4425 30438
rect 4449 30436 4505 30438
rect 4529 30436 4585 30438
rect 4526 29960 4582 30016
rect 4289 29402 4345 29404
rect 4369 29402 4425 29404
rect 4449 29402 4505 29404
rect 4529 29402 4585 29404
rect 4289 29350 4315 29402
rect 4315 29350 4345 29402
rect 4369 29350 4379 29402
rect 4379 29350 4425 29402
rect 4449 29350 4495 29402
rect 4495 29350 4505 29402
rect 4529 29350 4559 29402
rect 4559 29350 4585 29402
rect 4289 29348 4345 29350
rect 4369 29348 4425 29350
rect 4449 29348 4505 29350
rect 4529 29348 4585 29350
rect 4289 28314 4345 28316
rect 4369 28314 4425 28316
rect 4449 28314 4505 28316
rect 4529 28314 4585 28316
rect 4289 28262 4315 28314
rect 4315 28262 4345 28314
rect 4369 28262 4379 28314
rect 4379 28262 4425 28314
rect 4449 28262 4495 28314
rect 4495 28262 4505 28314
rect 4529 28262 4559 28314
rect 4559 28262 4585 28314
rect 4289 28260 4345 28262
rect 4369 28260 4425 28262
rect 4449 28260 4505 28262
rect 4529 28260 4585 28262
rect 4066 27376 4122 27432
rect 5262 37304 5318 37360
rect 5722 50904 5778 50960
rect 5538 49156 5594 49192
rect 5538 49136 5540 49156
rect 5540 49136 5592 49156
rect 5592 49136 5594 49156
rect 5538 49000 5594 49056
rect 5630 48864 5686 48920
rect 5630 46452 5632 46472
rect 5632 46452 5684 46472
rect 5684 46452 5686 46472
rect 5630 46416 5686 46452
rect 5630 44376 5686 44432
rect 5814 50768 5870 50824
rect 5814 48204 5870 48240
rect 5814 48184 5816 48204
rect 5816 48184 5868 48204
rect 5868 48184 5870 48204
rect 5814 47676 5816 47696
rect 5816 47676 5868 47696
rect 5868 47676 5870 47696
rect 5814 47640 5870 47676
rect 5722 41928 5778 41984
rect 5630 41384 5686 41440
rect 5630 41112 5686 41168
rect 5630 41012 5632 41032
rect 5632 41012 5684 41032
rect 5684 41012 5686 41032
rect 5630 40976 5686 41012
rect 5538 40840 5594 40896
rect 5446 29144 5502 29200
rect 4289 27226 4345 27228
rect 4369 27226 4425 27228
rect 4449 27226 4505 27228
rect 4529 27226 4585 27228
rect 4289 27174 4315 27226
rect 4315 27174 4345 27226
rect 4369 27174 4379 27226
rect 4379 27174 4425 27226
rect 4449 27174 4495 27226
rect 4495 27174 4505 27226
rect 4529 27174 4559 27226
rect 4559 27174 4585 27226
rect 4289 27172 4345 27174
rect 4369 27172 4425 27174
rect 4449 27172 4505 27174
rect 4529 27172 4585 27174
rect 4289 26138 4345 26140
rect 4369 26138 4425 26140
rect 4449 26138 4505 26140
rect 4529 26138 4585 26140
rect 4289 26086 4315 26138
rect 4315 26086 4345 26138
rect 4369 26086 4379 26138
rect 4379 26086 4425 26138
rect 4449 26086 4495 26138
rect 4495 26086 4505 26138
rect 4529 26086 4559 26138
rect 4559 26086 4585 26138
rect 4289 26084 4345 26086
rect 4369 26084 4425 26086
rect 4449 26084 4505 26086
rect 4529 26084 4585 26086
rect 4158 25200 4214 25256
rect 4066 23160 4122 23216
rect 4289 25050 4345 25052
rect 4369 25050 4425 25052
rect 4449 25050 4505 25052
rect 4529 25050 4585 25052
rect 4289 24998 4315 25050
rect 4315 24998 4345 25050
rect 4369 24998 4379 25050
rect 4379 24998 4425 25050
rect 4449 24998 4495 25050
rect 4495 24998 4505 25050
rect 4529 24998 4559 25050
rect 4559 24998 4585 25050
rect 4289 24996 4345 24998
rect 4369 24996 4425 24998
rect 4449 24996 4505 24998
rect 4529 24996 4585 24998
rect 5170 26560 5226 26616
rect 5170 24384 5226 24440
rect 4289 23962 4345 23964
rect 4369 23962 4425 23964
rect 4449 23962 4505 23964
rect 4529 23962 4585 23964
rect 4289 23910 4315 23962
rect 4315 23910 4345 23962
rect 4369 23910 4379 23962
rect 4379 23910 4425 23962
rect 4449 23910 4495 23962
rect 4495 23910 4505 23962
rect 4529 23910 4559 23962
rect 4559 23910 4585 23962
rect 4289 23908 4345 23910
rect 4369 23908 4425 23910
rect 4449 23908 4505 23910
rect 4529 23908 4585 23910
rect 4710 22888 4766 22944
rect 4289 22874 4345 22876
rect 4369 22874 4425 22876
rect 4449 22874 4505 22876
rect 4529 22874 4585 22876
rect 4289 22822 4315 22874
rect 4315 22822 4345 22874
rect 4369 22822 4379 22874
rect 4379 22822 4425 22874
rect 4449 22822 4495 22874
rect 4495 22822 4505 22874
rect 4529 22822 4559 22874
rect 4559 22822 4585 22874
rect 4289 22820 4345 22822
rect 4369 22820 4425 22822
rect 4449 22820 4505 22822
rect 4529 22820 4585 22822
rect 5078 23468 5080 23488
rect 5080 23468 5132 23488
rect 5132 23468 5134 23488
rect 5078 23432 5134 23468
rect 7194 71304 7250 71360
rect 6642 69400 6698 69456
rect 7102 68992 7158 69048
rect 6090 63280 6146 63336
rect 6274 60560 6330 60616
rect 6182 60036 6238 60072
rect 6182 60016 6184 60036
rect 6184 60016 6236 60036
rect 6236 60016 6238 60036
rect 6274 59336 6330 59392
rect 6274 55664 6330 55720
rect 6182 54068 6184 54088
rect 6184 54068 6236 54088
rect 6236 54068 6238 54088
rect 6182 54032 6238 54068
rect 6090 52672 6146 52728
rect 6182 52128 6238 52184
rect 6366 53896 6422 53952
rect 6642 59744 6698 59800
rect 7194 67124 7196 67144
rect 7196 67124 7248 67144
rect 7248 67124 7250 67144
rect 7194 67088 7250 67124
rect 10956 74010 11012 74012
rect 11036 74010 11092 74012
rect 11116 74010 11172 74012
rect 11196 74010 11252 74012
rect 10956 73958 10982 74010
rect 10982 73958 11012 74010
rect 11036 73958 11046 74010
rect 11046 73958 11092 74010
rect 11116 73958 11162 74010
rect 11162 73958 11172 74010
rect 11196 73958 11226 74010
rect 11226 73958 11252 74010
rect 10956 73956 11012 73958
rect 11036 73956 11092 73958
rect 11116 73956 11172 73958
rect 11196 73956 11252 73958
rect 17622 74010 17678 74012
rect 17702 74010 17758 74012
rect 17782 74010 17838 74012
rect 17862 74010 17918 74012
rect 17622 73958 17648 74010
rect 17648 73958 17678 74010
rect 17702 73958 17712 74010
rect 17712 73958 17758 74010
rect 17782 73958 17828 74010
rect 17828 73958 17838 74010
rect 17862 73958 17892 74010
rect 17892 73958 17918 74010
rect 17622 73956 17678 73958
rect 17702 73956 17758 73958
rect 17782 73956 17838 73958
rect 17862 73956 17918 73958
rect 8482 73344 8538 73400
rect 7622 72378 7678 72380
rect 7702 72378 7758 72380
rect 7782 72378 7838 72380
rect 7862 72378 7918 72380
rect 7622 72326 7648 72378
rect 7648 72326 7678 72378
rect 7702 72326 7712 72378
rect 7712 72326 7758 72378
rect 7782 72326 7828 72378
rect 7828 72326 7838 72378
rect 7862 72326 7892 72378
rect 7892 72326 7918 72378
rect 7622 72324 7678 72326
rect 7702 72324 7758 72326
rect 7782 72324 7838 72326
rect 7862 72324 7918 72326
rect 7622 71290 7678 71292
rect 7702 71290 7758 71292
rect 7782 71290 7838 71292
rect 7862 71290 7918 71292
rect 7622 71238 7648 71290
rect 7648 71238 7678 71290
rect 7702 71238 7712 71290
rect 7712 71238 7758 71290
rect 7782 71238 7828 71290
rect 7828 71238 7838 71290
rect 7862 71238 7892 71290
rect 7892 71238 7918 71290
rect 7622 71236 7678 71238
rect 7702 71236 7758 71238
rect 7782 71236 7838 71238
rect 7862 71236 7918 71238
rect 7470 70352 7526 70408
rect 7838 70352 7894 70408
rect 7622 70202 7678 70204
rect 7702 70202 7758 70204
rect 7782 70202 7838 70204
rect 7862 70202 7918 70204
rect 7622 70150 7648 70202
rect 7648 70150 7678 70202
rect 7702 70150 7712 70202
rect 7712 70150 7758 70202
rect 7782 70150 7828 70202
rect 7828 70150 7838 70202
rect 7862 70150 7892 70202
rect 7892 70150 7918 70202
rect 7622 70148 7678 70150
rect 7702 70148 7758 70150
rect 7782 70148 7838 70150
rect 7862 70148 7918 70150
rect 7622 69114 7678 69116
rect 7702 69114 7758 69116
rect 7782 69114 7838 69116
rect 7862 69114 7918 69116
rect 7622 69062 7648 69114
rect 7648 69062 7678 69114
rect 7702 69062 7712 69114
rect 7712 69062 7758 69114
rect 7782 69062 7828 69114
rect 7828 69062 7838 69114
rect 7862 69062 7892 69114
rect 7892 69062 7918 69114
rect 7622 69060 7678 69062
rect 7702 69060 7758 69062
rect 7782 69060 7838 69062
rect 7862 69060 7918 69062
rect 8022 68876 8078 68912
rect 8022 68856 8024 68876
rect 8024 68856 8076 68876
rect 8076 68856 8078 68876
rect 7194 64504 7250 64560
rect 7194 63552 7250 63608
rect 7194 62328 7250 62384
rect 7102 62056 7158 62112
rect 6642 58520 6698 58576
rect 6734 54304 6790 54360
rect 6734 54204 6736 54224
rect 6736 54204 6788 54224
rect 6788 54204 6790 54224
rect 6734 54168 6790 54204
rect 6734 54032 6790 54088
rect 6090 50224 6146 50280
rect 6090 49272 6146 49328
rect 5998 48592 6054 48648
rect 6090 48320 6146 48376
rect 6090 47912 6146 47968
rect 6550 51720 6606 51776
rect 6458 51176 6514 51232
rect 6458 50088 6514 50144
rect 6274 49544 6330 49600
rect 6182 45464 6238 45520
rect 6182 43016 6238 43072
rect 6182 42744 6238 42800
rect 5998 41676 6054 41712
rect 5998 41656 6000 41676
rect 6000 41656 6052 41676
rect 6052 41656 6054 41676
rect 5998 39480 6054 39536
rect 5814 36352 5870 36408
rect 5998 36216 6054 36272
rect 5722 33380 5778 33416
rect 5722 33360 5724 33380
rect 5724 33360 5776 33380
rect 5776 33360 5778 33380
rect 5814 31884 5870 31920
rect 5814 31864 5816 31884
rect 5816 31864 5868 31884
rect 5868 31864 5870 31884
rect 6274 41384 6330 41440
rect 6274 41248 6330 41304
rect 6182 40432 6238 40488
rect 6182 39908 6238 39944
rect 6182 39888 6184 39908
rect 6184 39888 6236 39908
rect 6236 39888 6238 39908
rect 6182 39752 6238 39808
rect 6274 36660 6276 36680
rect 6276 36660 6328 36680
rect 6328 36660 6330 36680
rect 6274 36624 6330 36660
rect 6182 33496 6238 33552
rect 7622 68026 7678 68028
rect 7702 68026 7758 68028
rect 7782 68026 7838 68028
rect 7862 68026 7918 68028
rect 7622 67974 7648 68026
rect 7648 67974 7678 68026
rect 7702 67974 7712 68026
rect 7712 67974 7758 68026
rect 7782 67974 7828 68026
rect 7828 67974 7838 68026
rect 7862 67974 7892 68026
rect 7892 67974 7918 68026
rect 7622 67972 7678 67974
rect 7702 67972 7758 67974
rect 7782 67972 7838 67974
rect 7862 67972 7918 67974
rect 8390 70388 8392 70408
rect 8392 70388 8444 70408
rect 8444 70388 8446 70408
rect 8390 70352 8446 70388
rect 8206 70216 8262 70272
rect 8482 69672 8538 69728
rect 8390 69400 8446 69456
rect 8206 69128 8262 69184
rect 7622 66938 7678 66940
rect 7702 66938 7758 66940
rect 7782 66938 7838 66940
rect 7862 66938 7918 66940
rect 7622 66886 7648 66938
rect 7648 66886 7678 66938
rect 7702 66886 7712 66938
rect 7712 66886 7758 66938
rect 7782 66886 7828 66938
rect 7828 66886 7838 66938
rect 7862 66886 7892 66938
rect 7892 66886 7918 66938
rect 7622 66884 7678 66886
rect 7702 66884 7758 66886
rect 7782 66884 7838 66886
rect 7862 66884 7918 66886
rect 7562 66136 7618 66192
rect 7622 65850 7678 65852
rect 7702 65850 7758 65852
rect 7782 65850 7838 65852
rect 7862 65850 7918 65852
rect 7622 65798 7648 65850
rect 7648 65798 7678 65850
rect 7702 65798 7712 65850
rect 7712 65798 7758 65850
rect 7782 65798 7828 65850
rect 7828 65798 7838 65850
rect 7862 65798 7892 65850
rect 7892 65798 7918 65850
rect 7622 65796 7678 65798
rect 7702 65796 7758 65798
rect 7782 65796 7838 65798
rect 7862 65796 7918 65798
rect 7622 64762 7678 64764
rect 7702 64762 7758 64764
rect 7782 64762 7838 64764
rect 7862 64762 7918 64764
rect 7622 64710 7648 64762
rect 7648 64710 7678 64762
rect 7702 64710 7712 64762
rect 7712 64710 7758 64762
rect 7782 64710 7828 64762
rect 7828 64710 7838 64762
rect 7862 64710 7892 64762
rect 7892 64710 7918 64762
rect 7622 64708 7678 64710
rect 7702 64708 7758 64710
rect 7782 64708 7838 64710
rect 7862 64708 7918 64710
rect 7930 63860 7932 63880
rect 7932 63860 7984 63880
rect 7984 63860 7986 63880
rect 7930 63824 7986 63860
rect 7622 63674 7678 63676
rect 7702 63674 7758 63676
rect 7782 63674 7838 63676
rect 7862 63674 7918 63676
rect 7622 63622 7648 63674
rect 7648 63622 7678 63674
rect 7702 63622 7712 63674
rect 7712 63622 7758 63674
rect 7782 63622 7828 63674
rect 7828 63622 7838 63674
rect 7862 63622 7892 63674
rect 7892 63622 7918 63674
rect 7622 63620 7678 63622
rect 7702 63620 7758 63622
rect 7782 63620 7838 63622
rect 7862 63620 7918 63622
rect 7746 63316 7748 63336
rect 7748 63316 7800 63336
rect 7800 63316 7802 63336
rect 7746 63280 7802 63316
rect 7286 59608 7342 59664
rect 7286 59336 7342 59392
rect 7010 55936 7066 55992
rect 7010 52536 7066 52592
rect 6826 51584 6882 51640
rect 6734 51040 6790 51096
rect 6826 50904 6882 50960
rect 6642 47640 6698 47696
rect 7010 51484 7012 51504
rect 7012 51484 7064 51504
rect 7064 51484 7066 51504
rect 7010 51448 7066 51484
rect 7010 50804 7012 50824
rect 7012 50804 7064 50824
rect 7064 50804 7066 50824
rect 7010 50768 7066 50804
rect 6366 33088 6422 33144
rect 6366 31728 6422 31784
rect 5170 22888 5226 22944
rect 4289 21786 4345 21788
rect 4369 21786 4425 21788
rect 4449 21786 4505 21788
rect 4529 21786 4585 21788
rect 4289 21734 4315 21786
rect 4315 21734 4345 21786
rect 4369 21734 4379 21786
rect 4379 21734 4425 21786
rect 4449 21734 4495 21786
rect 4495 21734 4505 21786
rect 4529 21734 4559 21786
rect 4559 21734 4585 21786
rect 4289 21732 4345 21734
rect 4369 21732 4425 21734
rect 4449 21732 4505 21734
rect 4529 21732 4585 21734
rect 4289 20698 4345 20700
rect 4369 20698 4425 20700
rect 4449 20698 4505 20700
rect 4529 20698 4585 20700
rect 4289 20646 4315 20698
rect 4315 20646 4345 20698
rect 4369 20646 4379 20698
rect 4379 20646 4425 20698
rect 4449 20646 4495 20698
rect 4495 20646 4505 20698
rect 4529 20646 4559 20698
rect 4559 20646 4585 20698
rect 4289 20644 4345 20646
rect 4369 20644 4425 20646
rect 4449 20644 4505 20646
rect 4529 20644 4585 20646
rect 4066 19236 4122 19272
rect 4066 19216 4068 19236
rect 4068 19216 4120 19236
rect 4120 19216 4122 19236
rect 4289 19610 4345 19612
rect 4369 19610 4425 19612
rect 4449 19610 4505 19612
rect 4529 19610 4585 19612
rect 4289 19558 4315 19610
rect 4315 19558 4345 19610
rect 4369 19558 4379 19610
rect 4379 19558 4425 19610
rect 4449 19558 4495 19610
rect 4495 19558 4505 19610
rect 4529 19558 4559 19610
rect 4559 19558 4585 19610
rect 4289 19556 4345 19558
rect 4369 19556 4425 19558
rect 4449 19556 4505 19558
rect 4529 19556 4585 19558
rect 4710 19352 4766 19408
rect 5906 23432 5962 23488
rect 6918 47776 6974 47832
rect 7010 45056 7066 45112
rect 7378 58928 7434 58984
rect 7746 62756 7802 62792
rect 7746 62736 7748 62756
rect 7748 62736 7800 62756
rect 7800 62736 7802 62756
rect 7622 62586 7678 62588
rect 7702 62586 7758 62588
rect 7782 62586 7838 62588
rect 7862 62586 7918 62588
rect 7622 62534 7648 62586
rect 7648 62534 7678 62586
rect 7702 62534 7712 62586
rect 7712 62534 7758 62586
rect 7782 62534 7828 62586
rect 7828 62534 7838 62586
rect 7862 62534 7892 62586
rect 7892 62534 7918 62586
rect 7622 62532 7678 62534
rect 7702 62532 7758 62534
rect 7782 62532 7838 62534
rect 7862 62532 7918 62534
rect 7622 61498 7678 61500
rect 7702 61498 7758 61500
rect 7782 61498 7838 61500
rect 7862 61498 7918 61500
rect 7622 61446 7648 61498
rect 7648 61446 7678 61498
rect 7702 61446 7712 61498
rect 7712 61446 7758 61498
rect 7782 61446 7828 61498
rect 7828 61446 7838 61498
rect 7862 61446 7892 61498
rect 7892 61446 7918 61498
rect 7622 61444 7678 61446
rect 7702 61444 7758 61446
rect 7782 61444 7838 61446
rect 7862 61444 7918 61446
rect 7562 60560 7618 60616
rect 7622 60410 7678 60412
rect 7702 60410 7758 60412
rect 7782 60410 7838 60412
rect 7862 60410 7918 60412
rect 7622 60358 7648 60410
rect 7648 60358 7678 60410
rect 7702 60358 7712 60410
rect 7712 60358 7758 60410
rect 7782 60358 7828 60410
rect 7828 60358 7838 60410
rect 7862 60358 7892 60410
rect 7892 60358 7918 60410
rect 7622 60356 7678 60358
rect 7702 60356 7758 60358
rect 7782 60356 7838 60358
rect 7862 60356 7918 60358
rect 7622 59322 7678 59324
rect 7702 59322 7758 59324
rect 7782 59322 7838 59324
rect 7862 59322 7918 59324
rect 7622 59270 7648 59322
rect 7648 59270 7678 59322
rect 7702 59270 7712 59322
rect 7712 59270 7758 59322
rect 7782 59270 7828 59322
rect 7828 59270 7838 59322
rect 7862 59270 7892 59322
rect 7892 59270 7918 59322
rect 7622 59268 7678 59270
rect 7702 59268 7758 59270
rect 7782 59268 7838 59270
rect 7862 59268 7918 59270
rect 7622 58234 7678 58236
rect 7702 58234 7758 58236
rect 7782 58234 7838 58236
rect 7862 58234 7918 58236
rect 7622 58182 7648 58234
rect 7648 58182 7678 58234
rect 7702 58182 7712 58234
rect 7712 58182 7758 58234
rect 7782 58182 7828 58234
rect 7828 58182 7838 58234
rect 7862 58182 7892 58234
rect 7892 58182 7918 58234
rect 7622 58180 7678 58182
rect 7702 58180 7758 58182
rect 7782 58180 7838 58182
rect 7862 58180 7918 58182
rect 7562 57976 7618 58032
rect 7838 57840 7894 57896
rect 7930 57296 7986 57352
rect 7622 57146 7678 57148
rect 7702 57146 7758 57148
rect 7782 57146 7838 57148
rect 7862 57146 7918 57148
rect 7622 57094 7648 57146
rect 7648 57094 7678 57146
rect 7702 57094 7712 57146
rect 7712 57094 7758 57146
rect 7782 57094 7828 57146
rect 7828 57094 7838 57146
rect 7862 57094 7892 57146
rect 7892 57094 7918 57146
rect 7622 57092 7678 57094
rect 7702 57092 7758 57094
rect 7782 57092 7838 57094
rect 7862 57092 7918 57094
rect 7622 56058 7678 56060
rect 7702 56058 7758 56060
rect 7782 56058 7838 56060
rect 7862 56058 7918 56060
rect 7622 56006 7648 56058
rect 7648 56006 7678 56058
rect 7702 56006 7712 56058
rect 7712 56006 7758 56058
rect 7782 56006 7828 56058
rect 7828 56006 7838 56058
rect 7862 56006 7892 56058
rect 7892 56006 7918 56058
rect 7622 56004 7678 56006
rect 7702 56004 7758 56006
rect 7782 56004 7838 56006
rect 7862 56004 7918 56006
rect 7286 55020 7288 55040
rect 7288 55020 7340 55040
rect 7340 55020 7342 55040
rect 7286 54984 7342 55020
rect 7378 53896 7434 53952
rect 7622 54970 7678 54972
rect 7702 54970 7758 54972
rect 7782 54970 7838 54972
rect 7862 54970 7918 54972
rect 7622 54918 7648 54970
rect 7648 54918 7678 54970
rect 7702 54918 7712 54970
rect 7712 54918 7758 54970
rect 7782 54918 7828 54970
rect 7828 54918 7838 54970
rect 7862 54918 7892 54970
rect 7892 54918 7918 54970
rect 7622 54916 7678 54918
rect 7702 54916 7758 54918
rect 7782 54916 7838 54918
rect 7862 54916 7918 54918
rect 7838 54712 7894 54768
rect 7622 53882 7678 53884
rect 7702 53882 7758 53884
rect 7782 53882 7838 53884
rect 7862 53882 7918 53884
rect 7622 53830 7648 53882
rect 7648 53830 7678 53882
rect 7702 53830 7712 53882
rect 7712 53830 7758 53882
rect 7782 53830 7828 53882
rect 7828 53830 7838 53882
rect 7862 53830 7892 53882
rect 7892 53830 7918 53882
rect 7622 53828 7678 53830
rect 7702 53828 7758 53830
rect 7782 53828 7838 53830
rect 7862 53828 7918 53830
rect 7622 52794 7678 52796
rect 7702 52794 7758 52796
rect 7782 52794 7838 52796
rect 7862 52794 7918 52796
rect 7622 52742 7648 52794
rect 7648 52742 7678 52794
rect 7702 52742 7712 52794
rect 7712 52742 7758 52794
rect 7782 52742 7828 52794
rect 7828 52742 7838 52794
rect 7862 52742 7892 52794
rect 7892 52742 7918 52794
rect 7622 52740 7678 52742
rect 7702 52740 7758 52742
rect 7782 52740 7838 52742
rect 7862 52740 7918 52742
rect 7622 51706 7678 51708
rect 7702 51706 7758 51708
rect 7782 51706 7838 51708
rect 7862 51706 7918 51708
rect 7622 51654 7648 51706
rect 7648 51654 7678 51706
rect 7702 51654 7712 51706
rect 7712 51654 7758 51706
rect 7782 51654 7828 51706
rect 7828 51654 7838 51706
rect 7862 51654 7892 51706
rect 7892 51654 7918 51706
rect 7622 51652 7678 51654
rect 7702 51652 7758 51654
rect 7782 51652 7838 51654
rect 7862 51652 7918 51654
rect 7930 51468 7986 51504
rect 7930 51448 7932 51468
rect 7932 51448 7984 51468
rect 7984 51448 7986 51468
rect 7746 51312 7802 51368
rect 7622 50618 7678 50620
rect 7702 50618 7758 50620
rect 7782 50618 7838 50620
rect 7862 50618 7918 50620
rect 7622 50566 7648 50618
rect 7648 50566 7678 50618
rect 7702 50566 7712 50618
rect 7712 50566 7758 50618
rect 7782 50566 7828 50618
rect 7828 50566 7838 50618
rect 7862 50566 7892 50618
rect 7892 50566 7918 50618
rect 7622 50564 7678 50566
rect 7702 50564 7758 50566
rect 7782 50564 7838 50566
rect 7862 50564 7918 50566
rect 8206 65456 8262 65512
rect 8298 64776 8354 64832
rect 8850 71032 8906 71088
rect 9402 71984 9458 72040
rect 9586 70624 9642 70680
rect 9678 70352 9734 70408
rect 9770 70216 9826 70272
rect 9586 69944 9642 70000
rect 9402 69264 9458 69320
rect 9770 69264 9826 69320
rect 9402 69128 9458 69184
rect 8666 64776 8722 64832
rect 8390 63416 8446 63472
rect 8574 63416 8630 63472
rect 8298 61260 8354 61296
rect 8298 61240 8300 61260
rect 8300 61240 8352 61260
rect 8352 61240 8354 61260
rect 8758 62872 8814 62928
rect 8390 60152 8446 60208
rect 8298 58828 8300 58848
rect 8300 58828 8352 58848
rect 8352 58828 8354 58848
rect 8298 58792 8354 58828
rect 8298 55956 8354 55992
rect 8298 55936 8300 55956
rect 8300 55936 8352 55956
rect 8352 55936 8354 55956
rect 8390 54440 8446 54496
rect 8114 52808 8170 52864
rect 8206 52672 8262 52728
rect 8114 52400 8170 52456
rect 7470 50088 7526 50144
rect 8022 50360 8078 50416
rect 7838 49816 7894 49872
rect 6918 43968 6974 44024
rect 7378 48340 7434 48376
rect 7378 48320 7380 48340
rect 7380 48320 7432 48340
rect 7432 48320 7434 48340
rect 7622 49530 7678 49532
rect 7702 49530 7758 49532
rect 7782 49530 7838 49532
rect 7862 49530 7918 49532
rect 7622 49478 7648 49530
rect 7648 49478 7678 49530
rect 7702 49478 7712 49530
rect 7712 49478 7758 49530
rect 7782 49478 7828 49530
rect 7828 49478 7838 49530
rect 7862 49478 7892 49530
rect 7892 49478 7918 49530
rect 7622 49476 7678 49478
rect 7702 49476 7758 49478
rect 7782 49476 7838 49478
rect 7862 49476 7918 49478
rect 7746 48628 7748 48648
rect 7748 48628 7800 48648
rect 7800 48628 7802 48648
rect 7746 48592 7802 48628
rect 7622 48442 7678 48444
rect 7702 48442 7758 48444
rect 7782 48442 7838 48444
rect 7862 48442 7918 48444
rect 7622 48390 7648 48442
rect 7648 48390 7678 48442
rect 7702 48390 7712 48442
rect 7712 48390 7758 48442
rect 7782 48390 7828 48442
rect 7828 48390 7838 48442
rect 7862 48390 7892 48442
rect 7892 48390 7918 48442
rect 7622 48388 7678 48390
rect 7702 48388 7758 48390
rect 7782 48388 7838 48390
rect 7862 48388 7918 48390
rect 7930 48184 7986 48240
rect 8298 51176 8354 51232
rect 8298 49136 8354 49192
rect 8114 48456 8170 48512
rect 8574 58520 8630 58576
rect 9126 65728 9182 65784
rect 9126 63960 9182 64016
rect 9126 63824 9182 63880
rect 10322 72120 10378 72176
rect 10690 73208 10746 73264
rect 10956 72922 11012 72924
rect 11036 72922 11092 72924
rect 11116 72922 11172 72924
rect 11196 72922 11252 72924
rect 10956 72870 10982 72922
rect 10982 72870 11012 72922
rect 11036 72870 11046 72922
rect 11046 72870 11092 72922
rect 11116 72870 11162 72922
rect 11162 72870 11172 72922
rect 11196 72870 11226 72922
rect 11226 72870 11252 72922
rect 10956 72868 11012 72870
rect 11036 72868 11092 72870
rect 11116 72868 11172 72870
rect 11196 72868 11252 72870
rect 14289 73466 14345 73468
rect 14369 73466 14425 73468
rect 14449 73466 14505 73468
rect 14529 73466 14585 73468
rect 14289 73414 14315 73466
rect 14315 73414 14345 73466
rect 14369 73414 14379 73466
rect 14379 73414 14425 73466
rect 14449 73414 14495 73466
rect 14495 73414 14505 73466
rect 14529 73414 14559 73466
rect 14559 73414 14585 73466
rect 14289 73412 14345 73414
rect 14369 73412 14425 73414
rect 14449 73412 14505 73414
rect 14529 73412 14585 73414
rect 17622 72922 17678 72924
rect 17702 72922 17758 72924
rect 17782 72922 17838 72924
rect 17862 72922 17918 72924
rect 17622 72870 17648 72922
rect 17648 72870 17678 72922
rect 17702 72870 17712 72922
rect 17712 72870 17758 72922
rect 17782 72870 17828 72922
rect 17828 72870 17838 72922
rect 17862 72870 17892 72922
rect 17892 72870 17918 72922
rect 17622 72868 17678 72870
rect 17702 72868 17758 72870
rect 17782 72868 17838 72870
rect 17862 72868 17918 72870
rect 16302 72664 16358 72720
rect 11794 72564 11796 72584
rect 11796 72564 11848 72584
rect 11848 72564 11850 72584
rect 10046 68856 10102 68912
rect 9678 67124 9680 67144
rect 9680 67124 9732 67144
rect 9732 67124 9734 67144
rect 9678 67088 9734 67124
rect 9402 65592 9458 65648
rect 9218 63416 9274 63472
rect 9218 62192 9274 62248
rect 9034 59764 9090 59800
rect 9034 59744 9036 59764
rect 9036 59744 9088 59764
rect 9088 59744 9090 59764
rect 8850 55800 8906 55856
rect 8850 54984 8906 55040
rect 8850 53644 8906 53680
rect 8850 53624 8852 53644
rect 8852 53624 8904 53644
rect 8904 53624 8906 53644
rect 8574 49952 8630 50008
rect 8114 48048 8170 48104
rect 8114 47912 8170 47968
rect 7622 47354 7678 47356
rect 7702 47354 7758 47356
rect 7782 47354 7838 47356
rect 7862 47354 7918 47356
rect 7622 47302 7648 47354
rect 7648 47302 7678 47354
rect 7702 47302 7712 47354
rect 7712 47302 7758 47354
rect 7782 47302 7828 47354
rect 7828 47302 7838 47354
rect 7862 47302 7892 47354
rect 7892 47302 7918 47354
rect 7622 47300 7678 47302
rect 7702 47300 7758 47302
rect 7782 47300 7838 47302
rect 7862 47300 7918 47302
rect 7622 46266 7678 46268
rect 7702 46266 7758 46268
rect 7782 46266 7838 46268
rect 7862 46266 7918 46268
rect 7622 46214 7648 46266
rect 7648 46214 7678 46266
rect 7702 46214 7712 46266
rect 7712 46214 7758 46266
rect 7782 46214 7828 46266
rect 7828 46214 7838 46266
rect 7862 46214 7892 46266
rect 7892 46214 7918 46266
rect 7622 46212 7678 46214
rect 7702 46212 7758 46214
rect 7782 46212 7838 46214
rect 7862 46212 7918 46214
rect 7930 45600 7986 45656
rect 7622 45178 7678 45180
rect 7702 45178 7758 45180
rect 7782 45178 7838 45180
rect 7862 45178 7918 45180
rect 7622 45126 7648 45178
rect 7648 45126 7678 45178
rect 7702 45126 7712 45178
rect 7712 45126 7758 45178
rect 7782 45126 7828 45178
rect 7828 45126 7838 45178
rect 7862 45126 7892 45178
rect 7892 45126 7918 45178
rect 7622 45124 7678 45126
rect 7702 45124 7758 45126
rect 7782 45124 7838 45126
rect 7862 45124 7918 45126
rect 7562 44920 7618 44976
rect 7010 43696 7066 43752
rect 6918 42200 6974 42256
rect 6918 42064 6974 42120
rect 7102 41520 7158 41576
rect 7010 41268 7066 41304
rect 7010 41248 7012 41268
rect 7012 41248 7064 41268
rect 7064 41248 7066 41268
rect 6734 37748 6736 37768
rect 6736 37748 6788 37768
rect 6788 37748 6790 37768
rect 6734 37712 6790 37748
rect 7286 40976 7342 41032
rect 7286 38120 7342 38176
rect 7622 44090 7678 44092
rect 7702 44090 7758 44092
rect 7782 44090 7838 44092
rect 7862 44090 7918 44092
rect 7622 44038 7648 44090
rect 7648 44038 7678 44090
rect 7702 44038 7712 44090
rect 7712 44038 7758 44090
rect 7782 44038 7828 44090
rect 7828 44038 7838 44090
rect 7862 44038 7892 44090
rect 7892 44038 7918 44090
rect 7622 44036 7678 44038
rect 7702 44036 7758 44038
rect 7782 44036 7838 44038
rect 7862 44036 7918 44038
rect 7622 43002 7678 43004
rect 7702 43002 7758 43004
rect 7782 43002 7838 43004
rect 7862 43002 7918 43004
rect 7622 42950 7648 43002
rect 7648 42950 7678 43002
rect 7702 42950 7712 43002
rect 7712 42950 7758 43002
rect 7782 42950 7828 43002
rect 7828 42950 7838 43002
rect 7862 42950 7892 43002
rect 7892 42950 7918 43002
rect 7622 42948 7678 42950
rect 7702 42948 7758 42950
rect 7782 42948 7838 42950
rect 7862 42948 7918 42950
rect 7562 42608 7618 42664
rect 7746 42220 7802 42256
rect 7746 42200 7748 42220
rect 7748 42200 7800 42220
rect 7800 42200 7802 42220
rect 7622 41914 7678 41916
rect 7702 41914 7758 41916
rect 7782 41914 7838 41916
rect 7862 41914 7918 41916
rect 7622 41862 7648 41914
rect 7648 41862 7678 41914
rect 7702 41862 7712 41914
rect 7712 41862 7758 41914
rect 7782 41862 7828 41914
rect 7828 41862 7838 41914
rect 7862 41862 7892 41914
rect 7892 41862 7918 41914
rect 7622 41860 7678 41862
rect 7702 41860 7758 41862
rect 7782 41860 7838 41862
rect 7862 41860 7918 41862
rect 7470 40976 7526 41032
rect 7622 40826 7678 40828
rect 7702 40826 7758 40828
rect 7782 40826 7838 40828
rect 7862 40826 7918 40828
rect 7622 40774 7648 40826
rect 7648 40774 7678 40826
rect 7702 40774 7712 40826
rect 7712 40774 7758 40826
rect 7782 40774 7828 40826
rect 7828 40774 7838 40826
rect 7862 40774 7892 40826
rect 7892 40774 7918 40826
rect 7622 40772 7678 40774
rect 7702 40772 7758 40774
rect 7782 40772 7838 40774
rect 7862 40772 7918 40774
rect 7622 39738 7678 39740
rect 7702 39738 7758 39740
rect 7782 39738 7838 39740
rect 7862 39738 7918 39740
rect 7622 39686 7648 39738
rect 7648 39686 7678 39738
rect 7702 39686 7712 39738
rect 7712 39686 7758 39738
rect 7782 39686 7828 39738
rect 7828 39686 7838 39738
rect 7862 39686 7892 39738
rect 7892 39686 7918 39738
rect 7622 39684 7678 39686
rect 7702 39684 7758 39686
rect 7782 39684 7838 39686
rect 7862 39684 7918 39686
rect 7562 39380 7564 39400
rect 7564 39380 7616 39400
rect 7616 39380 7618 39400
rect 7562 39344 7618 39380
rect 7654 38936 7710 38992
rect 6734 37032 6790 37088
rect 6826 36352 6882 36408
rect 6734 34040 6790 34096
rect 6826 33768 6882 33824
rect 6826 33652 6882 33688
rect 6826 33632 6828 33652
rect 6828 33632 6880 33652
rect 6880 33632 6882 33652
rect 6826 32952 6882 33008
rect 6826 32272 6882 32328
rect 6826 31728 6882 31784
rect 7622 38650 7678 38652
rect 7702 38650 7758 38652
rect 7782 38650 7838 38652
rect 7862 38650 7918 38652
rect 7622 38598 7648 38650
rect 7648 38598 7678 38650
rect 7702 38598 7712 38650
rect 7712 38598 7758 38650
rect 7782 38598 7828 38650
rect 7828 38598 7838 38650
rect 7862 38598 7892 38650
rect 7892 38598 7918 38650
rect 7622 38596 7678 38598
rect 7702 38596 7758 38598
rect 7782 38596 7838 38598
rect 7862 38596 7918 38598
rect 7378 37304 7434 37360
rect 7622 37562 7678 37564
rect 7702 37562 7758 37564
rect 7782 37562 7838 37564
rect 7862 37562 7918 37564
rect 7622 37510 7648 37562
rect 7648 37510 7678 37562
rect 7702 37510 7712 37562
rect 7712 37510 7758 37562
rect 7782 37510 7828 37562
rect 7828 37510 7838 37562
rect 7862 37510 7892 37562
rect 7892 37510 7918 37562
rect 7622 37508 7678 37510
rect 7702 37508 7758 37510
rect 7782 37508 7838 37510
rect 7862 37508 7918 37510
rect 7930 37032 7986 37088
rect 7622 36474 7678 36476
rect 7702 36474 7758 36476
rect 7782 36474 7838 36476
rect 7862 36474 7918 36476
rect 7622 36422 7648 36474
rect 7648 36422 7678 36474
rect 7702 36422 7712 36474
rect 7712 36422 7758 36474
rect 7782 36422 7828 36474
rect 7828 36422 7838 36474
rect 7862 36422 7892 36474
rect 7892 36422 7918 36474
rect 7622 36420 7678 36422
rect 7702 36420 7758 36422
rect 7782 36420 7838 36422
rect 7862 36420 7918 36422
rect 7622 35386 7678 35388
rect 7702 35386 7758 35388
rect 7782 35386 7838 35388
rect 7862 35386 7918 35388
rect 7622 35334 7648 35386
rect 7648 35334 7678 35386
rect 7702 35334 7712 35386
rect 7712 35334 7758 35386
rect 7782 35334 7828 35386
rect 7828 35334 7838 35386
rect 7862 35334 7892 35386
rect 7892 35334 7918 35386
rect 7622 35332 7678 35334
rect 7702 35332 7758 35334
rect 7782 35332 7838 35334
rect 7862 35332 7918 35334
rect 7930 34584 7986 34640
rect 7470 34448 7526 34504
rect 7622 34298 7678 34300
rect 7702 34298 7758 34300
rect 7782 34298 7838 34300
rect 7862 34298 7918 34300
rect 7622 34246 7648 34298
rect 7648 34246 7678 34298
rect 7702 34246 7712 34298
rect 7712 34246 7758 34298
rect 7782 34246 7828 34298
rect 7828 34246 7838 34298
rect 7862 34246 7892 34298
rect 7892 34246 7918 34298
rect 7622 34244 7678 34246
rect 7702 34244 7758 34246
rect 7782 34244 7838 34246
rect 7862 34244 7918 34246
rect 7622 33210 7678 33212
rect 7702 33210 7758 33212
rect 7782 33210 7838 33212
rect 7862 33210 7918 33212
rect 7622 33158 7648 33210
rect 7648 33158 7678 33210
rect 7702 33158 7712 33210
rect 7712 33158 7758 33210
rect 7782 33158 7828 33210
rect 7828 33158 7838 33210
rect 7862 33158 7892 33210
rect 7892 33158 7918 33210
rect 7622 33156 7678 33158
rect 7702 33156 7758 33158
rect 7782 33156 7838 33158
rect 7862 33156 7918 33158
rect 7378 32680 7434 32736
rect 8114 39616 8170 39672
rect 8022 32564 8078 32600
rect 8022 32544 8024 32564
rect 8024 32544 8076 32564
rect 8076 32544 8078 32564
rect 7622 32122 7678 32124
rect 7702 32122 7758 32124
rect 7782 32122 7838 32124
rect 7862 32122 7918 32124
rect 7622 32070 7648 32122
rect 7648 32070 7678 32122
rect 7702 32070 7712 32122
rect 7712 32070 7758 32122
rect 7782 32070 7828 32122
rect 7828 32070 7838 32122
rect 7862 32070 7892 32122
rect 7892 32070 7918 32122
rect 7622 32068 7678 32070
rect 7702 32068 7758 32070
rect 7782 32068 7838 32070
rect 7862 32068 7918 32070
rect 7194 29144 7250 29200
rect 7010 24384 7066 24440
rect 6642 24012 6644 24032
rect 6644 24012 6696 24032
rect 6696 24012 6698 24032
rect 6642 23976 6698 24012
rect 7622 31034 7678 31036
rect 7702 31034 7758 31036
rect 7782 31034 7838 31036
rect 7862 31034 7918 31036
rect 7622 30982 7648 31034
rect 7648 30982 7678 31034
rect 7702 30982 7712 31034
rect 7712 30982 7758 31034
rect 7782 30982 7828 31034
rect 7828 30982 7838 31034
rect 7862 30982 7892 31034
rect 7892 30982 7918 31034
rect 7622 30980 7678 30982
rect 7702 30980 7758 30982
rect 7782 30980 7838 30982
rect 7862 30980 7918 30982
rect 7654 30540 7656 30560
rect 7656 30540 7708 30560
rect 7708 30540 7710 30560
rect 7654 30504 7710 30540
rect 7622 29946 7678 29948
rect 7702 29946 7758 29948
rect 7782 29946 7838 29948
rect 7862 29946 7918 29948
rect 7622 29894 7648 29946
rect 7648 29894 7678 29946
rect 7702 29894 7712 29946
rect 7712 29894 7758 29946
rect 7782 29894 7828 29946
rect 7828 29894 7838 29946
rect 7862 29894 7892 29946
rect 7892 29894 7918 29946
rect 7622 29892 7678 29894
rect 7702 29892 7758 29894
rect 7782 29892 7838 29894
rect 7862 29892 7918 29894
rect 8114 29008 8170 29064
rect 7622 28858 7678 28860
rect 7702 28858 7758 28860
rect 7782 28858 7838 28860
rect 7862 28858 7918 28860
rect 7622 28806 7648 28858
rect 7648 28806 7678 28858
rect 7702 28806 7712 28858
rect 7712 28806 7758 28858
rect 7782 28806 7828 28858
rect 7828 28806 7838 28858
rect 7862 28806 7892 28858
rect 7892 28806 7918 28858
rect 7622 28804 7678 28806
rect 7702 28804 7758 28806
rect 7782 28804 7838 28806
rect 7862 28804 7918 28806
rect 8114 28600 8170 28656
rect 7622 27770 7678 27772
rect 7702 27770 7758 27772
rect 7782 27770 7838 27772
rect 7862 27770 7918 27772
rect 7622 27718 7648 27770
rect 7648 27718 7678 27770
rect 7702 27718 7712 27770
rect 7712 27718 7758 27770
rect 7782 27718 7828 27770
rect 7828 27718 7838 27770
rect 7862 27718 7892 27770
rect 7892 27718 7918 27770
rect 7622 27716 7678 27718
rect 7702 27716 7758 27718
rect 7782 27716 7838 27718
rect 7862 27716 7918 27718
rect 7622 26682 7678 26684
rect 7702 26682 7758 26684
rect 7782 26682 7838 26684
rect 7862 26682 7918 26684
rect 7622 26630 7648 26682
rect 7648 26630 7678 26682
rect 7702 26630 7712 26682
rect 7712 26630 7758 26682
rect 7782 26630 7828 26682
rect 7828 26630 7838 26682
rect 7862 26630 7892 26682
rect 7892 26630 7918 26682
rect 7622 26628 7678 26630
rect 7702 26628 7758 26630
rect 7782 26628 7838 26630
rect 7862 26628 7918 26630
rect 7622 25594 7678 25596
rect 7702 25594 7758 25596
rect 7782 25594 7838 25596
rect 7862 25594 7918 25596
rect 7622 25542 7648 25594
rect 7648 25542 7678 25594
rect 7702 25542 7712 25594
rect 7712 25542 7758 25594
rect 7782 25542 7828 25594
rect 7828 25542 7838 25594
rect 7862 25542 7892 25594
rect 7892 25542 7918 25594
rect 7622 25540 7678 25542
rect 7702 25540 7758 25542
rect 7782 25540 7838 25542
rect 7862 25540 7918 25542
rect 7622 24506 7678 24508
rect 7702 24506 7758 24508
rect 7782 24506 7838 24508
rect 7862 24506 7918 24508
rect 7622 24454 7648 24506
rect 7648 24454 7678 24506
rect 7702 24454 7712 24506
rect 7712 24454 7758 24506
rect 7782 24454 7828 24506
rect 7828 24454 7838 24506
rect 7862 24454 7892 24506
rect 7892 24454 7918 24506
rect 7622 24452 7678 24454
rect 7702 24452 7758 24454
rect 7782 24452 7838 24454
rect 7862 24452 7918 24454
rect 7470 23976 7526 24032
rect 7622 23418 7678 23420
rect 7702 23418 7758 23420
rect 7782 23418 7838 23420
rect 7862 23418 7918 23420
rect 7622 23366 7648 23418
rect 7648 23366 7678 23418
rect 7702 23366 7712 23418
rect 7712 23366 7758 23418
rect 7782 23366 7828 23418
rect 7828 23366 7838 23418
rect 7862 23366 7892 23418
rect 7892 23366 7918 23418
rect 7622 23364 7678 23366
rect 7702 23364 7758 23366
rect 7782 23364 7838 23366
rect 7862 23364 7918 23366
rect 7622 22330 7678 22332
rect 7702 22330 7758 22332
rect 7782 22330 7838 22332
rect 7862 22330 7918 22332
rect 7622 22278 7648 22330
rect 7648 22278 7678 22330
rect 7702 22278 7712 22330
rect 7712 22278 7758 22330
rect 7782 22278 7828 22330
rect 7828 22278 7838 22330
rect 7862 22278 7892 22330
rect 7892 22278 7918 22330
rect 7622 22276 7678 22278
rect 7702 22276 7758 22278
rect 7782 22276 7838 22278
rect 7862 22276 7918 22278
rect 8114 22208 8170 22264
rect 8390 46824 8446 46880
rect 8574 46144 8630 46200
rect 8758 50904 8814 50960
rect 8758 50632 8814 50688
rect 8942 51176 8998 51232
rect 8942 50904 8998 50960
rect 8298 42744 8354 42800
rect 8298 38528 8354 38584
rect 8298 38392 8354 38448
rect 8298 33768 8354 33824
rect 8298 32680 8354 32736
rect 10046 65900 10048 65920
rect 10048 65900 10100 65920
rect 10100 65900 10102 65920
rect 10046 65864 10102 65900
rect 9402 62892 9458 62928
rect 9402 62872 9404 62892
rect 9404 62872 9456 62892
rect 9456 62872 9458 62892
rect 9954 63960 10010 64016
rect 9218 54168 9274 54224
rect 9218 51720 9274 51776
rect 9218 49816 9274 49872
rect 8942 45600 8998 45656
rect 9034 44104 9090 44160
rect 8942 41656 8998 41712
rect 10414 67224 10470 67280
rect 10046 62872 10102 62928
rect 10046 61240 10102 61296
rect 9954 60696 10010 60752
rect 9862 59336 9918 59392
rect 9586 57976 9642 58032
rect 9494 56208 9550 56264
rect 9494 55664 9550 55720
rect 9678 57044 9734 57080
rect 9678 57024 9680 57044
rect 9680 57024 9732 57044
rect 9732 57024 9734 57044
rect 9678 55392 9734 55448
rect 9494 53896 9550 53952
rect 9862 56344 9918 56400
rect 10046 59336 10102 59392
rect 9678 52808 9734 52864
rect 9586 51584 9642 51640
rect 9678 51312 9734 51368
rect 9218 41520 9274 41576
rect 9034 40452 9090 40488
rect 9034 40432 9036 40452
rect 9036 40432 9088 40452
rect 9088 40432 9090 40452
rect 9034 38256 9090 38312
rect 9218 38936 9274 38992
rect 9218 38664 9274 38720
rect 9678 49952 9734 50008
rect 9586 48628 9588 48648
rect 9588 48628 9640 48648
rect 9640 48628 9642 48648
rect 9586 48592 9642 48628
rect 9954 54168 10010 54224
rect 9954 53080 10010 53136
rect 10956 71834 11012 71836
rect 11036 71834 11092 71836
rect 11116 71834 11172 71836
rect 11196 71834 11252 71836
rect 10956 71782 10982 71834
rect 10982 71782 11012 71834
rect 11036 71782 11046 71834
rect 11046 71782 11092 71834
rect 11116 71782 11162 71834
rect 11162 71782 11172 71834
rect 11196 71782 11226 71834
rect 11226 71782 11252 71834
rect 10956 71780 11012 71782
rect 11036 71780 11092 71782
rect 11116 71780 11172 71782
rect 11196 71780 11252 71782
rect 10956 70746 11012 70748
rect 11036 70746 11092 70748
rect 11116 70746 11172 70748
rect 11196 70746 11252 70748
rect 10956 70694 10982 70746
rect 10982 70694 11012 70746
rect 11036 70694 11046 70746
rect 11046 70694 11092 70746
rect 11116 70694 11162 70746
rect 11162 70694 11172 70746
rect 11196 70694 11226 70746
rect 11226 70694 11252 70746
rect 10956 70692 11012 70694
rect 11036 70692 11092 70694
rect 11116 70692 11172 70694
rect 11196 70692 11252 70694
rect 10956 69658 11012 69660
rect 11036 69658 11092 69660
rect 11116 69658 11172 69660
rect 11196 69658 11252 69660
rect 10956 69606 10982 69658
rect 10982 69606 11012 69658
rect 11036 69606 11046 69658
rect 11046 69606 11092 69658
rect 11116 69606 11162 69658
rect 11162 69606 11172 69658
rect 11196 69606 11226 69658
rect 11226 69606 11252 69658
rect 10956 69604 11012 69606
rect 11036 69604 11092 69606
rect 11116 69604 11172 69606
rect 11196 69604 11252 69606
rect 10598 65864 10654 65920
rect 10956 68570 11012 68572
rect 11036 68570 11092 68572
rect 11116 68570 11172 68572
rect 11196 68570 11252 68572
rect 10956 68518 10982 68570
rect 10982 68518 11012 68570
rect 11036 68518 11046 68570
rect 11046 68518 11092 68570
rect 11116 68518 11162 68570
rect 11162 68518 11172 68570
rect 11196 68518 11226 68570
rect 11226 68518 11252 68570
rect 10956 68516 11012 68518
rect 11036 68516 11092 68518
rect 11116 68516 11172 68518
rect 11196 68516 11252 68518
rect 11794 72528 11850 72564
rect 11610 70352 11666 70408
rect 11518 70080 11574 70136
rect 10956 67482 11012 67484
rect 11036 67482 11092 67484
rect 11116 67482 11172 67484
rect 11196 67482 11252 67484
rect 10956 67430 10982 67482
rect 10982 67430 11012 67482
rect 11036 67430 11046 67482
rect 11046 67430 11092 67482
rect 11116 67430 11162 67482
rect 11162 67430 11172 67482
rect 11196 67430 11226 67482
rect 11226 67430 11252 67482
rect 10956 67428 11012 67430
rect 11036 67428 11092 67430
rect 11116 67428 11172 67430
rect 11196 67428 11252 67430
rect 10956 66394 11012 66396
rect 11036 66394 11092 66396
rect 11116 66394 11172 66396
rect 11196 66394 11252 66396
rect 10956 66342 10982 66394
rect 10982 66342 11012 66394
rect 11036 66342 11046 66394
rect 11046 66342 11092 66394
rect 11116 66342 11162 66394
rect 11162 66342 11172 66394
rect 11196 66342 11226 66394
rect 11226 66342 11252 66394
rect 10956 66340 11012 66342
rect 11036 66340 11092 66342
rect 11116 66340 11172 66342
rect 11196 66340 11252 66342
rect 10782 65184 10838 65240
rect 10414 60152 10470 60208
rect 10414 59336 10470 59392
rect 10414 58384 10470 58440
rect 10414 56380 10416 56400
rect 10416 56380 10468 56400
rect 10468 56380 10470 56400
rect 10414 56344 10470 56380
rect 10230 53100 10286 53136
rect 10230 53080 10232 53100
rect 10232 53080 10284 53100
rect 10284 53080 10286 53100
rect 10138 52436 10140 52456
rect 10140 52436 10192 52456
rect 10192 52436 10194 52456
rect 10138 52400 10194 52436
rect 10138 51448 10194 51504
rect 10138 50768 10194 50824
rect 10138 49836 10194 49872
rect 10138 49816 10140 49836
rect 10140 49816 10192 49836
rect 10192 49816 10194 49836
rect 10322 51060 10378 51096
rect 10322 51040 10324 51060
rect 10324 51040 10376 51060
rect 10376 51040 10378 51060
rect 10322 50804 10324 50824
rect 10324 50804 10376 50824
rect 10376 50804 10378 50824
rect 10322 50768 10378 50804
rect 10230 49680 10286 49736
rect 9954 49136 10010 49192
rect 9862 45500 9864 45520
rect 9864 45500 9916 45520
rect 9916 45500 9918 45520
rect 9862 45464 9918 45500
rect 9954 45192 10010 45248
rect 9586 42608 9642 42664
rect 9862 43732 9864 43752
rect 9864 43732 9916 43752
rect 9916 43732 9918 43752
rect 9862 43696 9918 43732
rect 9494 41384 9550 41440
rect 9402 39516 9404 39536
rect 9404 39516 9456 39536
rect 9456 39516 9458 39536
rect 9402 39480 9458 39516
rect 9126 37848 9182 37904
rect 8942 34584 8998 34640
rect 8758 31728 8814 31784
rect 9678 38664 9734 38720
rect 9586 37712 9642 37768
rect 9954 38664 10010 38720
rect 9126 34040 9182 34096
rect 9310 32836 9366 32872
rect 9310 32816 9312 32836
rect 9312 32816 9364 32836
rect 9364 32816 9366 32836
rect 9034 25200 9090 25256
rect 7622 21242 7678 21244
rect 7702 21242 7758 21244
rect 7782 21242 7838 21244
rect 7862 21242 7918 21244
rect 7622 21190 7648 21242
rect 7648 21190 7678 21242
rect 7702 21190 7712 21242
rect 7712 21190 7758 21242
rect 7782 21190 7828 21242
rect 7828 21190 7838 21242
rect 7862 21190 7892 21242
rect 7892 21190 7918 21242
rect 7622 21188 7678 21190
rect 7702 21188 7758 21190
rect 7782 21188 7838 21190
rect 7862 21188 7918 21190
rect 7622 20154 7678 20156
rect 7702 20154 7758 20156
rect 7782 20154 7838 20156
rect 7862 20154 7918 20156
rect 7622 20102 7648 20154
rect 7648 20102 7678 20154
rect 7702 20102 7712 20154
rect 7712 20102 7758 20154
rect 7782 20102 7828 20154
rect 7828 20102 7838 20154
rect 7862 20102 7892 20154
rect 7892 20102 7918 20154
rect 7622 20100 7678 20102
rect 7702 20100 7758 20102
rect 7782 20100 7838 20102
rect 7862 20100 7918 20102
rect 4289 18522 4345 18524
rect 4369 18522 4425 18524
rect 4449 18522 4505 18524
rect 4529 18522 4585 18524
rect 4289 18470 4315 18522
rect 4315 18470 4345 18522
rect 4369 18470 4379 18522
rect 4379 18470 4425 18522
rect 4449 18470 4495 18522
rect 4495 18470 4505 18522
rect 4529 18470 4559 18522
rect 4559 18470 4585 18522
rect 4289 18468 4345 18470
rect 4369 18468 4425 18470
rect 4449 18468 4505 18470
rect 4529 18468 4585 18470
rect 4289 17434 4345 17436
rect 4369 17434 4425 17436
rect 4449 17434 4505 17436
rect 4529 17434 4585 17436
rect 4289 17382 4315 17434
rect 4315 17382 4345 17434
rect 4369 17382 4379 17434
rect 4379 17382 4425 17434
rect 4449 17382 4495 17434
rect 4495 17382 4505 17434
rect 4529 17382 4559 17434
rect 4559 17382 4585 17434
rect 4289 17380 4345 17382
rect 4369 17380 4425 17382
rect 4449 17380 4505 17382
rect 4529 17380 4585 17382
rect 4289 16346 4345 16348
rect 4369 16346 4425 16348
rect 4449 16346 4505 16348
rect 4529 16346 4585 16348
rect 4289 16294 4315 16346
rect 4315 16294 4345 16346
rect 4369 16294 4379 16346
rect 4379 16294 4425 16346
rect 4449 16294 4495 16346
rect 4495 16294 4505 16346
rect 4529 16294 4559 16346
rect 4559 16294 4585 16346
rect 4289 16292 4345 16294
rect 4369 16292 4425 16294
rect 4449 16292 4505 16294
rect 4529 16292 4585 16294
rect 4289 15258 4345 15260
rect 4369 15258 4425 15260
rect 4449 15258 4505 15260
rect 4529 15258 4585 15260
rect 4289 15206 4315 15258
rect 4315 15206 4345 15258
rect 4369 15206 4379 15258
rect 4379 15206 4425 15258
rect 4449 15206 4495 15258
rect 4495 15206 4505 15258
rect 4529 15206 4559 15258
rect 4559 15206 4585 15258
rect 4289 15204 4345 15206
rect 4369 15204 4425 15206
rect 4449 15204 4505 15206
rect 4529 15204 4585 15206
rect 3238 14592 3294 14648
rect 5078 14864 5134 14920
rect 3974 14356 3976 14376
rect 3976 14356 4028 14376
rect 4028 14356 4030 14376
rect 3974 14320 4030 14356
rect 4289 14170 4345 14172
rect 4369 14170 4425 14172
rect 4449 14170 4505 14172
rect 4529 14170 4585 14172
rect 4289 14118 4315 14170
rect 4315 14118 4345 14170
rect 4369 14118 4379 14170
rect 4379 14118 4425 14170
rect 4449 14118 4495 14170
rect 4495 14118 4505 14170
rect 4529 14118 4559 14170
rect 4559 14118 4585 14170
rect 4289 14116 4345 14118
rect 4369 14116 4425 14118
rect 4449 14116 4505 14118
rect 4529 14116 4585 14118
rect 3790 13776 3846 13832
rect 8482 19488 8538 19544
rect 7622 19066 7678 19068
rect 7702 19066 7758 19068
rect 7782 19066 7838 19068
rect 7862 19066 7918 19068
rect 7622 19014 7648 19066
rect 7648 19014 7678 19066
rect 7702 19014 7712 19066
rect 7712 19014 7758 19066
rect 7782 19014 7828 19066
rect 7828 19014 7838 19066
rect 7862 19014 7892 19066
rect 7892 19014 7918 19066
rect 7622 19012 7678 19014
rect 7702 19012 7758 19014
rect 7782 19012 7838 19014
rect 7862 19012 7918 19014
rect 7622 17978 7678 17980
rect 7702 17978 7758 17980
rect 7782 17978 7838 17980
rect 7862 17978 7918 17980
rect 7622 17926 7648 17978
rect 7648 17926 7678 17978
rect 7702 17926 7712 17978
rect 7712 17926 7758 17978
rect 7782 17926 7828 17978
rect 7828 17926 7838 17978
rect 7862 17926 7892 17978
rect 7892 17926 7918 17978
rect 7622 17924 7678 17926
rect 7702 17924 7758 17926
rect 7782 17924 7838 17926
rect 7862 17924 7918 17926
rect 8022 16940 8024 16960
rect 8024 16940 8076 16960
rect 8076 16940 8078 16960
rect 8022 16904 8078 16940
rect 7622 16890 7678 16892
rect 7702 16890 7758 16892
rect 7782 16890 7838 16892
rect 7862 16890 7918 16892
rect 7622 16838 7648 16890
rect 7648 16838 7678 16890
rect 7702 16838 7712 16890
rect 7712 16838 7758 16890
rect 7782 16838 7828 16890
rect 7828 16838 7838 16890
rect 7862 16838 7892 16890
rect 7892 16838 7918 16890
rect 7622 16836 7678 16838
rect 7702 16836 7758 16838
rect 7782 16836 7838 16838
rect 7862 16836 7918 16838
rect 6918 16632 6974 16688
rect 5906 16088 5962 16144
rect 4618 13268 4620 13288
rect 4620 13268 4672 13288
rect 4672 13268 4674 13288
rect 4618 13232 4674 13268
rect 4289 13082 4345 13084
rect 4369 13082 4425 13084
rect 4449 13082 4505 13084
rect 4529 13082 4585 13084
rect 4289 13030 4315 13082
rect 4315 13030 4345 13082
rect 4369 13030 4379 13082
rect 4379 13030 4425 13082
rect 4449 13030 4495 13082
rect 4495 13030 4505 13082
rect 4529 13030 4559 13082
rect 4559 13030 4585 13082
rect 4289 13028 4345 13030
rect 4369 13028 4425 13030
rect 4449 13028 4505 13030
rect 4529 13028 4585 13030
rect 3054 12824 3110 12880
rect 2962 12688 3018 12744
rect 5630 13096 5686 13152
rect 3790 12300 3846 12336
rect 3790 12280 3792 12300
rect 3792 12280 3844 12300
rect 3844 12280 3846 12300
rect 4289 11994 4345 11996
rect 4369 11994 4425 11996
rect 4449 11994 4505 11996
rect 4529 11994 4585 11996
rect 4289 11942 4315 11994
rect 4315 11942 4345 11994
rect 4369 11942 4379 11994
rect 4379 11942 4425 11994
rect 4449 11942 4495 11994
rect 4495 11942 4505 11994
rect 4529 11942 4559 11994
rect 4559 11942 4585 11994
rect 4289 11940 4345 11942
rect 4369 11940 4425 11942
rect 4449 11940 4505 11942
rect 4529 11940 4585 11942
rect 7622 15802 7678 15804
rect 7702 15802 7758 15804
rect 7782 15802 7838 15804
rect 7862 15802 7918 15804
rect 7622 15750 7648 15802
rect 7648 15750 7678 15802
rect 7702 15750 7712 15802
rect 7712 15750 7758 15802
rect 7782 15750 7828 15802
rect 7828 15750 7838 15802
rect 7862 15750 7892 15802
rect 7892 15750 7918 15802
rect 7622 15748 7678 15750
rect 7702 15748 7758 15750
rect 7782 15748 7838 15750
rect 7862 15748 7918 15750
rect 7286 14456 7342 14512
rect 7622 14714 7678 14716
rect 7702 14714 7758 14716
rect 7782 14714 7838 14716
rect 7862 14714 7918 14716
rect 7622 14662 7648 14714
rect 7648 14662 7678 14714
rect 7702 14662 7712 14714
rect 7712 14662 7758 14714
rect 7782 14662 7828 14714
rect 7828 14662 7838 14714
rect 7862 14662 7892 14714
rect 7892 14662 7918 14714
rect 7622 14660 7678 14662
rect 7702 14660 7758 14662
rect 7782 14660 7838 14662
rect 7862 14660 7918 14662
rect 8298 13912 8354 13968
rect 7622 13626 7678 13628
rect 7702 13626 7758 13628
rect 7782 13626 7838 13628
rect 7862 13626 7918 13628
rect 7622 13574 7648 13626
rect 7648 13574 7678 13626
rect 7702 13574 7712 13626
rect 7712 13574 7758 13626
rect 7782 13574 7828 13626
rect 7828 13574 7838 13626
rect 7862 13574 7892 13626
rect 7892 13574 7918 13626
rect 7622 13572 7678 13574
rect 7702 13572 7758 13574
rect 7782 13572 7838 13574
rect 7862 13572 7918 13574
rect 5814 11736 5870 11792
rect 3146 10140 3148 10160
rect 3148 10140 3200 10160
rect 3200 10140 3202 10160
rect 3146 10104 3202 10140
rect 3974 11056 4030 11112
rect 4289 10906 4345 10908
rect 4369 10906 4425 10908
rect 4449 10906 4505 10908
rect 4529 10906 4585 10908
rect 4289 10854 4315 10906
rect 4315 10854 4345 10906
rect 4369 10854 4379 10906
rect 4379 10854 4425 10906
rect 4449 10854 4495 10906
rect 4495 10854 4505 10906
rect 4529 10854 4559 10906
rect 4559 10854 4585 10906
rect 4289 10852 4345 10854
rect 4369 10852 4425 10854
rect 4449 10852 4505 10854
rect 4529 10852 4585 10854
rect 8298 12688 8354 12744
rect 7622 12538 7678 12540
rect 7702 12538 7758 12540
rect 7782 12538 7838 12540
rect 7862 12538 7918 12540
rect 7622 12486 7648 12538
rect 7648 12486 7678 12538
rect 7702 12486 7712 12538
rect 7712 12486 7758 12538
rect 7782 12486 7828 12538
rect 7828 12486 7838 12538
rect 7862 12486 7892 12538
rect 7892 12486 7918 12538
rect 7622 12484 7678 12486
rect 7702 12484 7758 12486
rect 7782 12484 7838 12486
rect 7862 12484 7918 12486
rect 9586 34448 9642 34504
rect 10230 45364 10232 45384
rect 10232 45364 10284 45384
rect 10284 45364 10286 45384
rect 10230 45328 10286 45364
rect 10690 64776 10746 64832
rect 11242 65728 11298 65784
rect 10956 65306 11012 65308
rect 11036 65306 11092 65308
rect 11116 65306 11172 65308
rect 11196 65306 11252 65308
rect 10956 65254 10982 65306
rect 10982 65254 11012 65306
rect 11036 65254 11046 65306
rect 11046 65254 11092 65306
rect 11116 65254 11162 65306
rect 11162 65254 11172 65306
rect 11196 65254 11226 65306
rect 11226 65254 11252 65306
rect 10956 65252 11012 65254
rect 11036 65252 11092 65254
rect 11116 65252 11172 65254
rect 11196 65252 11252 65254
rect 10956 64218 11012 64220
rect 11036 64218 11092 64220
rect 11116 64218 11172 64220
rect 11196 64218 11252 64220
rect 10956 64166 10982 64218
rect 10982 64166 11012 64218
rect 11036 64166 11046 64218
rect 11046 64166 11092 64218
rect 11116 64166 11162 64218
rect 11162 64166 11172 64218
rect 11196 64166 11226 64218
rect 11226 64166 11252 64218
rect 10956 64164 11012 64166
rect 11036 64164 11092 64166
rect 11116 64164 11172 64166
rect 11196 64164 11252 64166
rect 11150 63552 11206 63608
rect 10956 63130 11012 63132
rect 11036 63130 11092 63132
rect 11116 63130 11172 63132
rect 11196 63130 11252 63132
rect 10956 63078 10982 63130
rect 10982 63078 11012 63130
rect 11036 63078 11046 63130
rect 11046 63078 11092 63130
rect 11116 63078 11162 63130
rect 11162 63078 11172 63130
rect 11196 63078 11226 63130
rect 11226 63078 11252 63130
rect 10956 63076 11012 63078
rect 11036 63076 11092 63078
rect 11116 63076 11172 63078
rect 11196 63076 11252 63078
rect 10598 62192 10654 62248
rect 10782 62600 10838 62656
rect 11610 68176 11666 68232
rect 11518 62600 11574 62656
rect 10956 62042 11012 62044
rect 11036 62042 11092 62044
rect 11116 62042 11172 62044
rect 11196 62042 11252 62044
rect 10956 61990 10982 62042
rect 10982 61990 11012 62042
rect 11036 61990 11046 62042
rect 11046 61990 11092 62042
rect 11116 61990 11162 62042
rect 11162 61990 11172 62042
rect 11196 61990 11226 62042
rect 11226 61990 11252 62042
rect 10956 61988 11012 61990
rect 11036 61988 11092 61990
rect 11116 61988 11172 61990
rect 11196 61988 11252 61990
rect 11058 61260 11114 61296
rect 11058 61240 11060 61260
rect 11060 61240 11112 61260
rect 11112 61240 11114 61260
rect 10956 60954 11012 60956
rect 11036 60954 11092 60956
rect 11116 60954 11172 60956
rect 11196 60954 11252 60956
rect 10956 60902 10982 60954
rect 10982 60902 11012 60954
rect 11036 60902 11046 60954
rect 11046 60902 11092 60954
rect 11116 60902 11162 60954
rect 11162 60902 11172 60954
rect 11196 60902 11226 60954
rect 11226 60902 11252 60954
rect 10956 60900 11012 60902
rect 11036 60900 11092 60902
rect 11116 60900 11172 60902
rect 11196 60900 11252 60902
rect 10874 60696 10930 60752
rect 10782 59744 10838 59800
rect 10690 59508 10692 59528
rect 10692 59508 10744 59528
rect 10744 59508 10746 59528
rect 10690 59472 10746 59508
rect 10690 59064 10746 59120
rect 10690 56072 10746 56128
rect 10506 54032 10562 54088
rect 10598 53644 10654 53680
rect 10598 53624 10600 53644
rect 10600 53624 10652 53644
rect 10652 53624 10654 53644
rect 10598 52536 10654 52592
rect 10956 59866 11012 59868
rect 11036 59866 11092 59868
rect 11116 59866 11172 59868
rect 11196 59866 11252 59868
rect 10956 59814 10982 59866
rect 10982 59814 11012 59866
rect 11036 59814 11046 59866
rect 11046 59814 11092 59866
rect 11116 59814 11162 59866
rect 11162 59814 11172 59866
rect 11196 59814 11226 59866
rect 11226 59814 11252 59866
rect 10956 59812 11012 59814
rect 11036 59812 11092 59814
rect 11116 59812 11172 59814
rect 11196 59812 11252 59814
rect 10956 58778 11012 58780
rect 11036 58778 11092 58780
rect 11116 58778 11172 58780
rect 11196 58778 11252 58780
rect 10956 58726 10982 58778
rect 10982 58726 11012 58778
rect 11036 58726 11046 58778
rect 11046 58726 11092 58778
rect 11116 58726 11162 58778
rect 11162 58726 11172 58778
rect 11196 58726 11226 58778
rect 11226 58726 11252 58778
rect 10956 58724 11012 58726
rect 11036 58724 11092 58726
rect 11116 58724 11172 58726
rect 11196 58724 11252 58726
rect 11150 57840 11206 57896
rect 10956 57690 11012 57692
rect 11036 57690 11092 57692
rect 11116 57690 11172 57692
rect 11196 57690 11252 57692
rect 10956 57638 10982 57690
rect 10982 57638 11012 57690
rect 11036 57638 11046 57690
rect 11046 57638 11092 57690
rect 11116 57638 11162 57690
rect 11162 57638 11172 57690
rect 11196 57638 11226 57690
rect 11226 57638 11252 57690
rect 10956 57636 11012 57638
rect 11036 57636 11092 57638
rect 11116 57636 11172 57638
rect 11196 57636 11252 57638
rect 10966 57432 11022 57488
rect 10956 56602 11012 56604
rect 11036 56602 11092 56604
rect 11116 56602 11172 56604
rect 11196 56602 11252 56604
rect 10956 56550 10982 56602
rect 10982 56550 11012 56602
rect 11036 56550 11046 56602
rect 11046 56550 11092 56602
rect 11116 56550 11162 56602
rect 11162 56550 11172 56602
rect 11196 56550 11226 56602
rect 11226 56550 11252 56602
rect 10956 56548 11012 56550
rect 11036 56548 11092 56550
rect 11116 56548 11172 56550
rect 11196 56548 11252 56550
rect 10966 56072 11022 56128
rect 11150 55664 11206 55720
rect 10956 55514 11012 55516
rect 11036 55514 11092 55516
rect 11116 55514 11172 55516
rect 11196 55514 11252 55516
rect 10956 55462 10982 55514
rect 10982 55462 11012 55514
rect 11036 55462 11046 55514
rect 11046 55462 11092 55514
rect 11116 55462 11162 55514
rect 11162 55462 11172 55514
rect 11196 55462 11226 55514
rect 11226 55462 11252 55514
rect 10956 55460 11012 55462
rect 11036 55460 11092 55462
rect 11116 55460 11172 55462
rect 11196 55460 11252 55462
rect 10956 54426 11012 54428
rect 11036 54426 11092 54428
rect 11116 54426 11172 54428
rect 11196 54426 11252 54428
rect 10956 54374 10982 54426
rect 10982 54374 11012 54426
rect 11036 54374 11046 54426
rect 11046 54374 11092 54426
rect 11116 54374 11162 54426
rect 11162 54374 11172 54426
rect 11196 54374 11226 54426
rect 11226 54374 11252 54426
rect 10956 54372 11012 54374
rect 11036 54372 11092 54374
rect 11116 54372 11172 54374
rect 11196 54372 11252 54374
rect 10966 54168 11022 54224
rect 10956 53338 11012 53340
rect 11036 53338 11092 53340
rect 11116 53338 11172 53340
rect 11196 53338 11252 53340
rect 10956 53286 10982 53338
rect 10982 53286 11012 53338
rect 11036 53286 11046 53338
rect 11046 53286 11092 53338
rect 11116 53286 11162 53338
rect 11162 53286 11172 53338
rect 11196 53286 11226 53338
rect 11226 53286 11252 53338
rect 10956 53284 11012 53286
rect 11036 53284 11092 53286
rect 11116 53284 11172 53286
rect 11196 53284 11252 53286
rect 11518 60016 11574 60072
rect 11978 69944 12034 70000
rect 11610 59472 11666 59528
rect 11610 57704 11666 57760
rect 11518 55276 11574 55312
rect 11518 55256 11520 55276
rect 11520 55256 11572 55276
rect 11572 55256 11574 55276
rect 11702 56208 11758 56264
rect 11426 53896 11482 53952
rect 11978 68992 12034 69048
rect 12622 65864 12678 65920
rect 12438 65456 12494 65512
rect 12070 62056 12126 62112
rect 12070 56480 12126 56536
rect 12530 64776 12586 64832
rect 14289 72378 14345 72380
rect 14369 72378 14425 72380
rect 14449 72378 14505 72380
rect 14529 72378 14585 72380
rect 14289 72326 14315 72378
rect 14315 72326 14345 72378
rect 14369 72326 14379 72378
rect 14379 72326 14425 72378
rect 14449 72326 14495 72378
rect 14495 72326 14505 72378
rect 14529 72326 14559 72378
rect 14559 72326 14585 72378
rect 14289 72324 14345 72326
rect 14369 72324 14425 72326
rect 14449 72324 14505 72326
rect 14529 72324 14585 72326
rect 14289 71290 14345 71292
rect 14369 71290 14425 71292
rect 14449 71290 14505 71292
rect 14529 71290 14585 71292
rect 14289 71238 14315 71290
rect 14315 71238 14345 71290
rect 14369 71238 14379 71290
rect 14379 71238 14425 71290
rect 14449 71238 14495 71290
rect 14495 71238 14505 71290
rect 14529 71238 14559 71290
rect 14559 71238 14585 71290
rect 14289 71236 14345 71238
rect 14369 71236 14425 71238
rect 14449 71236 14505 71238
rect 14529 71236 14585 71238
rect 14289 70202 14345 70204
rect 14369 70202 14425 70204
rect 14449 70202 14505 70204
rect 14529 70202 14585 70204
rect 14289 70150 14315 70202
rect 14315 70150 14345 70202
rect 14369 70150 14379 70202
rect 14379 70150 14425 70202
rect 14449 70150 14495 70202
rect 14495 70150 14505 70202
rect 14529 70150 14559 70202
rect 14559 70150 14585 70202
rect 14289 70148 14345 70150
rect 14369 70148 14425 70150
rect 14449 70148 14505 70150
rect 14529 70148 14585 70150
rect 14289 69114 14345 69116
rect 14369 69114 14425 69116
rect 14449 69114 14505 69116
rect 14529 69114 14585 69116
rect 14289 69062 14315 69114
rect 14315 69062 14345 69114
rect 14369 69062 14379 69114
rect 14379 69062 14425 69114
rect 14449 69062 14495 69114
rect 14495 69062 14505 69114
rect 14529 69062 14559 69114
rect 14559 69062 14585 69114
rect 14289 69060 14345 69062
rect 14369 69060 14425 69062
rect 14449 69060 14505 69062
rect 14529 69060 14585 69062
rect 12438 62192 12494 62248
rect 12438 60832 12494 60888
rect 11886 55120 11942 55176
rect 11610 53352 11666 53408
rect 11426 52400 11482 52456
rect 10956 52250 11012 52252
rect 11036 52250 11092 52252
rect 11116 52250 11172 52252
rect 11196 52250 11252 52252
rect 10956 52198 10982 52250
rect 10982 52198 11012 52250
rect 11036 52198 11046 52250
rect 11046 52198 11092 52250
rect 11116 52198 11162 52250
rect 11162 52198 11172 52250
rect 11196 52198 11226 52250
rect 11226 52198 11252 52250
rect 10956 52196 11012 52198
rect 11036 52196 11092 52198
rect 11116 52196 11172 52198
rect 11196 52196 11252 52198
rect 11058 51448 11114 51504
rect 10966 51312 11022 51368
rect 11334 51468 11390 51504
rect 11334 51448 11336 51468
rect 11336 51448 11388 51468
rect 11388 51448 11390 51468
rect 10782 51040 10838 51096
rect 10690 50904 10746 50960
rect 10506 49680 10562 49736
rect 10598 49308 10600 49328
rect 10600 49308 10652 49328
rect 10652 49308 10654 49328
rect 10598 49272 10654 49308
rect 10322 43852 10378 43888
rect 10322 43832 10324 43852
rect 10324 43832 10376 43852
rect 10376 43832 10378 43852
rect 10230 42764 10286 42800
rect 10230 42744 10232 42764
rect 10232 42744 10284 42764
rect 10284 42744 10286 42764
rect 10230 42608 10286 42664
rect 10414 42880 10470 42936
rect 10322 40588 10378 40624
rect 10322 40568 10324 40588
rect 10324 40568 10376 40588
rect 10376 40568 10378 40588
rect 10322 39092 10378 39128
rect 10322 39072 10324 39092
rect 10324 39072 10376 39092
rect 10376 39072 10378 39092
rect 9862 32988 9864 33008
rect 9864 32988 9916 33008
rect 9916 32988 9918 33008
rect 9862 32952 9918 32988
rect 9494 31220 9496 31240
rect 9496 31220 9548 31240
rect 9548 31220 9550 31240
rect 9494 31184 9550 31220
rect 9310 26444 9366 26480
rect 9310 26424 9312 26444
rect 9312 26424 9364 26444
rect 9364 26424 9366 26444
rect 9494 25608 9550 25664
rect 9402 20476 9404 20496
rect 9404 20476 9456 20496
rect 9456 20476 9458 20496
rect 9402 20440 9458 20476
rect 9402 17720 9458 17776
rect 9494 13388 9550 13424
rect 9494 13368 9496 13388
rect 9496 13368 9548 13388
rect 9548 13368 9550 13388
rect 9494 12960 9550 13016
rect 7622 11450 7678 11452
rect 7702 11450 7758 11452
rect 7782 11450 7838 11452
rect 7862 11450 7918 11452
rect 7622 11398 7648 11450
rect 7648 11398 7678 11450
rect 7702 11398 7712 11450
rect 7712 11398 7758 11450
rect 7782 11398 7828 11450
rect 7828 11398 7838 11450
rect 7862 11398 7892 11450
rect 7892 11398 7918 11450
rect 7622 11396 7678 11398
rect 7702 11396 7758 11398
rect 7782 11396 7838 11398
rect 7862 11396 7918 11398
rect 8114 11348 8170 11384
rect 8114 11328 8116 11348
rect 8116 11328 8168 11348
rect 8168 11328 8170 11348
rect 7470 11056 7526 11112
rect 8758 10668 8814 10704
rect 8758 10648 8760 10668
rect 8760 10648 8812 10668
rect 8812 10648 8814 10668
rect 7622 10362 7678 10364
rect 7702 10362 7758 10364
rect 7782 10362 7838 10364
rect 7862 10362 7918 10364
rect 7622 10310 7648 10362
rect 7648 10310 7678 10362
rect 7702 10310 7712 10362
rect 7712 10310 7758 10362
rect 7782 10310 7828 10362
rect 7828 10310 7838 10362
rect 7862 10310 7892 10362
rect 7892 10310 7918 10362
rect 7622 10308 7678 10310
rect 7702 10308 7758 10310
rect 7782 10308 7838 10310
rect 7862 10308 7918 10310
rect 3974 9832 4030 9888
rect 8114 10240 8170 10296
rect 4289 9818 4345 9820
rect 4369 9818 4425 9820
rect 4449 9818 4505 9820
rect 4529 9818 4585 9820
rect 4289 9766 4315 9818
rect 4315 9766 4345 9818
rect 4369 9766 4379 9818
rect 4379 9766 4425 9818
rect 4449 9766 4495 9818
rect 4495 9766 4505 9818
rect 4529 9766 4559 9818
rect 4559 9766 4585 9818
rect 4289 9764 4345 9766
rect 4369 9764 4425 9766
rect 4449 9764 4505 9766
rect 4529 9764 4585 9766
rect 7838 9460 7840 9480
rect 7840 9460 7892 9480
rect 7892 9460 7894 9480
rect 7838 9424 7894 9460
rect 8482 10376 8538 10432
rect 8574 9324 8576 9344
rect 8576 9324 8628 9344
rect 8628 9324 8630 9344
rect 8574 9288 8630 9324
rect 7622 9274 7678 9276
rect 7702 9274 7758 9276
rect 7782 9274 7838 9276
rect 7862 9274 7918 9276
rect 7622 9222 7648 9274
rect 7648 9222 7678 9274
rect 7702 9222 7712 9274
rect 7712 9222 7758 9274
rect 7782 9222 7828 9274
rect 7828 9222 7838 9274
rect 7862 9222 7892 9274
rect 7892 9222 7918 9274
rect 7622 9220 7678 9222
rect 7702 9220 7758 9222
rect 7782 9220 7838 9222
rect 7862 9220 7918 9222
rect 4289 8730 4345 8732
rect 4369 8730 4425 8732
rect 4449 8730 4505 8732
rect 4529 8730 4585 8732
rect 4289 8678 4315 8730
rect 4315 8678 4345 8730
rect 4369 8678 4379 8730
rect 4379 8678 4425 8730
rect 4449 8678 4495 8730
rect 4495 8678 4505 8730
rect 4529 8678 4559 8730
rect 4559 8678 4585 8730
rect 4289 8676 4345 8678
rect 4369 8676 4425 8678
rect 4449 8676 4505 8678
rect 4529 8676 4585 8678
rect 7622 8186 7678 8188
rect 7702 8186 7758 8188
rect 7782 8186 7838 8188
rect 7862 8186 7918 8188
rect 7622 8134 7648 8186
rect 7648 8134 7678 8186
rect 7702 8134 7712 8186
rect 7712 8134 7758 8186
rect 7782 8134 7828 8186
rect 7828 8134 7838 8186
rect 7862 8134 7892 8186
rect 7892 8134 7918 8186
rect 7622 8132 7678 8134
rect 7702 8132 7758 8134
rect 7782 8132 7838 8134
rect 7862 8132 7918 8134
rect 4289 7642 4345 7644
rect 4369 7642 4425 7644
rect 4449 7642 4505 7644
rect 4529 7642 4585 7644
rect 4289 7590 4315 7642
rect 4315 7590 4345 7642
rect 4369 7590 4379 7642
rect 4379 7590 4425 7642
rect 4449 7590 4495 7642
rect 4495 7590 4505 7642
rect 4529 7590 4559 7642
rect 4559 7590 4585 7642
rect 4289 7588 4345 7590
rect 4369 7588 4425 7590
rect 4449 7588 4505 7590
rect 4529 7588 4585 7590
rect 8942 7792 8998 7848
rect 8758 7420 8760 7440
rect 8760 7420 8812 7440
rect 8812 7420 8814 7440
rect 8758 7384 8814 7420
rect 5722 7248 5778 7304
rect 4066 7112 4122 7168
rect 5538 7148 5540 7168
rect 5540 7148 5592 7168
rect 5592 7148 5594 7168
rect 5538 7112 5594 7148
rect 3422 6704 3478 6760
rect 7622 7098 7678 7100
rect 7702 7098 7758 7100
rect 7782 7098 7838 7100
rect 7862 7098 7918 7100
rect 7622 7046 7648 7098
rect 7648 7046 7678 7098
rect 7702 7046 7712 7098
rect 7712 7046 7758 7098
rect 7782 7046 7828 7098
rect 7828 7046 7838 7098
rect 7862 7046 7892 7098
rect 7892 7046 7918 7098
rect 7622 7044 7678 7046
rect 7702 7044 7758 7046
rect 7782 7044 7838 7046
rect 7862 7044 7918 7046
rect 7286 6704 7342 6760
rect 4289 6554 4345 6556
rect 4369 6554 4425 6556
rect 4449 6554 4505 6556
rect 4529 6554 4585 6556
rect 4289 6502 4315 6554
rect 4315 6502 4345 6554
rect 4369 6502 4379 6554
rect 4379 6502 4425 6554
rect 4449 6502 4495 6554
rect 4495 6502 4505 6554
rect 4529 6502 4559 6554
rect 4559 6502 4585 6554
rect 4289 6500 4345 6502
rect 4369 6500 4425 6502
rect 4449 6500 4505 6502
rect 4529 6500 4585 6502
rect 7622 6010 7678 6012
rect 7702 6010 7758 6012
rect 7782 6010 7838 6012
rect 7862 6010 7918 6012
rect 7622 5958 7648 6010
rect 7648 5958 7678 6010
rect 7702 5958 7712 6010
rect 7712 5958 7758 6010
rect 7782 5958 7828 6010
rect 7828 5958 7838 6010
rect 7862 5958 7892 6010
rect 7892 5958 7918 6010
rect 7622 5956 7678 5958
rect 7702 5956 7758 5958
rect 7782 5956 7838 5958
rect 7862 5956 7918 5958
rect 4066 5888 4122 5944
rect 3790 5772 3846 5808
rect 3790 5752 3792 5772
rect 3792 5752 3844 5772
rect 3844 5752 3846 5772
rect 4289 5466 4345 5468
rect 4369 5466 4425 5468
rect 4449 5466 4505 5468
rect 4529 5466 4585 5468
rect 4289 5414 4315 5466
rect 4315 5414 4345 5466
rect 4369 5414 4379 5466
rect 4379 5414 4425 5466
rect 4449 5414 4495 5466
rect 4495 5414 4505 5466
rect 4529 5414 4559 5466
rect 4559 5414 4585 5466
rect 4289 5412 4345 5414
rect 4369 5412 4425 5414
rect 4449 5412 4505 5414
rect 4529 5412 4585 5414
rect 2134 5108 2136 5128
rect 2136 5108 2188 5128
rect 2188 5108 2190 5128
rect 2134 5072 2190 5108
rect 4066 4664 4122 4720
rect 3054 4528 3110 4584
rect 1674 4256 1730 4312
rect 4289 4378 4345 4380
rect 4369 4378 4425 4380
rect 4449 4378 4505 4380
rect 4529 4378 4585 4380
rect 4289 4326 4315 4378
rect 4315 4326 4345 4378
rect 4369 4326 4379 4378
rect 4379 4326 4425 4378
rect 4449 4326 4495 4378
rect 4495 4326 4505 4378
rect 4529 4326 4559 4378
rect 4559 4326 4585 4378
rect 4289 4324 4345 4326
rect 4369 4324 4425 4326
rect 4449 4324 4505 4326
rect 4529 4324 4585 4326
rect 4066 3440 4122 3496
rect 4289 3290 4345 3292
rect 4369 3290 4425 3292
rect 4449 3290 4505 3292
rect 4529 3290 4585 3292
rect 4289 3238 4315 3290
rect 4315 3238 4345 3290
rect 4369 3238 4379 3290
rect 4379 3238 4425 3290
rect 4449 3238 4495 3290
rect 4495 3238 4505 3290
rect 4529 3238 4559 3290
rect 4559 3238 4585 3290
rect 4289 3236 4345 3238
rect 4369 3236 4425 3238
rect 4449 3236 4505 3238
rect 4529 3236 4585 3238
rect 7622 4922 7678 4924
rect 7702 4922 7758 4924
rect 7782 4922 7838 4924
rect 7862 4922 7918 4924
rect 7622 4870 7648 4922
rect 7648 4870 7678 4922
rect 7702 4870 7712 4922
rect 7712 4870 7758 4922
rect 7782 4870 7828 4922
rect 7828 4870 7838 4922
rect 7862 4870 7892 4922
rect 7892 4870 7918 4922
rect 7622 4868 7678 4870
rect 7702 4868 7758 4870
rect 7782 4868 7838 4870
rect 7862 4868 7918 4870
rect 7622 3834 7678 3836
rect 7702 3834 7758 3836
rect 7782 3834 7838 3836
rect 7862 3834 7918 3836
rect 7622 3782 7648 3834
rect 7648 3782 7678 3834
rect 7702 3782 7712 3834
rect 7712 3782 7758 3834
rect 7782 3782 7828 3834
rect 7828 3782 7838 3834
rect 7862 3782 7892 3834
rect 7892 3782 7918 3834
rect 7622 3780 7678 3782
rect 7702 3780 7758 3782
rect 7782 3780 7838 3782
rect 7862 3780 7918 3782
rect 7622 2746 7678 2748
rect 7702 2746 7758 2748
rect 7782 2746 7838 2748
rect 7862 2746 7918 2748
rect 7622 2694 7648 2746
rect 7648 2694 7678 2746
rect 7702 2694 7712 2746
rect 7712 2694 7758 2746
rect 7782 2694 7828 2746
rect 7828 2694 7838 2746
rect 7862 2694 7892 2746
rect 7892 2694 7918 2746
rect 7622 2692 7678 2694
rect 7702 2692 7758 2694
rect 7782 2692 7838 2694
rect 7862 2692 7918 2694
rect 7286 2624 7342 2680
rect 3422 2488 3478 2544
rect 4289 2202 4345 2204
rect 4369 2202 4425 2204
rect 4449 2202 4505 2204
rect 4529 2202 4585 2204
rect 4289 2150 4315 2202
rect 4315 2150 4345 2202
rect 4369 2150 4379 2202
rect 4379 2150 4425 2202
rect 4449 2150 4495 2202
rect 4495 2150 4505 2202
rect 4529 2150 4559 2202
rect 4559 2150 4585 2202
rect 4289 2148 4345 2150
rect 4369 2148 4425 2150
rect 4449 2148 4505 2150
rect 4529 2148 4585 2150
rect 3422 1808 3478 1864
rect 9402 10532 9458 10568
rect 9402 10512 9404 10532
rect 9404 10512 9456 10532
rect 9456 10512 9458 10532
rect 10046 32816 10102 32872
rect 9770 23976 9826 24032
rect 10690 46044 10692 46064
rect 10692 46044 10744 46064
rect 10744 46044 10746 46064
rect 10690 46008 10746 46044
rect 10956 51162 11012 51164
rect 11036 51162 11092 51164
rect 11116 51162 11172 51164
rect 11196 51162 11252 51164
rect 10956 51110 10982 51162
rect 10982 51110 11012 51162
rect 11036 51110 11046 51162
rect 11046 51110 11092 51162
rect 11116 51110 11162 51162
rect 11162 51110 11172 51162
rect 11196 51110 11226 51162
rect 11226 51110 11252 51162
rect 10956 51108 11012 51110
rect 11036 51108 11092 51110
rect 11116 51108 11172 51110
rect 11196 51108 11252 51110
rect 10966 50904 11022 50960
rect 10966 50380 11022 50416
rect 10966 50360 10968 50380
rect 10968 50360 11020 50380
rect 11020 50360 11022 50380
rect 10956 50074 11012 50076
rect 11036 50074 11092 50076
rect 11116 50074 11172 50076
rect 11196 50074 11252 50076
rect 10956 50022 10982 50074
rect 10982 50022 11012 50074
rect 11036 50022 11046 50074
rect 11046 50022 11092 50074
rect 11116 50022 11162 50074
rect 11162 50022 11172 50074
rect 11196 50022 11226 50074
rect 11226 50022 11252 50074
rect 10956 50020 11012 50022
rect 11036 50020 11092 50022
rect 11116 50020 11172 50022
rect 11196 50020 11252 50022
rect 10966 49816 11022 49872
rect 10956 48986 11012 48988
rect 11036 48986 11092 48988
rect 11116 48986 11172 48988
rect 11196 48986 11252 48988
rect 10956 48934 10982 48986
rect 10982 48934 11012 48986
rect 11036 48934 11046 48986
rect 11046 48934 11092 48986
rect 11116 48934 11162 48986
rect 11162 48934 11172 48986
rect 11196 48934 11226 48986
rect 11226 48934 11252 48986
rect 10956 48932 11012 48934
rect 11036 48932 11092 48934
rect 11116 48932 11172 48934
rect 11196 48932 11252 48934
rect 10966 48728 11022 48784
rect 11242 48628 11244 48648
rect 11244 48628 11296 48648
rect 11296 48628 11298 48648
rect 11242 48592 11298 48628
rect 10956 47898 11012 47900
rect 11036 47898 11092 47900
rect 11116 47898 11172 47900
rect 11196 47898 11252 47900
rect 10956 47846 10982 47898
rect 10982 47846 11012 47898
rect 11036 47846 11046 47898
rect 11046 47846 11092 47898
rect 11116 47846 11162 47898
rect 11162 47846 11172 47898
rect 11196 47846 11226 47898
rect 11226 47846 11252 47898
rect 10956 47844 11012 47846
rect 11036 47844 11092 47846
rect 11116 47844 11172 47846
rect 11196 47844 11252 47846
rect 10966 47640 11022 47696
rect 10956 46810 11012 46812
rect 11036 46810 11092 46812
rect 11116 46810 11172 46812
rect 11196 46810 11252 46812
rect 10956 46758 10982 46810
rect 10982 46758 11012 46810
rect 11036 46758 11046 46810
rect 11046 46758 11092 46810
rect 11116 46758 11162 46810
rect 11162 46758 11172 46810
rect 11196 46758 11226 46810
rect 11226 46758 11252 46810
rect 10956 46756 11012 46758
rect 11036 46756 11092 46758
rect 11116 46756 11172 46758
rect 11196 46756 11252 46758
rect 10956 45722 11012 45724
rect 11036 45722 11092 45724
rect 11116 45722 11172 45724
rect 11196 45722 11252 45724
rect 10956 45670 10982 45722
rect 10982 45670 11012 45722
rect 11036 45670 11046 45722
rect 11046 45670 11092 45722
rect 11116 45670 11162 45722
rect 11162 45670 11172 45722
rect 11196 45670 11226 45722
rect 11226 45670 11252 45722
rect 10956 45668 11012 45670
rect 11036 45668 11092 45670
rect 11116 45668 11172 45670
rect 11196 45668 11252 45670
rect 10874 45464 10930 45520
rect 10956 44634 11012 44636
rect 11036 44634 11092 44636
rect 11116 44634 11172 44636
rect 11196 44634 11252 44636
rect 10956 44582 10982 44634
rect 10982 44582 11012 44634
rect 11036 44582 11046 44634
rect 11046 44582 11092 44634
rect 11116 44582 11162 44634
rect 11162 44582 11172 44634
rect 11196 44582 11226 44634
rect 11226 44582 11252 44634
rect 10956 44580 11012 44582
rect 11036 44580 11092 44582
rect 11116 44580 11172 44582
rect 11196 44580 11252 44582
rect 10874 44376 10930 44432
rect 10956 43546 11012 43548
rect 11036 43546 11092 43548
rect 11116 43546 11172 43548
rect 11196 43546 11252 43548
rect 10956 43494 10982 43546
rect 10982 43494 11012 43546
rect 11036 43494 11046 43546
rect 11046 43494 11092 43546
rect 11116 43494 11162 43546
rect 11162 43494 11172 43546
rect 11196 43494 11226 43546
rect 11226 43494 11252 43546
rect 10956 43492 11012 43494
rect 11036 43492 11092 43494
rect 11116 43492 11172 43494
rect 11196 43492 11252 43494
rect 10782 42628 10838 42664
rect 10782 42608 10784 42628
rect 10784 42608 10836 42628
rect 10836 42608 10838 42628
rect 10966 42744 11022 42800
rect 10956 42458 11012 42460
rect 11036 42458 11092 42460
rect 11116 42458 11172 42460
rect 11196 42458 11252 42460
rect 10956 42406 10982 42458
rect 10982 42406 11012 42458
rect 11036 42406 11046 42458
rect 11046 42406 11092 42458
rect 11116 42406 11162 42458
rect 11162 42406 11172 42458
rect 11196 42406 11226 42458
rect 11226 42406 11252 42458
rect 10956 42404 11012 42406
rect 11036 42404 11092 42406
rect 11116 42404 11172 42406
rect 11196 42404 11252 42406
rect 10956 41370 11012 41372
rect 11036 41370 11092 41372
rect 11116 41370 11172 41372
rect 11196 41370 11252 41372
rect 10956 41318 10982 41370
rect 10982 41318 11012 41370
rect 11036 41318 11046 41370
rect 11046 41318 11092 41370
rect 11116 41318 11162 41370
rect 11162 41318 11172 41370
rect 11196 41318 11226 41370
rect 11226 41318 11252 41370
rect 10956 41316 11012 41318
rect 11036 41316 11092 41318
rect 11116 41316 11172 41318
rect 11196 41316 11252 41318
rect 10506 38664 10562 38720
rect 10506 38392 10562 38448
rect 10230 32972 10286 33008
rect 10230 32952 10232 32972
rect 10232 32952 10284 32972
rect 10284 32952 10286 32972
rect 10230 32308 10232 32328
rect 10232 32308 10284 32328
rect 10284 32308 10286 32328
rect 10230 32272 10286 32308
rect 10230 32136 10286 32192
rect 10230 30776 10286 30832
rect 10506 36760 10562 36816
rect 10874 40588 10930 40624
rect 10874 40568 10876 40588
rect 10876 40568 10928 40588
rect 10928 40568 10930 40588
rect 10956 40282 11012 40284
rect 11036 40282 11092 40284
rect 11116 40282 11172 40284
rect 11196 40282 11252 40284
rect 10956 40230 10982 40282
rect 10982 40230 11012 40282
rect 11036 40230 11046 40282
rect 11046 40230 11092 40282
rect 11116 40230 11162 40282
rect 11162 40230 11172 40282
rect 11196 40230 11226 40282
rect 11226 40230 11252 40282
rect 10956 40228 11012 40230
rect 11036 40228 11092 40230
rect 11116 40228 11172 40230
rect 11196 40228 11252 40230
rect 10874 39788 10876 39808
rect 10876 39788 10928 39808
rect 10928 39788 10930 39808
rect 10874 39752 10930 39788
rect 10956 39194 11012 39196
rect 11036 39194 11092 39196
rect 11116 39194 11172 39196
rect 11196 39194 11252 39196
rect 10956 39142 10982 39194
rect 10982 39142 11012 39194
rect 11036 39142 11046 39194
rect 11046 39142 11092 39194
rect 11116 39142 11162 39194
rect 11162 39142 11172 39194
rect 11196 39142 11226 39194
rect 11226 39142 11252 39194
rect 10956 39140 11012 39142
rect 11036 39140 11092 39142
rect 11116 39140 11172 39142
rect 11196 39140 11252 39142
rect 11058 38664 11114 38720
rect 11242 38664 11298 38720
rect 10956 38106 11012 38108
rect 11036 38106 11092 38108
rect 11116 38106 11172 38108
rect 11196 38106 11252 38108
rect 10956 38054 10982 38106
rect 10982 38054 11012 38106
rect 11036 38054 11046 38106
rect 11046 38054 11092 38106
rect 11116 38054 11162 38106
rect 11162 38054 11172 38106
rect 11196 38054 11226 38106
rect 11226 38054 11252 38106
rect 10956 38052 11012 38054
rect 11036 38052 11092 38054
rect 11116 38052 11172 38054
rect 11196 38052 11252 38054
rect 11242 37848 11298 37904
rect 10506 33224 10562 33280
rect 11794 53116 11796 53136
rect 11796 53116 11848 53136
rect 11848 53116 11850 53136
rect 11794 53080 11850 53116
rect 11610 51584 11666 51640
rect 11886 52672 11942 52728
rect 11794 51040 11850 51096
rect 11794 50904 11850 50960
rect 11702 50496 11758 50552
rect 11610 50224 11666 50280
rect 11426 48320 11482 48376
rect 11610 47640 11666 47696
rect 12438 56924 12440 56944
rect 12440 56924 12492 56944
rect 12492 56924 12494 56944
rect 12438 56888 12494 56924
rect 13450 68176 13506 68232
rect 13082 63860 13084 63880
rect 13084 63860 13136 63880
rect 13136 63860 13138 63880
rect 13082 63824 13138 63860
rect 13082 63688 13138 63744
rect 12898 63144 12954 63200
rect 12898 61104 12954 61160
rect 12714 56480 12770 56536
rect 12530 55936 12586 55992
rect 12346 54168 12402 54224
rect 11978 51176 12034 51232
rect 11886 50360 11942 50416
rect 11886 48728 11942 48784
rect 11702 47096 11758 47152
rect 11610 46960 11666 47016
rect 11518 45464 11574 45520
rect 11610 42200 11666 42256
rect 11518 41384 11574 41440
rect 11794 45464 11850 45520
rect 11702 39924 11704 39944
rect 11704 39924 11756 39944
rect 11756 39924 11758 39944
rect 11702 39888 11758 39924
rect 11702 39616 11758 39672
rect 11518 39344 11574 39400
rect 10956 37018 11012 37020
rect 11036 37018 11092 37020
rect 11116 37018 11172 37020
rect 11196 37018 11252 37020
rect 10956 36966 10982 37018
rect 10982 36966 11012 37018
rect 11036 36966 11046 37018
rect 11046 36966 11092 37018
rect 11116 36966 11162 37018
rect 11162 36966 11172 37018
rect 11196 36966 11226 37018
rect 11226 36966 11252 37018
rect 10956 36964 11012 36966
rect 11036 36964 11092 36966
rect 11116 36964 11172 36966
rect 11196 36964 11252 36966
rect 10782 34448 10838 34504
rect 10690 31864 10746 31920
rect 10956 35930 11012 35932
rect 11036 35930 11092 35932
rect 11116 35930 11172 35932
rect 11196 35930 11252 35932
rect 10956 35878 10982 35930
rect 10982 35878 11012 35930
rect 11036 35878 11046 35930
rect 11046 35878 11092 35930
rect 11116 35878 11162 35930
rect 11162 35878 11172 35930
rect 11196 35878 11226 35930
rect 11226 35878 11252 35930
rect 10956 35876 11012 35878
rect 11036 35876 11092 35878
rect 11116 35876 11172 35878
rect 11196 35876 11252 35878
rect 10956 34842 11012 34844
rect 11036 34842 11092 34844
rect 11116 34842 11172 34844
rect 11196 34842 11252 34844
rect 10956 34790 10982 34842
rect 10982 34790 11012 34842
rect 11036 34790 11046 34842
rect 11046 34790 11092 34842
rect 11116 34790 11162 34842
rect 11162 34790 11172 34842
rect 11196 34790 11226 34842
rect 11226 34790 11252 34842
rect 10956 34788 11012 34790
rect 11036 34788 11092 34790
rect 11116 34788 11172 34790
rect 11196 34788 11252 34790
rect 11426 34040 11482 34096
rect 10956 33754 11012 33756
rect 11036 33754 11092 33756
rect 11116 33754 11172 33756
rect 11196 33754 11252 33756
rect 10956 33702 10982 33754
rect 10982 33702 11012 33754
rect 11036 33702 11046 33754
rect 11046 33702 11092 33754
rect 11116 33702 11162 33754
rect 11162 33702 11172 33754
rect 11196 33702 11226 33754
rect 11226 33702 11252 33754
rect 10956 33700 11012 33702
rect 11036 33700 11092 33702
rect 11116 33700 11172 33702
rect 11196 33700 11252 33702
rect 10956 32666 11012 32668
rect 11036 32666 11092 32668
rect 11116 32666 11172 32668
rect 11196 32666 11252 32668
rect 10956 32614 10982 32666
rect 10982 32614 11012 32666
rect 11036 32614 11046 32666
rect 11046 32614 11092 32666
rect 11116 32614 11162 32666
rect 11162 32614 11172 32666
rect 11196 32614 11226 32666
rect 11226 32614 11252 32666
rect 10956 32612 11012 32614
rect 11036 32612 11092 32614
rect 11116 32612 11172 32614
rect 11196 32612 11252 32614
rect 11334 31728 11390 31784
rect 10956 31578 11012 31580
rect 11036 31578 11092 31580
rect 11116 31578 11172 31580
rect 11196 31578 11252 31580
rect 10956 31526 10982 31578
rect 10982 31526 11012 31578
rect 11036 31526 11046 31578
rect 11046 31526 11092 31578
rect 11116 31526 11162 31578
rect 11162 31526 11172 31578
rect 11196 31526 11226 31578
rect 11226 31526 11252 31578
rect 10956 31524 11012 31526
rect 11036 31524 11092 31526
rect 11116 31524 11172 31526
rect 11196 31524 11252 31526
rect 10782 31340 10838 31376
rect 10782 31320 10784 31340
rect 10784 31320 10836 31340
rect 10836 31320 10838 31340
rect 10598 30776 10654 30832
rect 10506 30232 10562 30288
rect 10506 26968 10562 27024
rect 10046 24268 10102 24304
rect 10046 24248 10048 24268
rect 10048 24248 10100 24268
rect 10100 24248 10102 24268
rect 10690 30504 10746 30560
rect 11334 30812 11336 30832
rect 11336 30812 11388 30832
rect 11388 30812 11390 30832
rect 11334 30776 11390 30812
rect 10956 30490 11012 30492
rect 11036 30490 11092 30492
rect 11116 30490 11172 30492
rect 11196 30490 11252 30492
rect 10956 30438 10982 30490
rect 10982 30438 11012 30490
rect 11036 30438 11046 30490
rect 11046 30438 11092 30490
rect 11116 30438 11162 30490
rect 11162 30438 11172 30490
rect 11196 30438 11226 30490
rect 11226 30438 11252 30490
rect 10956 30436 11012 30438
rect 11036 30436 11092 30438
rect 11116 30436 11172 30438
rect 11196 30436 11252 30438
rect 10966 29708 11022 29744
rect 10966 29688 10968 29708
rect 10968 29688 11020 29708
rect 11020 29688 11022 29708
rect 10956 29402 11012 29404
rect 11036 29402 11092 29404
rect 11116 29402 11172 29404
rect 11196 29402 11252 29404
rect 10956 29350 10982 29402
rect 10982 29350 11012 29402
rect 11036 29350 11046 29402
rect 11046 29350 11092 29402
rect 11116 29350 11162 29402
rect 11162 29350 11172 29402
rect 11196 29350 11226 29402
rect 11226 29350 11252 29402
rect 10956 29348 11012 29350
rect 11036 29348 11092 29350
rect 11116 29348 11172 29350
rect 11196 29348 11252 29350
rect 10956 28314 11012 28316
rect 11036 28314 11092 28316
rect 11116 28314 11172 28316
rect 11196 28314 11252 28316
rect 10956 28262 10982 28314
rect 10982 28262 11012 28314
rect 11036 28262 11046 28314
rect 11046 28262 11092 28314
rect 11116 28262 11162 28314
rect 11162 28262 11172 28314
rect 11196 28262 11226 28314
rect 11226 28262 11252 28314
rect 10956 28260 11012 28262
rect 11036 28260 11092 28262
rect 11116 28260 11172 28262
rect 11196 28260 11252 28262
rect 10956 27226 11012 27228
rect 11036 27226 11092 27228
rect 11116 27226 11172 27228
rect 11196 27226 11252 27228
rect 10956 27174 10982 27226
rect 10982 27174 11012 27226
rect 11036 27174 11046 27226
rect 11046 27174 11092 27226
rect 11116 27174 11162 27226
rect 11162 27174 11172 27226
rect 11196 27174 11226 27226
rect 11226 27174 11252 27226
rect 10956 27172 11012 27174
rect 11036 27172 11092 27174
rect 11116 27172 11172 27174
rect 11196 27172 11252 27174
rect 11518 33088 11574 33144
rect 11518 31184 11574 31240
rect 12070 48048 12126 48104
rect 12254 50088 12310 50144
rect 12622 54068 12624 54088
rect 12624 54068 12676 54088
rect 12676 54068 12678 54088
rect 12622 54032 12678 54068
rect 13910 68076 13912 68096
rect 13912 68076 13964 68096
rect 13964 68076 13966 68096
rect 13910 68040 13966 68076
rect 14289 68026 14345 68028
rect 14369 68026 14425 68028
rect 14449 68026 14505 68028
rect 14529 68026 14585 68028
rect 14289 67974 14315 68026
rect 14315 67974 14345 68026
rect 14369 67974 14379 68026
rect 14379 67974 14425 68026
rect 14449 67974 14495 68026
rect 14495 67974 14505 68026
rect 14529 67974 14559 68026
rect 14559 67974 14585 68026
rect 14289 67972 14345 67974
rect 14369 67972 14425 67974
rect 14449 67972 14505 67974
rect 14529 67972 14585 67974
rect 14094 67768 14150 67824
rect 13910 65864 13966 65920
rect 13450 64368 13506 64424
rect 13450 63688 13506 63744
rect 13266 60832 13322 60888
rect 12990 57296 13046 57352
rect 12898 52944 12954 53000
rect 12898 52672 12954 52728
rect 12898 51484 12900 51504
rect 12900 51484 12952 51504
rect 12952 51484 12954 51504
rect 12898 51448 12954 51484
rect 12990 50904 13046 50960
rect 12898 49544 12954 49600
rect 12622 48728 12678 48784
rect 12346 47368 12402 47424
rect 12346 47232 12402 47288
rect 12622 48456 12678 48512
rect 12714 47776 12770 47832
rect 12070 44648 12126 44704
rect 12070 44376 12126 44432
rect 11978 38836 11980 38856
rect 11980 38836 12032 38856
rect 12032 38836 12034 38856
rect 11978 38800 12034 38836
rect 11978 38120 12034 38176
rect 12254 41112 12310 41168
rect 11978 31864 12034 31920
rect 11886 31728 11942 31784
rect 11886 30232 11942 30288
rect 11518 28872 11574 28928
rect 11518 27920 11574 27976
rect 12806 47504 12862 47560
rect 14370 67260 14372 67280
rect 14372 67260 14424 67280
rect 14424 67260 14426 67280
rect 14370 67224 14426 67260
rect 14289 66938 14345 66940
rect 14369 66938 14425 66940
rect 14449 66938 14505 66940
rect 14529 66938 14585 66940
rect 14289 66886 14315 66938
rect 14315 66886 14345 66938
rect 14369 66886 14379 66938
rect 14379 66886 14425 66938
rect 14449 66886 14495 66938
rect 14495 66886 14505 66938
rect 14529 66886 14559 66938
rect 14559 66886 14585 66938
rect 14289 66884 14345 66886
rect 14369 66884 14425 66886
rect 14449 66884 14505 66886
rect 14529 66884 14585 66886
rect 14738 65900 14740 65920
rect 14740 65900 14792 65920
rect 14792 65900 14794 65920
rect 14738 65864 14794 65900
rect 14289 65850 14345 65852
rect 14369 65850 14425 65852
rect 14449 65850 14505 65852
rect 14529 65850 14585 65852
rect 14289 65798 14315 65850
rect 14315 65798 14345 65850
rect 14369 65798 14379 65850
rect 14379 65798 14425 65850
rect 14449 65798 14495 65850
rect 14495 65798 14505 65850
rect 14529 65798 14559 65850
rect 14559 65798 14585 65850
rect 14289 65796 14345 65798
rect 14369 65796 14425 65798
rect 14449 65796 14505 65798
rect 14529 65796 14585 65798
rect 14289 64762 14345 64764
rect 14369 64762 14425 64764
rect 14449 64762 14505 64764
rect 14529 64762 14585 64764
rect 14289 64710 14315 64762
rect 14315 64710 14345 64762
rect 14369 64710 14379 64762
rect 14379 64710 14425 64762
rect 14449 64710 14495 64762
rect 14495 64710 14505 64762
rect 14529 64710 14559 64762
rect 14559 64710 14585 64762
rect 14289 64708 14345 64710
rect 14369 64708 14425 64710
rect 14449 64708 14505 64710
rect 14529 64708 14585 64710
rect 14370 64504 14426 64560
rect 14289 63674 14345 63676
rect 14369 63674 14425 63676
rect 14449 63674 14505 63676
rect 14529 63674 14585 63676
rect 14289 63622 14315 63674
rect 14315 63622 14345 63674
rect 14369 63622 14379 63674
rect 14379 63622 14425 63674
rect 14449 63622 14495 63674
rect 14495 63622 14505 63674
rect 14529 63622 14559 63674
rect 14559 63622 14585 63674
rect 14289 63620 14345 63622
rect 14369 63620 14425 63622
rect 14449 63620 14505 63622
rect 14529 63620 14585 63622
rect 14289 62586 14345 62588
rect 14369 62586 14425 62588
rect 14449 62586 14505 62588
rect 14529 62586 14585 62588
rect 14289 62534 14315 62586
rect 14315 62534 14345 62586
rect 14369 62534 14379 62586
rect 14379 62534 14425 62586
rect 14449 62534 14495 62586
rect 14495 62534 14505 62586
rect 14529 62534 14559 62586
rect 14559 62534 14585 62586
rect 14289 62532 14345 62534
rect 14369 62532 14425 62534
rect 14449 62532 14505 62534
rect 14529 62532 14585 62534
rect 14289 61498 14345 61500
rect 14369 61498 14425 61500
rect 14449 61498 14505 61500
rect 14529 61498 14585 61500
rect 14289 61446 14315 61498
rect 14315 61446 14345 61498
rect 14369 61446 14379 61498
rect 14379 61446 14425 61498
rect 14449 61446 14495 61498
rect 14495 61446 14505 61498
rect 14529 61446 14559 61498
rect 14559 61446 14585 61498
rect 14289 61444 14345 61446
rect 14369 61444 14425 61446
rect 14449 61444 14505 61446
rect 14529 61444 14585 61446
rect 14738 60968 14794 61024
rect 14094 60696 14150 60752
rect 14738 60696 14794 60752
rect 14289 60410 14345 60412
rect 14369 60410 14425 60412
rect 14449 60410 14505 60412
rect 14529 60410 14585 60412
rect 14289 60358 14315 60410
rect 14315 60358 14345 60410
rect 14369 60358 14379 60410
rect 14379 60358 14425 60410
rect 14449 60358 14495 60410
rect 14495 60358 14505 60410
rect 14529 60358 14559 60410
rect 14559 60358 14585 60410
rect 14289 60356 14345 60358
rect 14369 60356 14425 60358
rect 14449 60356 14505 60358
rect 14529 60356 14585 60358
rect 14738 60308 14794 60344
rect 14738 60288 14740 60308
rect 14740 60288 14792 60308
rect 14792 60288 14794 60308
rect 14186 60152 14242 60208
rect 14094 60016 14150 60072
rect 14002 59472 14058 59528
rect 13358 51040 13414 51096
rect 13450 50904 13506 50960
rect 13358 50768 13414 50824
rect 13174 50224 13230 50280
rect 13358 49816 13414 49872
rect 13266 48084 13268 48104
rect 13268 48084 13320 48104
rect 13320 48084 13322 48104
rect 13266 48048 13322 48084
rect 13174 46824 13230 46880
rect 13266 46552 13322 46608
rect 12530 43288 12586 43344
rect 12346 40432 12402 40488
rect 12346 38256 12402 38312
rect 13266 46008 13322 46064
rect 13174 42608 13230 42664
rect 12990 42220 13046 42256
rect 12990 42200 12992 42220
rect 12992 42200 13044 42220
rect 13044 42200 13046 42220
rect 13174 41556 13176 41576
rect 13176 41556 13228 41576
rect 13228 41556 13230 41576
rect 13174 41520 13230 41556
rect 13082 39788 13084 39808
rect 13084 39788 13136 39808
rect 13136 39788 13138 39808
rect 13082 39752 13138 39788
rect 12714 38120 12770 38176
rect 12898 37304 12954 37360
rect 13082 36236 13138 36272
rect 13082 36216 13084 36236
rect 13084 36216 13136 36236
rect 13136 36216 13138 36236
rect 12806 33496 12862 33552
rect 12622 33224 12678 33280
rect 12162 28464 12218 28520
rect 11978 28056 12034 28112
rect 11150 26308 11206 26344
rect 11150 26288 11152 26308
rect 11152 26288 11204 26308
rect 11204 26288 11206 26308
rect 10956 26138 11012 26140
rect 11036 26138 11092 26140
rect 11116 26138 11172 26140
rect 11196 26138 11252 26140
rect 10956 26086 10982 26138
rect 10982 26086 11012 26138
rect 11036 26086 11046 26138
rect 11046 26086 11092 26138
rect 11116 26086 11162 26138
rect 11162 26086 11172 26138
rect 11196 26086 11226 26138
rect 11226 26086 11252 26138
rect 10956 26084 11012 26086
rect 11036 26084 11092 26086
rect 11116 26084 11172 26086
rect 11196 26084 11252 26086
rect 10956 25050 11012 25052
rect 11036 25050 11092 25052
rect 11116 25050 11172 25052
rect 11196 25050 11252 25052
rect 10956 24998 10982 25050
rect 10982 24998 11012 25050
rect 11036 24998 11046 25050
rect 11046 24998 11092 25050
rect 11116 24998 11162 25050
rect 11162 24998 11172 25050
rect 11196 24998 11226 25050
rect 11226 24998 11252 25050
rect 10956 24996 11012 24998
rect 11036 24996 11092 24998
rect 11116 24996 11172 24998
rect 11196 24996 11252 24998
rect 11426 24928 11482 24984
rect 10956 23962 11012 23964
rect 11036 23962 11092 23964
rect 11116 23962 11172 23964
rect 11196 23962 11252 23964
rect 10956 23910 10982 23962
rect 10982 23910 11012 23962
rect 11036 23910 11046 23962
rect 11046 23910 11092 23962
rect 11116 23910 11162 23962
rect 11162 23910 11172 23962
rect 11196 23910 11226 23962
rect 11226 23910 11252 23962
rect 10956 23908 11012 23910
rect 11036 23908 11092 23910
rect 11116 23908 11172 23910
rect 11196 23908 11252 23910
rect 10230 22888 10286 22944
rect 10956 22874 11012 22876
rect 11036 22874 11092 22876
rect 11116 22874 11172 22876
rect 11196 22874 11252 22876
rect 10956 22822 10982 22874
rect 10982 22822 11012 22874
rect 11036 22822 11046 22874
rect 11046 22822 11092 22874
rect 11116 22822 11162 22874
rect 11162 22822 11172 22874
rect 11196 22822 11226 22874
rect 11226 22822 11252 22874
rect 10956 22820 11012 22822
rect 11036 22820 11092 22822
rect 11116 22820 11172 22822
rect 11196 22820 11252 22822
rect 9678 22108 9680 22128
rect 9680 22108 9732 22128
rect 9732 22108 9734 22128
rect 9678 22072 9734 22108
rect 9862 22208 9918 22264
rect 9770 19488 9826 19544
rect 9770 16904 9826 16960
rect 10506 22072 10562 22128
rect 11426 22616 11482 22672
rect 10956 21786 11012 21788
rect 11036 21786 11092 21788
rect 11116 21786 11172 21788
rect 11196 21786 11252 21788
rect 10956 21734 10982 21786
rect 10982 21734 11012 21786
rect 11036 21734 11046 21786
rect 11046 21734 11092 21786
rect 11116 21734 11162 21786
rect 11162 21734 11172 21786
rect 11196 21734 11226 21786
rect 11226 21734 11252 21786
rect 10956 21732 11012 21734
rect 11036 21732 11092 21734
rect 11116 21732 11172 21734
rect 11196 21732 11252 21734
rect 10956 20698 11012 20700
rect 11036 20698 11092 20700
rect 11116 20698 11172 20700
rect 11196 20698 11252 20700
rect 10956 20646 10982 20698
rect 10982 20646 11012 20698
rect 11036 20646 11046 20698
rect 11046 20646 11092 20698
rect 11116 20646 11162 20698
rect 11162 20646 11172 20698
rect 11196 20646 11226 20698
rect 11226 20646 11252 20698
rect 10956 20644 11012 20646
rect 11036 20644 11092 20646
rect 11116 20644 11172 20646
rect 11196 20644 11252 20646
rect 10956 19610 11012 19612
rect 11036 19610 11092 19612
rect 11116 19610 11172 19612
rect 11196 19610 11252 19612
rect 10956 19558 10982 19610
rect 10982 19558 11012 19610
rect 11036 19558 11046 19610
rect 11046 19558 11092 19610
rect 11116 19558 11162 19610
rect 11162 19558 11172 19610
rect 11196 19558 11226 19610
rect 11226 19558 11252 19610
rect 10956 19556 11012 19558
rect 11036 19556 11092 19558
rect 11116 19556 11172 19558
rect 11196 19556 11252 19558
rect 9678 16652 9734 16688
rect 9678 16632 9680 16652
rect 9680 16632 9732 16652
rect 9732 16632 9734 16652
rect 10782 18828 10838 18864
rect 10782 18808 10784 18828
rect 10784 18808 10836 18828
rect 10836 18808 10838 18828
rect 11242 18808 11298 18864
rect 10956 18522 11012 18524
rect 11036 18522 11092 18524
rect 11116 18522 11172 18524
rect 11196 18522 11252 18524
rect 10956 18470 10982 18522
rect 10982 18470 11012 18522
rect 11036 18470 11046 18522
rect 11046 18470 11092 18522
rect 11116 18470 11162 18522
rect 11162 18470 11172 18522
rect 11196 18470 11226 18522
rect 11226 18470 11252 18522
rect 10956 18468 11012 18470
rect 11036 18468 11092 18470
rect 11116 18468 11172 18470
rect 11196 18468 11252 18470
rect 10956 17434 11012 17436
rect 11036 17434 11092 17436
rect 11116 17434 11172 17436
rect 11196 17434 11252 17436
rect 10956 17382 10982 17434
rect 10982 17382 11012 17434
rect 11036 17382 11046 17434
rect 11046 17382 11092 17434
rect 11116 17382 11162 17434
rect 11162 17382 11172 17434
rect 11196 17382 11226 17434
rect 11226 17382 11252 17434
rect 10956 17380 11012 17382
rect 11036 17380 11092 17382
rect 11116 17380 11172 17382
rect 11196 17380 11252 17382
rect 11334 16632 11390 16688
rect 10956 16346 11012 16348
rect 11036 16346 11092 16348
rect 11116 16346 11172 16348
rect 11196 16346 11252 16348
rect 10956 16294 10982 16346
rect 10982 16294 11012 16346
rect 11036 16294 11046 16346
rect 11046 16294 11092 16346
rect 11116 16294 11162 16346
rect 11162 16294 11172 16346
rect 11196 16294 11226 16346
rect 11226 16294 11252 16346
rect 10956 16292 11012 16294
rect 11036 16292 11092 16294
rect 11116 16292 11172 16294
rect 11196 16292 11252 16294
rect 12070 25780 12072 25800
rect 12072 25780 12124 25800
rect 12124 25780 12126 25800
rect 12070 25744 12126 25780
rect 12162 25644 12164 25664
rect 12164 25644 12216 25664
rect 12216 25644 12218 25664
rect 12162 25608 12218 25644
rect 11978 25200 12034 25256
rect 11978 23704 12034 23760
rect 10956 15258 11012 15260
rect 11036 15258 11092 15260
rect 11116 15258 11172 15260
rect 11196 15258 11252 15260
rect 10956 15206 10982 15258
rect 10982 15206 11012 15258
rect 11036 15206 11046 15258
rect 11046 15206 11092 15258
rect 11116 15206 11162 15258
rect 11162 15206 11172 15258
rect 11196 15206 11226 15258
rect 11226 15206 11252 15258
rect 10956 15204 11012 15206
rect 11036 15204 11092 15206
rect 11116 15204 11172 15206
rect 11196 15204 11252 15206
rect 9862 14456 9918 14512
rect 9770 13132 9772 13152
rect 9772 13132 9824 13152
rect 9824 13132 9826 13152
rect 9770 13096 9826 13132
rect 10322 13232 10378 13288
rect 10230 12960 10286 13016
rect 9586 11600 9642 11656
rect 10956 14170 11012 14172
rect 11036 14170 11092 14172
rect 11116 14170 11172 14172
rect 11196 14170 11252 14172
rect 10956 14118 10982 14170
rect 10982 14118 11012 14170
rect 11036 14118 11046 14170
rect 11046 14118 11092 14170
rect 11116 14118 11162 14170
rect 11162 14118 11172 14170
rect 11196 14118 11226 14170
rect 11226 14118 11252 14170
rect 10956 14116 11012 14118
rect 11036 14116 11092 14118
rect 11116 14116 11172 14118
rect 11196 14116 11252 14118
rect 10956 13082 11012 13084
rect 11036 13082 11092 13084
rect 11116 13082 11172 13084
rect 11196 13082 11252 13084
rect 10956 13030 10982 13082
rect 10982 13030 11012 13082
rect 11036 13030 11046 13082
rect 11046 13030 11092 13082
rect 11116 13030 11162 13082
rect 11162 13030 11172 13082
rect 11196 13030 11226 13082
rect 11226 13030 11252 13082
rect 10956 13028 11012 13030
rect 11036 13028 11092 13030
rect 11116 13028 11172 13030
rect 11196 13028 11252 13030
rect 11794 19116 11796 19136
rect 11796 19116 11848 19136
rect 11848 19116 11850 19136
rect 11794 19080 11850 19116
rect 10956 11994 11012 11996
rect 11036 11994 11092 11996
rect 11116 11994 11172 11996
rect 11196 11994 11252 11996
rect 10956 11942 10982 11994
rect 10982 11942 11012 11994
rect 11036 11942 11046 11994
rect 11046 11942 11092 11994
rect 11116 11942 11162 11994
rect 11162 11942 11172 11994
rect 11196 11942 11226 11994
rect 11226 11942 11252 11994
rect 10956 11940 11012 11942
rect 11036 11940 11092 11942
rect 11116 11940 11172 11942
rect 11196 11940 11252 11942
rect 11794 17584 11850 17640
rect 11058 11328 11114 11384
rect 12162 19352 12218 19408
rect 12070 18400 12126 18456
rect 13542 50088 13598 50144
rect 13726 56752 13782 56808
rect 13726 56228 13782 56264
rect 13726 56208 13728 56228
rect 13728 56208 13780 56228
rect 13780 56208 13782 56228
rect 13726 55392 13782 55448
rect 14094 57976 14150 58032
rect 15198 63280 15254 63336
rect 15198 62328 15254 62384
rect 15382 63824 15438 63880
rect 15382 62464 15438 62520
rect 14922 60968 14978 61024
rect 14289 59322 14345 59324
rect 14369 59322 14425 59324
rect 14449 59322 14505 59324
rect 14529 59322 14585 59324
rect 14289 59270 14315 59322
rect 14315 59270 14345 59322
rect 14369 59270 14379 59322
rect 14379 59270 14425 59322
rect 14449 59270 14495 59322
rect 14495 59270 14505 59322
rect 14529 59270 14559 59322
rect 14559 59270 14585 59322
rect 14289 59268 14345 59270
rect 14369 59268 14425 59270
rect 14449 59268 14505 59270
rect 14529 59268 14585 59270
rect 14830 59064 14886 59120
rect 14289 58234 14345 58236
rect 14369 58234 14425 58236
rect 14449 58234 14505 58236
rect 14529 58234 14585 58236
rect 14289 58182 14315 58234
rect 14315 58182 14345 58234
rect 14369 58182 14379 58234
rect 14379 58182 14425 58234
rect 14449 58182 14495 58234
rect 14495 58182 14505 58234
rect 14529 58182 14559 58234
rect 14559 58182 14585 58234
rect 14289 58180 14345 58182
rect 14369 58180 14425 58182
rect 14449 58180 14505 58182
rect 14529 58180 14585 58182
rect 14830 57976 14886 58032
rect 14289 57146 14345 57148
rect 14369 57146 14425 57148
rect 14449 57146 14505 57148
rect 14529 57146 14585 57148
rect 14289 57094 14315 57146
rect 14315 57094 14345 57146
rect 14369 57094 14379 57146
rect 14379 57094 14425 57146
rect 14449 57094 14495 57146
rect 14495 57094 14505 57146
rect 14529 57094 14559 57146
rect 14559 57094 14585 57146
rect 14289 57092 14345 57094
rect 14369 57092 14425 57094
rect 14449 57092 14505 57094
rect 14529 57092 14585 57094
rect 14289 56058 14345 56060
rect 14369 56058 14425 56060
rect 14449 56058 14505 56060
rect 14529 56058 14585 56060
rect 14289 56006 14315 56058
rect 14315 56006 14345 56058
rect 14369 56006 14379 56058
rect 14379 56006 14425 56058
rect 14449 56006 14495 56058
rect 14495 56006 14505 56058
rect 14529 56006 14559 56058
rect 14559 56006 14585 56058
rect 14289 56004 14345 56006
rect 14369 56004 14425 56006
rect 14449 56004 14505 56006
rect 14529 56004 14585 56006
rect 14370 55392 14426 55448
rect 14186 55292 14188 55312
rect 14188 55292 14240 55312
rect 14240 55292 14242 55312
rect 14186 55256 14242 55292
rect 14289 54970 14345 54972
rect 14369 54970 14425 54972
rect 14449 54970 14505 54972
rect 14529 54970 14585 54972
rect 14289 54918 14315 54970
rect 14315 54918 14345 54970
rect 14369 54918 14379 54970
rect 14379 54918 14425 54970
rect 14449 54918 14495 54970
rect 14495 54918 14505 54970
rect 14529 54918 14559 54970
rect 14559 54918 14585 54970
rect 14289 54916 14345 54918
rect 14369 54916 14425 54918
rect 14449 54916 14505 54918
rect 14529 54916 14585 54918
rect 14646 54712 14702 54768
rect 13910 52400 13966 52456
rect 14289 53882 14345 53884
rect 14369 53882 14425 53884
rect 14449 53882 14505 53884
rect 14529 53882 14585 53884
rect 14289 53830 14315 53882
rect 14315 53830 14345 53882
rect 14369 53830 14379 53882
rect 14379 53830 14425 53882
rect 14449 53830 14495 53882
rect 14495 53830 14505 53882
rect 14529 53830 14559 53882
rect 14559 53830 14585 53882
rect 14289 53828 14345 53830
rect 14369 53828 14425 53830
rect 14449 53828 14505 53830
rect 14529 53828 14585 53830
rect 14738 53624 14794 53680
rect 13726 51992 13782 52048
rect 13726 51876 13782 51912
rect 13726 51856 13728 51876
rect 13728 51856 13780 51876
rect 13780 51856 13782 51876
rect 13726 50904 13782 50960
rect 13726 49136 13782 49192
rect 13542 48728 13598 48784
rect 13634 47096 13690 47152
rect 13542 46824 13598 46880
rect 13542 46416 13598 46472
rect 13542 45328 13598 45384
rect 13542 44376 13598 44432
rect 14002 50224 14058 50280
rect 13818 43968 13874 44024
rect 13818 43288 13874 43344
rect 13358 38120 13414 38176
rect 13818 40588 13874 40624
rect 13818 40568 13820 40588
rect 13820 40568 13872 40588
rect 13872 40568 13874 40588
rect 13726 38548 13782 38584
rect 13726 38528 13728 38548
rect 13728 38528 13780 38548
rect 13780 38528 13782 38548
rect 13174 31728 13230 31784
rect 12530 21528 12586 21584
rect 12898 23604 12900 23624
rect 12900 23604 12952 23624
rect 12952 23604 12954 23624
rect 12898 23568 12954 23604
rect 12898 23180 12954 23216
rect 12898 23160 12900 23180
rect 12900 23160 12952 23180
rect 12952 23160 12954 23180
rect 12622 19352 12678 19408
rect 10956 10906 11012 10908
rect 11036 10906 11092 10908
rect 11116 10906 11172 10908
rect 11196 10906 11252 10908
rect 10956 10854 10982 10906
rect 10982 10854 11012 10906
rect 11036 10854 11046 10906
rect 11046 10854 11092 10906
rect 11116 10854 11162 10906
rect 11162 10854 11172 10906
rect 11196 10854 11226 10906
rect 11226 10854 11252 10906
rect 10956 10852 11012 10854
rect 11036 10852 11092 10854
rect 11116 10852 11172 10854
rect 11196 10852 11252 10854
rect 10138 10240 10194 10296
rect 9770 9036 9826 9072
rect 9770 9016 9772 9036
rect 9772 9016 9824 9036
rect 9824 9016 9826 9036
rect 9678 7248 9734 7304
rect 10598 8880 10654 8936
rect 10506 8472 10562 8528
rect 10138 7928 10194 7984
rect 10782 10376 10838 10432
rect 10956 9818 11012 9820
rect 11036 9818 11092 9820
rect 11116 9818 11172 9820
rect 11196 9818 11252 9820
rect 10956 9766 10982 9818
rect 10982 9766 11012 9818
rect 11036 9766 11046 9818
rect 11046 9766 11092 9818
rect 11116 9766 11162 9818
rect 11162 9766 11172 9818
rect 11196 9766 11226 9818
rect 11226 9766 11252 9818
rect 10956 9764 11012 9766
rect 11036 9764 11092 9766
rect 11116 9764 11172 9766
rect 11196 9764 11252 9766
rect 11610 10648 11666 10704
rect 11150 9560 11206 9616
rect 10956 8730 11012 8732
rect 11036 8730 11092 8732
rect 11116 8730 11172 8732
rect 11196 8730 11252 8732
rect 10956 8678 10982 8730
rect 10982 8678 11012 8730
rect 11036 8678 11046 8730
rect 11046 8678 11092 8730
rect 11116 8678 11162 8730
rect 11162 8678 11172 8730
rect 11196 8678 11226 8730
rect 11226 8678 11252 8730
rect 10956 8676 11012 8678
rect 11036 8676 11092 8678
rect 11116 8676 11172 8678
rect 11196 8676 11252 8678
rect 11518 9288 11574 9344
rect 10874 8336 10930 8392
rect 10956 7642 11012 7644
rect 11036 7642 11092 7644
rect 11116 7642 11172 7644
rect 11196 7642 11252 7644
rect 10956 7590 10982 7642
rect 10982 7590 11012 7642
rect 11036 7590 11046 7642
rect 11046 7590 11092 7642
rect 11116 7590 11162 7642
rect 11162 7590 11172 7642
rect 11196 7590 11226 7642
rect 11226 7590 11252 7642
rect 10956 7588 11012 7590
rect 11036 7588 11092 7590
rect 11116 7588 11172 7590
rect 11196 7588 11252 7590
rect 11794 10648 11850 10704
rect 11702 9288 11758 9344
rect 11610 7928 11666 7984
rect 10956 6554 11012 6556
rect 11036 6554 11092 6556
rect 11116 6554 11172 6556
rect 11196 6554 11252 6556
rect 10956 6502 10982 6554
rect 10982 6502 11012 6554
rect 11036 6502 11046 6554
rect 11046 6502 11092 6554
rect 11116 6502 11162 6554
rect 11162 6502 11172 6554
rect 11196 6502 11226 6554
rect 11226 6502 11252 6554
rect 10956 6500 11012 6502
rect 11036 6500 11092 6502
rect 11116 6500 11172 6502
rect 11196 6500 11252 6502
rect 11978 8472 12034 8528
rect 12530 16088 12586 16144
rect 12346 13776 12402 13832
rect 12254 12316 12256 12336
rect 12256 12316 12308 12336
rect 12308 12316 12310 12336
rect 12254 12280 12310 12316
rect 12254 11600 12310 11656
rect 12254 10512 12310 10568
rect 12438 9288 12494 9344
rect 11886 7792 11942 7848
rect 11794 6160 11850 6216
rect 11426 5652 11428 5672
rect 11428 5652 11480 5672
rect 11480 5652 11482 5672
rect 11426 5616 11482 5652
rect 10956 5466 11012 5468
rect 11036 5466 11092 5468
rect 11116 5466 11172 5468
rect 11196 5466 11252 5468
rect 10956 5414 10982 5466
rect 10982 5414 11012 5466
rect 11036 5414 11046 5466
rect 11046 5414 11092 5466
rect 11116 5414 11162 5466
rect 11162 5414 11172 5466
rect 11196 5414 11226 5466
rect 11226 5414 11252 5466
rect 10956 5412 11012 5414
rect 11036 5412 11092 5414
rect 11116 5412 11172 5414
rect 11196 5412 11252 5414
rect 9862 4664 9918 4720
rect 10046 4664 10102 4720
rect 10956 4378 11012 4380
rect 11036 4378 11092 4380
rect 11116 4378 11172 4380
rect 11196 4378 11252 4380
rect 10956 4326 10982 4378
rect 10982 4326 11012 4378
rect 11036 4326 11046 4378
rect 11046 4326 11092 4378
rect 11116 4326 11162 4378
rect 11162 4326 11172 4378
rect 11196 4326 11226 4378
rect 11226 4326 11252 4378
rect 10956 4324 11012 4326
rect 11036 4324 11092 4326
rect 11116 4324 11172 4326
rect 11196 4324 11252 4326
rect 10956 3290 11012 3292
rect 11036 3290 11092 3292
rect 11116 3290 11172 3292
rect 11196 3290 11252 3292
rect 10956 3238 10982 3290
rect 10982 3238 11012 3290
rect 11036 3238 11046 3290
rect 11046 3238 11092 3290
rect 11116 3238 11162 3290
rect 11162 3238 11172 3290
rect 11196 3238 11226 3290
rect 11226 3238 11252 3290
rect 10956 3236 11012 3238
rect 11036 3236 11092 3238
rect 11116 3236 11172 3238
rect 11196 3236 11252 3238
rect 10046 2488 10102 2544
rect 13634 33904 13690 33960
rect 14094 49952 14150 50008
rect 14289 52794 14345 52796
rect 14369 52794 14425 52796
rect 14449 52794 14505 52796
rect 14529 52794 14585 52796
rect 14289 52742 14315 52794
rect 14315 52742 14345 52794
rect 14369 52742 14379 52794
rect 14379 52742 14425 52794
rect 14449 52742 14495 52794
rect 14495 52742 14505 52794
rect 14529 52742 14559 52794
rect 14559 52742 14585 52794
rect 14289 52740 14345 52742
rect 14369 52740 14425 52742
rect 14449 52740 14505 52742
rect 14529 52740 14585 52742
rect 14289 51706 14345 51708
rect 14369 51706 14425 51708
rect 14449 51706 14505 51708
rect 14529 51706 14585 51708
rect 14289 51654 14315 51706
rect 14315 51654 14345 51706
rect 14369 51654 14379 51706
rect 14379 51654 14425 51706
rect 14449 51654 14495 51706
rect 14495 51654 14505 51706
rect 14529 51654 14559 51706
rect 14559 51654 14585 51706
rect 14289 51652 14345 51654
rect 14369 51652 14425 51654
rect 14449 51652 14505 51654
rect 14529 51652 14585 51654
rect 14289 50618 14345 50620
rect 14369 50618 14425 50620
rect 14449 50618 14505 50620
rect 14529 50618 14585 50620
rect 14289 50566 14315 50618
rect 14315 50566 14345 50618
rect 14369 50566 14379 50618
rect 14379 50566 14425 50618
rect 14449 50566 14495 50618
rect 14495 50566 14505 50618
rect 14529 50566 14559 50618
rect 14559 50566 14585 50618
rect 14289 50564 14345 50566
rect 14369 50564 14425 50566
rect 14449 50564 14505 50566
rect 14529 50564 14585 50566
rect 14289 49530 14345 49532
rect 14369 49530 14425 49532
rect 14449 49530 14505 49532
rect 14529 49530 14585 49532
rect 14289 49478 14315 49530
rect 14315 49478 14345 49530
rect 14369 49478 14379 49530
rect 14379 49478 14425 49530
rect 14449 49478 14495 49530
rect 14495 49478 14505 49530
rect 14529 49478 14559 49530
rect 14559 49478 14585 49530
rect 14289 49476 14345 49478
rect 14369 49476 14425 49478
rect 14449 49476 14505 49478
rect 14529 49476 14585 49478
rect 14186 48864 14242 48920
rect 14094 47252 14150 47288
rect 14094 47232 14096 47252
rect 14096 47232 14148 47252
rect 14148 47232 14150 47252
rect 14002 41420 14004 41440
rect 14004 41420 14056 41440
rect 14056 41420 14058 41440
rect 14002 41384 14058 41420
rect 14289 48442 14345 48444
rect 14369 48442 14425 48444
rect 14449 48442 14505 48444
rect 14529 48442 14585 48444
rect 14289 48390 14315 48442
rect 14315 48390 14345 48442
rect 14369 48390 14379 48442
rect 14379 48390 14425 48442
rect 14449 48390 14495 48442
rect 14495 48390 14505 48442
rect 14529 48390 14559 48442
rect 14559 48390 14585 48442
rect 14289 48388 14345 48390
rect 14369 48388 14425 48390
rect 14449 48388 14505 48390
rect 14529 48388 14585 48390
rect 14289 47354 14345 47356
rect 14369 47354 14425 47356
rect 14449 47354 14505 47356
rect 14529 47354 14585 47356
rect 14289 47302 14315 47354
rect 14315 47302 14345 47354
rect 14369 47302 14379 47354
rect 14379 47302 14425 47354
rect 14449 47302 14495 47354
rect 14495 47302 14505 47354
rect 14529 47302 14559 47354
rect 14559 47302 14585 47354
rect 14289 47300 14345 47302
rect 14369 47300 14425 47302
rect 14449 47300 14505 47302
rect 14529 47300 14585 47302
rect 14289 46266 14345 46268
rect 14369 46266 14425 46268
rect 14449 46266 14505 46268
rect 14529 46266 14585 46268
rect 14289 46214 14315 46266
rect 14315 46214 14345 46266
rect 14369 46214 14379 46266
rect 14379 46214 14425 46266
rect 14449 46214 14495 46266
rect 14495 46214 14505 46266
rect 14529 46214 14559 46266
rect 14559 46214 14585 46266
rect 14289 46212 14345 46214
rect 14369 46212 14425 46214
rect 14449 46212 14505 46214
rect 14529 46212 14585 46214
rect 14922 56752 14978 56808
rect 14830 50904 14886 50960
rect 14830 49136 14886 49192
rect 14289 45178 14345 45180
rect 14369 45178 14425 45180
rect 14449 45178 14505 45180
rect 14529 45178 14585 45180
rect 14289 45126 14315 45178
rect 14315 45126 14345 45178
rect 14369 45126 14379 45178
rect 14379 45126 14425 45178
rect 14449 45126 14495 45178
rect 14495 45126 14505 45178
rect 14529 45126 14559 45178
rect 14559 45126 14585 45178
rect 14289 45124 14345 45126
rect 14369 45124 14425 45126
rect 14449 45124 14505 45126
rect 14529 45124 14585 45126
rect 14554 44684 14556 44704
rect 14556 44684 14608 44704
rect 14608 44684 14610 44704
rect 14554 44648 14610 44684
rect 14289 44090 14345 44092
rect 14369 44090 14425 44092
rect 14449 44090 14505 44092
rect 14529 44090 14585 44092
rect 14289 44038 14315 44090
rect 14315 44038 14345 44090
rect 14369 44038 14379 44090
rect 14379 44038 14425 44090
rect 14449 44038 14495 44090
rect 14495 44038 14505 44090
rect 14529 44038 14559 44090
rect 14559 44038 14585 44090
rect 14289 44036 14345 44038
rect 14369 44036 14425 44038
rect 14449 44036 14505 44038
rect 14529 44036 14585 44038
rect 14289 43002 14345 43004
rect 14369 43002 14425 43004
rect 14449 43002 14505 43004
rect 14529 43002 14585 43004
rect 14289 42950 14315 43002
rect 14315 42950 14345 43002
rect 14369 42950 14379 43002
rect 14379 42950 14425 43002
rect 14449 42950 14495 43002
rect 14495 42950 14505 43002
rect 14529 42950 14559 43002
rect 14559 42950 14585 43002
rect 14289 42948 14345 42950
rect 14369 42948 14425 42950
rect 14449 42948 14505 42950
rect 14529 42948 14585 42950
rect 14289 41914 14345 41916
rect 14369 41914 14425 41916
rect 14449 41914 14505 41916
rect 14529 41914 14585 41916
rect 14289 41862 14315 41914
rect 14315 41862 14345 41914
rect 14369 41862 14379 41914
rect 14379 41862 14425 41914
rect 14449 41862 14495 41914
rect 14495 41862 14505 41914
rect 14529 41862 14559 41914
rect 14559 41862 14585 41914
rect 14289 41860 14345 41862
rect 14369 41860 14425 41862
rect 14449 41860 14505 41862
rect 14529 41860 14585 41862
rect 14554 40976 14610 41032
rect 14289 40826 14345 40828
rect 14369 40826 14425 40828
rect 14449 40826 14505 40828
rect 14529 40826 14585 40828
rect 14289 40774 14315 40826
rect 14315 40774 14345 40826
rect 14369 40774 14379 40826
rect 14379 40774 14425 40826
rect 14449 40774 14495 40826
rect 14495 40774 14505 40826
rect 14529 40774 14559 40826
rect 14559 40774 14585 40826
rect 14289 40772 14345 40774
rect 14369 40772 14425 40774
rect 14449 40772 14505 40774
rect 14529 40772 14585 40774
rect 14830 45600 14886 45656
rect 15014 54984 15070 55040
rect 15106 50224 15162 50280
rect 15014 49680 15070 49736
rect 15106 45872 15162 45928
rect 15014 43832 15070 43888
rect 14289 39738 14345 39740
rect 14369 39738 14425 39740
rect 14449 39738 14505 39740
rect 14529 39738 14585 39740
rect 14289 39686 14315 39738
rect 14315 39686 14345 39738
rect 14369 39686 14379 39738
rect 14379 39686 14425 39738
rect 14449 39686 14495 39738
rect 14495 39686 14505 39738
rect 14529 39686 14559 39738
rect 14559 39686 14585 39738
rect 14289 39684 14345 39686
rect 14369 39684 14425 39686
rect 14449 39684 14505 39686
rect 14529 39684 14585 39686
rect 14646 39480 14702 39536
rect 14289 38650 14345 38652
rect 14369 38650 14425 38652
rect 14449 38650 14505 38652
rect 14529 38650 14585 38652
rect 14289 38598 14315 38650
rect 14315 38598 14345 38650
rect 14369 38598 14379 38650
rect 14379 38598 14425 38650
rect 14449 38598 14495 38650
rect 14495 38598 14505 38650
rect 14529 38598 14559 38650
rect 14559 38598 14585 38650
rect 14289 38596 14345 38598
rect 14369 38596 14425 38598
rect 14449 38596 14505 38598
rect 14529 38596 14585 38598
rect 14922 41248 14978 41304
rect 15106 43288 15162 43344
rect 15106 43152 15162 43208
rect 14646 38256 14702 38312
rect 14289 37562 14345 37564
rect 14369 37562 14425 37564
rect 14449 37562 14505 37564
rect 14529 37562 14585 37564
rect 14289 37510 14315 37562
rect 14315 37510 14345 37562
rect 14369 37510 14379 37562
rect 14379 37510 14425 37562
rect 14449 37510 14495 37562
rect 14495 37510 14505 37562
rect 14529 37510 14559 37562
rect 14559 37510 14585 37562
rect 14289 37508 14345 37510
rect 14369 37508 14425 37510
rect 14449 37508 14505 37510
rect 14529 37508 14585 37510
rect 13818 31184 13874 31240
rect 13542 26968 13598 27024
rect 13266 23060 13268 23080
rect 13268 23060 13320 23080
rect 13320 23060 13322 23080
rect 13266 23024 13322 23060
rect 13450 24928 13506 24984
rect 13634 22480 13690 22536
rect 14289 36474 14345 36476
rect 14369 36474 14425 36476
rect 14449 36474 14505 36476
rect 14529 36474 14585 36476
rect 14289 36422 14315 36474
rect 14315 36422 14345 36474
rect 14369 36422 14379 36474
rect 14379 36422 14425 36474
rect 14449 36422 14495 36474
rect 14495 36422 14505 36474
rect 14529 36422 14559 36474
rect 14559 36422 14585 36474
rect 14289 36420 14345 36422
rect 14369 36420 14425 36422
rect 14449 36420 14505 36422
rect 14529 36420 14585 36422
rect 14289 35386 14345 35388
rect 14369 35386 14425 35388
rect 14449 35386 14505 35388
rect 14529 35386 14585 35388
rect 14289 35334 14315 35386
rect 14315 35334 14345 35386
rect 14369 35334 14379 35386
rect 14379 35334 14425 35386
rect 14449 35334 14495 35386
rect 14495 35334 14505 35386
rect 14529 35334 14559 35386
rect 14559 35334 14585 35386
rect 14289 35332 14345 35334
rect 14369 35332 14425 35334
rect 14449 35332 14505 35334
rect 14529 35332 14585 35334
rect 14094 34448 14150 34504
rect 14289 34298 14345 34300
rect 14369 34298 14425 34300
rect 14449 34298 14505 34300
rect 14529 34298 14585 34300
rect 14289 34246 14315 34298
rect 14315 34246 14345 34298
rect 14369 34246 14379 34298
rect 14379 34246 14425 34298
rect 14449 34246 14495 34298
rect 14495 34246 14505 34298
rect 14529 34246 14559 34298
rect 14559 34246 14585 34298
rect 14289 34244 14345 34246
rect 14369 34244 14425 34246
rect 14449 34244 14505 34246
rect 14529 34244 14585 34246
rect 14289 33210 14345 33212
rect 14369 33210 14425 33212
rect 14449 33210 14505 33212
rect 14529 33210 14585 33212
rect 14289 33158 14315 33210
rect 14315 33158 14345 33210
rect 14369 33158 14379 33210
rect 14379 33158 14425 33210
rect 14449 33158 14495 33210
rect 14495 33158 14505 33210
rect 14529 33158 14559 33210
rect 14559 33158 14585 33210
rect 14289 33156 14345 33158
rect 14369 33156 14425 33158
rect 14449 33156 14505 33158
rect 14529 33156 14585 33158
rect 14289 32122 14345 32124
rect 14369 32122 14425 32124
rect 14449 32122 14505 32124
rect 14529 32122 14585 32124
rect 14289 32070 14315 32122
rect 14315 32070 14345 32122
rect 14369 32070 14379 32122
rect 14379 32070 14425 32122
rect 14449 32070 14495 32122
rect 14495 32070 14505 32122
rect 14529 32070 14559 32122
rect 14559 32070 14585 32122
rect 14289 32068 14345 32070
rect 14369 32068 14425 32070
rect 14449 32068 14505 32070
rect 14529 32068 14585 32070
rect 14289 31034 14345 31036
rect 14369 31034 14425 31036
rect 14449 31034 14505 31036
rect 14529 31034 14585 31036
rect 14289 30982 14315 31034
rect 14315 30982 14345 31034
rect 14369 30982 14379 31034
rect 14379 30982 14425 31034
rect 14449 30982 14495 31034
rect 14495 30982 14505 31034
rect 14529 30982 14559 31034
rect 14559 30982 14585 31034
rect 14289 30980 14345 30982
rect 14369 30980 14425 30982
rect 14449 30980 14505 30982
rect 14529 30980 14585 30982
rect 14186 30232 14242 30288
rect 14289 29946 14345 29948
rect 14369 29946 14425 29948
rect 14449 29946 14505 29948
rect 14529 29946 14585 29948
rect 14289 29894 14315 29946
rect 14315 29894 14345 29946
rect 14369 29894 14379 29946
rect 14379 29894 14425 29946
rect 14449 29894 14495 29946
rect 14495 29894 14505 29946
rect 14529 29894 14559 29946
rect 14559 29894 14585 29946
rect 14289 29892 14345 29894
rect 14369 29892 14425 29894
rect 14449 29892 14505 29894
rect 14529 29892 14585 29894
rect 14289 28858 14345 28860
rect 14369 28858 14425 28860
rect 14449 28858 14505 28860
rect 14529 28858 14585 28860
rect 14289 28806 14315 28858
rect 14315 28806 14345 28858
rect 14369 28806 14379 28858
rect 14379 28806 14425 28858
rect 14449 28806 14495 28858
rect 14495 28806 14505 28858
rect 14529 28806 14559 28858
rect 14559 28806 14585 28858
rect 14289 28804 14345 28806
rect 14369 28804 14425 28806
rect 14449 28804 14505 28806
rect 14529 28804 14585 28806
rect 15382 61104 15438 61160
rect 15382 60968 15438 61024
rect 15382 60016 15438 60072
rect 15566 62228 15568 62248
rect 15568 62228 15620 62248
rect 15620 62228 15622 62248
rect 15566 62192 15622 62228
rect 16210 63180 16212 63200
rect 16212 63180 16264 63200
rect 16264 63180 16266 63200
rect 16210 63144 16266 63180
rect 16118 60832 16174 60888
rect 16026 60424 16082 60480
rect 15474 57024 15530 57080
rect 15290 55120 15346 55176
rect 15382 54984 15438 55040
rect 15566 54576 15622 54632
rect 15474 53352 15530 53408
rect 15382 52400 15438 52456
rect 15290 52264 15346 52320
rect 15290 50904 15346 50960
rect 15842 57840 15898 57896
rect 17498 72528 17554 72584
rect 17622 71834 17678 71836
rect 17702 71834 17758 71836
rect 17782 71834 17838 71836
rect 17862 71834 17918 71836
rect 17622 71782 17648 71834
rect 17648 71782 17678 71834
rect 17702 71782 17712 71834
rect 17712 71782 17758 71834
rect 17782 71782 17828 71834
rect 17828 71782 17838 71834
rect 17862 71782 17892 71834
rect 17892 71782 17918 71834
rect 17622 71780 17678 71782
rect 17702 71780 17758 71782
rect 17782 71780 17838 71782
rect 17862 71780 17918 71782
rect 17622 70746 17678 70748
rect 17702 70746 17758 70748
rect 17782 70746 17838 70748
rect 17862 70746 17918 70748
rect 17622 70694 17648 70746
rect 17648 70694 17678 70746
rect 17702 70694 17712 70746
rect 17712 70694 17758 70746
rect 17782 70694 17828 70746
rect 17828 70694 17838 70746
rect 17862 70694 17892 70746
rect 17892 70694 17918 70746
rect 17622 70692 17678 70694
rect 17702 70692 17758 70694
rect 17782 70692 17838 70694
rect 17862 70692 17918 70694
rect 17622 69658 17678 69660
rect 17702 69658 17758 69660
rect 17782 69658 17838 69660
rect 17862 69658 17918 69660
rect 17622 69606 17648 69658
rect 17648 69606 17678 69658
rect 17702 69606 17712 69658
rect 17712 69606 17758 69658
rect 17782 69606 17828 69658
rect 17828 69606 17838 69658
rect 17862 69606 17892 69658
rect 17892 69606 17918 69658
rect 17622 69604 17678 69606
rect 17702 69604 17758 69606
rect 17782 69604 17838 69606
rect 17862 69604 17918 69606
rect 17498 68720 17554 68776
rect 17622 68570 17678 68572
rect 17702 68570 17758 68572
rect 17782 68570 17838 68572
rect 17862 68570 17918 68572
rect 17622 68518 17648 68570
rect 17648 68518 17678 68570
rect 17702 68518 17712 68570
rect 17712 68518 17758 68570
rect 17782 68518 17828 68570
rect 17828 68518 17838 68570
rect 17862 68518 17892 68570
rect 17892 68518 17918 68570
rect 17622 68516 17678 68518
rect 17702 68516 17758 68518
rect 17782 68516 17838 68518
rect 17862 68516 17918 68518
rect 17622 67482 17678 67484
rect 17702 67482 17758 67484
rect 17782 67482 17838 67484
rect 17862 67482 17918 67484
rect 17622 67430 17648 67482
rect 17648 67430 17678 67482
rect 17702 67430 17712 67482
rect 17712 67430 17758 67482
rect 17782 67430 17828 67482
rect 17828 67430 17838 67482
rect 17862 67430 17892 67482
rect 17892 67430 17918 67482
rect 17622 67428 17678 67430
rect 17702 67428 17758 67430
rect 17782 67428 17838 67430
rect 17862 67428 17918 67430
rect 17130 67224 17186 67280
rect 16394 65456 16450 65512
rect 17498 67088 17554 67144
rect 16670 66580 16672 66600
rect 16672 66580 16724 66600
rect 16724 66580 16726 66600
rect 16670 66544 16726 66580
rect 17622 66394 17678 66396
rect 17702 66394 17758 66396
rect 17782 66394 17838 66396
rect 17862 66394 17918 66396
rect 17622 66342 17648 66394
rect 17648 66342 17678 66394
rect 17702 66342 17712 66394
rect 17712 66342 17758 66394
rect 17782 66342 17828 66394
rect 17828 66342 17838 66394
rect 17862 66342 17892 66394
rect 17892 66342 17918 66394
rect 17622 66340 17678 66342
rect 17702 66340 17758 66342
rect 17782 66340 17838 66342
rect 17862 66340 17918 66342
rect 16486 64504 16542 64560
rect 16394 63824 16450 63880
rect 16486 61784 16542 61840
rect 16946 65864 17002 65920
rect 16854 64404 16856 64424
rect 16856 64404 16908 64424
rect 16908 64404 16910 64424
rect 16854 64368 16910 64404
rect 17498 65592 17554 65648
rect 17622 65306 17678 65308
rect 17702 65306 17758 65308
rect 17782 65306 17838 65308
rect 17862 65306 17918 65308
rect 17622 65254 17648 65306
rect 17648 65254 17678 65306
rect 17702 65254 17712 65306
rect 17712 65254 17758 65306
rect 17782 65254 17828 65306
rect 17828 65254 17838 65306
rect 17862 65254 17892 65306
rect 17892 65254 17918 65306
rect 17622 65252 17678 65254
rect 17702 65252 17758 65254
rect 17782 65252 17838 65254
rect 17862 65252 17918 65254
rect 17622 64218 17678 64220
rect 17702 64218 17758 64220
rect 17782 64218 17838 64220
rect 17862 64218 17918 64220
rect 17622 64166 17648 64218
rect 17648 64166 17678 64218
rect 17702 64166 17712 64218
rect 17712 64166 17758 64218
rect 17782 64166 17828 64218
rect 17828 64166 17838 64218
rect 17862 64166 17892 64218
rect 17892 64166 17918 64218
rect 17622 64164 17678 64166
rect 17702 64164 17758 64166
rect 17782 64164 17838 64166
rect 17862 64164 17918 64166
rect 17622 63130 17678 63132
rect 17702 63130 17758 63132
rect 17782 63130 17838 63132
rect 17862 63130 17918 63132
rect 17622 63078 17648 63130
rect 17648 63078 17678 63130
rect 17702 63078 17712 63130
rect 17712 63078 17758 63130
rect 17782 63078 17828 63130
rect 17828 63078 17838 63130
rect 17862 63078 17892 63130
rect 17892 63078 17918 63130
rect 17622 63076 17678 63078
rect 17702 63076 17758 63078
rect 17782 63076 17838 63078
rect 17862 63076 17918 63078
rect 17498 62736 17554 62792
rect 17622 62042 17678 62044
rect 17702 62042 17758 62044
rect 17782 62042 17838 62044
rect 17862 62042 17918 62044
rect 17622 61990 17648 62042
rect 17648 61990 17678 62042
rect 17702 61990 17712 62042
rect 17712 61990 17758 62042
rect 17782 61990 17828 62042
rect 17828 61990 17838 62042
rect 17862 61990 17892 62042
rect 17892 61990 17918 62042
rect 17622 61988 17678 61990
rect 17702 61988 17758 61990
rect 17782 61988 17838 61990
rect 17862 61988 17918 61990
rect 17622 60954 17678 60956
rect 17702 60954 17758 60956
rect 17782 60954 17838 60956
rect 17862 60954 17918 60956
rect 17622 60902 17648 60954
rect 17648 60902 17678 60954
rect 17702 60902 17712 60954
rect 17712 60902 17758 60954
rect 17782 60902 17828 60954
rect 17828 60902 17838 60954
rect 17862 60902 17892 60954
rect 17892 60902 17918 60954
rect 17622 60900 17678 60902
rect 17702 60900 17758 60902
rect 17782 60900 17838 60902
rect 17862 60900 17918 60902
rect 17498 60560 17554 60616
rect 16670 60288 16726 60344
rect 16578 60152 16634 60208
rect 17622 59866 17678 59868
rect 17702 59866 17758 59868
rect 17782 59866 17838 59868
rect 17862 59866 17918 59868
rect 17622 59814 17648 59866
rect 17648 59814 17678 59866
rect 17702 59814 17712 59866
rect 17712 59814 17758 59866
rect 17782 59814 17828 59866
rect 17828 59814 17838 59866
rect 17862 59814 17892 59866
rect 17892 59814 17918 59866
rect 17622 59812 17678 59814
rect 17702 59812 17758 59814
rect 17782 59812 17838 59814
rect 17862 59812 17918 59814
rect 16486 59064 16542 59120
rect 17622 58778 17678 58780
rect 17702 58778 17758 58780
rect 17782 58778 17838 58780
rect 17862 58778 17918 58780
rect 17622 58726 17648 58778
rect 17648 58726 17678 58778
rect 17702 58726 17712 58778
rect 17712 58726 17758 58778
rect 17782 58726 17828 58778
rect 17828 58726 17838 58778
rect 17862 58726 17892 58778
rect 17892 58726 17918 58778
rect 17622 58724 17678 58726
rect 17702 58724 17758 58726
rect 17782 58724 17838 58726
rect 17862 58724 17918 58726
rect 16394 58384 16450 58440
rect 16302 57976 16358 58032
rect 17622 57690 17678 57692
rect 17702 57690 17758 57692
rect 17782 57690 17838 57692
rect 17862 57690 17918 57692
rect 17622 57638 17648 57690
rect 17648 57638 17678 57690
rect 17702 57638 17712 57690
rect 17712 57638 17758 57690
rect 17782 57638 17828 57690
rect 17828 57638 17838 57690
rect 17862 57638 17892 57690
rect 17892 57638 17918 57690
rect 17622 57636 17678 57638
rect 17702 57636 17758 57638
rect 17782 57636 17838 57638
rect 17862 57636 17918 57638
rect 16026 57296 16082 57352
rect 15750 52808 15806 52864
rect 16670 56652 16672 56672
rect 16672 56652 16724 56672
rect 16724 56652 16726 56672
rect 16670 56616 16726 56652
rect 16210 56344 16266 56400
rect 17622 56602 17678 56604
rect 17702 56602 17758 56604
rect 17782 56602 17838 56604
rect 17862 56602 17918 56604
rect 17622 56550 17648 56602
rect 17648 56550 17678 56602
rect 17702 56550 17712 56602
rect 17712 56550 17758 56602
rect 17782 56550 17828 56602
rect 17828 56550 17838 56602
rect 17862 56550 17892 56602
rect 17892 56550 17918 56602
rect 17622 56548 17678 56550
rect 17702 56548 17758 56550
rect 17782 56548 17838 56550
rect 17862 56548 17918 56550
rect 17498 55800 17554 55856
rect 16394 55664 16450 55720
rect 17130 55412 17186 55448
rect 17130 55392 17132 55412
rect 17132 55392 17184 55412
rect 17184 55392 17186 55412
rect 16026 54168 16082 54224
rect 15658 49408 15714 49464
rect 15658 49272 15714 49328
rect 15566 47132 15568 47152
rect 15568 47132 15620 47152
rect 15620 47132 15622 47152
rect 15566 47096 15622 47132
rect 15290 42200 15346 42256
rect 15198 40704 15254 40760
rect 15106 39344 15162 39400
rect 17622 55514 17678 55516
rect 17702 55514 17758 55516
rect 17782 55514 17838 55516
rect 17862 55514 17918 55516
rect 17622 55462 17648 55514
rect 17648 55462 17678 55514
rect 17702 55462 17712 55514
rect 17712 55462 17758 55514
rect 17782 55462 17828 55514
rect 17828 55462 17838 55514
rect 17862 55462 17892 55514
rect 17892 55462 17918 55514
rect 17622 55460 17678 55462
rect 17702 55460 17758 55462
rect 17782 55460 17838 55462
rect 17862 55460 17918 55462
rect 16118 51176 16174 51232
rect 16118 50904 16174 50960
rect 16026 49816 16082 49872
rect 15934 45056 15990 45112
rect 15658 43968 15714 44024
rect 15566 41656 15622 41712
rect 15474 41520 15530 41576
rect 14830 34060 14886 34096
rect 14830 34040 14832 34060
rect 14832 34040 14884 34060
rect 14884 34040 14886 34060
rect 14830 30232 14886 30288
rect 14289 27770 14345 27772
rect 14369 27770 14425 27772
rect 14449 27770 14505 27772
rect 14529 27770 14585 27772
rect 14289 27718 14315 27770
rect 14315 27718 14345 27770
rect 14369 27718 14379 27770
rect 14379 27718 14425 27770
rect 14449 27718 14495 27770
rect 14495 27718 14505 27770
rect 14529 27718 14559 27770
rect 14559 27718 14585 27770
rect 14289 27716 14345 27718
rect 14369 27716 14425 27718
rect 14449 27716 14505 27718
rect 14529 27716 14585 27718
rect 14289 26682 14345 26684
rect 14369 26682 14425 26684
rect 14449 26682 14505 26684
rect 14529 26682 14585 26684
rect 14289 26630 14315 26682
rect 14315 26630 14345 26682
rect 14369 26630 14379 26682
rect 14379 26630 14425 26682
rect 14449 26630 14495 26682
rect 14495 26630 14505 26682
rect 14529 26630 14559 26682
rect 14559 26630 14585 26682
rect 14289 26628 14345 26630
rect 14369 26628 14425 26630
rect 14449 26628 14505 26630
rect 14529 26628 14585 26630
rect 14289 25594 14345 25596
rect 14369 25594 14425 25596
rect 14449 25594 14505 25596
rect 14529 25594 14585 25596
rect 14289 25542 14315 25594
rect 14315 25542 14345 25594
rect 14369 25542 14379 25594
rect 14379 25542 14425 25594
rect 14449 25542 14495 25594
rect 14495 25542 14505 25594
rect 14529 25542 14559 25594
rect 14559 25542 14585 25594
rect 14289 25540 14345 25542
rect 14369 25540 14425 25542
rect 14449 25540 14505 25542
rect 14529 25540 14585 25542
rect 14002 24792 14058 24848
rect 14289 24506 14345 24508
rect 14369 24506 14425 24508
rect 14449 24506 14505 24508
rect 14529 24506 14585 24508
rect 14289 24454 14315 24506
rect 14315 24454 14345 24506
rect 14369 24454 14379 24506
rect 14379 24454 14425 24506
rect 14449 24454 14495 24506
rect 14495 24454 14505 24506
rect 14529 24454 14559 24506
rect 14559 24454 14585 24506
rect 14289 24452 14345 24454
rect 14369 24452 14425 24454
rect 14449 24452 14505 24454
rect 14529 24452 14585 24454
rect 15106 37848 15162 37904
rect 15566 41248 15622 41304
rect 15382 37460 15438 37496
rect 15382 37440 15384 37460
rect 15384 37440 15436 37460
rect 15436 37440 15438 37460
rect 15382 37168 15438 37224
rect 15106 32816 15162 32872
rect 16578 53388 16580 53408
rect 16580 53388 16632 53408
rect 16632 53388 16634 53408
rect 16578 53352 16634 53388
rect 16854 53080 16910 53136
rect 16762 52944 16818 53000
rect 16302 49816 16358 49872
rect 16670 49680 16726 49736
rect 16670 49172 16672 49192
rect 16672 49172 16724 49192
rect 16724 49172 16726 49192
rect 16670 49136 16726 49172
rect 16394 47096 16450 47152
rect 16302 46960 16358 47016
rect 15842 43424 15898 43480
rect 16026 42744 16082 42800
rect 15934 42336 15990 42392
rect 15750 41692 15752 41712
rect 15752 41692 15804 41712
rect 15804 41692 15806 41712
rect 15750 41656 15806 41692
rect 15658 39208 15714 39264
rect 15934 39500 15990 39536
rect 15934 39480 15936 39500
rect 15936 39480 15988 39500
rect 15988 39480 15990 39500
rect 15658 35672 15714 35728
rect 15566 34448 15622 34504
rect 15566 33496 15622 33552
rect 15290 31184 15346 31240
rect 14646 23704 14702 23760
rect 13818 22752 13874 22808
rect 13542 19080 13598 19136
rect 13818 19896 13874 19952
rect 12990 10376 13046 10432
rect 13634 18300 13636 18320
rect 13636 18300 13688 18320
rect 13688 18300 13690 18320
rect 13634 18264 13690 18300
rect 13818 13912 13874 13968
rect 13726 12708 13782 12744
rect 13726 12688 13728 12708
rect 13728 12688 13780 12708
rect 13780 12688 13782 12708
rect 13634 11772 13636 11792
rect 13636 11772 13688 11792
rect 13688 11772 13690 11792
rect 13634 11736 13690 11772
rect 14289 23418 14345 23420
rect 14369 23418 14425 23420
rect 14449 23418 14505 23420
rect 14529 23418 14585 23420
rect 14289 23366 14315 23418
rect 14315 23366 14345 23418
rect 14369 23366 14379 23418
rect 14379 23366 14425 23418
rect 14449 23366 14495 23418
rect 14495 23366 14505 23418
rect 14529 23366 14559 23418
rect 14559 23366 14585 23418
rect 14289 23364 14345 23366
rect 14369 23364 14425 23366
rect 14449 23364 14505 23366
rect 14529 23364 14585 23366
rect 14289 22330 14345 22332
rect 14369 22330 14425 22332
rect 14449 22330 14505 22332
rect 14529 22330 14585 22332
rect 14289 22278 14315 22330
rect 14315 22278 14345 22330
rect 14369 22278 14379 22330
rect 14379 22278 14425 22330
rect 14449 22278 14495 22330
rect 14495 22278 14505 22330
rect 14529 22278 14559 22330
rect 14559 22278 14585 22330
rect 14289 22276 14345 22278
rect 14369 22276 14425 22278
rect 14449 22276 14505 22278
rect 14529 22276 14585 22278
rect 14370 22072 14426 22128
rect 15014 23568 15070 23624
rect 14289 21242 14345 21244
rect 14369 21242 14425 21244
rect 14449 21242 14505 21244
rect 14529 21242 14585 21244
rect 14289 21190 14315 21242
rect 14315 21190 14345 21242
rect 14369 21190 14379 21242
rect 14379 21190 14425 21242
rect 14449 21190 14495 21242
rect 14495 21190 14505 21242
rect 14529 21190 14559 21242
rect 14559 21190 14585 21242
rect 14289 21188 14345 21190
rect 14369 21188 14425 21190
rect 14449 21188 14505 21190
rect 14529 21188 14585 21190
rect 15198 22480 15254 22536
rect 14289 20154 14345 20156
rect 14369 20154 14425 20156
rect 14449 20154 14505 20156
rect 14529 20154 14585 20156
rect 14289 20102 14315 20154
rect 14315 20102 14345 20154
rect 14369 20102 14379 20154
rect 14379 20102 14425 20154
rect 14449 20102 14495 20154
rect 14495 20102 14505 20154
rect 14529 20102 14559 20154
rect 14559 20102 14585 20154
rect 14289 20100 14345 20102
rect 14369 20100 14425 20102
rect 14449 20100 14505 20102
rect 14529 20100 14585 20102
rect 14738 19780 14794 19816
rect 14738 19760 14740 19780
rect 14740 19760 14792 19780
rect 14792 19760 14794 19780
rect 14186 19216 14242 19272
rect 14289 19066 14345 19068
rect 14369 19066 14425 19068
rect 14449 19066 14505 19068
rect 14529 19066 14585 19068
rect 14289 19014 14315 19066
rect 14315 19014 14345 19066
rect 14369 19014 14379 19066
rect 14379 19014 14425 19066
rect 14449 19014 14495 19066
rect 14495 19014 14505 19066
rect 14529 19014 14559 19066
rect 14559 19014 14585 19066
rect 14289 19012 14345 19014
rect 14369 19012 14425 19014
rect 14449 19012 14505 19014
rect 14529 19012 14585 19014
rect 14646 18420 14702 18456
rect 14646 18400 14648 18420
rect 14648 18400 14700 18420
rect 14700 18400 14702 18420
rect 14289 17978 14345 17980
rect 14369 17978 14425 17980
rect 14449 17978 14505 17980
rect 14529 17978 14585 17980
rect 14289 17926 14315 17978
rect 14315 17926 14345 17978
rect 14369 17926 14379 17978
rect 14379 17926 14425 17978
rect 14449 17926 14495 17978
rect 14495 17926 14505 17978
rect 14529 17926 14559 17978
rect 14559 17926 14585 17978
rect 14289 17924 14345 17926
rect 14369 17924 14425 17926
rect 14449 17924 14505 17926
rect 14529 17924 14585 17926
rect 14289 16890 14345 16892
rect 14369 16890 14425 16892
rect 14449 16890 14505 16892
rect 14529 16890 14585 16892
rect 14289 16838 14315 16890
rect 14315 16838 14345 16890
rect 14369 16838 14379 16890
rect 14379 16838 14425 16890
rect 14449 16838 14495 16890
rect 14495 16838 14505 16890
rect 14529 16838 14559 16890
rect 14559 16838 14585 16890
rect 14289 16836 14345 16838
rect 14369 16836 14425 16838
rect 14449 16836 14505 16838
rect 14529 16836 14585 16838
rect 14289 15802 14345 15804
rect 14369 15802 14425 15804
rect 14449 15802 14505 15804
rect 14529 15802 14585 15804
rect 14289 15750 14315 15802
rect 14315 15750 14345 15802
rect 14369 15750 14379 15802
rect 14379 15750 14425 15802
rect 14449 15750 14495 15802
rect 14495 15750 14505 15802
rect 14529 15750 14559 15802
rect 14559 15750 14585 15802
rect 14289 15748 14345 15750
rect 14369 15748 14425 15750
rect 14449 15748 14505 15750
rect 14529 15748 14585 15750
rect 14278 15272 14334 15328
rect 14289 14714 14345 14716
rect 14369 14714 14425 14716
rect 14449 14714 14505 14716
rect 14529 14714 14585 14716
rect 14289 14662 14315 14714
rect 14315 14662 14345 14714
rect 14369 14662 14379 14714
rect 14379 14662 14425 14714
rect 14449 14662 14495 14714
rect 14495 14662 14505 14714
rect 14529 14662 14559 14714
rect 14559 14662 14585 14714
rect 14289 14660 14345 14662
rect 14369 14660 14425 14662
rect 14449 14660 14505 14662
rect 14529 14660 14585 14662
rect 14289 13626 14345 13628
rect 14369 13626 14425 13628
rect 14449 13626 14505 13628
rect 14529 13626 14585 13628
rect 14289 13574 14315 13626
rect 14315 13574 14345 13626
rect 14369 13574 14379 13626
rect 14379 13574 14425 13626
rect 14449 13574 14495 13626
rect 14495 13574 14505 13626
rect 14529 13574 14559 13626
rect 14559 13574 14585 13626
rect 14289 13572 14345 13574
rect 14369 13572 14425 13574
rect 14449 13572 14505 13574
rect 14529 13572 14585 13574
rect 14289 12538 14345 12540
rect 14369 12538 14425 12540
rect 14449 12538 14505 12540
rect 14529 12538 14585 12540
rect 14289 12486 14315 12538
rect 14315 12486 14345 12538
rect 14369 12486 14379 12538
rect 14379 12486 14425 12538
rect 14449 12486 14495 12538
rect 14495 12486 14505 12538
rect 14529 12486 14559 12538
rect 14559 12486 14585 12538
rect 14289 12484 14345 12486
rect 14369 12484 14425 12486
rect 14449 12484 14505 12486
rect 14529 12484 14585 12486
rect 14186 12300 14242 12336
rect 14186 12280 14188 12300
rect 14188 12280 14240 12300
rect 14240 12280 14242 12300
rect 14186 11872 14242 11928
rect 14278 11636 14280 11656
rect 14280 11636 14332 11656
rect 14332 11636 14334 11656
rect 14278 11600 14334 11636
rect 14289 11450 14345 11452
rect 14369 11450 14425 11452
rect 14449 11450 14505 11452
rect 14529 11450 14585 11452
rect 14289 11398 14315 11450
rect 14315 11398 14345 11450
rect 14369 11398 14379 11450
rect 14379 11398 14425 11450
rect 14449 11398 14495 11450
rect 14495 11398 14505 11450
rect 14529 11398 14559 11450
rect 14559 11398 14585 11450
rect 14289 11396 14345 11398
rect 14369 11396 14425 11398
rect 14449 11396 14505 11398
rect 14529 11396 14585 11398
rect 13818 10548 13820 10568
rect 13820 10548 13872 10568
rect 13872 10548 13874 10568
rect 13818 10512 13874 10548
rect 13174 9424 13230 9480
rect 12990 8880 13046 8936
rect 14002 9560 14058 9616
rect 14289 10362 14345 10364
rect 14369 10362 14425 10364
rect 14449 10362 14505 10364
rect 14529 10362 14585 10364
rect 14289 10310 14315 10362
rect 14315 10310 14345 10362
rect 14369 10310 14379 10362
rect 14379 10310 14425 10362
rect 14449 10310 14495 10362
rect 14495 10310 14505 10362
rect 14529 10310 14559 10362
rect 14559 10310 14585 10362
rect 14289 10308 14345 10310
rect 14369 10308 14425 10310
rect 14449 10308 14505 10310
rect 14529 10308 14585 10310
rect 14186 9424 14242 9480
rect 14289 9274 14345 9276
rect 14369 9274 14425 9276
rect 14449 9274 14505 9276
rect 14529 9274 14585 9276
rect 14289 9222 14315 9274
rect 14315 9222 14345 9274
rect 14369 9222 14379 9274
rect 14379 9222 14425 9274
rect 14449 9222 14495 9274
rect 14495 9222 14505 9274
rect 14529 9222 14559 9274
rect 14559 9222 14585 9274
rect 14289 9220 14345 9222
rect 14369 9220 14425 9222
rect 14449 9220 14505 9222
rect 14529 9220 14585 9222
rect 13634 6332 13636 6352
rect 13636 6332 13688 6352
rect 13688 6332 13690 6352
rect 13634 6296 13690 6332
rect 14186 8336 14242 8392
rect 14289 8186 14345 8188
rect 14369 8186 14425 8188
rect 14449 8186 14505 8188
rect 14529 8186 14585 8188
rect 14289 8134 14315 8186
rect 14315 8134 14345 8186
rect 14369 8134 14379 8186
rect 14379 8134 14425 8186
rect 14449 8134 14495 8186
rect 14495 8134 14505 8186
rect 14529 8134 14559 8186
rect 14559 8134 14585 8186
rect 14289 8132 14345 8134
rect 14369 8132 14425 8134
rect 14449 8132 14505 8134
rect 14529 8132 14585 8134
rect 14289 7098 14345 7100
rect 14369 7098 14425 7100
rect 14449 7098 14505 7100
rect 14529 7098 14585 7100
rect 14289 7046 14315 7098
rect 14315 7046 14345 7098
rect 14369 7046 14379 7098
rect 14379 7046 14425 7098
rect 14449 7046 14495 7098
rect 14495 7046 14505 7098
rect 14529 7046 14559 7098
rect 14559 7046 14585 7098
rect 14289 7044 14345 7046
rect 14369 7044 14425 7046
rect 14449 7044 14505 7046
rect 14529 7044 14585 7046
rect 15566 25880 15622 25936
rect 15842 30268 15844 30288
rect 15844 30268 15896 30288
rect 15896 30268 15898 30288
rect 15842 30232 15898 30268
rect 16394 43696 16450 43752
rect 16394 42744 16450 42800
rect 16394 41520 16450 41576
rect 16302 41112 16358 41168
rect 16210 40568 16266 40624
rect 16302 39500 16358 39536
rect 16302 39480 16304 39500
rect 16304 39480 16356 39500
rect 16356 39480 16358 39500
rect 16486 39888 16542 39944
rect 17622 54426 17678 54428
rect 17702 54426 17758 54428
rect 17782 54426 17838 54428
rect 17862 54426 17918 54428
rect 17622 54374 17648 54426
rect 17648 54374 17678 54426
rect 17702 54374 17712 54426
rect 17712 54374 17758 54426
rect 17782 54374 17828 54426
rect 17828 54374 17838 54426
rect 17862 54374 17892 54426
rect 17892 54374 17918 54426
rect 17622 54372 17678 54374
rect 17702 54372 17758 54374
rect 17782 54372 17838 54374
rect 17862 54372 17918 54374
rect 17406 53352 17462 53408
rect 17622 53338 17678 53340
rect 17702 53338 17758 53340
rect 17782 53338 17838 53340
rect 17862 53338 17918 53340
rect 17622 53286 17648 53338
rect 17648 53286 17678 53338
rect 17702 53286 17712 53338
rect 17712 53286 17758 53338
rect 17782 53286 17828 53338
rect 17828 53286 17838 53338
rect 17862 53286 17892 53338
rect 17892 53286 17918 53338
rect 17622 53284 17678 53286
rect 17702 53284 17758 53286
rect 17782 53284 17838 53286
rect 17862 53284 17918 53286
rect 17958 52980 17960 53000
rect 17960 52980 18012 53000
rect 18012 52980 18014 53000
rect 17958 52944 18014 52980
rect 17622 52250 17678 52252
rect 17702 52250 17758 52252
rect 17782 52250 17838 52252
rect 17862 52250 17918 52252
rect 17622 52198 17648 52250
rect 17648 52198 17678 52250
rect 17702 52198 17712 52250
rect 17712 52198 17758 52250
rect 17782 52198 17828 52250
rect 17828 52198 17838 52250
rect 17862 52198 17892 52250
rect 17892 52198 17918 52250
rect 17622 52196 17678 52198
rect 17702 52196 17758 52198
rect 17782 52196 17838 52198
rect 17862 52196 17918 52198
rect 17498 51856 17554 51912
rect 17038 47096 17094 47152
rect 16946 46960 17002 47016
rect 16762 41676 16818 41712
rect 16762 41656 16764 41676
rect 16764 41656 16816 41676
rect 16816 41656 16818 41676
rect 15658 24928 15714 24984
rect 15658 24792 15714 24848
rect 16302 27940 16358 27976
rect 16302 27920 16304 27940
rect 16304 27920 16356 27940
rect 16356 27920 16358 27940
rect 17222 46416 17278 46472
rect 17038 41384 17094 41440
rect 17038 41248 17094 41304
rect 17622 51162 17678 51164
rect 17702 51162 17758 51164
rect 17782 51162 17838 51164
rect 17862 51162 17918 51164
rect 17622 51110 17648 51162
rect 17648 51110 17678 51162
rect 17702 51110 17712 51162
rect 17712 51110 17758 51162
rect 17782 51110 17828 51162
rect 17828 51110 17838 51162
rect 17862 51110 17892 51162
rect 17892 51110 17918 51162
rect 17622 51108 17678 51110
rect 17702 51108 17758 51110
rect 17782 51108 17838 51110
rect 17862 51108 17918 51110
rect 18142 50088 18198 50144
rect 17622 50074 17678 50076
rect 17702 50074 17758 50076
rect 17782 50074 17838 50076
rect 17862 50074 17918 50076
rect 17622 50022 17648 50074
rect 17648 50022 17678 50074
rect 17702 50022 17712 50074
rect 17712 50022 17758 50074
rect 17782 50022 17828 50074
rect 17828 50022 17838 50074
rect 17862 50022 17892 50074
rect 17892 50022 17918 50074
rect 17622 50020 17678 50022
rect 17702 50020 17758 50022
rect 17782 50020 17838 50022
rect 17862 50020 17918 50022
rect 17622 48986 17678 48988
rect 17702 48986 17758 48988
rect 17782 48986 17838 48988
rect 17862 48986 17918 48988
rect 17622 48934 17648 48986
rect 17648 48934 17678 48986
rect 17702 48934 17712 48986
rect 17712 48934 17758 48986
rect 17782 48934 17828 48986
rect 17828 48934 17838 48986
rect 17862 48934 17892 48986
rect 17892 48934 17918 48986
rect 17622 48932 17678 48934
rect 17702 48932 17758 48934
rect 17782 48932 17838 48934
rect 17862 48932 17918 48934
rect 17622 47898 17678 47900
rect 17702 47898 17758 47900
rect 17782 47898 17838 47900
rect 17862 47898 17918 47900
rect 17622 47846 17648 47898
rect 17648 47846 17678 47898
rect 17702 47846 17712 47898
rect 17712 47846 17758 47898
rect 17782 47846 17828 47898
rect 17828 47846 17838 47898
rect 17862 47846 17892 47898
rect 17892 47846 17918 47898
rect 17622 47844 17678 47846
rect 17702 47844 17758 47846
rect 17782 47844 17838 47846
rect 17862 47844 17918 47846
rect 17622 46810 17678 46812
rect 17702 46810 17758 46812
rect 17782 46810 17838 46812
rect 17862 46810 17918 46812
rect 17622 46758 17648 46810
rect 17648 46758 17678 46810
rect 17702 46758 17712 46810
rect 17712 46758 17758 46810
rect 17782 46758 17828 46810
rect 17828 46758 17838 46810
rect 17862 46758 17892 46810
rect 17892 46758 17918 46810
rect 17622 46756 17678 46758
rect 17702 46756 17758 46758
rect 17782 46756 17838 46758
rect 17862 46756 17918 46758
rect 17622 45722 17678 45724
rect 17702 45722 17758 45724
rect 17782 45722 17838 45724
rect 17862 45722 17918 45724
rect 17622 45670 17648 45722
rect 17648 45670 17678 45722
rect 17702 45670 17712 45722
rect 17712 45670 17758 45722
rect 17782 45670 17828 45722
rect 17828 45670 17838 45722
rect 17862 45670 17892 45722
rect 17892 45670 17918 45722
rect 17622 45668 17678 45670
rect 17702 45668 17758 45670
rect 17782 45668 17838 45670
rect 17862 45668 17918 45670
rect 17622 44634 17678 44636
rect 17702 44634 17758 44636
rect 17782 44634 17838 44636
rect 17862 44634 17918 44636
rect 17622 44582 17648 44634
rect 17648 44582 17678 44634
rect 17702 44582 17712 44634
rect 17712 44582 17758 44634
rect 17782 44582 17828 44634
rect 17828 44582 17838 44634
rect 17862 44582 17892 44634
rect 17892 44582 17918 44634
rect 17622 44580 17678 44582
rect 17702 44580 17758 44582
rect 17782 44580 17838 44582
rect 17862 44580 17918 44582
rect 17622 43546 17678 43548
rect 17702 43546 17758 43548
rect 17782 43546 17838 43548
rect 17862 43546 17918 43548
rect 17622 43494 17648 43546
rect 17648 43494 17678 43546
rect 17702 43494 17712 43546
rect 17712 43494 17758 43546
rect 17782 43494 17828 43546
rect 17828 43494 17838 43546
rect 17862 43494 17892 43546
rect 17892 43494 17918 43546
rect 17622 43492 17678 43494
rect 17702 43492 17758 43494
rect 17782 43492 17838 43494
rect 17862 43492 17918 43494
rect 17622 42458 17678 42460
rect 17702 42458 17758 42460
rect 17782 42458 17838 42460
rect 17862 42458 17918 42460
rect 17622 42406 17648 42458
rect 17648 42406 17678 42458
rect 17702 42406 17712 42458
rect 17712 42406 17758 42458
rect 17782 42406 17828 42458
rect 17828 42406 17838 42458
rect 17862 42406 17892 42458
rect 17892 42406 17918 42458
rect 17622 42404 17678 42406
rect 17702 42404 17758 42406
rect 17782 42404 17838 42406
rect 17862 42404 17918 42406
rect 17958 42064 18014 42120
rect 17774 41792 17830 41848
rect 17222 40296 17278 40352
rect 17222 40024 17278 40080
rect 16118 24928 16174 24984
rect 15198 21392 15254 21448
rect 15106 21256 15162 21312
rect 16118 22772 16174 22808
rect 16118 22752 16120 22772
rect 16120 22752 16172 22772
rect 16172 22752 16174 22772
rect 16026 22616 16082 22672
rect 15934 21256 15990 21312
rect 16394 25472 16450 25528
rect 17130 36488 17186 36544
rect 17130 34448 17186 34504
rect 17130 33940 17132 33960
rect 17132 33940 17184 33960
rect 17184 33940 17186 33960
rect 17130 33904 17186 33940
rect 17038 33496 17094 33552
rect 17130 33088 17186 33144
rect 17130 32816 17186 32872
rect 17622 41370 17678 41372
rect 17702 41370 17758 41372
rect 17782 41370 17838 41372
rect 17862 41370 17918 41372
rect 17622 41318 17648 41370
rect 17648 41318 17678 41370
rect 17702 41318 17712 41370
rect 17712 41318 17758 41370
rect 17782 41318 17828 41370
rect 17828 41318 17838 41370
rect 17862 41318 17892 41370
rect 17892 41318 17918 41370
rect 17622 41316 17678 41318
rect 17702 41316 17758 41318
rect 17782 41316 17838 41318
rect 17862 41316 17918 41318
rect 17622 40282 17678 40284
rect 17702 40282 17758 40284
rect 17782 40282 17838 40284
rect 17862 40282 17918 40284
rect 17622 40230 17648 40282
rect 17648 40230 17678 40282
rect 17702 40230 17712 40282
rect 17712 40230 17758 40282
rect 17782 40230 17828 40282
rect 17828 40230 17838 40282
rect 17862 40230 17892 40282
rect 17892 40230 17918 40282
rect 17622 40228 17678 40230
rect 17702 40228 17758 40230
rect 17782 40228 17838 40230
rect 17862 40228 17918 40230
rect 17622 39194 17678 39196
rect 17702 39194 17758 39196
rect 17782 39194 17838 39196
rect 17862 39194 17918 39196
rect 17622 39142 17648 39194
rect 17648 39142 17678 39194
rect 17702 39142 17712 39194
rect 17712 39142 17758 39194
rect 17782 39142 17828 39194
rect 17828 39142 17838 39194
rect 17862 39142 17892 39194
rect 17892 39142 17918 39194
rect 17622 39140 17678 39142
rect 17702 39140 17758 39142
rect 17782 39140 17838 39142
rect 17862 39140 17918 39142
rect 18234 42608 18290 42664
rect 18234 39480 18290 39536
rect 17622 38106 17678 38108
rect 17702 38106 17758 38108
rect 17782 38106 17838 38108
rect 17862 38106 17918 38108
rect 17622 38054 17648 38106
rect 17648 38054 17678 38106
rect 17702 38054 17712 38106
rect 17712 38054 17758 38106
rect 17782 38054 17828 38106
rect 17828 38054 17838 38106
rect 17862 38054 17892 38106
rect 17892 38054 17918 38106
rect 17622 38052 17678 38054
rect 17702 38052 17758 38054
rect 17782 38052 17838 38054
rect 17862 38052 17918 38054
rect 17498 37168 17554 37224
rect 17622 37018 17678 37020
rect 17702 37018 17758 37020
rect 17782 37018 17838 37020
rect 17862 37018 17918 37020
rect 17622 36966 17648 37018
rect 17648 36966 17678 37018
rect 17702 36966 17712 37018
rect 17712 36966 17758 37018
rect 17782 36966 17828 37018
rect 17828 36966 17838 37018
rect 17862 36966 17892 37018
rect 17892 36966 17918 37018
rect 17622 36964 17678 36966
rect 17702 36964 17758 36966
rect 17782 36964 17838 36966
rect 17862 36964 17918 36966
rect 17622 35930 17678 35932
rect 17702 35930 17758 35932
rect 17782 35930 17838 35932
rect 17862 35930 17918 35932
rect 17622 35878 17648 35930
rect 17648 35878 17678 35930
rect 17702 35878 17712 35930
rect 17712 35878 17758 35930
rect 17782 35878 17828 35930
rect 17828 35878 17838 35930
rect 17862 35878 17892 35930
rect 17892 35878 17918 35930
rect 17622 35876 17678 35878
rect 17702 35876 17758 35878
rect 17782 35876 17838 35878
rect 17862 35876 17918 35878
rect 17498 35128 17554 35184
rect 17622 34842 17678 34844
rect 17702 34842 17758 34844
rect 17782 34842 17838 34844
rect 17862 34842 17918 34844
rect 17622 34790 17648 34842
rect 17648 34790 17678 34842
rect 17702 34790 17712 34842
rect 17712 34790 17758 34842
rect 17782 34790 17828 34842
rect 17828 34790 17838 34842
rect 17862 34790 17892 34842
rect 17892 34790 17918 34842
rect 17622 34788 17678 34790
rect 17702 34788 17758 34790
rect 17782 34788 17838 34790
rect 17862 34788 17918 34790
rect 17622 33754 17678 33756
rect 17702 33754 17758 33756
rect 17782 33754 17838 33756
rect 17862 33754 17918 33756
rect 17622 33702 17648 33754
rect 17648 33702 17678 33754
rect 17702 33702 17712 33754
rect 17712 33702 17758 33754
rect 17782 33702 17828 33754
rect 17828 33702 17838 33754
rect 17862 33702 17892 33754
rect 17892 33702 17918 33754
rect 17622 33700 17678 33702
rect 17702 33700 17758 33702
rect 17782 33700 17838 33702
rect 17862 33700 17918 33702
rect 17406 32988 17408 33008
rect 17408 32988 17460 33008
rect 17460 32988 17462 33008
rect 17406 32952 17462 32988
rect 17622 32666 17678 32668
rect 17702 32666 17758 32668
rect 17782 32666 17838 32668
rect 17862 32666 17918 32668
rect 17622 32614 17648 32666
rect 17648 32614 17678 32666
rect 17702 32614 17712 32666
rect 17712 32614 17758 32666
rect 17782 32614 17828 32666
rect 17828 32614 17838 32666
rect 17862 32614 17892 32666
rect 17892 32614 17918 32666
rect 17622 32612 17678 32614
rect 17702 32612 17758 32614
rect 17782 32612 17838 32614
rect 17862 32612 17918 32614
rect 17498 32408 17554 32464
rect 17222 29688 17278 29744
rect 18050 35808 18106 35864
rect 17774 31728 17830 31784
rect 17622 31578 17678 31580
rect 17702 31578 17758 31580
rect 17782 31578 17838 31580
rect 17862 31578 17918 31580
rect 17622 31526 17648 31578
rect 17648 31526 17678 31578
rect 17702 31526 17712 31578
rect 17712 31526 17758 31578
rect 17782 31526 17828 31578
rect 17828 31526 17838 31578
rect 17862 31526 17892 31578
rect 17892 31526 17918 31578
rect 17622 31524 17678 31526
rect 17702 31524 17758 31526
rect 17782 31524 17838 31526
rect 17862 31524 17918 31526
rect 17774 31048 17830 31104
rect 17622 30490 17678 30492
rect 17702 30490 17758 30492
rect 17782 30490 17838 30492
rect 17862 30490 17918 30492
rect 17622 30438 17648 30490
rect 17648 30438 17678 30490
rect 17702 30438 17712 30490
rect 17712 30438 17758 30490
rect 17782 30438 17828 30490
rect 17828 30438 17838 30490
rect 17862 30438 17892 30490
rect 17892 30438 17918 30490
rect 17622 30436 17678 30438
rect 17702 30436 17758 30438
rect 17782 30436 17838 30438
rect 17862 30436 17918 30438
rect 17866 30252 17922 30288
rect 17866 30232 17868 30252
rect 17868 30232 17920 30252
rect 17920 30232 17922 30252
rect 17622 29402 17678 29404
rect 17702 29402 17758 29404
rect 17782 29402 17838 29404
rect 17862 29402 17918 29404
rect 17622 29350 17648 29402
rect 17648 29350 17678 29402
rect 17702 29350 17712 29402
rect 17712 29350 17758 29402
rect 17782 29350 17828 29402
rect 17828 29350 17838 29402
rect 17862 29350 17892 29402
rect 17892 29350 17918 29402
rect 17622 29348 17678 29350
rect 17702 29348 17758 29350
rect 17782 29348 17838 29350
rect 17862 29348 17918 29350
rect 17774 29044 17776 29064
rect 17776 29044 17828 29064
rect 17828 29044 17830 29064
rect 17774 29008 17830 29044
rect 17622 28314 17678 28316
rect 17702 28314 17758 28316
rect 17782 28314 17838 28316
rect 17862 28314 17918 28316
rect 17622 28262 17648 28314
rect 17648 28262 17678 28314
rect 17702 28262 17712 28314
rect 17712 28262 17758 28314
rect 17782 28262 17828 28314
rect 17828 28262 17838 28314
rect 17862 28262 17892 28314
rect 17892 28262 17918 28314
rect 17622 28260 17678 28262
rect 17702 28260 17758 28262
rect 17782 28260 17838 28262
rect 17862 28260 17918 28262
rect 17774 28076 17830 28112
rect 17774 28056 17776 28076
rect 17776 28056 17828 28076
rect 17828 28056 17830 28076
rect 17498 27648 17554 27704
rect 17038 25880 17094 25936
rect 16670 24928 16726 24984
rect 16394 24112 16450 24168
rect 15474 20848 15530 20904
rect 15382 20032 15438 20088
rect 15198 18672 15254 18728
rect 15014 18400 15070 18456
rect 15198 18264 15254 18320
rect 15106 17992 15162 18048
rect 15198 17584 15254 17640
rect 16578 21292 16580 21312
rect 16580 21292 16632 21312
rect 16632 21292 16634 21312
rect 16578 21256 16634 21292
rect 15934 19896 15990 19952
rect 15382 14864 15438 14920
rect 15198 13776 15254 13832
rect 15014 10512 15070 10568
rect 14289 6010 14345 6012
rect 14369 6010 14425 6012
rect 14449 6010 14505 6012
rect 14529 6010 14585 6012
rect 14289 5958 14315 6010
rect 14315 5958 14345 6010
rect 14369 5958 14379 6010
rect 14379 5958 14425 6010
rect 14449 5958 14495 6010
rect 14495 5958 14505 6010
rect 14529 5958 14559 6010
rect 14559 5958 14585 6010
rect 14289 5956 14345 5958
rect 14369 5956 14425 5958
rect 14449 5956 14505 5958
rect 14529 5956 14585 5958
rect 14094 5752 14150 5808
rect 14646 5772 14702 5808
rect 14646 5752 14648 5772
rect 14648 5752 14700 5772
rect 14700 5752 14702 5772
rect 14289 4922 14345 4924
rect 14369 4922 14425 4924
rect 14449 4922 14505 4924
rect 14529 4922 14585 4924
rect 14289 4870 14315 4922
rect 14315 4870 14345 4922
rect 14369 4870 14379 4922
rect 14379 4870 14425 4922
rect 14449 4870 14495 4922
rect 14495 4870 14505 4922
rect 14529 4870 14559 4922
rect 14559 4870 14585 4922
rect 14289 4868 14345 4870
rect 14369 4868 14425 4870
rect 14449 4868 14505 4870
rect 14529 4868 14585 4870
rect 14646 4664 14702 4720
rect 15198 11192 15254 11248
rect 15382 11736 15438 11792
rect 15566 15952 15622 16008
rect 15566 13912 15622 13968
rect 15658 13368 15714 13424
rect 17622 27226 17678 27228
rect 17702 27226 17758 27228
rect 17782 27226 17838 27228
rect 17862 27226 17918 27228
rect 17622 27174 17648 27226
rect 17648 27174 17678 27226
rect 17702 27174 17712 27226
rect 17712 27174 17758 27226
rect 17782 27174 17828 27226
rect 17828 27174 17838 27226
rect 17862 27174 17892 27226
rect 17892 27174 17918 27226
rect 17622 27172 17678 27174
rect 17702 27172 17758 27174
rect 17782 27172 17838 27174
rect 17862 27172 17918 27174
rect 17590 26968 17646 27024
rect 17622 26138 17678 26140
rect 17702 26138 17758 26140
rect 17782 26138 17838 26140
rect 17862 26138 17918 26140
rect 17622 26086 17648 26138
rect 17648 26086 17678 26138
rect 17702 26086 17712 26138
rect 17712 26086 17758 26138
rect 17782 26086 17828 26138
rect 17828 26086 17838 26138
rect 17862 26086 17892 26138
rect 17892 26086 17918 26138
rect 17622 26084 17678 26086
rect 17702 26084 17758 26086
rect 17782 26084 17838 26086
rect 17862 26084 17918 26086
rect 17590 25880 17646 25936
rect 17622 25050 17678 25052
rect 17702 25050 17758 25052
rect 17782 25050 17838 25052
rect 17862 25050 17918 25052
rect 17622 24998 17648 25050
rect 17648 24998 17678 25050
rect 17702 24998 17712 25050
rect 17712 24998 17758 25050
rect 17782 24998 17828 25050
rect 17828 24998 17838 25050
rect 17862 24998 17892 25050
rect 17892 24998 17918 25050
rect 17622 24996 17678 24998
rect 17702 24996 17758 24998
rect 17782 24996 17838 24998
rect 17862 24996 17918 24998
rect 17590 24792 17646 24848
rect 17130 23432 17186 23488
rect 17622 23962 17678 23964
rect 17702 23962 17758 23964
rect 17782 23962 17838 23964
rect 17862 23962 17918 23964
rect 17622 23910 17648 23962
rect 17648 23910 17678 23962
rect 17702 23910 17712 23962
rect 17712 23910 17758 23962
rect 17782 23910 17828 23962
rect 17828 23910 17838 23962
rect 17862 23910 17892 23962
rect 17892 23910 17918 23962
rect 17622 23908 17678 23910
rect 17702 23908 17758 23910
rect 17782 23908 17838 23910
rect 17862 23908 17918 23910
rect 17622 22874 17678 22876
rect 17702 22874 17758 22876
rect 17782 22874 17838 22876
rect 17862 22874 17918 22876
rect 17622 22822 17648 22874
rect 17648 22822 17678 22874
rect 17702 22822 17712 22874
rect 17712 22822 17758 22874
rect 17782 22822 17828 22874
rect 17828 22822 17838 22874
rect 17862 22822 17892 22874
rect 17892 22822 17918 22874
rect 17622 22820 17678 22822
rect 17702 22820 17758 22822
rect 17782 22820 17838 22822
rect 17862 22820 17918 22822
rect 17622 21786 17678 21788
rect 17702 21786 17758 21788
rect 17782 21786 17838 21788
rect 17862 21786 17918 21788
rect 17622 21734 17648 21786
rect 17648 21734 17678 21786
rect 17702 21734 17712 21786
rect 17712 21734 17758 21786
rect 17782 21734 17828 21786
rect 17828 21734 17838 21786
rect 17862 21734 17892 21786
rect 17892 21734 17918 21786
rect 17622 21732 17678 21734
rect 17702 21732 17758 21734
rect 17782 21732 17838 21734
rect 17862 21732 17918 21734
rect 17622 20698 17678 20700
rect 17702 20698 17758 20700
rect 17782 20698 17838 20700
rect 17862 20698 17918 20700
rect 17622 20646 17648 20698
rect 17648 20646 17678 20698
rect 17702 20646 17712 20698
rect 17712 20646 17758 20698
rect 17782 20646 17828 20698
rect 17828 20646 17838 20698
rect 17862 20646 17892 20698
rect 17892 20646 17918 20698
rect 17622 20644 17678 20646
rect 17702 20644 17758 20646
rect 17782 20644 17838 20646
rect 17862 20644 17918 20646
rect 17622 19610 17678 19612
rect 17702 19610 17758 19612
rect 17782 19610 17838 19612
rect 17862 19610 17918 19612
rect 17622 19558 17648 19610
rect 17648 19558 17678 19610
rect 17702 19558 17712 19610
rect 17712 19558 17758 19610
rect 17782 19558 17828 19610
rect 17828 19558 17838 19610
rect 17862 19558 17892 19610
rect 17892 19558 17918 19610
rect 17622 19556 17678 19558
rect 17702 19556 17758 19558
rect 17782 19556 17838 19558
rect 17862 19556 17918 19558
rect 15382 9968 15438 10024
rect 15198 9560 15254 9616
rect 15198 7112 15254 7168
rect 15566 9152 15622 9208
rect 15658 8356 15714 8392
rect 15658 8336 15660 8356
rect 15660 8336 15712 8356
rect 15712 8336 15714 8356
rect 15658 7828 15660 7848
rect 15660 7828 15712 7848
rect 15712 7828 15714 7848
rect 15658 7792 15714 7828
rect 14289 3834 14345 3836
rect 14369 3834 14425 3836
rect 14449 3834 14505 3836
rect 14529 3834 14585 3836
rect 14289 3782 14315 3834
rect 14315 3782 14345 3834
rect 14369 3782 14379 3834
rect 14379 3782 14425 3834
rect 14449 3782 14495 3834
rect 14495 3782 14505 3834
rect 14529 3782 14559 3834
rect 14559 3782 14585 3834
rect 14289 3780 14345 3782
rect 14369 3780 14425 3782
rect 14449 3780 14505 3782
rect 14529 3780 14585 3782
rect 14289 2746 14345 2748
rect 14369 2746 14425 2748
rect 14449 2746 14505 2748
rect 14529 2746 14585 2748
rect 14289 2694 14315 2746
rect 14315 2694 14345 2746
rect 14369 2694 14379 2746
rect 14379 2694 14425 2746
rect 14449 2694 14495 2746
rect 14495 2694 14505 2746
rect 14529 2694 14559 2746
rect 14559 2694 14585 2746
rect 14289 2692 14345 2694
rect 14369 2692 14425 2694
rect 14449 2692 14505 2694
rect 14529 2692 14585 2694
rect 10956 2202 11012 2204
rect 11036 2202 11092 2204
rect 11116 2202 11172 2204
rect 11196 2202 11252 2204
rect 10956 2150 10982 2202
rect 10982 2150 11012 2202
rect 11036 2150 11046 2202
rect 11046 2150 11092 2202
rect 11116 2150 11162 2202
rect 11162 2150 11172 2202
rect 11196 2150 11226 2202
rect 11226 2150 11252 2202
rect 10956 2148 11012 2150
rect 11036 2148 11092 2150
rect 11116 2148 11172 2150
rect 11196 2148 11252 2150
rect 9494 1400 9550 1456
rect 16394 15408 16450 15464
rect 16026 15272 16082 15328
rect 16210 14592 16266 14648
rect 17622 18522 17678 18524
rect 17702 18522 17758 18524
rect 17782 18522 17838 18524
rect 17862 18522 17918 18524
rect 17622 18470 17648 18522
rect 17648 18470 17678 18522
rect 17702 18470 17712 18522
rect 17712 18470 17758 18522
rect 17782 18470 17828 18522
rect 17828 18470 17838 18522
rect 17862 18470 17892 18522
rect 17892 18470 17918 18522
rect 17622 18468 17678 18470
rect 17702 18468 17758 18470
rect 17782 18468 17838 18470
rect 17862 18468 17918 18470
rect 16854 18400 16910 18456
rect 17622 17434 17678 17436
rect 17702 17434 17758 17436
rect 17782 17434 17838 17436
rect 17862 17434 17918 17436
rect 17622 17382 17648 17434
rect 17648 17382 17678 17434
rect 17702 17382 17712 17434
rect 17712 17382 17758 17434
rect 17782 17382 17828 17434
rect 17828 17382 17838 17434
rect 17862 17382 17892 17434
rect 17892 17382 17918 17434
rect 17622 17380 17678 17382
rect 17702 17380 17758 17382
rect 17782 17380 17838 17382
rect 17862 17380 17918 17382
rect 17622 16346 17678 16348
rect 17702 16346 17758 16348
rect 17782 16346 17838 16348
rect 17862 16346 17918 16348
rect 17622 16294 17648 16346
rect 17648 16294 17678 16346
rect 17702 16294 17712 16346
rect 17712 16294 17758 16346
rect 17782 16294 17828 16346
rect 17828 16294 17838 16346
rect 17862 16294 17892 16346
rect 17892 16294 17918 16346
rect 17622 16292 17678 16294
rect 17702 16292 17758 16294
rect 17782 16292 17838 16294
rect 17862 16292 17918 16294
rect 16946 15816 17002 15872
rect 16118 12824 16174 12880
rect 16394 12552 16450 12608
rect 16026 7792 16082 7848
rect 15934 6704 15990 6760
rect 16026 5616 16082 5672
rect 16854 14320 16910 14376
rect 16762 13232 16818 13288
rect 16762 11872 16818 11928
rect 17622 15258 17678 15260
rect 17702 15258 17758 15260
rect 17782 15258 17838 15260
rect 17862 15258 17918 15260
rect 17622 15206 17648 15258
rect 17648 15206 17678 15258
rect 17702 15206 17712 15258
rect 17712 15206 17758 15258
rect 17782 15206 17828 15258
rect 17828 15206 17838 15258
rect 17862 15206 17892 15258
rect 17892 15206 17918 15258
rect 17622 15204 17678 15206
rect 17702 15204 17758 15206
rect 17782 15204 17838 15206
rect 17862 15204 17918 15206
rect 17622 14170 17678 14172
rect 17702 14170 17758 14172
rect 17782 14170 17838 14172
rect 17862 14170 17918 14172
rect 17622 14118 17648 14170
rect 17648 14118 17678 14170
rect 17702 14118 17712 14170
rect 17712 14118 17758 14170
rect 17782 14118 17828 14170
rect 17828 14118 17838 14170
rect 17862 14118 17892 14170
rect 17892 14118 17918 14170
rect 17622 14116 17678 14118
rect 17702 14116 17758 14118
rect 17782 14116 17838 14118
rect 17862 14116 17918 14118
rect 16302 6024 16358 6080
rect 16118 5072 16174 5128
rect 15566 3032 15622 3088
rect 16394 3712 16450 3768
rect 17314 10104 17370 10160
rect 16670 6024 16726 6080
rect 17622 13082 17678 13084
rect 17702 13082 17758 13084
rect 17782 13082 17838 13084
rect 17862 13082 17918 13084
rect 17622 13030 17648 13082
rect 17648 13030 17678 13082
rect 17702 13030 17712 13082
rect 17712 13030 17758 13082
rect 17782 13030 17828 13082
rect 17828 13030 17838 13082
rect 17862 13030 17892 13082
rect 17892 13030 17918 13082
rect 17622 13028 17678 13030
rect 17702 13028 17758 13030
rect 17782 13028 17838 13030
rect 17862 13028 17918 13030
rect 17622 11994 17678 11996
rect 17702 11994 17758 11996
rect 17782 11994 17838 11996
rect 17862 11994 17918 11996
rect 17622 11942 17648 11994
rect 17648 11942 17678 11994
rect 17702 11942 17712 11994
rect 17712 11942 17758 11994
rect 17782 11942 17828 11994
rect 17828 11942 17838 11994
rect 17862 11942 17892 11994
rect 17892 11942 17918 11994
rect 17622 11940 17678 11942
rect 17702 11940 17758 11942
rect 17782 11940 17838 11942
rect 17862 11940 17918 11942
rect 17622 10906 17678 10908
rect 17702 10906 17758 10908
rect 17782 10906 17838 10908
rect 17862 10906 17918 10908
rect 17622 10854 17648 10906
rect 17648 10854 17678 10906
rect 17702 10854 17712 10906
rect 17712 10854 17758 10906
rect 17782 10854 17828 10906
rect 17828 10854 17838 10906
rect 17862 10854 17892 10906
rect 17892 10854 17918 10906
rect 17622 10852 17678 10854
rect 17702 10852 17758 10854
rect 17782 10852 17838 10854
rect 17862 10852 17918 10854
rect 17622 9818 17678 9820
rect 17702 9818 17758 9820
rect 17782 9818 17838 9820
rect 17862 9818 17918 9820
rect 17622 9766 17648 9818
rect 17648 9766 17678 9818
rect 17702 9766 17712 9818
rect 17712 9766 17758 9818
rect 17782 9766 17828 9818
rect 17828 9766 17838 9818
rect 17862 9766 17892 9818
rect 17892 9766 17918 9818
rect 17622 9764 17678 9766
rect 17702 9764 17758 9766
rect 17782 9764 17838 9766
rect 17862 9764 17918 9766
rect 17622 8730 17678 8732
rect 17702 8730 17758 8732
rect 17782 8730 17838 8732
rect 17862 8730 17918 8732
rect 17622 8678 17648 8730
rect 17648 8678 17678 8730
rect 17702 8678 17712 8730
rect 17712 8678 17758 8730
rect 17782 8678 17828 8730
rect 17828 8678 17838 8730
rect 17862 8678 17892 8730
rect 17892 8678 17918 8730
rect 17622 8676 17678 8678
rect 17702 8676 17758 8678
rect 17782 8676 17838 8678
rect 17862 8676 17918 8678
rect 17622 7642 17678 7644
rect 17702 7642 17758 7644
rect 17782 7642 17838 7644
rect 17862 7642 17918 7644
rect 17622 7590 17648 7642
rect 17648 7590 17678 7642
rect 17702 7590 17712 7642
rect 17712 7590 17758 7642
rect 17782 7590 17828 7642
rect 17828 7590 17838 7642
rect 17862 7590 17892 7642
rect 17892 7590 17918 7642
rect 17622 7588 17678 7590
rect 17702 7588 17758 7590
rect 17782 7588 17838 7590
rect 17862 7588 17918 7590
rect 17406 6724 17462 6760
rect 17406 6704 17408 6724
rect 17408 6704 17460 6724
rect 17460 6704 17462 6724
rect 17622 6554 17678 6556
rect 17702 6554 17758 6556
rect 17782 6554 17838 6556
rect 17862 6554 17918 6556
rect 17622 6502 17648 6554
rect 17648 6502 17678 6554
rect 17702 6502 17712 6554
rect 17712 6502 17758 6554
rect 17782 6502 17828 6554
rect 17828 6502 17838 6554
rect 17862 6502 17892 6554
rect 17892 6502 17918 6554
rect 17622 6500 17678 6502
rect 17702 6500 17758 6502
rect 17782 6500 17838 6502
rect 17862 6500 17918 6502
rect 17622 5466 17678 5468
rect 17702 5466 17758 5468
rect 17782 5466 17838 5468
rect 17862 5466 17918 5468
rect 17622 5414 17648 5466
rect 17648 5414 17678 5466
rect 17702 5414 17712 5466
rect 17712 5414 17758 5466
rect 17782 5414 17828 5466
rect 17828 5414 17838 5466
rect 17862 5414 17892 5466
rect 17892 5414 17918 5466
rect 17622 5412 17678 5414
rect 17702 5412 17758 5414
rect 17782 5412 17838 5414
rect 17862 5412 17918 5414
rect 17038 4528 17094 4584
rect 17622 4378 17678 4380
rect 17702 4378 17758 4380
rect 17782 4378 17838 4380
rect 17862 4378 17918 4380
rect 17622 4326 17648 4378
rect 17648 4326 17678 4378
rect 17702 4326 17712 4378
rect 17712 4326 17758 4378
rect 17782 4326 17828 4378
rect 17828 4326 17838 4378
rect 17862 4326 17892 4378
rect 17892 4326 17918 4378
rect 17622 4324 17678 4326
rect 17702 4324 17758 4326
rect 17782 4324 17838 4326
rect 17862 4324 17918 4326
rect 17622 3290 17678 3292
rect 17702 3290 17758 3292
rect 17782 3290 17838 3292
rect 17862 3290 17918 3292
rect 17622 3238 17648 3290
rect 17648 3238 17678 3290
rect 17702 3238 17712 3290
rect 17712 3238 17758 3290
rect 17782 3238 17828 3290
rect 17828 3238 17838 3290
rect 17862 3238 17892 3290
rect 17892 3238 17918 3290
rect 17622 3236 17678 3238
rect 17702 3236 17758 3238
rect 17782 3236 17838 3238
rect 17862 3236 17918 3238
rect 16486 2352 16542 2408
rect 17622 2202 17678 2204
rect 17702 2202 17758 2204
rect 17782 2202 17838 2204
rect 17862 2202 17918 2204
rect 17622 2150 17648 2202
rect 17648 2150 17678 2202
rect 17702 2150 17712 2202
rect 17712 2150 17758 2202
rect 17782 2150 17828 2202
rect 17828 2150 17838 2202
rect 17862 2150 17892 2202
rect 17892 2150 17918 2202
rect 17622 2148 17678 2150
rect 17702 2148 17758 2150
rect 17782 2148 17838 2150
rect 17862 2148 17918 2150
rect 16302 1672 16358 1728
rect 15198 992 15254 1048
rect 9310 312 9366 368
rect 11334 312 11390 368
<< metal3 >>
rect 5390 79596 5396 79660
rect 5460 79658 5466 79660
rect 5460 79598 19442 79658
rect 5460 79596 5466 79598
rect 0 79522 480 79552
rect 3601 79522 3667 79525
rect 0 79520 3667 79522
rect 0 79464 3606 79520
rect 3662 79464 3667 79520
rect 0 79462 3667 79464
rect 19382 79522 19442 79598
rect 19520 79522 20000 79552
rect 19382 79462 20000 79522
rect 0 79432 480 79462
rect 3601 79459 3667 79462
rect 19520 79432 20000 79462
rect 16021 78842 16087 78845
rect 19520 78842 20000 78872
rect 16021 78840 20000 78842
rect 16021 78784 16026 78840
rect 16082 78784 20000 78840
rect 16021 78782 20000 78784
rect 16021 78779 16087 78782
rect 19520 78752 20000 78782
rect 0 78706 480 78736
rect 3785 78706 3851 78709
rect 0 78704 3851 78706
rect 0 78648 3790 78704
rect 3846 78648 3851 78704
rect 0 78646 3851 78648
rect 0 78616 480 78646
rect 3785 78643 3851 78646
rect 15929 78162 15995 78165
rect 19520 78162 20000 78192
rect 15929 78160 20000 78162
rect 15929 78104 15934 78160
rect 15990 78104 20000 78160
rect 15929 78102 20000 78104
rect 15929 78099 15995 78102
rect 19520 78072 20000 78102
rect 0 77890 480 77920
rect 2865 77890 2931 77893
rect 0 77888 2931 77890
rect 0 77832 2870 77888
rect 2926 77832 2931 77888
rect 0 77830 2931 77832
rect 0 77800 480 77830
rect 2865 77827 2931 77830
rect 7610 77824 7930 77825
rect 7610 77760 7618 77824
rect 7682 77760 7698 77824
rect 7762 77760 7778 77824
rect 7842 77760 7858 77824
rect 7922 77760 7930 77824
rect 7610 77759 7930 77760
rect 14277 77824 14597 77825
rect 14277 77760 14285 77824
rect 14349 77760 14365 77824
rect 14429 77760 14445 77824
rect 14509 77760 14525 77824
rect 14589 77760 14597 77824
rect 14277 77759 14597 77760
rect 14958 77420 14964 77484
rect 15028 77482 15034 77484
rect 19520 77482 20000 77512
rect 15028 77422 20000 77482
rect 15028 77420 15034 77422
rect 19520 77392 20000 77422
rect 4277 77280 4597 77281
rect 4277 77216 4285 77280
rect 4349 77216 4365 77280
rect 4429 77216 4445 77280
rect 4509 77216 4525 77280
rect 4589 77216 4597 77280
rect 4277 77215 4597 77216
rect 10944 77280 11264 77281
rect 10944 77216 10952 77280
rect 11016 77216 11032 77280
rect 11096 77216 11112 77280
rect 11176 77216 11192 77280
rect 11256 77216 11264 77280
rect 10944 77215 11264 77216
rect 17610 77280 17930 77281
rect 17610 77216 17618 77280
rect 17682 77216 17698 77280
rect 17762 77216 17778 77280
rect 17842 77216 17858 77280
rect 17922 77216 17930 77280
rect 17610 77215 17930 77216
rect 0 77074 480 77104
rect 2129 77074 2195 77077
rect 0 77072 2195 77074
rect 0 77016 2134 77072
rect 2190 77016 2195 77072
rect 0 77014 2195 77016
rect 0 76984 480 77014
rect 2129 77011 2195 77014
rect 19520 76802 20000 76832
rect 15886 76742 20000 76802
rect 7610 76736 7930 76737
rect 7610 76672 7618 76736
rect 7682 76672 7698 76736
rect 7762 76672 7778 76736
rect 7842 76672 7858 76736
rect 7922 76672 7930 76736
rect 7610 76671 7930 76672
rect 14277 76736 14597 76737
rect 14277 76672 14285 76736
rect 14349 76672 14365 76736
rect 14429 76672 14445 76736
rect 14509 76672 14525 76736
rect 14589 76672 14597 76736
rect 14277 76671 14597 76672
rect 5206 76332 5212 76396
rect 5276 76394 5282 76396
rect 15886 76394 15946 76742
rect 19520 76712 20000 76742
rect 5276 76334 15946 76394
rect 5276 76332 5282 76334
rect 0 76258 480 76288
rect 4061 76258 4127 76261
rect 0 76256 4127 76258
rect 0 76200 4066 76256
rect 4122 76200 4127 76256
rect 0 76198 4127 76200
rect 0 76168 480 76198
rect 4061 76195 4127 76198
rect 4277 76192 4597 76193
rect 4277 76128 4285 76192
rect 4349 76128 4365 76192
rect 4429 76128 4445 76192
rect 4509 76128 4525 76192
rect 4589 76128 4597 76192
rect 4277 76127 4597 76128
rect 10944 76192 11264 76193
rect 10944 76128 10952 76192
rect 11016 76128 11032 76192
rect 11096 76128 11112 76192
rect 11176 76128 11192 76192
rect 11256 76128 11264 76192
rect 10944 76127 11264 76128
rect 17610 76192 17930 76193
rect 17610 76128 17618 76192
rect 17682 76128 17698 76192
rect 17762 76128 17778 76192
rect 17842 76128 17858 76192
rect 17922 76128 17930 76192
rect 17610 76127 17930 76128
rect 19520 76122 20000 76152
rect 18094 76062 20000 76122
rect 4838 75924 4844 75988
rect 4908 75986 4914 75988
rect 18094 75986 18154 76062
rect 19520 76032 20000 76062
rect 4908 75926 18154 75986
rect 4908 75924 4914 75926
rect 7610 75648 7930 75649
rect 7610 75584 7618 75648
rect 7682 75584 7698 75648
rect 7762 75584 7778 75648
rect 7842 75584 7858 75648
rect 7922 75584 7930 75648
rect 7610 75583 7930 75584
rect 14277 75648 14597 75649
rect 14277 75584 14285 75648
rect 14349 75584 14365 75648
rect 14429 75584 14445 75648
rect 14509 75584 14525 75648
rect 14589 75584 14597 75648
rect 14277 75583 14597 75584
rect 0 75442 480 75472
rect 3417 75442 3483 75445
rect 0 75440 3483 75442
rect 0 75384 3422 75440
rect 3478 75384 3483 75440
rect 0 75382 3483 75384
rect 0 75352 480 75382
rect 3417 75379 3483 75382
rect 5022 75380 5028 75444
rect 5092 75442 5098 75444
rect 19520 75442 20000 75472
rect 5092 75382 20000 75442
rect 5092 75380 5098 75382
rect 19520 75352 20000 75382
rect 4889 75306 4955 75309
rect 7005 75306 7071 75309
rect 4889 75304 7071 75306
rect 4889 75248 4894 75304
rect 4950 75248 7010 75304
rect 7066 75248 7071 75304
rect 4889 75246 7071 75248
rect 4889 75243 4955 75246
rect 7005 75243 7071 75246
rect 4277 75104 4597 75105
rect 4277 75040 4285 75104
rect 4349 75040 4365 75104
rect 4429 75040 4445 75104
rect 4509 75040 4525 75104
rect 4589 75040 4597 75104
rect 4277 75039 4597 75040
rect 10944 75104 11264 75105
rect 10944 75040 10952 75104
rect 11016 75040 11032 75104
rect 11096 75040 11112 75104
rect 11176 75040 11192 75104
rect 11256 75040 11264 75104
rect 10944 75039 11264 75040
rect 17610 75104 17930 75105
rect 17610 75040 17618 75104
rect 17682 75040 17698 75104
rect 17762 75040 17778 75104
rect 17842 75040 17858 75104
rect 17922 75040 17930 75104
rect 17610 75039 17930 75040
rect 2446 74700 2452 74764
rect 2516 74762 2522 74764
rect 19520 74762 20000 74792
rect 2516 74702 20000 74762
rect 2516 74700 2522 74702
rect 19520 74672 20000 74702
rect 0 74626 480 74656
rect 4613 74626 4679 74629
rect 0 74624 4679 74626
rect 0 74568 4618 74624
rect 4674 74568 4679 74624
rect 0 74566 4679 74568
rect 0 74536 480 74566
rect 4613 74563 4679 74566
rect 7610 74560 7930 74561
rect 7610 74496 7618 74560
rect 7682 74496 7698 74560
rect 7762 74496 7778 74560
rect 7842 74496 7858 74560
rect 7922 74496 7930 74560
rect 7610 74495 7930 74496
rect 14277 74560 14597 74561
rect 14277 74496 14285 74560
rect 14349 74496 14365 74560
rect 14429 74496 14445 74560
rect 14509 74496 14525 74560
rect 14589 74496 14597 74560
rect 14277 74495 14597 74496
rect 19520 74082 20000 74112
rect 18094 74022 20000 74082
rect 4277 74016 4597 74017
rect 4277 73952 4285 74016
rect 4349 73952 4365 74016
rect 4429 73952 4445 74016
rect 4509 73952 4525 74016
rect 4589 73952 4597 74016
rect 4277 73951 4597 73952
rect 10944 74016 11264 74017
rect 10944 73952 10952 74016
rect 11016 73952 11032 74016
rect 11096 73952 11112 74016
rect 11176 73952 11192 74016
rect 11256 73952 11264 74016
rect 10944 73951 11264 73952
rect 17610 74016 17930 74017
rect 17610 73952 17618 74016
rect 17682 73952 17698 74016
rect 17762 73952 17778 74016
rect 17842 73952 17858 74016
rect 17922 73952 17930 74016
rect 17610 73951 17930 73952
rect 0 73810 480 73840
rect 4797 73810 4863 73813
rect 0 73808 4863 73810
rect 0 73752 4802 73808
rect 4858 73752 4863 73808
rect 0 73750 4863 73752
rect 0 73720 480 73750
rect 4797 73747 4863 73750
rect 7230 73748 7236 73812
rect 7300 73810 7306 73812
rect 18094 73810 18154 74022
rect 19520 73992 20000 74022
rect 7300 73750 18154 73810
rect 7300 73748 7306 73750
rect 5073 73674 5139 73677
rect 7005 73674 7071 73677
rect 5073 73672 7071 73674
rect 5073 73616 5078 73672
rect 5134 73616 7010 73672
rect 7066 73616 7071 73672
rect 5073 73614 7071 73616
rect 5073 73611 5139 73614
rect 7005 73611 7071 73614
rect 7610 73472 7930 73473
rect 7610 73408 7618 73472
rect 7682 73408 7698 73472
rect 7762 73408 7778 73472
rect 7842 73408 7858 73472
rect 7922 73408 7930 73472
rect 7610 73407 7930 73408
rect 14277 73472 14597 73473
rect 14277 73408 14285 73472
rect 14349 73408 14365 73472
rect 14429 73408 14445 73472
rect 14509 73408 14525 73472
rect 14589 73408 14597 73472
rect 14277 73407 14597 73408
rect 3877 73402 3943 73405
rect 5993 73402 6059 73405
rect 3877 73400 6059 73402
rect 3877 73344 3882 73400
rect 3938 73344 5998 73400
rect 6054 73344 6059 73400
rect 3877 73342 6059 73344
rect 3877 73339 3943 73342
rect 5993 73339 6059 73342
rect 8477 73402 8543 73405
rect 19520 73402 20000 73432
rect 8477 73400 10978 73402
rect 8477 73344 8482 73400
rect 8538 73344 10978 73400
rect 8477 73342 10978 73344
rect 8477 73339 8543 73342
rect 4337 73266 4403 73269
rect 6913 73266 6979 73269
rect 4337 73264 6979 73266
rect 4337 73208 4342 73264
rect 4398 73208 6918 73264
rect 6974 73208 6979 73264
rect 4337 73206 6979 73208
rect 4337 73203 4403 73206
rect 6913 73203 6979 73206
rect 10685 73268 10751 73269
rect 10685 73264 10732 73268
rect 10796 73266 10802 73268
rect 10918 73266 10978 73342
rect 15886 73342 20000 73402
rect 15886 73266 15946 73342
rect 19520 73312 20000 73342
rect 10685 73208 10690 73264
rect 10685 73204 10732 73208
rect 10796 73206 10842 73266
rect 10918 73206 15946 73266
rect 10796 73204 10802 73206
rect 10685 73203 10751 73204
rect 0 73130 480 73160
rect 4245 73130 4311 73133
rect 0 73128 4311 73130
rect 0 73072 4250 73128
rect 4306 73072 4311 73128
rect 0 73070 4311 73072
rect 0 73040 480 73070
rect 4245 73067 4311 73070
rect 4277 72928 4597 72929
rect 4277 72864 4285 72928
rect 4349 72864 4365 72928
rect 4429 72864 4445 72928
rect 4509 72864 4525 72928
rect 4589 72864 4597 72928
rect 4277 72863 4597 72864
rect 10944 72928 11264 72929
rect 10944 72864 10952 72928
rect 11016 72864 11032 72928
rect 11096 72864 11112 72928
rect 11176 72864 11192 72928
rect 11256 72864 11264 72928
rect 10944 72863 11264 72864
rect 17610 72928 17930 72929
rect 17610 72864 17618 72928
rect 17682 72864 17698 72928
rect 17762 72864 17778 72928
rect 17842 72864 17858 72928
rect 17922 72864 17930 72928
rect 17610 72863 17930 72864
rect 16297 72722 16363 72725
rect 19520 72722 20000 72752
rect 16297 72720 20000 72722
rect 16297 72664 16302 72720
rect 16358 72664 20000 72720
rect 16297 72662 20000 72664
rect 16297 72659 16363 72662
rect 19520 72632 20000 72662
rect 11789 72586 11855 72589
rect 17493 72586 17559 72589
rect 11789 72584 17559 72586
rect 11789 72528 11794 72584
rect 11850 72528 17498 72584
rect 17554 72528 17559 72584
rect 11789 72526 17559 72528
rect 11789 72523 11855 72526
rect 17493 72523 17559 72526
rect 7610 72384 7930 72385
rect 0 72314 480 72344
rect 7610 72320 7618 72384
rect 7682 72320 7698 72384
rect 7762 72320 7778 72384
rect 7842 72320 7858 72384
rect 7922 72320 7930 72384
rect 7610 72319 7930 72320
rect 14277 72384 14597 72385
rect 14277 72320 14285 72384
rect 14349 72320 14365 72384
rect 14429 72320 14445 72384
rect 14509 72320 14525 72384
rect 14589 72320 14597 72384
rect 14277 72319 14597 72320
rect 2865 72314 2931 72317
rect 0 72312 2931 72314
rect 0 72256 2870 72312
rect 2926 72256 2931 72312
rect 0 72254 2931 72256
rect 0 72224 480 72254
rect 2865 72251 2931 72254
rect 7097 72178 7163 72181
rect 10317 72178 10383 72181
rect 7097 72176 10383 72178
rect 7097 72120 7102 72176
rect 7158 72120 10322 72176
rect 10378 72120 10383 72176
rect 7097 72118 10383 72120
rect 7097 72115 7163 72118
rect 10317 72115 10383 72118
rect 9397 72042 9463 72045
rect 19520 72042 20000 72072
rect 9397 72040 20000 72042
rect 9397 71984 9402 72040
rect 9458 71984 20000 72040
rect 9397 71982 20000 71984
rect 9397 71979 9463 71982
rect 19520 71952 20000 71982
rect 4277 71840 4597 71841
rect 4277 71776 4285 71840
rect 4349 71776 4365 71840
rect 4429 71776 4445 71840
rect 4509 71776 4525 71840
rect 4589 71776 4597 71840
rect 4277 71775 4597 71776
rect 10944 71840 11264 71841
rect 10944 71776 10952 71840
rect 11016 71776 11032 71840
rect 11096 71776 11112 71840
rect 11176 71776 11192 71840
rect 11256 71776 11264 71840
rect 10944 71775 11264 71776
rect 17610 71840 17930 71841
rect 17610 71776 17618 71840
rect 17682 71776 17698 71840
rect 17762 71776 17778 71840
rect 17842 71776 17858 71840
rect 17922 71776 17930 71840
rect 17610 71775 17930 71776
rect 0 71498 480 71528
rect 4102 71498 4108 71500
rect 0 71438 4108 71498
rect 0 71408 480 71438
rect 4102 71436 4108 71438
rect 4172 71436 4178 71500
rect 3693 71362 3759 71365
rect 7189 71362 7255 71365
rect 3693 71360 7255 71362
rect 3693 71304 3698 71360
rect 3754 71304 7194 71360
rect 7250 71304 7255 71360
rect 3693 71302 7255 71304
rect 3693 71299 3759 71302
rect 7189 71299 7255 71302
rect 16614 71300 16620 71364
rect 16684 71362 16690 71364
rect 19520 71362 20000 71392
rect 16684 71302 20000 71362
rect 16684 71300 16690 71302
rect 7610 71296 7930 71297
rect 7610 71232 7618 71296
rect 7682 71232 7698 71296
rect 7762 71232 7778 71296
rect 7842 71232 7858 71296
rect 7922 71232 7930 71296
rect 7610 71231 7930 71232
rect 14277 71296 14597 71297
rect 14277 71232 14285 71296
rect 14349 71232 14365 71296
rect 14429 71232 14445 71296
rect 14509 71232 14525 71296
rect 14589 71232 14597 71296
rect 19520 71272 20000 71302
rect 14277 71231 14597 71232
rect 8845 71090 8911 71093
rect 8845 71088 18154 71090
rect 8845 71032 8850 71088
rect 8906 71032 18154 71088
rect 8845 71030 18154 71032
rect 8845 71027 8911 71030
rect 4277 70752 4597 70753
rect 0 70682 480 70712
rect 4277 70688 4285 70752
rect 4349 70688 4365 70752
rect 4429 70688 4445 70752
rect 4509 70688 4525 70752
rect 4589 70688 4597 70752
rect 4277 70687 4597 70688
rect 10944 70752 11264 70753
rect 10944 70688 10952 70752
rect 11016 70688 11032 70752
rect 11096 70688 11112 70752
rect 11176 70688 11192 70752
rect 11256 70688 11264 70752
rect 10944 70687 11264 70688
rect 17610 70752 17930 70753
rect 17610 70688 17618 70752
rect 17682 70688 17698 70752
rect 17762 70688 17778 70752
rect 17842 70688 17858 70752
rect 17922 70688 17930 70752
rect 17610 70687 17930 70688
rect 9581 70684 9647 70685
rect 0 70622 3802 70682
rect 0 70592 480 70622
rect 3742 70546 3802 70622
rect 9581 70680 9628 70684
rect 9692 70682 9698 70684
rect 18094 70682 18154 71030
rect 19520 70682 20000 70712
rect 9581 70624 9586 70680
rect 9581 70620 9628 70624
rect 9692 70622 9738 70682
rect 18094 70622 20000 70682
rect 9692 70620 9698 70622
rect 9581 70619 9647 70620
rect 19520 70592 20000 70622
rect 4654 70546 4660 70548
rect 3742 70486 4660 70546
rect 4654 70484 4660 70486
rect 4724 70484 4730 70548
rect 4705 70410 4771 70413
rect 7465 70410 7531 70413
rect 4705 70408 7531 70410
rect 4705 70352 4710 70408
rect 4766 70352 7470 70408
rect 7526 70352 7531 70408
rect 4705 70350 7531 70352
rect 4705 70347 4771 70350
rect 7465 70347 7531 70350
rect 7833 70410 7899 70413
rect 8150 70410 8156 70412
rect 7833 70408 8156 70410
rect 7833 70352 7838 70408
rect 7894 70352 8156 70408
rect 7833 70350 8156 70352
rect 7833 70347 7899 70350
rect 8150 70348 8156 70350
rect 8220 70348 8226 70412
rect 8385 70410 8451 70413
rect 9673 70410 9739 70413
rect 8385 70408 9739 70410
rect 8385 70352 8390 70408
rect 8446 70352 9678 70408
rect 9734 70352 9739 70408
rect 8385 70350 9739 70352
rect 8385 70347 8451 70350
rect 9673 70347 9739 70350
rect 11605 70410 11671 70413
rect 11605 70408 11714 70410
rect 11605 70352 11610 70408
rect 11666 70352 11714 70408
rect 11605 70347 11714 70352
rect 8201 70274 8267 70277
rect 9765 70274 9831 70277
rect 8201 70272 9831 70274
rect 8201 70216 8206 70272
rect 8262 70216 9770 70272
rect 9826 70216 9831 70272
rect 8201 70214 9831 70216
rect 8201 70211 8267 70214
rect 9765 70211 9831 70214
rect 7610 70208 7930 70209
rect 7610 70144 7618 70208
rect 7682 70144 7698 70208
rect 7762 70144 7778 70208
rect 7842 70144 7858 70208
rect 7922 70144 7930 70208
rect 7610 70143 7930 70144
rect 11513 70138 11579 70141
rect 11654 70138 11714 70347
rect 14277 70208 14597 70209
rect 14277 70144 14285 70208
rect 14349 70144 14365 70208
rect 14429 70144 14445 70208
rect 14509 70144 14525 70208
rect 14589 70144 14597 70208
rect 14277 70143 14597 70144
rect 11513 70136 11714 70138
rect 11513 70080 11518 70136
rect 11574 70080 11714 70136
rect 11513 70078 11714 70080
rect 11513 70075 11579 70078
rect 9581 70002 9647 70005
rect 11973 70002 12039 70005
rect 19520 70002 20000 70032
rect 9581 70000 12039 70002
rect 9581 69944 9586 70000
rect 9642 69944 11978 70000
rect 12034 69944 12039 70000
rect 9581 69942 12039 69944
rect 9581 69939 9647 69942
rect 11973 69939 12039 69942
rect 19382 69942 20000 70002
rect 0 69866 480 69896
rect 3969 69866 4035 69869
rect 0 69864 4035 69866
rect 0 69808 3974 69864
rect 4030 69808 4035 69864
rect 0 69806 4035 69808
rect 0 69776 480 69806
rect 3969 69803 4035 69806
rect 6862 69668 6868 69732
rect 6932 69730 6938 69732
rect 8477 69730 8543 69733
rect 6932 69728 8543 69730
rect 6932 69672 8482 69728
rect 8538 69672 8543 69728
rect 6932 69670 8543 69672
rect 6932 69668 6938 69670
rect 8477 69667 8543 69670
rect 4277 69664 4597 69665
rect 4277 69600 4285 69664
rect 4349 69600 4365 69664
rect 4429 69600 4445 69664
rect 4509 69600 4525 69664
rect 4589 69600 4597 69664
rect 4277 69599 4597 69600
rect 10944 69664 11264 69665
rect 10944 69600 10952 69664
rect 11016 69600 11032 69664
rect 11096 69600 11112 69664
rect 11176 69600 11192 69664
rect 11256 69600 11264 69664
rect 10944 69599 11264 69600
rect 17610 69664 17930 69665
rect 17610 69600 17618 69664
rect 17682 69600 17698 69664
rect 17762 69600 17778 69664
rect 17842 69600 17858 69664
rect 17922 69600 17930 69664
rect 17610 69599 17930 69600
rect 4705 69594 4771 69597
rect 4705 69592 10794 69594
rect 4705 69536 4710 69592
rect 4766 69536 10794 69592
rect 4705 69534 10794 69536
rect 4705 69531 4771 69534
rect 2865 69458 2931 69461
rect 5809 69458 5875 69461
rect 2865 69456 5875 69458
rect 2865 69400 2870 69456
rect 2926 69400 5814 69456
rect 5870 69400 5875 69456
rect 2865 69398 5875 69400
rect 2865 69395 2931 69398
rect 5809 69395 5875 69398
rect 6637 69458 6703 69461
rect 8385 69458 8451 69461
rect 6637 69456 8451 69458
rect 6637 69400 6642 69456
rect 6698 69400 8390 69456
rect 8446 69400 8451 69456
rect 6637 69398 8451 69400
rect 10734 69458 10794 69534
rect 19382 69458 19442 69942
rect 19520 69912 20000 69942
rect 10734 69398 19442 69458
rect 6637 69395 6703 69398
rect 8385 69395 8451 69398
rect 2957 69322 3023 69325
rect 9397 69322 9463 69325
rect 2957 69320 9463 69322
rect 2957 69264 2962 69320
rect 3018 69264 9402 69320
rect 9458 69264 9463 69320
rect 2957 69262 9463 69264
rect 2957 69259 3023 69262
rect 9397 69259 9463 69262
rect 9765 69322 9831 69325
rect 19520 69322 20000 69352
rect 9765 69320 20000 69322
rect 9765 69264 9770 69320
rect 9826 69264 20000 69320
rect 9765 69262 20000 69264
rect 9765 69259 9831 69262
rect 19520 69232 20000 69262
rect 3049 69186 3115 69189
rect 5349 69186 5415 69189
rect 3049 69184 5415 69186
rect 3049 69128 3054 69184
rect 3110 69128 5354 69184
rect 5410 69128 5415 69184
rect 3049 69126 5415 69128
rect 3049 69123 3115 69126
rect 5349 69123 5415 69126
rect 8201 69186 8267 69189
rect 9397 69186 9463 69189
rect 8201 69184 9463 69186
rect 8201 69128 8206 69184
rect 8262 69128 9402 69184
rect 9458 69128 9463 69184
rect 8201 69126 9463 69128
rect 8201 69123 8267 69126
rect 9397 69123 9463 69126
rect 7610 69120 7930 69121
rect 0 69050 480 69080
rect 7610 69056 7618 69120
rect 7682 69056 7698 69120
rect 7762 69056 7778 69120
rect 7842 69056 7858 69120
rect 7922 69056 7930 69120
rect 7610 69055 7930 69056
rect 14277 69120 14597 69121
rect 14277 69056 14285 69120
rect 14349 69056 14365 69120
rect 14429 69056 14445 69120
rect 14509 69056 14525 69120
rect 14589 69056 14597 69120
rect 14277 69055 14597 69056
rect 2037 69050 2103 69053
rect 0 69048 2103 69050
rect 0 68992 2042 69048
rect 2098 68992 2103 69048
rect 0 68990 2103 68992
rect 0 68960 480 68990
rect 2037 68987 2103 68990
rect 3601 69050 3667 69053
rect 7097 69050 7163 69053
rect 11973 69052 12039 69053
rect 11973 69050 12020 69052
rect 3601 69048 7163 69050
rect 3601 68992 3606 69048
rect 3662 68992 7102 69048
rect 7158 68992 7163 69048
rect 3601 68990 7163 68992
rect 11928 69048 12020 69050
rect 11928 68992 11978 69048
rect 11928 68990 12020 68992
rect 3601 68987 3667 68990
rect 7097 68987 7163 68990
rect 11973 68988 12020 68990
rect 12084 68988 12090 69052
rect 11973 68987 12039 68988
rect 8017 68914 8083 68917
rect 10041 68914 10107 68917
rect 8017 68912 10107 68914
rect 8017 68856 8022 68912
rect 8078 68856 10046 68912
rect 10102 68856 10107 68912
rect 8017 68854 10107 68856
rect 8017 68851 8083 68854
rect 10041 68851 10107 68854
rect 2630 68716 2636 68780
rect 2700 68778 2706 68780
rect 4705 68778 4771 68781
rect 2700 68776 4771 68778
rect 2700 68720 4710 68776
rect 4766 68720 4771 68776
rect 2700 68718 4771 68720
rect 2700 68716 2706 68718
rect 4705 68715 4771 68718
rect 5073 68778 5139 68781
rect 17493 68778 17559 68781
rect 5073 68776 17559 68778
rect 5073 68720 5078 68776
rect 5134 68720 17498 68776
rect 17554 68720 17559 68776
rect 5073 68718 17559 68720
rect 5073 68715 5139 68718
rect 17493 68715 17559 68718
rect 19520 68642 20000 68672
rect 18094 68582 20000 68642
rect 4277 68576 4597 68577
rect 4277 68512 4285 68576
rect 4349 68512 4365 68576
rect 4429 68512 4445 68576
rect 4509 68512 4525 68576
rect 4589 68512 4597 68576
rect 4277 68511 4597 68512
rect 10944 68576 11264 68577
rect 10944 68512 10952 68576
rect 11016 68512 11032 68576
rect 11096 68512 11112 68576
rect 11176 68512 11192 68576
rect 11256 68512 11264 68576
rect 10944 68511 11264 68512
rect 17610 68576 17930 68577
rect 17610 68512 17618 68576
rect 17682 68512 17698 68576
rect 17762 68512 17778 68576
rect 17842 68512 17858 68576
rect 17922 68512 17930 68576
rect 17610 68511 17930 68512
rect 14038 68308 14044 68372
rect 14108 68370 14114 68372
rect 18094 68370 18154 68582
rect 19520 68552 20000 68582
rect 14108 68310 18154 68370
rect 14108 68308 14114 68310
rect 0 68234 480 68264
rect 4153 68234 4219 68237
rect 0 68232 4219 68234
rect 0 68176 4158 68232
rect 4214 68176 4219 68232
rect 0 68174 4219 68176
rect 0 68144 480 68174
rect 4153 68171 4219 68174
rect 11605 68234 11671 68237
rect 13445 68234 13511 68237
rect 11605 68232 13511 68234
rect 11605 68176 11610 68232
rect 11666 68176 13450 68232
rect 13506 68176 13511 68232
rect 11605 68174 13511 68176
rect 11605 68171 11671 68174
rect 13445 68171 13511 68174
rect 13905 68100 13971 68101
rect 13854 68036 13860 68100
rect 13924 68098 13971 68100
rect 13924 68096 14016 68098
rect 13966 68040 14016 68096
rect 13924 68038 14016 68040
rect 13924 68036 13971 68038
rect 13905 68035 13971 68036
rect 7610 68032 7930 68033
rect 7610 67968 7618 68032
rect 7682 67968 7698 68032
rect 7762 67968 7778 68032
rect 7842 67968 7858 68032
rect 7922 67968 7930 68032
rect 7610 67967 7930 67968
rect 14277 68032 14597 68033
rect 14277 67968 14285 68032
rect 14349 67968 14365 68032
rect 14429 67968 14445 68032
rect 14509 67968 14525 68032
rect 14589 67968 14597 68032
rect 14277 67967 14597 67968
rect 19520 67962 20000 67992
rect 14736 67902 20000 67962
rect 14089 67826 14155 67829
rect 14736 67826 14796 67902
rect 19520 67872 20000 67902
rect 14089 67824 14796 67826
rect 14089 67768 14094 67824
rect 14150 67768 14796 67824
rect 14089 67766 14796 67768
rect 14089 67763 14155 67766
rect 4277 67488 4597 67489
rect 0 67418 480 67448
rect 4277 67424 4285 67488
rect 4349 67424 4365 67488
rect 4429 67424 4445 67488
rect 4509 67424 4525 67488
rect 4589 67424 4597 67488
rect 4277 67423 4597 67424
rect 10944 67488 11264 67489
rect 10944 67424 10952 67488
rect 11016 67424 11032 67488
rect 11096 67424 11112 67488
rect 11176 67424 11192 67488
rect 11256 67424 11264 67488
rect 10944 67423 11264 67424
rect 17610 67488 17930 67489
rect 17610 67424 17618 67488
rect 17682 67424 17698 67488
rect 17762 67424 17778 67488
rect 17842 67424 17858 67488
rect 17922 67424 17930 67488
rect 17610 67423 17930 67424
rect 1301 67418 1367 67421
rect 0 67416 1367 67418
rect 0 67360 1306 67416
rect 1362 67360 1367 67416
rect 0 67358 1367 67360
rect 0 67328 480 67358
rect 1301 67355 1367 67358
rect 10409 67282 10475 67285
rect 14365 67282 14431 67285
rect 10409 67280 14431 67282
rect 10409 67224 10414 67280
rect 10470 67224 14370 67280
rect 14426 67224 14431 67280
rect 10409 67222 14431 67224
rect 10409 67219 10475 67222
rect 14365 67219 14431 67222
rect 17125 67282 17191 67285
rect 19520 67282 20000 67312
rect 17125 67280 20000 67282
rect 17125 67224 17130 67280
rect 17186 67224 20000 67280
rect 17125 67222 20000 67224
rect 17125 67219 17191 67222
rect 19520 67192 20000 67222
rect 5257 67146 5323 67149
rect 7189 67146 7255 67149
rect 5257 67144 7255 67146
rect 5257 67088 5262 67144
rect 5318 67088 7194 67144
rect 7250 67088 7255 67144
rect 5257 67086 7255 67088
rect 5257 67083 5323 67086
rect 7189 67083 7255 67086
rect 9673 67146 9739 67149
rect 17493 67146 17559 67149
rect 9673 67144 17559 67146
rect 9673 67088 9678 67144
rect 9734 67088 17498 67144
rect 17554 67088 17559 67144
rect 9673 67086 17559 67088
rect 9673 67083 9739 67086
rect 17493 67083 17559 67086
rect 7610 66944 7930 66945
rect 7610 66880 7618 66944
rect 7682 66880 7698 66944
rect 7762 66880 7778 66944
rect 7842 66880 7858 66944
rect 7922 66880 7930 66944
rect 7610 66879 7930 66880
rect 14277 66944 14597 66945
rect 14277 66880 14285 66944
rect 14349 66880 14365 66944
rect 14429 66880 14445 66944
rect 14509 66880 14525 66944
rect 14589 66880 14597 66944
rect 14277 66879 14597 66880
rect 0 66738 480 66768
rect 1669 66738 1735 66741
rect 0 66736 1735 66738
rect 0 66680 1674 66736
rect 1730 66680 1735 66736
rect 0 66678 1735 66680
rect 0 66648 480 66678
rect 1669 66675 1735 66678
rect 16665 66602 16731 66605
rect 19520 66602 20000 66632
rect 16665 66600 20000 66602
rect 16665 66544 16670 66600
rect 16726 66544 20000 66600
rect 16665 66542 20000 66544
rect 16665 66539 16731 66542
rect 19520 66512 20000 66542
rect 4277 66400 4597 66401
rect 4277 66336 4285 66400
rect 4349 66336 4365 66400
rect 4429 66336 4445 66400
rect 4509 66336 4525 66400
rect 4589 66336 4597 66400
rect 4277 66335 4597 66336
rect 10944 66400 11264 66401
rect 10944 66336 10952 66400
rect 11016 66336 11032 66400
rect 11096 66336 11112 66400
rect 11176 66336 11192 66400
rect 11256 66336 11264 66400
rect 10944 66335 11264 66336
rect 17610 66400 17930 66401
rect 17610 66336 17618 66400
rect 17682 66336 17698 66400
rect 17762 66336 17778 66400
rect 17842 66336 17858 66400
rect 17922 66336 17930 66400
rect 17610 66335 17930 66336
rect 5441 66194 5507 66197
rect 7557 66194 7623 66197
rect 5441 66192 7623 66194
rect 5441 66136 5446 66192
rect 5502 66136 7562 66192
rect 7618 66136 7623 66192
rect 5441 66134 7623 66136
rect 5441 66131 5507 66134
rect 7557 66131 7623 66134
rect 0 65922 480 65952
rect 3509 65922 3575 65925
rect 0 65920 3575 65922
rect 0 65864 3514 65920
rect 3570 65864 3575 65920
rect 0 65862 3575 65864
rect 0 65832 480 65862
rect 3509 65859 3575 65862
rect 10041 65922 10107 65925
rect 10358 65922 10364 65924
rect 10041 65920 10364 65922
rect 10041 65864 10046 65920
rect 10102 65864 10364 65920
rect 10041 65862 10364 65864
rect 10041 65859 10107 65862
rect 10358 65860 10364 65862
rect 10428 65860 10434 65924
rect 10593 65922 10659 65925
rect 12617 65922 12683 65925
rect 13905 65922 13971 65925
rect 14733 65924 14799 65925
rect 14733 65922 14780 65924
rect 10593 65920 13971 65922
rect 10593 65864 10598 65920
rect 10654 65864 12622 65920
rect 12678 65864 13910 65920
rect 13966 65864 13971 65920
rect 10593 65862 13971 65864
rect 14688 65920 14780 65922
rect 14688 65864 14738 65920
rect 14688 65862 14780 65864
rect 10593 65859 10659 65862
rect 12617 65859 12683 65862
rect 13905 65859 13971 65862
rect 14733 65860 14780 65862
rect 14844 65860 14850 65924
rect 16941 65922 17007 65925
rect 19520 65922 20000 65952
rect 16941 65920 20000 65922
rect 16941 65864 16946 65920
rect 17002 65864 20000 65920
rect 16941 65862 20000 65864
rect 14733 65859 14799 65860
rect 16941 65859 17007 65862
rect 7610 65856 7930 65857
rect 7610 65792 7618 65856
rect 7682 65792 7698 65856
rect 7762 65792 7778 65856
rect 7842 65792 7858 65856
rect 7922 65792 7930 65856
rect 7610 65791 7930 65792
rect 14277 65856 14597 65857
rect 14277 65792 14285 65856
rect 14349 65792 14365 65856
rect 14429 65792 14445 65856
rect 14509 65792 14525 65856
rect 14589 65792 14597 65856
rect 19520 65832 20000 65862
rect 14277 65791 14597 65792
rect 9121 65786 9187 65789
rect 11237 65786 11303 65789
rect 11462 65786 11468 65788
rect 9121 65784 11468 65786
rect 9121 65728 9126 65784
rect 9182 65728 11242 65784
rect 11298 65728 11468 65784
rect 9121 65726 11468 65728
rect 9121 65723 9187 65726
rect 11237 65723 11303 65726
rect 11462 65724 11468 65726
rect 11532 65724 11538 65788
rect 9397 65650 9463 65653
rect 17493 65650 17559 65653
rect 9397 65648 17559 65650
rect 9397 65592 9402 65648
rect 9458 65592 17498 65648
rect 17554 65592 17559 65648
rect 9397 65590 17559 65592
rect 9397 65587 9463 65590
rect 17493 65587 17559 65590
rect 8201 65514 8267 65517
rect 12433 65514 12499 65517
rect 8201 65512 12499 65514
rect 8201 65456 8206 65512
rect 8262 65456 12438 65512
rect 12494 65456 12499 65512
rect 8201 65454 12499 65456
rect 8201 65451 8267 65454
rect 12433 65451 12499 65454
rect 16389 65514 16455 65517
rect 16389 65512 18154 65514
rect 16389 65456 16394 65512
rect 16450 65456 18154 65512
rect 16389 65454 18154 65456
rect 16389 65451 16455 65454
rect 4277 65312 4597 65313
rect 4277 65248 4285 65312
rect 4349 65248 4365 65312
rect 4429 65248 4445 65312
rect 4509 65248 4525 65312
rect 4589 65248 4597 65312
rect 4277 65247 4597 65248
rect 10944 65312 11264 65313
rect 10944 65248 10952 65312
rect 11016 65248 11032 65312
rect 11096 65248 11112 65312
rect 11176 65248 11192 65312
rect 11256 65248 11264 65312
rect 10944 65247 11264 65248
rect 17610 65312 17930 65313
rect 17610 65248 17618 65312
rect 17682 65248 17698 65312
rect 17762 65248 17778 65312
rect 17842 65248 17858 65312
rect 17922 65248 17930 65312
rect 17610 65247 17930 65248
rect 10542 65180 10548 65244
rect 10612 65242 10618 65244
rect 10777 65242 10843 65245
rect 10612 65240 10843 65242
rect 10612 65184 10782 65240
rect 10838 65184 10843 65240
rect 10612 65182 10843 65184
rect 18094 65242 18154 65454
rect 19520 65242 20000 65272
rect 18094 65182 20000 65242
rect 10612 65180 10618 65182
rect 10777 65179 10843 65182
rect 19520 65152 20000 65182
rect 0 65106 480 65136
rect 1761 65106 1827 65109
rect 0 65104 1827 65106
rect 0 65048 1766 65104
rect 1822 65048 1827 65104
rect 0 65046 1827 65048
rect 0 65016 480 65046
rect 1761 65043 1827 65046
rect 8293 64834 8359 64837
rect 8661 64834 8727 64837
rect 8293 64832 8727 64834
rect 8293 64776 8298 64832
rect 8354 64776 8666 64832
rect 8722 64776 8727 64832
rect 8293 64774 8727 64776
rect 8293 64771 8359 64774
rect 8661 64771 8727 64774
rect 10685 64834 10751 64837
rect 12525 64834 12591 64837
rect 10685 64832 12591 64834
rect 10685 64776 10690 64832
rect 10746 64776 12530 64832
rect 12586 64776 12591 64832
rect 10685 64774 12591 64776
rect 10685 64771 10751 64774
rect 12525 64771 12591 64774
rect 7610 64768 7930 64769
rect 7610 64704 7618 64768
rect 7682 64704 7698 64768
rect 7762 64704 7778 64768
rect 7842 64704 7858 64768
rect 7922 64704 7930 64768
rect 7610 64703 7930 64704
rect 14277 64768 14597 64769
rect 14277 64704 14285 64768
rect 14349 64704 14365 64768
rect 14429 64704 14445 64768
rect 14509 64704 14525 64768
rect 14589 64704 14597 64768
rect 14277 64703 14597 64704
rect 7189 64562 7255 64565
rect 7414 64562 7420 64564
rect 7189 64560 7420 64562
rect 7189 64504 7194 64560
rect 7250 64504 7420 64560
rect 7189 64502 7420 64504
rect 7189 64499 7255 64502
rect 7414 64500 7420 64502
rect 7484 64562 7490 64564
rect 14365 64562 14431 64565
rect 7484 64560 14431 64562
rect 7484 64504 14370 64560
rect 14426 64504 14431 64560
rect 7484 64502 14431 64504
rect 7484 64500 7490 64502
rect 14365 64499 14431 64502
rect 16481 64562 16547 64565
rect 19520 64562 20000 64592
rect 16481 64560 20000 64562
rect 16481 64504 16486 64560
rect 16542 64504 20000 64560
rect 16481 64502 20000 64504
rect 16481 64499 16547 64502
rect 19520 64472 20000 64502
rect 13445 64426 13511 64429
rect 16849 64426 16915 64429
rect 13445 64424 16915 64426
rect 13445 64368 13450 64424
rect 13506 64368 16854 64424
rect 16910 64368 16915 64424
rect 13445 64366 16915 64368
rect 13445 64363 13511 64366
rect 16849 64363 16915 64366
rect 0 64290 480 64320
rect 2865 64290 2931 64293
rect 0 64288 2931 64290
rect 0 64232 2870 64288
rect 2926 64232 2931 64288
rect 0 64230 2931 64232
rect 0 64200 480 64230
rect 2865 64227 2931 64230
rect 4277 64224 4597 64225
rect 4277 64160 4285 64224
rect 4349 64160 4365 64224
rect 4429 64160 4445 64224
rect 4509 64160 4525 64224
rect 4589 64160 4597 64224
rect 4277 64159 4597 64160
rect 10944 64224 11264 64225
rect 10944 64160 10952 64224
rect 11016 64160 11032 64224
rect 11096 64160 11112 64224
rect 11176 64160 11192 64224
rect 11256 64160 11264 64224
rect 10944 64159 11264 64160
rect 17610 64224 17930 64225
rect 17610 64160 17618 64224
rect 17682 64160 17698 64224
rect 17762 64160 17778 64224
rect 17842 64160 17858 64224
rect 17922 64160 17930 64224
rect 17610 64159 17930 64160
rect 4061 64018 4127 64021
rect 5441 64018 5507 64021
rect 9121 64018 9187 64021
rect 4061 64016 5507 64018
rect 4061 63960 4066 64016
rect 4122 63960 5446 64016
rect 5502 63960 5507 64016
rect 4061 63958 5507 63960
rect 4061 63955 4127 63958
rect 5441 63955 5507 63958
rect 7790 64016 9187 64018
rect 7790 63960 9126 64016
rect 9182 63960 9187 64016
rect 7790 63958 9187 63960
rect 2681 63882 2747 63885
rect 4153 63882 4219 63885
rect 7790 63882 7850 63958
rect 9121 63955 9187 63958
rect 9806 63956 9812 64020
rect 9876 64018 9882 64020
rect 9949 64018 10015 64021
rect 9876 64016 10015 64018
rect 9876 63960 9954 64016
rect 10010 63960 10015 64016
rect 9876 63958 10015 63960
rect 9876 63956 9882 63958
rect 9949 63955 10015 63958
rect 2681 63880 4219 63882
rect 2681 63824 2686 63880
rect 2742 63824 4158 63880
rect 4214 63824 4219 63880
rect 2681 63822 4219 63824
rect 2681 63819 2747 63822
rect 4153 63819 4219 63822
rect 7468 63822 7850 63882
rect 7925 63882 7991 63885
rect 9121 63882 9187 63885
rect 7925 63880 9187 63882
rect 7925 63824 7930 63880
rect 7986 63824 9126 63880
rect 9182 63824 9187 63880
rect 7925 63822 9187 63824
rect 7468 63746 7528 63822
rect 7925 63819 7991 63822
rect 9121 63819 9187 63822
rect 13077 63882 13143 63885
rect 15377 63882 15443 63885
rect 13077 63880 15443 63882
rect 13077 63824 13082 63880
rect 13138 63824 15382 63880
rect 15438 63824 15443 63880
rect 13077 63822 15443 63824
rect 13077 63819 13143 63822
rect 15377 63819 15443 63822
rect 16389 63882 16455 63885
rect 19520 63882 20000 63912
rect 16389 63880 20000 63882
rect 16389 63824 16394 63880
rect 16450 63824 20000 63880
rect 16389 63822 20000 63824
rect 16389 63819 16455 63822
rect 19520 63792 20000 63822
rect 2270 63686 7528 63746
rect 0 63474 480 63504
rect 2129 63474 2195 63477
rect 0 63472 2195 63474
rect 0 63416 2134 63472
rect 2190 63416 2195 63472
rect 0 63414 2195 63416
rect 0 63384 480 63414
rect 2129 63411 2195 63414
rect 2270 63338 2330 63686
rect 7046 63548 7052 63612
rect 7116 63610 7122 63612
rect 7189 63610 7255 63613
rect 7116 63608 7255 63610
rect 7116 63552 7194 63608
rect 7250 63552 7255 63608
rect 7116 63550 7255 63552
rect 7116 63548 7122 63550
rect 7189 63547 7255 63550
rect 2497 63474 2563 63477
rect 5625 63474 5691 63477
rect 2497 63472 5691 63474
rect 2497 63416 2502 63472
rect 2558 63416 5630 63472
rect 5686 63416 5691 63472
rect 2497 63414 5691 63416
rect 7468 63474 7528 63686
rect 13077 63746 13143 63749
rect 13445 63746 13511 63749
rect 13077 63744 13511 63746
rect 13077 63688 13082 63744
rect 13138 63688 13450 63744
rect 13506 63688 13511 63744
rect 13077 63686 13511 63688
rect 13077 63683 13143 63686
rect 13445 63683 13511 63686
rect 7610 63680 7930 63681
rect 7610 63616 7618 63680
rect 7682 63616 7698 63680
rect 7762 63616 7778 63680
rect 7842 63616 7858 63680
rect 7922 63616 7930 63680
rect 7610 63615 7930 63616
rect 14277 63680 14597 63681
rect 14277 63616 14285 63680
rect 14349 63616 14365 63680
rect 14429 63616 14445 63680
rect 14509 63616 14525 63680
rect 14589 63616 14597 63680
rect 14277 63615 14597 63616
rect 11145 63610 11211 63613
rect 11102 63608 11211 63610
rect 11102 63552 11150 63608
rect 11206 63552 11211 63608
rect 11102 63547 11211 63552
rect 8385 63474 8451 63477
rect 7468 63472 8451 63474
rect 7468 63416 8390 63472
rect 8446 63416 8451 63472
rect 7468 63414 8451 63416
rect 2497 63411 2563 63414
rect 5625 63411 5691 63414
rect 8385 63411 8451 63414
rect 8569 63474 8635 63477
rect 9213 63474 9279 63477
rect 11102 63474 11162 63547
rect 8569 63472 11162 63474
rect 8569 63416 8574 63472
rect 8630 63416 9218 63472
rect 9274 63416 11162 63472
rect 8569 63414 11162 63416
rect 8569 63411 8635 63414
rect 9213 63411 9279 63414
rect 2497 63338 2563 63341
rect 2270 63336 2563 63338
rect 2270 63280 2502 63336
rect 2558 63280 2563 63336
rect 2270 63278 2563 63280
rect 2497 63275 2563 63278
rect 4521 63338 4587 63341
rect 6085 63338 6151 63341
rect 7741 63338 7807 63341
rect 4521 63336 7807 63338
rect 4521 63280 4526 63336
rect 4582 63280 6090 63336
rect 6146 63280 7746 63336
rect 7802 63280 7807 63336
rect 4521 63278 7807 63280
rect 4521 63275 4587 63278
rect 6085 63275 6151 63278
rect 7741 63275 7807 63278
rect 15193 63338 15259 63341
rect 15193 63336 18154 63338
rect 15193 63280 15198 63336
rect 15254 63280 18154 63336
rect 15193 63278 18154 63280
rect 15193 63275 15259 63278
rect 12893 63202 12959 63205
rect 16205 63202 16271 63205
rect 12893 63200 16271 63202
rect 12893 63144 12898 63200
rect 12954 63144 16210 63200
rect 16266 63144 16271 63200
rect 12893 63142 16271 63144
rect 18094 63202 18154 63278
rect 19520 63202 20000 63232
rect 18094 63142 20000 63202
rect 12893 63139 12959 63142
rect 16205 63139 16271 63142
rect 4277 63136 4597 63137
rect 4277 63072 4285 63136
rect 4349 63072 4365 63136
rect 4429 63072 4445 63136
rect 4509 63072 4525 63136
rect 4589 63072 4597 63136
rect 4277 63071 4597 63072
rect 10944 63136 11264 63137
rect 10944 63072 10952 63136
rect 11016 63072 11032 63136
rect 11096 63072 11112 63136
rect 11176 63072 11192 63136
rect 11256 63072 11264 63136
rect 10944 63071 11264 63072
rect 17610 63136 17930 63137
rect 17610 63072 17618 63136
rect 17682 63072 17698 63136
rect 17762 63072 17778 63136
rect 17842 63072 17858 63136
rect 17922 63072 17930 63136
rect 19520 63112 20000 63142
rect 17610 63071 17930 63072
rect 7230 63004 7236 63068
rect 7300 63066 7306 63068
rect 8334 63066 8340 63068
rect 7300 63006 8340 63066
rect 7300 63004 7306 63006
rect 8334 63004 8340 63006
rect 8404 63004 8410 63068
rect 3366 62868 3372 62932
rect 3436 62930 3442 62932
rect 8753 62930 8819 62933
rect 3436 62928 8819 62930
rect 3436 62872 8758 62928
rect 8814 62872 8819 62928
rect 3436 62870 8819 62872
rect 3436 62868 3442 62870
rect 8753 62867 8819 62870
rect 9397 62930 9463 62933
rect 10041 62930 10107 62933
rect 9397 62928 10107 62930
rect 9397 62872 9402 62928
rect 9458 62872 10046 62928
rect 10102 62872 10107 62928
rect 9397 62870 10107 62872
rect 9397 62867 9463 62870
rect 10041 62867 10107 62870
rect 7741 62794 7807 62797
rect 17493 62794 17559 62797
rect 7741 62792 17559 62794
rect 7741 62736 7746 62792
rect 7802 62736 17498 62792
rect 17554 62736 17559 62792
rect 7741 62734 17559 62736
rect 7741 62731 7807 62734
rect 17493 62731 17559 62734
rect 0 62658 480 62688
rect 1485 62658 1551 62661
rect 0 62656 1551 62658
rect 0 62600 1490 62656
rect 1546 62600 1551 62656
rect 0 62598 1551 62600
rect 0 62568 480 62598
rect 1485 62595 1551 62598
rect 10777 62658 10843 62661
rect 11513 62658 11579 62661
rect 10777 62656 11579 62658
rect 10777 62600 10782 62656
rect 10838 62600 11518 62656
rect 11574 62600 11579 62656
rect 10777 62598 11579 62600
rect 10777 62595 10843 62598
rect 11513 62595 11579 62598
rect 7610 62592 7930 62593
rect 7610 62528 7618 62592
rect 7682 62528 7698 62592
rect 7762 62528 7778 62592
rect 7842 62528 7858 62592
rect 7922 62528 7930 62592
rect 7610 62527 7930 62528
rect 14277 62592 14597 62593
rect 14277 62528 14285 62592
rect 14349 62528 14365 62592
rect 14429 62528 14445 62592
rect 14509 62528 14525 62592
rect 14589 62528 14597 62592
rect 14277 62527 14597 62528
rect 15377 62522 15443 62525
rect 19520 62522 20000 62552
rect 15377 62520 20000 62522
rect 15377 62464 15382 62520
rect 15438 62464 20000 62520
rect 15377 62462 20000 62464
rect 15377 62459 15443 62462
rect 19520 62432 20000 62462
rect 7189 62386 7255 62389
rect 12014 62386 12020 62388
rect 7189 62384 12020 62386
rect 7189 62328 7194 62384
rect 7250 62328 12020 62384
rect 7189 62326 12020 62328
rect 7189 62323 7255 62326
rect 12014 62324 12020 62326
rect 12084 62386 12090 62388
rect 15193 62386 15259 62389
rect 12084 62384 15259 62386
rect 12084 62328 15198 62384
rect 15254 62328 15259 62384
rect 12084 62326 15259 62328
rect 12084 62324 12090 62326
rect 15193 62323 15259 62326
rect 9213 62250 9279 62253
rect 9990 62250 9996 62252
rect 9213 62248 9996 62250
rect 9213 62192 9218 62248
rect 9274 62192 9996 62248
rect 9213 62190 9996 62192
rect 9213 62187 9279 62190
rect 9990 62188 9996 62190
rect 10060 62188 10066 62252
rect 10593 62250 10659 62253
rect 10593 62248 12082 62250
rect 10593 62192 10598 62248
rect 10654 62192 12082 62248
rect 10593 62190 12082 62192
rect 10593 62187 10659 62190
rect 12022 62117 12082 62190
rect 12198 62188 12204 62252
rect 12268 62250 12274 62252
rect 12433 62250 12499 62253
rect 15561 62250 15627 62253
rect 12268 62248 12499 62250
rect 12268 62192 12438 62248
rect 12494 62192 12499 62248
rect 12268 62190 12499 62192
rect 12268 62188 12274 62190
rect 12433 62187 12499 62190
rect 12574 62248 15627 62250
rect 12574 62192 15566 62248
rect 15622 62192 15627 62248
rect 12574 62190 15627 62192
rect 7097 62114 7163 62117
rect 10174 62114 10180 62116
rect 7097 62112 10180 62114
rect 7097 62056 7102 62112
rect 7158 62056 10180 62112
rect 7097 62054 10180 62056
rect 7097 62051 7163 62054
rect 10174 62052 10180 62054
rect 10244 62052 10250 62116
rect 12022 62114 12131 62117
rect 12574 62114 12634 62190
rect 15561 62187 15627 62190
rect 11938 62112 12634 62114
rect 11938 62056 12070 62112
rect 12126 62056 12634 62112
rect 11938 62054 12634 62056
rect 12065 62051 12131 62054
rect 4277 62048 4597 62049
rect 4277 61984 4285 62048
rect 4349 61984 4365 62048
rect 4429 61984 4445 62048
rect 4509 61984 4525 62048
rect 4589 61984 4597 62048
rect 4277 61983 4597 61984
rect 10944 62048 11264 62049
rect 10944 61984 10952 62048
rect 11016 61984 11032 62048
rect 11096 61984 11112 62048
rect 11176 61984 11192 62048
rect 11256 61984 11264 62048
rect 10944 61983 11264 61984
rect 17610 62048 17930 62049
rect 17610 61984 17618 62048
rect 17682 61984 17698 62048
rect 17762 61984 17778 62048
rect 17842 61984 17858 62048
rect 17922 61984 17930 62048
rect 17610 61983 17930 61984
rect 0 61842 480 61872
rect 1945 61842 2011 61845
rect 0 61840 2011 61842
rect 0 61784 1950 61840
rect 2006 61784 2011 61840
rect 0 61782 2011 61784
rect 0 61752 480 61782
rect 1945 61779 2011 61782
rect 16481 61842 16547 61845
rect 19520 61842 20000 61872
rect 16481 61840 20000 61842
rect 16481 61784 16486 61840
rect 16542 61784 20000 61840
rect 16481 61782 20000 61784
rect 16481 61779 16547 61782
rect 19520 61752 20000 61782
rect 7610 61504 7930 61505
rect 7610 61440 7618 61504
rect 7682 61440 7698 61504
rect 7762 61440 7778 61504
rect 7842 61440 7858 61504
rect 7922 61440 7930 61504
rect 7610 61439 7930 61440
rect 14277 61504 14597 61505
rect 14277 61440 14285 61504
rect 14349 61440 14365 61504
rect 14429 61440 14445 61504
rect 14509 61440 14525 61504
rect 14589 61440 14597 61504
rect 14277 61439 14597 61440
rect 8293 61298 8359 61301
rect 10041 61298 10107 61301
rect 8293 61296 10107 61298
rect 8293 61240 8298 61296
rect 8354 61240 10046 61296
rect 10102 61240 10107 61296
rect 8293 61238 10107 61240
rect 8293 61235 8359 61238
rect 10041 61235 10107 61238
rect 10542 61236 10548 61300
rect 10612 61298 10618 61300
rect 11053 61298 11119 61301
rect 10612 61296 11119 61298
rect 10612 61240 11058 61296
rect 11114 61240 11119 61296
rect 10612 61238 11119 61240
rect 10612 61236 10618 61238
rect 11053 61235 11119 61238
rect 14774 61236 14780 61300
rect 14844 61298 14850 61300
rect 15326 61298 15332 61300
rect 14844 61238 15332 61298
rect 14844 61236 14850 61238
rect 15326 61236 15332 61238
rect 15396 61236 15402 61300
rect 3141 61162 3207 61165
rect 3785 61162 3851 61165
rect 3141 61160 3851 61162
rect 3141 61104 3146 61160
rect 3202 61104 3790 61160
rect 3846 61104 3851 61160
rect 3141 61102 3851 61104
rect 3141 61099 3207 61102
rect 3785 61099 3851 61102
rect 10542 61100 10548 61164
rect 10612 61162 10618 61164
rect 12893 61162 12959 61165
rect 10612 61160 12959 61162
rect 10612 61104 12898 61160
rect 12954 61104 12959 61160
rect 10612 61102 12959 61104
rect 10612 61100 10618 61102
rect 12893 61099 12959 61102
rect 15377 61162 15443 61165
rect 19520 61162 20000 61192
rect 15377 61160 20000 61162
rect 15377 61104 15382 61160
rect 15438 61104 20000 61160
rect 15377 61102 20000 61104
rect 15377 61099 15443 61102
rect 19520 61072 20000 61102
rect 0 61026 480 61056
rect 1485 61026 1551 61029
rect 0 61024 1551 61026
rect 0 60968 1490 61024
rect 1546 60968 1551 61024
rect 0 60966 1551 60968
rect 0 60936 480 60966
rect 1485 60963 1551 60966
rect 14038 60964 14044 61028
rect 14108 61026 14114 61028
rect 14733 61026 14799 61029
rect 14108 61024 14799 61026
rect 14108 60968 14738 61024
rect 14794 60968 14799 61024
rect 14108 60966 14799 60968
rect 14108 60964 14114 60966
rect 14733 60963 14799 60966
rect 14917 61026 14983 61029
rect 15377 61026 15443 61029
rect 14917 61024 15443 61026
rect 14917 60968 14922 61024
rect 14978 60968 15382 61024
rect 15438 60968 15443 61024
rect 14917 60966 15443 60968
rect 14917 60963 14983 60966
rect 15377 60963 15443 60966
rect 4277 60960 4597 60961
rect 4277 60896 4285 60960
rect 4349 60896 4365 60960
rect 4429 60896 4445 60960
rect 4509 60896 4525 60960
rect 4589 60896 4597 60960
rect 4277 60895 4597 60896
rect 10944 60960 11264 60961
rect 10944 60896 10952 60960
rect 11016 60896 11032 60960
rect 11096 60896 11112 60960
rect 11176 60896 11192 60960
rect 11256 60896 11264 60960
rect 10944 60895 11264 60896
rect 17610 60960 17930 60961
rect 17610 60896 17618 60960
rect 17682 60896 17698 60960
rect 17762 60896 17778 60960
rect 17842 60896 17858 60960
rect 17922 60896 17930 60960
rect 17610 60895 17930 60896
rect 12433 60890 12499 60893
rect 13261 60890 13327 60893
rect 16113 60890 16179 60893
rect 12433 60888 16179 60890
rect 12433 60832 12438 60888
rect 12494 60832 13266 60888
rect 13322 60832 16118 60888
rect 16174 60832 16179 60888
rect 12433 60830 16179 60832
rect 12433 60827 12499 60830
rect 13261 60827 13327 60830
rect 16113 60827 16179 60830
rect 9806 60754 9812 60756
rect 4110 60694 9812 60754
rect 3325 60620 3391 60621
rect 3325 60618 3372 60620
rect 3280 60616 3372 60618
rect 3280 60560 3330 60616
rect 3280 60558 3372 60560
rect 3325 60556 3372 60558
rect 3436 60556 3442 60620
rect 3785 60618 3851 60621
rect 4110 60618 4170 60694
rect 9806 60692 9812 60694
rect 9876 60692 9882 60756
rect 9949 60754 10015 60757
rect 10869 60754 10935 60757
rect 14089 60756 14155 60757
rect 14038 60754 14044 60756
rect 9949 60752 10935 60754
rect 9949 60696 9954 60752
rect 10010 60696 10874 60752
rect 10930 60696 10935 60752
rect 9949 60694 10935 60696
rect 13998 60694 14044 60754
rect 14108 60752 14155 60756
rect 14150 60696 14155 60752
rect 9949 60691 10015 60694
rect 10869 60691 10935 60694
rect 14038 60692 14044 60694
rect 14108 60692 14155 60696
rect 14089 60691 14155 60692
rect 14733 60756 14799 60757
rect 14733 60752 14780 60756
rect 14844 60754 14850 60756
rect 14733 60696 14738 60752
rect 14733 60692 14780 60696
rect 14844 60694 14890 60754
rect 14844 60692 14850 60694
rect 14733 60691 14799 60692
rect 3785 60616 4170 60618
rect 3785 60560 3790 60616
rect 3846 60560 4170 60616
rect 3785 60558 4170 60560
rect 4981 60618 5047 60621
rect 6269 60618 6335 60621
rect 7557 60618 7623 60621
rect 17493 60618 17559 60621
rect 4981 60616 5090 60618
rect 4981 60560 4986 60616
rect 5042 60560 5090 60616
rect 3325 60555 3391 60556
rect 3785 60555 3851 60558
rect 4981 60555 5090 60560
rect 6269 60616 17559 60618
rect 6269 60560 6274 60616
rect 6330 60560 7562 60616
rect 7618 60560 17498 60616
rect 17554 60560 17559 60616
rect 6269 60558 17559 60560
rect 6269 60555 6335 60558
rect 7557 60555 7623 60558
rect 17493 60555 17559 60558
rect 2681 60482 2747 60485
rect 4337 60482 4403 60485
rect 2681 60480 4403 60482
rect 2681 60424 2686 60480
rect 2742 60424 4342 60480
rect 4398 60424 4403 60480
rect 2681 60422 4403 60424
rect 5030 60482 5090 60555
rect 5349 60482 5415 60485
rect 5030 60480 5415 60482
rect 5030 60424 5354 60480
rect 5410 60424 5415 60480
rect 5030 60422 5415 60424
rect 2681 60419 2747 60422
rect 4337 60419 4403 60422
rect 5349 60419 5415 60422
rect 16021 60482 16087 60485
rect 19520 60482 20000 60512
rect 16021 60480 20000 60482
rect 16021 60424 16026 60480
rect 16082 60424 20000 60480
rect 16021 60422 20000 60424
rect 16021 60419 16087 60422
rect 7610 60416 7930 60417
rect 0 60346 480 60376
rect 7610 60352 7618 60416
rect 7682 60352 7698 60416
rect 7762 60352 7778 60416
rect 7842 60352 7858 60416
rect 7922 60352 7930 60416
rect 7610 60351 7930 60352
rect 14277 60416 14597 60417
rect 14277 60352 14285 60416
rect 14349 60352 14365 60416
rect 14429 60352 14445 60416
rect 14509 60352 14525 60416
rect 14589 60352 14597 60416
rect 19520 60392 20000 60422
rect 14277 60351 14597 60352
rect 1577 60346 1643 60349
rect 0 60344 1643 60346
rect 0 60288 1582 60344
rect 1638 60288 1643 60344
rect 0 60286 1643 60288
rect 0 60256 480 60286
rect 1577 60283 1643 60286
rect 14733 60346 14799 60349
rect 16665 60346 16731 60349
rect 14733 60344 16731 60346
rect 14733 60288 14738 60344
rect 14794 60288 16670 60344
rect 16726 60288 16731 60344
rect 14733 60286 16731 60288
rect 14733 60283 14799 60286
rect 16665 60283 16731 60286
rect 2497 60210 2563 60213
rect 8385 60210 8451 60213
rect 2497 60208 8451 60210
rect 2497 60152 2502 60208
rect 2558 60152 8390 60208
rect 8446 60152 8451 60208
rect 2497 60150 8451 60152
rect 2497 60147 2563 60150
rect 8385 60147 8451 60150
rect 10409 60210 10475 60213
rect 14181 60210 14247 60213
rect 16573 60210 16639 60213
rect 10409 60208 16639 60210
rect 10409 60152 10414 60208
rect 10470 60152 14186 60208
rect 14242 60152 16578 60208
rect 16634 60152 16639 60208
rect 10409 60150 16639 60152
rect 10409 60147 10475 60150
rect 14181 60147 14247 60150
rect 16573 60147 16639 60150
rect 3693 60074 3759 60077
rect 6177 60074 6243 60077
rect 3693 60072 6243 60074
rect 3693 60016 3698 60072
rect 3754 60016 6182 60072
rect 6238 60016 6243 60072
rect 3693 60014 6243 60016
rect 3693 60011 3759 60014
rect 6177 60011 6243 60014
rect 9254 60012 9260 60076
rect 9324 60074 9330 60076
rect 11513 60074 11579 60077
rect 14089 60074 14155 60077
rect 9324 60072 14155 60074
rect 9324 60016 11518 60072
rect 11574 60016 14094 60072
rect 14150 60016 14155 60072
rect 9324 60014 14155 60016
rect 9324 60012 9330 60014
rect 11513 60011 11579 60014
rect 14089 60011 14155 60014
rect 15377 60074 15443 60077
rect 15377 60072 18154 60074
rect 15377 60016 15382 60072
rect 15438 60016 18154 60072
rect 15377 60014 18154 60016
rect 15377 60011 15443 60014
rect 4277 59872 4597 59873
rect 4277 59808 4285 59872
rect 4349 59808 4365 59872
rect 4429 59808 4445 59872
rect 4509 59808 4525 59872
rect 4589 59808 4597 59872
rect 4277 59807 4597 59808
rect 10944 59872 11264 59873
rect 10944 59808 10952 59872
rect 11016 59808 11032 59872
rect 11096 59808 11112 59872
rect 11176 59808 11192 59872
rect 11256 59808 11264 59872
rect 10944 59807 11264 59808
rect 17610 59872 17930 59873
rect 17610 59808 17618 59872
rect 17682 59808 17698 59872
rect 17762 59808 17778 59872
rect 17842 59808 17858 59872
rect 17922 59808 17930 59872
rect 17610 59807 17930 59808
rect 6637 59802 6703 59805
rect 9029 59802 9095 59805
rect 10777 59802 10843 59805
rect 6637 59800 9095 59802
rect 6637 59744 6642 59800
rect 6698 59744 9034 59800
rect 9090 59744 9095 59800
rect 6637 59742 9095 59744
rect 6637 59739 6703 59742
rect 9029 59739 9095 59742
rect 10550 59800 10843 59802
rect 10550 59744 10782 59800
rect 10838 59744 10843 59800
rect 10550 59742 10843 59744
rect 18094 59802 18154 60014
rect 19520 59802 20000 59832
rect 18094 59742 20000 59802
rect 2589 59666 2655 59669
rect 7281 59666 7347 59669
rect 2589 59664 10472 59666
rect 2589 59608 2594 59664
rect 2650 59608 7286 59664
rect 7342 59608 10472 59664
rect 2589 59606 10472 59608
rect 2589 59603 2655 59606
rect 7281 59603 7347 59606
rect 0 59530 480 59560
rect 1393 59530 1459 59533
rect 0 59528 1459 59530
rect 0 59472 1398 59528
rect 1454 59472 1459 59528
rect 0 59470 1459 59472
rect 0 59440 480 59470
rect 1393 59467 1459 59470
rect 10412 59397 10472 59606
rect 3417 59396 3483 59397
rect 3366 59332 3372 59396
rect 3436 59394 3483 59396
rect 6269 59394 6335 59397
rect 7281 59394 7347 59397
rect 3436 59392 3528 59394
rect 3478 59336 3528 59392
rect 3436 59334 3528 59336
rect 6269 59392 7347 59394
rect 6269 59336 6274 59392
rect 6330 59336 7286 59392
rect 7342 59336 7347 59392
rect 6269 59334 7347 59336
rect 3436 59332 3483 59334
rect 3417 59331 3483 59332
rect 6269 59331 6335 59334
rect 7281 59331 7347 59334
rect 9857 59394 9923 59397
rect 10041 59394 10107 59397
rect 9857 59392 10107 59394
rect 9857 59336 9862 59392
rect 9918 59336 10046 59392
rect 10102 59336 10107 59392
rect 9857 59334 10107 59336
rect 9857 59331 9923 59334
rect 10041 59331 10107 59334
rect 10409 59392 10475 59397
rect 10409 59336 10414 59392
rect 10470 59336 10475 59392
rect 10409 59331 10475 59336
rect 7610 59328 7930 59329
rect 7610 59264 7618 59328
rect 7682 59264 7698 59328
rect 7762 59264 7778 59328
rect 7842 59264 7858 59328
rect 7922 59264 7930 59328
rect 7610 59263 7930 59264
rect 4613 59258 4679 59261
rect 5441 59258 5507 59261
rect 4613 59256 5507 59258
rect 4613 59200 4618 59256
rect 4674 59200 5446 59256
rect 5502 59200 5507 59256
rect 4613 59198 5507 59200
rect 4613 59195 4679 59198
rect 5441 59195 5507 59198
rect 7230 58924 7236 58988
rect 7300 58986 7306 58988
rect 7373 58986 7439 58989
rect 7300 58984 7439 58986
rect 7300 58928 7378 58984
rect 7434 58928 7439 58984
rect 7300 58926 7439 58928
rect 7300 58924 7306 58926
rect 7373 58923 7439 58926
rect 4981 58850 5047 58853
rect 8293 58850 8359 58853
rect 4981 58848 8359 58850
rect 4981 58792 4986 58848
rect 5042 58792 8298 58848
rect 8354 58792 8359 58848
rect 4981 58790 8359 58792
rect 4981 58787 5047 58790
rect 8293 58787 8359 58790
rect 4277 58784 4597 58785
rect 0 58714 480 58744
rect 4277 58720 4285 58784
rect 4349 58720 4365 58784
rect 4429 58720 4445 58784
rect 4509 58720 4525 58784
rect 4589 58720 4597 58784
rect 4277 58719 4597 58720
rect 3550 58714 3556 58716
rect 0 58654 3556 58714
rect 0 58624 480 58654
rect 3550 58652 3556 58654
rect 3620 58652 3626 58716
rect 10550 58714 10610 59742
rect 10777 59739 10843 59742
rect 19520 59712 20000 59742
rect 10685 59530 10751 59533
rect 11605 59530 11671 59533
rect 13997 59530 14063 59533
rect 10685 59528 14063 59530
rect 10685 59472 10690 59528
rect 10746 59472 11610 59528
rect 11666 59472 14002 59528
rect 14058 59472 14063 59528
rect 10685 59470 14063 59472
rect 10685 59467 10751 59470
rect 11605 59467 11671 59470
rect 13997 59467 14063 59470
rect 14277 59328 14597 59329
rect 14277 59264 14285 59328
rect 14349 59264 14365 59328
rect 14429 59264 14445 59328
rect 14509 59264 14525 59328
rect 14589 59264 14597 59328
rect 14277 59263 14597 59264
rect 10685 59122 10751 59125
rect 14825 59122 14891 59125
rect 10685 59120 14891 59122
rect 10685 59064 10690 59120
rect 10746 59064 14830 59120
rect 14886 59064 14891 59120
rect 10685 59062 14891 59064
rect 10685 59059 10751 59062
rect 14825 59059 14891 59062
rect 16481 59122 16547 59125
rect 19520 59122 20000 59152
rect 16481 59120 20000 59122
rect 16481 59064 16486 59120
rect 16542 59064 20000 59120
rect 16481 59062 20000 59064
rect 16481 59059 16547 59062
rect 19520 59032 20000 59062
rect 10944 58784 11264 58785
rect 10944 58720 10952 58784
rect 11016 58720 11032 58784
rect 11096 58720 11112 58784
rect 11176 58720 11192 58784
rect 11256 58720 11264 58784
rect 10944 58719 11264 58720
rect 17610 58784 17930 58785
rect 17610 58720 17618 58784
rect 17682 58720 17698 58784
rect 17762 58720 17778 58784
rect 17842 58720 17858 58784
rect 17922 58720 17930 58784
rect 17610 58719 17930 58720
rect 10412 58654 10610 58714
rect 6637 58578 6703 58581
rect 8569 58578 8635 58581
rect 6637 58576 8635 58578
rect 6637 58520 6642 58576
rect 6698 58520 8574 58576
rect 8630 58520 8635 58576
rect 6637 58518 8635 58520
rect 6637 58515 6703 58518
rect 8569 58515 8635 58518
rect 10412 58445 10472 58654
rect 10409 58440 10475 58445
rect 10409 58384 10414 58440
rect 10470 58384 10475 58440
rect 10409 58379 10475 58384
rect 16389 58442 16455 58445
rect 19520 58442 20000 58472
rect 16389 58440 20000 58442
rect 16389 58384 16394 58440
rect 16450 58384 20000 58440
rect 16389 58382 20000 58384
rect 16389 58379 16455 58382
rect 19520 58352 20000 58382
rect 7610 58240 7930 58241
rect 7610 58176 7618 58240
rect 7682 58176 7698 58240
rect 7762 58176 7778 58240
rect 7842 58176 7858 58240
rect 7922 58176 7930 58240
rect 7610 58175 7930 58176
rect 14277 58240 14597 58241
rect 14277 58176 14285 58240
rect 14349 58176 14365 58240
rect 14429 58176 14445 58240
rect 14509 58176 14525 58240
rect 14589 58176 14597 58240
rect 14277 58175 14597 58176
rect 2313 58170 2379 58173
rect 5533 58170 5599 58173
rect 2313 58168 5599 58170
rect 2313 58112 2318 58168
rect 2374 58112 5538 58168
rect 5594 58112 5599 58168
rect 2313 58110 5599 58112
rect 2313 58107 2379 58110
rect 5533 58107 5599 58110
rect 7557 58034 7623 58037
rect 9581 58034 9647 58037
rect 14089 58034 14155 58037
rect 7557 58032 14155 58034
rect 7557 57976 7562 58032
rect 7618 57976 9586 58032
rect 9642 57976 14094 58032
rect 14150 57976 14155 58032
rect 7557 57974 14155 57976
rect 7557 57971 7623 57974
rect 9581 57971 9647 57974
rect 14089 57971 14155 57974
rect 14825 58034 14891 58037
rect 16297 58034 16363 58037
rect 14825 58032 16363 58034
rect 14825 57976 14830 58032
rect 14886 57976 16302 58032
rect 16358 57976 16363 58032
rect 14825 57974 16363 57976
rect 14825 57971 14891 57974
rect 16297 57971 16363 57974
rect 0 57898 480 57928
rect 3969 57898 4035 57901
rect 0 57896 4035 57898
rect 0 57840 3974 57896
rect 4030 57840 4035 57896
rect 0 57838 4035 57840
rect 0 57808 480 57838
rect 3969 57835 4035 57838
rect 7833 57898 7899 57901
rect 11145 57898 11211 57901
rect 7833 57896 11211 57898
rect 7833 57840 7838 57896
rect 7894 57840 11150 57896
rect 11206 57840 11211 57896
rect 7833 57838 11211 57840
rect 7833 57835 7899 57838
rect 11145 57835 11211 57838
rect 15837 57898 15903 57901
rect 15837 57896 18154 57898
rect 15837 57840 15842 57896
rect 15898 57840 18154 57896
rect 15837 57838 18154 57840
rect 15837 57835 15903 57838
rect 11605 57762 11671 57765
rect 11830 57762 11836 57764
rect 11605 57760 11836 57762
rect 11605 57704 11610 57760
rect 11666 57704 11836 57760
rect 11605 57702 11836 57704
rect 11605 57699 11671 57702
rect 11830 57700 11836 57702
rect 11900 57700 11906 57764
rect 18094 57762 18154 57838
rect 19520 57762 20000 57792
rect 18094 57702 20000 57762
rect 4277 57696 4597 57697
rect 4277 57632 4285 57696
rect 4349 57632 4365 57696
rect 4429 57632 4445 57696
rect 4509 57632 4525 57696
rect 4589 57632 4597 57696
rect 4277 57631 4597 57632
rect 10944 57696 11264 57697
rect 10944 57632 10952 57696
rect 11016 57632 11032 57696
rect 11096 57632 11112 57696
rect 11176 57632 11192 57696
rect 11256 57632 11264 57696
rect 10944 57631 11264 57632
rect 17610 57696 17930 57697
rect 17610 57632 17618 57696
rect 17682 57632 17698 57696
rect 17762 57632 17778 57696
rect 17842 57632 17858 57696
rect 17922 57632 17930 57696
rect 19520 57672 20000 57702
rect 17610 57631 17930 57632
rect 10358 57428 10364 57492
rect 10428 57490 10434 57492
rect 10961 57490 11027 57493
rect 10428 57488 11027 57490
rect 10428 57432 10966 57488
rect 11022 57432 11027 57488
rect 10428 57430 11027 57432
rect 10428 57428 10434 57430
rect 10961 57427 11027 57430
rect 3049 57354 3115 57357
rect 5625 57354 5691 57357
rect 3049 57352 5691 57354
rect 3049 57296 3054 57352
rect 3110 57296 5630 57352
rect 5686 57296 5691 57352
rect 3049 57294 5691 57296
rect 3049 57291 3115 57294
rect 5625 57291 5691 57294
rect 7925 57354 7991 57357
rect 9438 57354 9444 57356
rect 7925 57352 9444 57354
rect 7925 57296 7930 57352
rect 7986 57296 9444 57352
rect 7925 57294 9444 57296
rect 7925 57291 7991 57294
rect 9438 57292 9444 57294
rect 9508 57292 9514 57356
rect 12985 57354 13051 57357
rect 16021 57354 16087 57357
rect 12985 57352 16087 57354
rect 12985 57296 12990 57352
rect 13046 57296 16026 57352
rect 16082 57296 16087 57352
rect 12985 57294 16087 57296
rect 12985 57291 13051 57294
rect 16021 57291 16087 57294
rect 7610 57152 7930 57153
rect 0 57082 480 57112
rect 7610 57088 7618 57152
rect 7682 57088 7698 57152
rect 7762 57088 7778 57152
rect 7842 57088 7858 57152
rect 7922 57088 7930 57152
rect 7610 57087 7930 57088
rect 14277 57152 14597 57153
rect 14277 57088 14285 57152
rect 14349 57088 14365 57152
rect 14429 57088 14445 57152
rect 14509 57088 14525 57152
rect 14589 57088 14597 57152
rect 14277 57087 14597 57088
rect 1577 57082 1643 57085
rect 0 57080 1643 57082
rect 0 57024 1582 57080
rect 1638 57024 1643 57080
rect 0 57022 1643 57024
rect 0 56992 480 57022
rect 1577 57019 1643 57022
rect 9673 57080 9739 57085
rect 9673 57024 9678 57080
rect 9734 57024 9739 57080
rect 9673 57019 9739 57024
rect 15469 57082 15535 57085
rect 19520 57082 20000 57112
rect 15469 57080 20000 57082
rect 15469 57024 15474 57080
rect 15530 57024 20000 57080
rect 15469 57022 20000 57024
rect 15469 57019 15535 57022
rect 9676 56946 9736 57019
rect 19520 56992 20000 57022
rect 12433 56946 12499 56949
rect 9676 56944 12499 56946
rect 9676 56888 12438 56944
rect 12494 56888 12499 56944
rect 9676 56886 12499 56888
rect 12433 56883 12499 56886
rect 13721 56810 13787 56813
rect 14917 56810 14983 56813
rect 13721 56808 14983 56810
rect 13721 56752 13726 56808
rect 13782 56752 14922 56808
rect 14978 56752 14983 56808
rect 13721 56750 14983 56752
rect 13721 56747 13787 56750
rect 14917 56747 14983 56750
rect 12566 56612 12572 56676
rect 12636 56674 12642 56676
rect 16665 56674 16731 56677
rect 12636 56672 16731 56674
rect 12636 56616 16670 56672
rect 16726 56616 16731 56672
rect 12636 56614 16731 56616
rect 12636 56612 12642 56614
rect 16665 56611 16731 56614
rect 4277 56608 4597 56609
rect 4277 56544 4285 56608
rect 4349 56544 4365 56608
rect 4429 56544 4445 56608
rect 4509 56544 4525 56608
rect 4589 56544 4597 56608
rect 4277 56543 4597 56544
rect 10944 56608 11264 56609
rect 10944 56544 10952 56608
rect 11016 56544 11032 56608
rect 11096 56544 11112 56608
rect 11176 56544 11192 56608
rect 11256 56544 11264 56608
rect 10944 56543 11264 56544
rect 17610 56608 17930 56609
rect 17610 56544 17618 56608
rect 17682 56544 17698 56608
rect 17762 56544 17778 56608
rect 17842 56544 17858 56608
rect 17922 56544 17930 56608
rect 17610 56543 17930 56544
rect 12065 56538 12131 56541
rect 12382 56538 12388 56540
rect 12065 56536 12388 56538
rect 12065 56480 12070 56536
rect 12126 56480 12388 56536
rect 12065 56478 12388 56480
rect 12065 56475 12131 56478
rect 12382 56476 12388 56478
rect 12452 56538 12458 56540
rect 12709 56538 12775 56541
rect 12452 56536 12775 56538
rect 12452 56480 12714 56536
rect 12770 56480 12775 56536
rect 12452 56478 12775 56480
rect 12452 56476 12458 56478
rect 12709 56475 12775 56478
rect 9070 56340 9076 56404
rect 9140 56402 9146 56404
rect 9857 56402 9923 56405
rect 10409 56404 10475 56405
rect 9140 56400 9923 56402
rect 9140 56344 9862 56400
rect 9918 56344 9923 56400
rect 9140 56342 9923 56344
rect 9140 56340 9146 56342
rect 9857 56339 9923 56342
rect 10358 56340 10364 56404
rect 10428 56402 10475 56404
rect 16205 56402 16271 56405
rect 19520 56402 20000 56432
rect 10428 56400 10520 56402
rect 10470 56344 10520 56400
rect 10428 56342 10520 56344
rect 16205 56400 20000 56402
rect 16205 56344 16210 56400
rect 16266 56344 20000 56400
rect 16205 56342 20000 56344
rect 10428 56340 10475 56342
rect 10409 56339 10475 56340
rect 16205 56339 16271 56342
rect 19520 56312 20000 56342
rect 0 56266 480 56296
rect 3693 56266 3759 56269
rect 0 56264 3759 56266
rect 0 56208 3698 56264
rect 3754 56208 3759 56264
rect 0 56206 3759 56208
rect 0 56176 480 56206
rect 3693 56203 3759 56206
rect 4797 56266 4863 56269
rect 8886 56266 8892 56268
rect 4797 56264 8892 56266
rect 4797 56208 4802 56264
rect 4858 56208 8892 56264
rect 4797 56206 8892 56208
rect 4797 56203 4863 56206
rect 8886 56204 8892 56206
rect 8956 56204 8962 56268
rect 9489 56266 9555 56269
rect 11697 56266 11763 56269
rect 13721 56266 13787 56269
rect 9489 56264 13787 56266
rect 9489 56208 9494 56264
rect 9550 56208 11702 56264
rect 11758 56208 13726 56264
rect 13782 56208 13787 56264
rect 9489 56206 13787 56208
rect 9489 56203 9555 56206
rect 11697 56203 11763 56206
rect 13721 56203 13787 56206
rect 5073 56130 5139 56133
rect 5574 56130 5580 56132
rect 5073 56128 5580 56130
rect 5073 56072 5078 56128
rect 5134 56072 5580 56128
rect 5073 56070 5580 56072
rect 5073 56067 5139 56070
rect 5574 56068 5580 56070
rect 5644 56068 5650 56132
rect 10685 56130 10751 56133
rect 10961 56130 11027 56133
rect 10685 56128 11027 56130
rect 10685 56072 10690 56128
rect 10746 56072 10966 56128
rect 11022 56072 11027 56128
rect 10685 56070 11027 56072
rect 10685 56067 10751 56070
rect 10961 56067 11027 56070
rect 7610 56064 7930 56065
rect 7610 56000 7618 56064
rect 7682 56000 7698 56064
rect 7762 56000 7778 56064
rect 7842 56000 7858 56064
rect 7922 56000 7930 56064
rect 7610 55999 7930 56000
rect 14277 56064 14597 56065
rect 14277 56000 14285 56064
rect 14349 56000 14365 56064
rect 14429 56000 14445 56064
rect 14509 56000 14525 56064
rect 14589 56000 14597 56064
rect 14277 55999 14597 56000
rect 3182 55932 3188 55996
rect 3252 55994 3258 55996
rect 7005 55994 7071 55997
rect 3252 55992 7071 55994
rect 3252 55936 7010 55992
rect 7066 55936 7071 55992
rect 3252 55934 7071 55936
rect 3252 55932 3258 55934
rect 7005 55931 7071 55934
rect 8293 55994 8359 55997
rect 12525 55994 12591 55997
rect 8293 55992 12591 55994
rect 8293 55936 8298 55992
rect 8354 55936 12530 55992
rect 12586 55936 12591 55992
rect 8293 55934 12591 55936
rect 8293 55931 8359 55934
rect 12525 55931 12591 55934
rect 8518 55796 8524 55860
rect 8588 55858 8594 55860
rect 8845 55858 8911 55861
rect 17493 55858 17559 55861
rect 8588 55856 17559 55858
rect 8588 55800 8850 55856
rect 8906 55800 17498 55856
rect 17554 55800 17559 55856
rect 8588 55798 17559 55800
rect 8588 55796 8594 55798
rect 8845 55795 8911 55798
rect 17493 55795 17559 55798
rect 3734 55660 3740 55724
rect 3804 55722 3810 55724
rect 5206 55722 5212 55724
rect 3804 55662 5212 55722
rect 3804 55660 3810 55662
rect 5206 55660 5212 55662
rect 5276 55660 5282 55724
rect 5942 55660 5948 55724
rect 6012 55722 6018 55724
rect 6269 55722 6335 55725
rect 6012 55720 6335 55722
rect 6012 55664 6274 55720
rect 6330 55664 6335 55720
rect 6012 55662 6335 55664
rect 6012 55660 6018 55662
rect 6269 55659 6335 55662
rect 9489 55722 9555 55725
rect 11145 55722 11211 55725
rect 9489 55720 11211 55722
rect 9489 55664 9494 55720
rect 9550 55664 11150 55720
rect 11206 55664 11211 55720
rect 9489 55662 11211 55664
rect 9489 55659 9555 55662
rect 11145 55659 11211 55662
rect 16389 55722 16455 55725
rect 19520 55722 20000 55752
rect 16389 55720 20000 55722
rect 16389 55664 16394 55720
rect 16450 55664 20000 55720
rect 16389 55662 20000 55664
rect 16389 55659 16455 55662
rect 19520 55632 20000 55662
rect 4277 55520 4597 55521
rect 0 55450 480 55480
rect 4277 55456 4285 55520
rect 4349 55456 4365 55520
rect 4429 55456 4445 55520
rect 4509 55456 4525 55520
rect 4589 55456 4597 55520
rect 4277 55455 4597 55456
rect 10944 55520 11264 55521
rect 10944 55456 10952 55520
rect 11016 55456 11032 55520
rect 11096 55456 11112 55520
rect 11176 55456 11192 55520
rect 11256 55456 11264 55520
rect 10944 55455 11264 55456
rect 17610 55520 17930 55521
rect 17610 55456 17618 55520
rect 17682 55456 17698 55520
rect 17762 55456 17778 55520
rect 17842 55456 17858 55520
rect 17922 55456 17930 55520
rect 17610 55455 17930 55456
rect 3918 55450 3924 55452
rect 0 55390 3924 55450
rect 0 55360 480 55390
rect 3918 55388 3924 55390
rect 3988 55388 3994 55452
rect 8702 55388 8708 55452
rect 8772 55450 8778 55452
rect 9673 55450 9739 55453
rect 8772 55448 9739 55450
rect 8772 55392 9678 55448
rect 9734 55392 9739 55448
rect 8772 55390 9739 55392
rect 8772 55388 8778 55390
rect 9673 55387 9739 55390
rect 13721 55450 13787 55453
rect 14365 55450 14431 55453
rect 17125 55450 17191 55453
rect 13721 55448 17191 55450
rect 13721 55392 13726 55448
rect 13782 55392 14370 55448
rect 14426 55392 17130 55448
rect 17186 55392 17191 55448
rect 13721 55390 17191 55392
rect 13721 55387 13787 55390
rect 14365 55387 14431 55390
rect 17125 55387 17191 55390
rect 11513 55314 11579 55317
rect 11646 55314 11652 55316
rect 11513 55312 11652 55314
rect 11513 55256 11518 55312
rect 11574 55256 11652 55312
rect 11513 55254 11652 55256
rect 11513 55251 11579 55254
rect 11646 55252 11652 55254
rect 11716 55252 11722 55316
rect 14181 55314 14247 55317
rect 14181 55312 15578 55314
rect 14181 55256 14186 55312
rect 14242 55256 15578 55312
rect 14181 55254 15578 55256
rect 14181 55251 14247 55254
rect 8886 55116 8892 55180
rect 8956 55178 8962 55180
rect 11881 55178 11947 55181
rect 8956 55176 11947 55178
rect 8956 55120 11886 55176
rect 11942 55120 11947 55176
rect 8956 55118 11947 55120
rect 8956 55116 8962 55118
rect 11838 55115 11947 55118
rect 12014 55116 12020 55180
rect 12084 55178 12090 55180
rect 12566 55178 12572 55180
rect 12084 55118 12572 55178
rect 12084 55116 12090 55118
rect 12566 55116 12572 55118
rect 12636 55116 12642 55180
rect 15285 55178 15351 55181
rect 13678 55176 15351 55178
rect 13678 55120 15290 55176
rect 15346 55120 15351 55176
rect 13678 55118 15351 55120
rect 2998 54980 3004 55044
rect 3068 55042 3074 55044
rect 4429 55042 4495 55045
rect 3068 55040 4495 55042
rect 3068 54984 4434 55040
rect 4490 54984 4495 55040
rect 3068 54982 4495 54984
rect 3068 54980 3074 54982
rect 4429 54979 4495 54982
rect 6126 54980 6132 55044
rect 6196 55042 6202 55044
rect 7281 55042 7347 55045
rect 6196 55040 7347 55042
rect 6196 54984 7286 55040
rect 7342 54984 7347 55040
rect 6196 54982 7347 54984
rect 6196 54980 6202 54982
rect 7281 54979 7347 54982
rect 8845 55042 8911 55045
rect 9254 55042 9260 55044
rect 8845 55040 9260 55042
rect 8845 54984 8850 55040
rect 8906 54984 9260 55040
rect 8845 54982 9260 54984
rect 8845 54979 8911 54982
rect 9254 54980 9260 54982
rect 9324 54980 9330 55044
rect 11838 55042 11898 55115
rect 13678 55042 13738 55118
rect 15285 55115 15351 55118
rect 11838 54982 13738 55042
rect 15009 55042 15075 55045
rect 15377 55042 15443 55045
rect 15009 55040 15443 55042
rect 15009 54984 15014 55040
rect 15070 54984 15382 55040
rect 15438 54984 15443 55040
rect 15009 54982 15443 54984
rect 15518 55042 15578 55254
rect 19520 55042 20000 55072
rect 15518 54982 20000 55042
rect 15009 54979 15075 54982
rect 15377 54979 15443 54982
rect 7610 54976 7930 54977
rect 7610 54912 7618 54976
rect 7682 54912 7698 54976
rect 7762 54912 7778 54976
rect 7842 54912 7858 54976
rect 7922 54912 7930 54976
rect 7610 54911 7930 54912
rect 14277 54976 14597 54977
rect 14277 54912 14285 54976
rect 14349 54912 14365 54976
rect 14429 54912 14445 54976
rect 14509 54912 14525 54976
rect 14589 54912 14597 54976
rect 19520 54952 20000 54982
rect 14277 54911 14597 54912
rect 9806 54844 9812 54908
rect 9876 54906 9882 54908
rect 12382 54906 12388 54908
rect 9876 54846 12388 54906
rect 9876 54844 9882 54846
rect 12382 54844 12388 54846
rect 12452 54844 12458 54908
rect 7833 54770 7899 54773
rect 14641 54770 14707 54773
rect 7833 54768 14707 54770
rect 7833 54712 7838 54768
rect 7894 54712 14646 54768
rect 14702 54712 14707 54768
rect 7833 54710 14707 54712
rect 7833 54707 7899 54710
rect 14641 54707 14707 54710
rect 0 54634 480 54664
rect 2313 54634 2379 54637
rect 0 54632 2379 54634
rect 0 54576 2318 54632
rect 2374 54576 2379 54632
rect 0 54574 2379 54576
rect 0 54544 480 54574
rect 2313 54571 2379 54574
rect 15561 54634 15627 54637
rect 15561 54632 18154 54634
rect 15561 54576 15566 54632
rect 15622 54576 18154 54632
rect 15561 54574 18154 54576
rect 15561 54571 15627 54574
rect 8385 54498 8451 54501
rect 6502 54496 8451 54498
rect 6502 54440 8390 54496
rect 8446 54440 8451 54496
rect 6502 54438 8451 54440
rect 4277 54432 4597 54433
rect 4277 54368 4285 54432
rect 4349 54368 4365 54432
rect 4429 54368 4445 54432
rect 4509 54368 4525 54432
rect 4589 54368 4597 54432
rect 4277 54367 4597 54368
rect 5758 54028 5764 54092
rect 5828 54090 5834 54092
rect 6177 54090 6243 54093
rect 6502 54090 6562 54438
rect 8385 54435 8451 54438
rect 10944 54432 11264 54433
rect 10944 54368 10952 54432
rect 11016 54368 11032 54432
rect 11096 54368 11112 54432
rect 11176 54368 11192 54432
rect 11256 54368 11264 54432
rect 10944 54367 11264 54368
rect 17610 54432 17930 54433
rect 17610 54368 17618 54432
rect 17682 54368 17698 54432
rect 17762 54368 17778 54432
rect 17842 54368 17858 54432
rect 17922 54368 17930 54432
rect 17610 54367 17930 54368
rect 6729 54364 6795 54365
rect 6678 54300 6684 54364
rect 6748 54362 6795 54364
rect 18094 54362 18154 54574
rect 19520 54362 20000 54392
rect 6748 54360 6840 54362
rect 6790 54304 6840 54360
rect 6748 54302 6840 54304
rect 18094 54302 20000 54362
rect 6748 54300 6795 54302
rect 6729 54299 6795 54300
rect 19520 54272 20000 54302
rect 6729 54226 6795 54229
rect 9213 54226 9279 54229
rect 9949 54226 10015 54229
rect 6729 54224 10015 54226
rect 6729 54168 6734 54224
rect 6790 54168 9218 54224
rect 9274 54168 9954 54224
rect 10010 54168 10015 54224
rect 6729 54166 10015 54168
rect 6729 54163 6795 54166
rect 9213 54163 9279 54166
rect 9949 54163 10015 54166
rect 10961 54226 11027 54229
rect 12341 54228 12407 54229
rect 11830 54226 11836 54228
rect 10961 54224 11836 54226
rect 10961 54168 10966 54224
rect 11022 54168 11836 54224
rect 10961 54166 11836 54168
rect 10961 54163 11027 54166
rect 11830 54164 11836 54166
rect 11900 54164 11906 54228
rect 12341 54226 12388 54228
rect 12300 54224 12388 54226
rect 12300 54168 12346 54224
rect 12300 54166 12388 54168
rect 12341 54164 12388 54166
rect 12452 54164 12458 54228
rect 16021 54226 16087 54229
rect 16021 54224 16130 54226
rect 16021 54168 16026 54224
rect 16082 54168 16130 54224
rect 12341 54163 12407 54164
rect 16021 54163 16130 54168
rect 5828 54088 6562 54090
rect 5828 54032 6182 54088
rect 6238 54032 6562 54088
rect 5828 54030 6562 54032
rect 6729 54090 6795 54093
rect 7230 54090 7236 54092
rect 6729 54088 7236 54090
rect 6729 54032 6734 54088
rect 6790 54032 7236 54088
rect 6729 54030 7236 54032
rect 5828 54028 5834 54030
rect 6177 54027 6243 54030
rect 6729 54027 6795 54030
rect 7230 54028 7236 54030
rect 7300 54028 7306 54092
rect 10501 54090 10567 54093
rect 12617 54090 12683 54093
rect 10501 54088 12683 54090
rect 10501 54032 10506 54088
rect 10562 54032 12622 54088
rect 12678 54032 12683 54088
rect 10501 54030 12683 54032
rect 10501 54027 10567 54030
rect 12617 54027 12683 54030
rect 6361 53954 6427 53957
rect 6494 53954 6500 53956
rect 6361 53952 6500 53954
rect 6361 53896 6366 53952
rect 6422 53896 6500 53952
rect 6361 53894 6500 53896
rect 6361 53891 6427 53894
rect 6494 53892 6500 53894
rect 6564 53892 6570 53956
rect 7230 53892 7236 53956
rect 7300 53954 7306 53956
rect 7373 53954 7439 53957
rect 7300 53952 7439 53954
rect 7300 53896 7378 53952
rect 7434 53896 7439 53952
rect 7300 53894 7439 53896
rect 7300 53892 7306 53894
rect 7373 53891 7439 53894
rect 9489 53954 9555 53957
rect 11421 53954 11487 53957
rect 11830 53954 11836 53956
rect 9489 53952 9828 53954
rect 9489 53896 9494 53952
rect 9550 53896 9828 53952
rect 9489 53894 9828 53896
rect 9489 53891 9555 53894
rect 7610 53888 7930 53889
rect 0 53818 480 53848
rect 7610 53824 7618 53888
rect 7682 53824 7698 53888
rect 7762 53824 7778 53888
rect 7842 53824 7858 53888
rect 7922 53824 7930 53888
rect 7610 53823 7930 53824
rect 1853 53818 1919 53821
rect 0 53816 1919 53818
rect 0 53760 1858 53816
rect 1914 53760 1919 53816
rect 0 53758 1919 53760
rect 9768 53818 9828 53894
rect 11421 53952 11836 53954
rect 11421 53896 11426 53952
rect 11482 53896 11836 53952
rect 11421 53894 11836 53896
rect 11421 53891 11487 53894
rect 11830 53892 11836 53894
rect 11900 53892 11906 53956
rect 14277 53888 14597 53889
rect 14277 53824 14285 53888
rect 14349 53824 14365 53888
rect 14429 53824 14445 53888
rect 14509 53824 14525 53888
rect 14589 53824 14597 53888
rect 14277 53823 14597 53824
rect 13118 53818 13124 53820
rect 9768 53758 13124 53818
rect 0 53728 480 53758
rect 1853 53755 1919 53758
rect 13118 53756 13124 53758
rect 13188 53756 13194 53820
rect 16070 53818 16130 54163
rect 16070 53758 16176 53818
rect 8845 53682 8911 53685
rect 9438 53682 9444 53684
rect 8845 53680 9444 53682
rect 8845 53624 8850 53680
rect 8906 53624 9444 53680
rect 8845 53622 9444 53624
rect 8845 53619 8911 53622
rect 9438 53620 9444 53622
rect 9508 53620 9514 53684
rect 10593 53682 10659 53685
rect 14733 53682 14799 53685
rect 10593 53680 14799 53682
rect 10593 53624 10598 53680
rect 10654 53624 14738 53680
rect 14794 53624 14799 53680
rect 10593 53622 14799 53624
rect 16116 53682 16176 53758
rect 19520 53682 20000 53712
rect 16116 53622 20000 53682
rect 10593 53619 10659 53622
rect 14733 53619 14799 53622
rect 19520 53592 20000 53622
rect 4337 53546 4403 53549
rect 4337 53544 4722 53546
rect 4337 53488 4342 53544
rect 4398 53488 4722 53544
rect 4337 53486 4722 53488
rect 4337 53483 4403 53486
rect 4277 53344 4597 53345
rect 4277 53280 4285 53344
rect 4349 53280 4365 53344
rect 4429 53280 4445 53344
rect 4509 53280 4525 53344
rect 4589 53280 4597 53344
rect 4277 53279 4597 53280
rect 0 53138 480 53168
rect 2865 53138 2931 53141
rect 0 53136 2931 53138
rect 0 53080 2870 53136
rect 2926 53080 2931 53136
rect 0 53078 2931 53080
rect 0 53048 480 53078
rect 2865 53075 2931 53078
rect 4521 53138 4587 53141
rect 4662 53138 4722 53486
rect 11605 53410 11671 53413
rect 15469 53410 15535 53413
rect 16573 53410 16639 53413
rect 17166 53410 17172 53412
rect 11605 53408 15535 53410
rect 11605 53352 11610 53408
rect 11666 53352 15474 53408
rect 15530 53352 15535 53408
rect 11605 53350 15535 53352
rect 11605 53347 11671 53350
rect 15469 53347 15535 53350
rect 15702 53408 17172 53410
rect 15702 53352 16578 53408
rect 16634 53352 17172 53408
rect 15702 53350 17172 53352
rect 10944 53344 11264 53345
rect 10944 53280 10952 53344
rect 11016 53280 11032 53344
rect 11096 53280 11112 53344
rect 11176 53280 11192 53344
rect 11256 53280 11264 53344
rect 10944 53279 11264 53280
rect 15702 53274 15762 53350
rect 16573 53347 16639 53350
rect 17166 53348 17172 53350
rect 17236 53410 17242 53412
rect 17401 53410 17467 53413
rect 17236 53408 17467 53410
rect 17236 53352 17406 53408
rect 17462 53352 17467 53408
rect 17236 53350 17467 53352
rect 17236 53348 17242 53350
rect 17401 53347 17467 53350
rect 17610 53344 17930 53345
rect 17610 53280 17618 53344
rect 17682 53280 17698 53344
rect 17762 53280 17778 53344
rect 17842 53280 17858 53344
rect 17922 53280 17930 53344
rect 17610 53279 17930 53280
rect 11470 53214 15762 53274
rect 4521 53136 4722 53138
rect 4521 53080 4526 53136
rect 4582 53080 4722 53136
rect 4521 53078 4722 53080
rect 4521 53075 4587 53078
rect 5942 53076 5948 53140
rect 6012 53138 6018 53140
rect 9949 53138 10015 53141
rect 6012 53136 10015 53138
rect 6012 53080 9954 53136
rect 10010 53080 10015 53136
rect 6012 53078 10015 53080
rect 6012 53076 6018 53078
rect 9949 53075 10015 53078
rect 10225 53138 10291 53141
rect 11470 53138 11530 53214
rect 10225 53136 11530 53138
rect 10225 53080 10230 53136
rect 10286 53080 11530 53136
rect 10225 53078 11530 53080
rect 11789 53138 11855 53141
rect 16849 53138 16915 53141
rect 11789 53136 16915 53138
rect 11789 53080 11794 53136
rect 11850 53080 16854 53136
rect 16910 53080 16915 53136
rect 11789 53078 16915 53080
rect 10225 53075 10291 53078
rect 11789 53075 11855 53078
rect 16849 53075 16915 53078
rect 5625 53002 5691 53005
rect 6310 53002 6316 53004
rect 5625 53000 6316 53002
rect 5625 52944 5630 53000
rect 5686 52944 6316 53000
rect 5625 52942 6316 52944
rect 5625 52939 5691 52942
rect 6310 52940 6316 52942
rect 6380 52940 6386 53004
rect 12893 53002 12959 53005
rect 16757 53002 16823 53005
rect 17953 53002 18019 53005
rect 12893 53000 18019 53002
rect 12893 52944 12898 53000
rect 12954 52944 16762 53000
rect 16818 52944 17958 53000
rect 18014 52944 18019 53000
rect 12893 52942 18019 52944
rect 12893 52939 12959 52942
rect 16757 52939 16823 52942
rect 17953 52939 18019 52942
rect 8109 52866 8175 52869
rect 9673 52866 9739 52869
rect 10358 52866 10364 52868
rect 8109 52864 10364 52866
rect 8109 52808 8114 52864
rect 8170 52808 9678 52864
rect 9734 52808 10364 52864
rect 8109 52806 10364 52808
rect 8109 52803 8175 52806
rect 9673 52803 9739 52806
rect 10358 52804 10364 52806
rect 10428 52804 10434 52868
rect 14958 52804 14964 52868
rect 15028 52866 15034 52868
rect 15326 52866 15332 52868
rect 15028 52806 15332 52866
rect 15028 52804 15034 52806
rect 15326 52804 15332 52806
rect 15396 52804 15402 52868
rect 15745 52866 15811 52869
rect 19520 52866 20000 52896
rect 15745 52864 20000 52866
rect 15745 52808 15750 52864
rect 15806 52808 20000 52864
rect 15745 52806 20000 52808
rect 15745 52803 15811 52806
rect 7610 52800 7930 52801
rect 7610 52736 7618 52800
rect 7682 52736 7698 52800
rect 7762 52736 7778 52800
rect 7842 52736 7858 52800
rect 7922 52736 7930 52800
rect 7610 52735 7930 52736
rect 14277 52800 14597 52801
rect 14277 52736 14285 52800
rect 14349 52736 14365 52800
rect 14429 52736 14445 52800
rect 14509 52736 14525 52800
rect 14589 52736 14597 52800
rect 19520 52776 20000 52806
rect 14277 52735 14597 52736
rect 3141 52730 3207 52733
rect 6085 52730 6151 52733
rect 3141 52728 6151 52730
rect 3141 52672 3146 52728
rect 3202 52672 6090 52728
rect 6146 52672 6151 52728
rect 3141 52670 6151 52672
rect 3141 52667 3207 52670
rect 6085 52667 6151 52670
rect 8201 52730 8267 52733
rect 8518 52730 8524 52732
rect 8201 52728 8524 52730
rect 8201 52672 8206 52728
rect 8262 52672 8524 52728
rect 8201 52670 8524 52672
rect 8201 52667 8267 52670
rect 8518 52668 8524 52670
rect 8588 52668 8594 52732
rect 11881 52730 11947 52733
rect 12566 52730 12572 52732
rect 11881 52728 12572 52730
rect 11881 52672 11886 52728
rect 11942 52672 12572 52728
rect 11881 52670 12572 52672
rect 11881 52667 11947 52670
rect 12566 52668 12572 52670
rect 12636 52668 12642 52732
rect 12893 52730 12959 52733
rect 13486 52730 13492 52732
rect 12893 52728 13492 52730
rect 12893 52672 12898 52728
rect 12954 52672 13492 52728
rect 12893 52670 13492 52672
rect 12893 52667 12959 52670
rect 13486 52668 13492 52670
rect 13556 52668 13562 52732
rect 1669 52594 1735 52597
rect 7005 52594 7071 52597
rect 1669 52592 7071 52594
rect 1669 52536 1674 52592
rect 1730 52536 7010 52592
rect 7066 52536 7071 52592
rect 1669 52534 7071 52536
rect 1669 52531 1735 52534
rect 7005 52531 7071 52534
rect 10358 52532 10364 52596
rect 10428 52594 10434 52596
rect 10593 52594 10659 52597
rect 10428 52592 10659 52594
rect 10428 52536 10598 52592
rect 10654 52536 10659 52592
rect 10428 52534 10659 52536
rect 10428 52532 10434 52534
rect 10593 52531 10659 52534
rect 8109 52458 8175 52461
rect 10133 52458 10199 52461
rect 11421 52458 11487 52461
rect 8109 52456 11487 52458
rect 8109 52400 8114 52456
rect 8170 52400 10138 52456
rect 10194 52400 11426 52456
rect 11482 52400 11487 52456
rect 8109 52398 11487 52400
rect 8109 52395 8175 52398
rect 10133 52395 10199 52398
rect 11421 52395 11487 52398
rect 13302 52396 13308 52460
rect 13372 52458 13378 52460
rect 13905 52458 13971 52461
rect 13372 52456 13971 52458
rect 13372 52400 13910 52456
rect 13966 52400 13971 52456
rect 13372 52398 13971 52400
rect 13372 52396 13378 52398
rect 13905 52395 13971 52398
rect 15377 52458 15443 52461
rect 15377 52456 18154 52458
rect 15377 52400 15382 52456
rect 15438 52400 18154 52456
rect 15377 52398 18154 52400
rect 15377 52395 15443 52398
rect 0 52322 480 52352
rect 1853 52322 1919 52325
rect 0 52320 1919 52322
rect 0 52264 1858 52320
rect 1914 52264 1919 52320
rect 0 52262 1919 52264
rect 0 52232 480 52262
rect 1853 52259 1919 52262
rect 15285 52322 15351 52325
rect 17350 52322 17356 52324
rect 15285 52320 17356 52322
rect 15285 52264 15290 52320
rect 15346 52264 17356 52320
rect 15285 52262 17356 52264
rect 15285 52259 15351 52262
rect 17350 52260 17356 52262
rect 17420 52260 17426 52324
rect 4277 52256 4597 52257
rect 4277 52192 4285 52256
rect 4349 52192 4365 52256
rect 4429 52192 4445 52256
rect 4509 52192 4525 52256
rect 4589 52192 4597 52256
rect 4277 52191 4597 52192
rect 10944 52256 11264 52257
rect 10944 52192 10952 52256
rect 11016 52192 11032 52256
rect 11096 52192 11112 52256
rect 11176 52192 11192 52256
rect 11256 52192 11264 52256
rect 10944 52191 11264 52192
rect 17610 52256 17930 52257
rect 17610 52192 17618 52256
rect 17682 52192 17698 52256
rect 17762 52192 17778 52256
rect 17842 52192 17858 52256
rect 17922 52192 17930 52256
rect 17610 52191 17930 52192
rect 5165 52186 5231 52189
rect 5574 52186 5580 52188
rect 5165 52184 5580 52186
rect 5165 52128 5170 52184
rect 5226 52128 5580 52184
rect 5165 52126 5580 52128
rect 5165 52123 5231 52126
rect 5574 52124 5580 52126
rect 5644 52124 5650 52188
rect 6177 52186 6243 52189
rect 18094 52186 18154 52398
rect 19520 52186 20000 52216
rect 6177 52184 6562 52186
rect 6177 52128 6182 52184
rect 6238 52128 6562 52184
rect 6177 52126 6562 52128
rect 18094 52126 20000 52186
rect 6177 52123 6243 52126
rect 6502 51781 6562 52126
rect 19520 52096 20000 52126
rect 13721 52050 13787 52053
rect 13721 52048 17786 52050
rect 13721 51992 13726 52048
rect 13782 51992 17786 52048
rect 13721 51990 17786 51992
rect 13721 51987 13787 51990
rect 13721 51914 13787 51917
rect 17493 51914 17559 51917
rect 13721 51912 17559 51914
rect 13721 51856 13726 51912
rect 13782 51856 17498 51912
rect 17554 51856 17559 51912
rect 13721 51854 17559 51856
rect 13721 51851 13787 51854
rect 17493 51851 17559 51854
rect 2773 51778 2839 51781
rect 3509 51778 3575 51781
rect 5533 51778 5599 51781
rect 2773 51776 5599 51778
rect 2773 51720 2778 51776
rect 2834 51720 3514 51776
rect 3570 51720 5538 51776
rect 5594 51720 5599 51776
rect 2773 51718 5599 51720
rect 6502 51776 6611 51781
rect 6502 51720 6550 51776
rect 6606 51720 6611 51776
rect 6502 51718 6611 51720
rect 2773 51715 2839 51718
rect 3509 51715 3575 51718
rect 5533 51715 5599 51718
rect 6545 51715 6611 51718
rect 9213 51778 9279 51781
rect 10542 51778 10548 51780
rect 9213 51776 10548 51778
rect 9213 51720 9218 51776
rect 9274 51720 10548 51776
rect 9213 51718 10548 51720
rect 9213 51715 9279 51718
rect 10542 51716 10548 51718
rect 10612 51716 10618 51780
rect 7610 51712 7930 51713
rect 7610 51648 7618 51712
rect 7682 51648 7698 51712
rect 7762 51648 7778 51712
rect 7842 51648 7858 51712
rect 7922 51648 7930 51712
rect 7610 51647 7930 51648
rect 14277 51712 14597 51713
rect 14277 51648 14285 51712
rect 14349 51648 14365 51712
rect 14429 51648 14445 51712
rect 14509 51648 14525 51712
rect 14589 51648 14597 51712
rect 14277 51647 14597 51648
rect 3550 51580 3556 51644
rect 3620 51642 3626 51644
rect 5257 51642 5323 51645
rect 3620 51640 5323 51642
rect 3620 51584 5262 51640
rect 5318 51584 5323 51640
rect 3620 51582 5323 51584
rect 3620 51580 3626 51582
rect 5257 51579 5323 51582
rect 6678 51580 6684 51644
rect 6748 51642 6754 51644
rect 6821 51642 6887 51645
rect 6748 51640 6887 51642
rect 6748 51584 6826 51640
rect 6882 51584 6887 51640
rect 6748 51582 6887 51584
rect 6748 51580 6754 51582
rect 6821 51579 6887 51582
rect 9581 51642 9647 51645
rect 11605 51642 11671 51645
rect 9581 51640 11671 51642
rect 9581 51584 9586 51640
rect 9642 51584 11610 51640
rect 11666 51584 11671 51640
rect 9581 51582 11671 51584
rect 9581 51579 9647 51582
rect 11605 51579 11671 51582
rect 0 51506 480 51536
rect 1485 51506 1551 51509
rect 0 51504 1551 51506
rect 0 51448 1490 51504
rect 1546 51448 1551 51504
rect 0 51446 1551 51448
rect 0 51416 480 51446
rect 1485 51443 1551 51446
rect 3366 51444 3372 51508
rect 3436 51506 3442 51508
rect 3436 51446 5458 51506
rect 3436 51444 3442 51446
rect 2998 51308 3004 51372
rect 3068 51370 3074 51372
rect 3601 51370 3667 51373
rect 3068 51368 3667 51370
rect 3068 51312 3606 51368
rect 3662 51312 3667 51368
rect 3068 51310 3667 51312
rect 3068 51308 3074 51310
rect 3601 51307 3667 51310
rect 3918 51308 3924 51372
rect 3988 51370 3994 51372
rect 3988 51310 5274 51370
rect 3988 51308 3994 51310
rect 5214 51236 5274 51310
rect 5398 51237 5458 51446
rect 5942 51444 5948 51508
rect 6012 51506 6018 51508
rect 7005 51506 7071 51509
rect 6012 51504 7071 51506
rect 6012 51448 7010 51504
rect 7066 51448 7071 51504
rect 6012 51446 7071 51448
rect 6012 51444 6018 51446
rect 5950 51370 6010 51444
rect 7005 51443 7071 51446
rect 7925 51506 7991 51509
rect 10133 51506 10199 51509
rect 7925 51504 10199 51506
rect 7925 51448 7930 51504
rect 7986 51448 10138 51504
rect 10194 51448 10199 51504
rect 7925 51446 10199 51448
rect 7925 51443 7991 51446
rect 10133 51443 10199 51446
rect 11053 51506 11119 51509
rect 11329 51506 11395 51509
rect 11053 51504 11395 51506
rect 11053 51448 11058 51504
rect 11114 51448 11334 51504
rect 11390 51448 11395 51504
rect 11053 51446 11395 51448
rect 11053 51443 11119 51446
rect 11329 51443 11395 51446
rect 12750 51444 12756 51508
rect 12820 51506 12826 51508
rect 12893 51506 12959 51509
rect 12820 51504 12959 51506
rect 12820 51448 12898 51504
rect 12954 51448 12959 51504
rect 12820 51446 12959 51448
rect 17726 51506 17786 51990
rect 19520 51506 20000 51536
rect 17726 51446 20000 51506
rect 12820 51444 12826 51446
rect 12893 51443 12959 51446
rect 19520 51416 20000 51446
rect 5582 51310 6010 51370
rect 5206 51172 5212 51236
rect 5276 51172 5282 51236
rect 5398 51232 5507 51237
rect 5398 51176 5446 51232
rect 5502 51176 5507 51232
rect 5398 51174 5507 51176
rect 5441 51171 5507 51174
rect 4277 51168 4597 51169
rect 4277 51104 4285 51168
rect 4349 51104 4365 51168
rect 4429 51104 4445 51168
rect 4509 51104 4525 51168
rect 4589 51104 4597 51168
rect 4277 51103 4597 51104
rect 4705 51098 4771 51101
rect 4889 51098 4955 51101
rect 5582 51098 5642 51310
rect 6678 51308 6684 51372
rect 6748 51370 6754 51372
rect 7046 51370 7052 51372
rect 6748 51310 7052 51370
rect 6748 51308 6754 51310
rect 7046 51308 7052 51310
rect 7116 51308 7122 51372
rect 7741 51370 7807 51373
rect 8334 51370 8340 51372
rect 7741 51368 8340 51370
rect 7741 51312 7746 51368
rect 7802 51312 8340 51368
rect 7741 51310 8340 51312
rect 7741 51307 7807 51310
rect 8334 51308 8340 51310
rect 8404 51308 8410 51372
rect 9673 51370 9739 51373
rect 10961 51370 11027 51373
rect 9673 51368 11027 51370
rect 9673 51312 9678 51368
rect 9734 51312 10966 51368
rect 11022 51312 11027 51368
rect 9673 51310 11027 51312
rect 9673 51307 9739 51310
rect 5942 51172 5948 51236
rect 6012 51234 6018 51236
rect 6453 51234 6519 51237
rect 6012 51232 6519 51234
rect 6012 51176 6458 51232
rect 6514 51176 6519 51232
rect 6012 51174 6519 51176
rect 6012 51172 6018 51174
rect 6453 51171 6519 51174
rect 7046 51172 7052 51236
rect 7116 51234 7122 51236
rect 7414 51234 7420 51236
rect 7116 51174 7420 51234
rect 7116 51172 7122 51174
rect 7414 51172 7420 51174
rect 7484 51172 7490 51236
rect 8293 51234 8359 51237
rect 8702 51234 8708 51236
rect 8293 51232 8708 51234
rect 8293 51176 8298 51232
rect 8354 51176 8708 51232
rect 8293 51174 8708 51176
rect 8293 51171 8359 51174
rect 8702 51172 8708 51174
rect 8772 51172 8778 51236
rect 8937 51234 9003 51237
rect 9254 51234 9260 51236
rect 8937 51232 9260 51234
rect 8937 51176 8942 51232
rect 8998 51176 9260 51232
rect 8937 51174 9260 51176
rect 8937 51171 9003 51174
rect 9254 51172 9260 51174
rect 9324 51172 9330 51236
rect 10780 51101 10840 51310
rect 10961 51307 11027 51310
rect 11973 51234 12039 51237
rect 16113 51234 16179 51237
rect 11516 51232 12039 51234
rect 11516 51176 11978 51232
rect 12034 51176 12039 51232
rect 11516 51174 12039 51176
rect 10944 51168 11264 51169
rect 10944 51104 10952 51168
rect 11016 51104 11032 51168
rect 11096 51104 11112 51168
rect 11176 51104 11192 51168
rect 11256 51104 11264 51168
rect 10944 51103 11264 51104
rect 4705 51096 5642 51098
rect 4705 51040 4710 51096
rect 4766 51040 4894 51096
rect 4950 51040 5642 51096
rect 4705 51038 5642 51040
rect 6729 51098 6795 51101
rect 7414 51098 7420 51100
rect 6729 51096 7420 51098
rect 6729 51040 6734 51096
rect 6790 51040 7420 51096
rect 6729 51038 7420 51040
rect 4705 51035 4771 51038
rect 4889 51035 4955 51038
rect 6729 51035 6795 51038
rect 7414 51036 7420 51038
rect 7484 51036 7490 51100
rect 9070 51098 9076 51100
rect 8342 51038 9076 51098
rect 5717 50964 5783 50965
rect 5717 50962 5764 50964
rect 5672 50960 5764 50962
rect 5672 50904 5722 50960
rect 5672 50902 5764 50904
rect 5717 50900 5764 50902
rect 5828 50900 5834 50964
rect 6821 50962 6887 50965
rect 8342 50962 8402 51038
rect 9070 51036 9076 51038
rect 9140 51098 9146 51100
rect 10317 51098 10383 51101
rect 9140 51096 10383 51098
rect 9140 51040 10322 51096
rect 10378 51040 10383 51096
rect 9140 51038 10383 51040
rect 9140 51036 9146 51038
rect 10317 51035 10383 51038
rect 10777 51096 10843 51101
rect 10777 51040 10782 51096
rect 10838 51040 10843 51096
rect 10777 51035 10843 51040
rect 6821 50960 8402 50962
rect 6821 50904 6826 50960
rect 6882 50904 8402 50960
rect 6821 50902 8402 50904
rect 8753 50962 8819 50965
rect 8937 50962 9003 50965
rect 8753 50960 9003 50962
rect 8753 50904 8758 50960
rect 8814 50904 8942 50960
rect 8998 50904 9003 50960
rect 8753 50902 9003 50904
rect 5717 50899 5783 50900
rect 6821 50899 6887 50902
rect 8753 50899 8819 50902
rect 8937 50899 9003 50902
rect 9438 50900 9444 50964
rect 9508 50962 9514 50964
rect 9508 50902 10426 50962
rect 9508 50900 9514 50902
rect 10366 50829 10426 50902
rect 10542 50900 10548 50964
rect 10612 50962 10618 50964
rect 10685 50962 10751 50965
rect 10612 50960 10751 50962
rect 10612 50904 10690 50960
rect 10746 50904 10751 50960
rect 10612 50902 10751 50904
rect 10612 50900 10618 50902
rect 10685 50899 10751 50902
rect 10961 50962 11027 50965
rect 11516 50962 11576 51174
rect 11973 51171 12039 51174
rect 16070 51232 16179 51234
rect 16070 51176 16118 51232
rect 16174 51176 16179 51232
rect 16070 51171 16179 51176
rect 11789 51098 11855 51101
rect 12934 51098 12940 51100
rect 11789 51096 12940 51098
rect 11789 51040 11794 51096
rect 11850 51040 12940 51096
rect 11789 51038 12940 51040
rect 11789 51035 11855 51038
rect 12934 51036 12940 51038
rect 13004 51036 13010 51100
rect 13353 51098 13419 51101
rect 13126 51096 13419 51098
rect 13126 51040 13358 51096
rect 13414 51040 13419 51096
rect 13126 51038 13419 51040
rect 10961 50960 11576 50962
rect 10961 50904 10966 50960
rect 11022 50904 11576 50960
rect 10961 50902 11576 50904
rect 11789 50962 11855 50965
rect 12985 50962 13051 50965
rect 11789 50960 13051 50962
rect 11789 50904 11794 50960
rect 11850 50904 12990 50960
rect 13046 50904 13051 50960
rect 11789 50902 13051 50904
rect 10961 50899 11027 50902
rect 11789 50899 11855 50902
rect 12985 50899 13051 50902
rect 5809 50826 5875 50829
rect 5942 50826 5948 50828
rect 5809 50824 5948 50826
rect 5809 50768 5814 50824
rect 5870 50768 5948 50824
rect 5809 50766 5948 50768
rect 5809 50763 5875 50766
rect 5942 50764 5948 50766
rect 6012 50764 6018 50828
rect 6862 50764 6868 50828
rect 6932 50764 6938 50828
rect 7005 50826 7071 50829
rect 10133 50826 10199 50829
rect 7005 50824 10199 50826
rect 7005 50768 7010 50824
rect 7066 50768 10138 50824
rect 10194 50768 10199 50824
rect 7005 50766 10199 50768
rect 0 50690 480 50720
rect 1710 50690 1716 50692
rect 0 50630 1716 50690
rect 0 50600 480 50630
rect 1710 50628 1716 50630
rect 1780 50628 1786 50692
rect 6678 50492 6684 50556
rect 6748 50554 6754 50556
rect 6870 50554 6930 50764
rect 7005 50763 7071 50766
rect 10133 50763 10199 50766
rect 10317 50824 10426 50829
rect 10317 50768 10322 50824
rect 10378 50768 10426 50824
rect 10317 50766 10426 50768
rect 10317 50763 10383 50766
rect 11646 50764 11652 50828
rect 11716 50764 11722 50828
rect 8753 50690 8819 50693
rect 9070 50690 9076 50692
rect 8753 50688 9076 50690
rect 8753 50632 8758 50688
rect 8814 50632 9076 50688
rect 8753 50630 9076 50632
rect 8753 50627 8819 50630
rect 9070 50628 9076 50630
rect 9140 50628 9146 50692
rect 9438 50628 9444 50692
rect 9508 50690 9514 50692
rect 11654 50690 11714 50764
rect 9508 50630 11714 50690
rect 13126 50690 13186 51038
rect 13353 51035 13419 51038
rect 14774 51036 14780 51100
rect 14844 51098 14850 51100
rect 15142 51098 15148 51100
rect 14844 51038 15148 51098
rect 14844 51036 14850 51038
rect 15142 51036 15148 51038
rect 15212 51036 15218 51100
rect 16070 50965 16130 51171
rect 17610 51168 17930 51169
rect 17610 51104 17618 51168
rect 17682 51104 17698 51168
rect 17762 51104 17778 51168
rect 17842 51104 17858 51168
rect 17922 51104 17930 51168
rect 17610 51103 17930 51104
rect 13445 50964 13511 50965
rect 13721 50964 13787 50965
rect 14825 50964 14891 50965
rect 13445 50962 13492 50964
rect 13400 50960 13492 50962
rect 13400 50904 13450 50960
rect 13400 50902 13492 50904
rect 13445 50900 13492 50902
rect 13556 50900 13562 50964
rect 13670 50900 13676 50964
rect 13740 50962 13787 50964
rect 14774 50962 14780 50964
rect 13740 50960 13832 50962
rect 13782 50904 13832 50960
rect 13740 50902 13832 50904
rect 14734 50902 14780 50962
rect 14844 50960 14891 50964
rect 14886 50904 14891 50960
rect 13740 50900 13787 50902
rect 14774 50900 14780 50902
rect 14844 50900 14891 50904
rect 13445 50899 13511 50900
rect 13721 50899 13787 50900
rect 14825 50899 14891 50900
rect 15285 50962 15351 50965
rect 16070 50962 16179 50965
rect 15285 50960 16179 50962
rect 15285 50904 15290 50960
rect 15346 50904 16118 50960
rect 16174 50904 16179 50960
rect 15285 50902 16179 50904
rect 15285 50899 15351 50902
rect 16113 50899 16179 50902
rect 13353 50826 13419 50829
rect 19520 50826 20000 50856
rect 13353 50824 20000 50826
rect 13353 50768 13358 50824
rect 13414 50768 20000 50824
rect 13353 50766 20000 50768
rect 13353 50763 13419 50766
rect 19520 50736 20000 50766
rect 13486 50690 13492 50692
rect 13126 50630 13492 50690
rect 9508 50628 9514 50630
rect 13486 50628 13492 50630
rect 13556 50628 13562 50692
rect 7610 50624 7930 50625
rect 7610 50560 7618 50624
rect 7682 50560 7698 50624
rect 7762 50560 7778 50624
rect 7842 50560 7858 50624
rect 7922 50560 7930 50624
rect 7610 50559 7930 50560
rect 14277 50624 14597 50625
rect 14277 50560 14285 50624
rect 14349 50560 14365 50624
rect 14429 50560 14445 50624
rect 14509 50560 14525 50624
rect 14589 50560 14597 50624
rect 14277 50559 14597 50560
rect 6748 50494 6930 50554
rect 6748 50492 6754 50494
rect 11462 50492 11468 50556
rect 11532 50554 11538 50556
rect 11697 50554 11763 50557
rect 11532 50552 11763 50554
rect 11532 50496 11702 50552
rect 11758 50496 11763 50552
rect 11532 50494 11763 50496
rect 11532 50492 11538 50494
rect 11697 50491 11763 50494
rect 6126 50356 6132 50420
rect 6196 50418 6202 50420
rect 8017 50418 8083 50421
rect 6196 50416 8083 50418
rect 6196 50360 8022 50416
rect 8078 50360 8083 50416
rect 6196 50358 8083 50360
rect 6196 50356 6202 50358
rect 8017 50355 8083 50358
rect 10961 50418 11027 50421
rect 10961 50416 11530 50418
rect 10961 50360 10966 50416
rect 11022 50360 11530 50416
rect 10961 50358 11530 50360
rect 10961 50355 11027 50358
rect 4061 50282 4127 50285
rect 6085 50282 6151 50285
rect 4061 50280 6151 50282
rect 4061 50224 4066 50280
rect 4122 50224 6090 50280
rect 6146 50224 6151 50280
rect 4061 50222 6151 50224
rect 11470 50282 11530 50358
rect 11881 50416 11947 50421
rect 11881 50360 11886 50416
rect 11942 50360 11947 50416
rect 11881 50355 11947 50360
rect 11605 50282 11671 50285
rect 11470 50280 11671 50282
rect 11470 50224 11610 50280
rect 11666 50224 11671 50280
rect 11470 50222 11671 50224
rect 4061 50219 4127 50222
rect 6085 50219 6151 50222
rect 11605 50219 11671 50222
rect 6126 50084 6132 50148
rect 6196 50146 6202 50148
rect 6453 50146 6519 50149
rect 6196 50144 6519 50146
rect 6196 50088 6458 50144
rect 6514 50088 6519 50144
rect 6196 50086 6519 50088
rect 6196 50084 6202 50086
rect 6453 50083 6519 50086
rect 7465 50146 7531 50149
rect 8334 50146 8340 50148
rect 7465 50144 8340 50146
rect 7465 50088 7470 50144
rect 7526 50088 8340 50144
rect 7465 50086 8340 50088
rect 7465 50083 7531 50086
rect 8334 50084 8340 50086
rect 8404 50084 8410 50148
rect 11884 50146 11944 50355
rect 13169 50282 13235 50285
rect 13302 50282 13308 50284
rect 13169 50280 13308 50282
rect 13169 50224 13174 50280
rect 13230 50224 13308 50280
rect 13169 50222 13308 50224
rect 13169 50219 13235 50222
rect 13302 50220 13308 50222
rect 13372 50220 13378 50284
rect 13997 50282 14063 50285
rect 15101 50282 15167 50285
rect 13997 50280 15167 50282
rect 13997 50224 14002 50280
rect 14058 50224 15106 50280
rect 15162 50224 15167 50280
rect 13997 50222 15167 50224
rect 13997 50219 14063 50222
rect 15101 50219 15167 50222
rect 12249 50146 12315 50149
rect 11884 50144 12315 50146
rect 11884 50088 12254 50144
rect 12310 50088 12315 50144
rect 11884 50086 12315 50088
rect 12249 50083 12315 50086
rect 13302 50084 13308 50148
rect 13372 50146 13378 50148
rect 13537 50146 13603 50149
rect 13372 50144 13603 50146
rect 13372 50088 13542 50144
rect 13598 50088 13603 50144
rect 13372 50086 13603 50088
rect 13372 50084 13378 50086
rect 13537 50083 13603 50086
rect 18137 50146 18203 50149
rect 19520 50146 20000 50176
rect 18137 50144 20000 50146
rect 18137 50088 18142 50144
rect 18198 50088 20000 50144
rect 18137 50086 20000 50088
rect 18137 50083 18203 50086
rect 4277 50080 4597 50081
rect 4277 50016 4285 50080
rect 4349 50016 4365 50080
rect 4429 50016 4445 50080
rect 4509 50016 4525 50080
rect 4589 50016 4597 50080
rect 4277 50015 4597 50016
rect 10944 50080 11264 50081
rect 10944 50016 10952 50080
rect 11016 50016 11032 50080
rect 11096 50016 11112 50080
rect 11176 50016 11192 50080
rect 11256 50016 11264 50080
rect 10944 50015 11264 50016
rect 17610 50080 17930 50081
rect 17610 50016 17618 50080
rect 17682 50016 17698 50080
rect 17762 50016 17778 50080
rect 17842 50016 17858 50080
rect 17922 50016 17930 50080
rect 19520 50056 20000 50086
rect 17610 50015 17930 50016
rect 2262 49948 2268 50012
rect 2332 50010 2338 50012
rect 2497 50010 2563 50013
rect 2332 50008 2563 50010
rect 2332 49952 2502 50008
rect 2558 49952 2563 50008
rect 2332 49950 2563 49952
rect 2332 49948 2338 49950
rect 2497 49947 2563 49950
rect 8569 50010 8635 50013
rect 9673 50012 9739 50013
rect 8569 50008 9506 50010
rect 8569 49952 8574 50008
rect 8630 49952 9506 50008
rect 8569 49950 9506 49952
rect 8569 49947 8635 49950
rect 0 49874 480 49904
rect 3049 49874 3115 49877
rect 0 49872 3115 49874
rect 0 49816 3054 49872
rect 3110 49816 3115 49872
rect 0 49814 3115 49816
rect 0 49784 480 49814
rect 3049 49811 3115 49814
rect 6862 49812 6868 49876
rect 6932 49874 6938 49876
rect 7833 49874 7899 49877
rect 6932 49872 7899 49874
rect 6932 49816 7838 49872
rect 7894 49816 7899 49872
rect 6932 49814 7899 49816
rect 6932 49812 6938 49814
rect 7833 49811 7899 49814
rect 9213 49876 9279 49877
rect 9213 49872 9260 49876
rect 9324 49874 9330 49876
rect 9213 49816 9218 49872
rect 9213 49812 9260 49816
rect 9324 49814 9370 49874
rect 9324 49812 9330 49814
rect 9213 49811 9279 49812
rect 2221 49738 2287 49741
rect 2865 49738 2931 49741
rect 2221 49736 2931 49738
rect 2221 49680 2226 49736
rect 2282 49680 2870 49736
rect 2926 49680 2931 49736
rect 2221 49678 2931 49680
rect 2221 49675 2287 49678
rect 2865 49675 2931 49678
rect 6269 49602 6335 49605
rect 6862 49602 6868 49604
rect 6269 49600 6868 49602
rect 6269 49544 6274 49600
rect 6330 49544 6868 49600
rect 6269 49542 6868 49544
rect 6269 49539 6335 49542
rect 6862 49540 6868 49542
rect 6932 49540 6938 49604
rect 7610 49536 7930 49537
rect 7610 49472 7618 49536
rect 7682 49472 7698 49536
rect 7762 49472 7778 49536
rect 7842 49472 7858 49536
rect 7922 49472 7930 49536
rect 7610 49471 7930 49472
rect 9254 49404 9260 49468
rect 9324 49466 9330 49468
rect 9446 49466 9506 49950
rect 9622 49948 9628 50012
rect 9692 50010 9739 50012
rect 14089 50010 14155 50013
rect 9692 50008 9784 50010
rect 9734 49952 9784 50008
rect 9692 49950 9784 49952
rect 13356 50008 14155 50010
rect 13356 49952 14094 50008
rect 14150 49952 14155 50008
rect 13356 49950 14155 49952
rect 9692 49948 9739 49950
rect 9673 49947 9739 49948
rect 13356 49877 13416 49950
rect 14089 49947 14155 49950
rect 9622 49812 9628 49876
rect 9692 49874 9698 49876
rect 10133 49874 10199 49877
rect 9692 49872 10199 49874
rect 9692 49816 10138 49872
rect 10194 49816 10199 49872
rect 9692 49814 10199 49816
rect 9692 49812 9698 49814
rect 10133 49811 10199 49814
rect 10542 49812 10548 49876
rect 10612 49874 10618 49876
rect 10961 49874 11027 49877
rect 10612 49872 11027 49874
rect 10612 49816 10966 49872
rect 11022 49816 11027 49872
rect 10612 49814 11027 49816
rect 10612 49812 10618 49814
rect 10961 49811 11027 49814
rect 13353 49872 13419 49877
rect 13353 49816 13358 49872
rect 13414 49816 13419 49872
rect 13353 49811 13419 49816
rect 16021 49874 16087 49877
rect 16297 49874 16363 49877
rect 16021 49872 16363 49874
rect 16021 49816 16026 49872
rect 16082 49816 16302 49872
rect 16358 49816 16363 49872
rect 16021 49814 16363 49816
rect 16021 49811 16087 49814
rect 16297 49811 16363 49814
rect 10225 49736 10291 49741
rect 10501 49740 10567 49741
rect 10501 49738 10548 49740
rect 10225 49680 10230 49736
rect 10286 49680 10291 49736
rect 10225 49675 10291 49680
rect 10456 49736 10548 49738
rect 10456 49680 10506 49736
rect 10456 49678 10548 49680
rect 10501 49676 10548 49678
rect 10612 49676 10618 49740
rect 15009 49738 15075 49741
rect 16665 49738 16731 49741
rect 15009 49736 16731 49738
rect 15009 49680 15014 49736
rect 15070 49680 16670 49736
rect 16726 49680 16731 49736
rect 15009 49678 16731 49680
rect 10501 49675 10567 49676
rect 15009 49675 15075 49678
rect 16665 49675 16731 49678
rect 10228 49602 10288 49675
rect 12893 49602 12959 49605
rect 10228 49600 12959 49602
rect 10228 49544 12898 49600
rect 12954 49544 12959 49600
rect 10228 49542 12959 49544
rect 12893 49539 12959 49542
rect 14277 49536 14597 49537
rect 14277 49472 14285 49536
rect 14349 49472 14365 49536
rect 14429 49472 14445 49536
rect 14509 49472 14525 49536
rect 14589 49472 14597 49536
rect 14277 49471 14597 49472
rect 9324 49406 9506 49466
rect 15653 49466 15719 49469
rect 19520 49466 20000 49496
rect 15653 49464 20000 49466
rect 15653 49408 15658 49464
rect 15714 49408 20000 49464
rect 15653 49406 20000 49408
rect 9324 49404 9330 49406
rect 15653 49403 15719 49406
rect 19520 49376 20000 49406
rect 6085 49330 6151 49333
rect 10593 49330 10659 49333
rect 6085 49328 10659 49330
rect 6085 49272 6090 49328
rect 6146 49272 10598 49328
rect 10654 49272 10659 49328
rect 6085 49270 10659 49272
rect 6085 49267 6151 49270
rect 10593 49267 10659 49270
rect 12566 49268 12572 49332
rect 12636 49330 12642 49332
rect 15653 49330 15719 49333
rect 12636 49328 15719 49330
rect 12636 49272 15658 49328
rect 15714 49272 15719 49328
rect 12636 49270 15719 49272
rect 12636 49268 12642 49270
rect 15653 49267 15719 49270
rect 3233 49194 3299 49197
rect 5390 49194 5396 49196
rect 3233 49192 5396 49194
rect 3233 49136 3238 49192
rect 3294 49136 5396 49192
rect 3233 49134 5396 49136
rect 3233 49131 3299 49134
rect 5390 49132 5396 49134
rect 5460 49132 5466 49196
rect 5533 49194 5599 49197
rect 8293 49194 8359 49197
rect 8886 49194 8892 49196
rect 5533 49192 8892 49194
rect 5533 49136 5538 49192
rect 5594 49136 8298 49192
rect 8354 49136 8892 49192
rect 5533 49134 8892 49136
rect 5533 49131 5599 49134
rect 8293 49131 8359 49134
rect 8886 49132 8892 49134
rect 8956 49132 8962 49196
rect 9949 49194 10015 49197
rect 13118 49194 13124 49196
rect 9949 49192 13124 49194
rect 9949 49136 9954 49192
rect 10010 49136 13124 49192
rect 9949 49134 13124 49136
rect 9949 49131 10015 49134
rect 13118 49132 13124 49134
rect 13188 49132 13194 49196
rect 13486 49132 13492 49196
rect 13556 49194 13562 49196
rect 13721 49194 13787 49197
rect 13556 49192 13787 49194
rect 13556 49136 13726 49192
rect 13782 49136 13787 49192
rect 13556 49134 13787 49136
rect 13556 49132 13562 49134
rect 13721 49131 13787 49134
rect 14825 49194 14891 49197
rect 16665 49194 16731 49197
rect 14825 49192 16731 49194
rect 14825 49136 14830 49192
rect 14886 49136 16670 49192
rect 16726 49136 16731 49192
rect 14825 49134 16731 49136
rect 14825 49131 14891 49134
rect 16665 49131 16731 49134
rect 0 49058 480 49088
rect 1945 49058 2011 49061
rect 0 49056 2011 49058
rect 0 49000 1950 49056
rect 2006 49000 2011 49056
rect 0 48998 2011 49000
rect 0 48968 480 48998
rect 1945 48995 2011 48998
rect 5349 49058 5415 49061
rect 5533 49058 5599 49061
rect 5349 49056 5599 49058
rect 5349 49000 5354 49056
rect 5410 49000 5538 49056
rect 5594 49000 5599 49056
rect 5349 48998 5599 49000
rect 5349 48995 5415 48998
rect 5533 48995 5599 48998
rect 4277 48992 4597 48993
rect 4277 48928 4285 48992
rect 4349 48928 4365 48992
rect 4429 48928 4445 48992
rect 4509 48928 4525 48992
rect 4589 48928 4597 48992
rect 4277 48927 4597 48928
rect 10944 48992 11264 48993
rect 10944 48928 10952 48992
rect 11016 48928 11032 48992
rect 11096 48928 11112 48992
rect 11176 48928 11192 48992
rect 11256 48928 11264 48992
rect 10944 48927 11264 48928
rect 17610 48992 17930 48993
rect 17610 48928 17618 48992
rect 17682 48928 17698 48992
rect 17762 48928 17778 48992
rect 17842 48928 17858 48992
rect 17922 48928 17930 48992
rect 17610 48927 17930 48928
rect 5390 48860 5396 48924
rect 5460 48922 5466 48924
rect 5625 48922 5691 48925
rect 14181 48922 14247 48925
rect 5460 48920 5691 48922
rect 5460 48864 5630 48920
rect 5686 48864 5691 48920
rect 5460 48862 5691 48864
rect 5460 48860 5466 48862
rect 5625 48859 5691 48862
rect 12022 48920 14247 48922
rect 12022 48864 14186 48920
rect 14242 48864 14247 48920
rect 12022 48862 14247 48864
rect 10961 48786 11027 48789
rect 11881 48786 11947 48789
rect 10961 48784 11947 48786
rect 10961 48728 10966 48784
rect 11022 48728 11886 48784
rect 11942 48728 11947 48784
rect 10961 48726 11947 48728
rect 10961 48723 11027 48726
rect 11881 48723 11947 48726
rect 2129 48650 2195 48653
rect 5993 48650 6059 48653
rect 7741 48650 7807 48653
rect 2129 48648 6059 48650
rect 2129 48592 2134 48648
rect 2190 48592 5998 48648
rect 6054 48592 6059 48648
rect 2129 48590 6059 48592
rect 2129 48587 2195 48590
rect 5993 48587 6059 48590
rect 7376 48648 7807 48650
rect 7376 48592 7746 48648
rect 7802 48592 7807 48648
rect 7376 48590 7807 48592
rect 7376 48381 7436 48590
rect 7741 48587 7807 48590
rect 9581 48650 9647 48653
rect 11237 48650 11303 48653
rect 12022 48650 12082 48862
rect 14181 48859 14247 48862
rect 12617 48786 12683 48789
rect 12750 48786 12756 48788
rect 12617 48784 12756 48786
rect 12617 48728 12622 48784
rect 12678 48728 12756 48784
rect 12617 48726 12756 48728
rect 12617 48723 12683 48726
rect 12750 48724 12756 48726
rect 12820 48724 12826 48788
rect 13537 48786 13603 48789
rect 19520 48786 20000 48816
rect 13537 48784 20000 48786
rect 13537 48728 13542 48784
rect 13598 48728 20000 48784
rect 13537 48726 20000 48728
rect 13537 48723 13603 48726
rect 19520 48696 20000 48726
rect 9581 48648 12082 48650
rect 9581 48592 9586 48648
rect 9642 48592 11242 48648
rect 11298 48592 12082 48648
rect 9581 48590 12082 48592
rect 9581 48587 9647 48590
rect 11237 48587 11303 48590
rect 8109 48514 8175 48517
rect 12617 48514 12683 48517
rect 8109 48512 12683 48514
rect 8109 48456 8114 48512
rect 8170 48456 12622 48512
rect 12678 48456 12683 48512
rect 8109 48454 12683 48456
rect 8109 48451 8175 48454
rect 12617 48451 12683 48454
rect 7610 48448 7930 48449
rect 7610 48384 7618 48448
rect 7682 48384 7698 48448
rect 7762 48384 7778 48448
rect 7842 48384 7858 48448
rect 7922 48384 7930 48448
rect 7610 48383 7930 48384
rect 14277 48448 14597 48449
rect 14277 48384 14285 48448
rect 14349 48384 14365 48448
rect 14429 48384 14445 48448
rect 14509 48384 14525 48448
rect 14589 48384 14597 48448
rect 14277 48383 14597 48384
rect 5758 48316 5764 48380
rect 5828 48378 5834 48380
rect 6085 48378 6151 48381
rect 5828 48376 6151 48378
rect 5828 48320 6090 48376
rect 6146 48320 6151 48376
rect 5828 48318 6151 48320
rect 5828 48316 5834 48318
rect 6085 48315 6151 48318
rect 7373 48376 7439 48381
rect 7373 48320 7378 48376
rect 7434 48320 7439 48376
rect 7373 48315 7439 48320
rect 8702 48316 8708 48380
rect 8772 48316 8778 48380
rect 11421 48378 11487 48381
rect 12934 48378 12940 48380
rect 11421 48376 12940 48378
rect 11421 48320 11426 48376
rect 11482 48320 12940 48376
rect 11421 48318 12940 48320
rect 0 48242 480 48272
rect 2773 48242 2839 48245
rect 0 48240 2839 48242
rect 0 48184 2778 48240
rect 2834 48184 2839 48240
rect 0 48182 2839 48184
rect 0 48152 480 48182
rect 2773 48179 2839 48182
rect 3417 48242 3483 48245
rect 3734 48242 3740 48244
rect 3417 48240 3740 48242
rect 3417 48184 3422 48240
rect 3478 48184 3740 48240
rect 3417 48182 3740 48184
rect 3417 48179 3483 48182
rect 3734 48180 3740 48182
rect 3804 48180 3810 48244
rect 5809 48242 5875 48245
rect 7925 48242 7991 48245
rect 8710 48242 8770 48316
rect 11421 48315 11487 48318
rect 12934 48316 12940 48318
rect 13004 48316 13010 48380
rect 5809 48240 8770 48242
rect 5809 48184 5814 48240
rect 5870 48184 7930 48240
rect 7986 48184 8770 48240
rect 5809 48182 8770 48184
rect 5809 48179 5875 48182
rect 7925 48179 7991 48182
rect 8109 48106 8175 48109
rect 12065 48106 12131 48109
rect 8109 48104 12131 48106
rect 8109 48048 8114 48104
rect 8170 48048 12070 48104
rect 12126 48048 12131 48104
rect 8109 48046 12131 48048
rect 8109 48043 8175 48046
rect 12065 48043 12131 48046
rect 13261 48106 13327 48109
rect 19520 48106 20000 48136
rect 13261 48104 20000 48106
rect 13261 48048 13266 48104
rect 13322 48048 20000 48104
rect 13261 48046 20000 48048
rect 13261 48043 13327 48046
rect 19520 48016 20000 48046
rect 6085 47970 6151 47973
rect 8109 47970 8175 47973
rect 6085 47968 8175 47970
rect 6085 47912 6090 47968
rect 6146 47912 8114 47968
rect 8170 47912 8175 47968
rect 6085 47910 8175 47912
rect 6085 47907 6151 47910
rect 8109 47907 8175 47910
rect 4277 47904 4597 47905
rect 4277 47840 4285 47904
rect 4349 47840 4365 47904
rect 4429 47840 4445 47904
rect 4509 47840 4525 47904
rect 4589 47840 4597 47904
rect 4277 47839 4597 47840
rect 10944 47904 11264 47905
rect 10944 47840 10952 47904
rect 11016 47840 11032 47904
rect 11096 47840 11112 47904
rect 11176 47840 11192 47904
rect 11256 47840 11264 47904
rect 10944 47839 11264 47840
rect 17610 47904 17930 47905
rect 17610 47840 17618 47904
rect 17682 47840 17698 47904
rect 17762 47840 17778 47904
rect 17842 47840 17858 47904
rect 17922 47840 17930 47904
rect 17610 47839 17930 47840
rect 6678 47772 6684 47836
rect 6748 47834 6754 47836
rect 6913 47834 6979 47837
rect 12709 47834 12775 47837
rect 6748 47832 6979 47834
rect 6748 47776 6918 47832
rect 6974 47776 6979 47832
rect 6748 47774 6979 47776
rect 6748 47772 6754 47774
rect 6913 47771 6979 47774
rect 11470 47832 12775 47834
rect 11470 47776 12714 47832
rect 12770 47776 12775 47832
rect 11470 47774 12775 47776
rect 5809 47698 5875 47701
rect 6310 47698 6316 47700
rect 5809 47696 6316 47698
rect 5809 47640 5814 47696
rect 5870 47640 6316 47696
rect 5809 47638 6316 47640
rect 5809 47635 5875 47638
rect 6310 47636 6316 47638
rect 6380 47698 6386 47700
rect 6637 47698 6703 47701
rect 6380 47696 6703 47698
rect 6380 47640 6642 47696
rect 6698 47640 6703 47696
rect 6380 47638 6703 47640
rect 6380 47636 6386 47638
rect 6637 47635 6703 47638
rect 10961 47698 11027 47701
rect 11470 47698 11530 47774
rect 12709 47771 12775 47774
rect 10961 47696 11530 47698
rect 10961 47640 10966 47696
rect 11022 47640 11530 47696
rect 10961 47638 11530 47640
rect 11605 47698 11671 47701
rect 12382 47698 12388 47700
rect 11605 47696 12388 47698
rect 11605 47640 11610 47696
rect 11666 47640 12388 47696
rect 11605 47638 12388 47640
rect 10961 47635 11027 47638
rect 11605 47635 11671 47638
rect 12382 47636 12388 47638
rect 12452 47636 12458 47700
rect 3918 47500 3924 47564
rect 3988 47562 3994 47564
rect 4153 47562 4219 47565
rect 3988 47560 4219 47562
rect 3988 47504 4158 47560
rect 4214 47504 4219 47560
rect 3988 47502 4219 47504
rect 3988 47500 3994 47502
rect 4153 47499 4219 47502
rect 12801 47562 12867 47565
rect 12801 47560 14842 47562
rect 12801 47504 12806 47560
rect 12862 47504 14842 47560
rect 12801 47502 14842 47504
rect 12801 47499 12867 47502
rect 0 47426 480 47456
rect 1301 47426 1367 47429
rect 0 47424 1367 47426
rect 0 47368 1306 47424
rect 1362 47368 1367 47424
rect 0 47366 1367 47368
rect 0 47336 480 47366
rect 1301 47363 1367 47366
rect 12341 47426 12407 47429
rect 12750 47426 12756 47428
rect 12341 47424 12756 47426
rect 12341 47368 12346 47424
rect 12402 47368 12756 47424
rect 12341 47366 12756 47368
rect 12341 47363 12407 47366
rect 12750 47364 12756 47366
rect 12820 47364 12826 47428
rect 14782 47426 14842 47502
rect 19520 47426 20000 47456
rect 14782 47366 20000 47426
rect 7610 47360 7930 47361
rect 7610 47296 7618 47360
rect 7682 47296 7698 47360
rect 7762 47296 7778 47360
rect 7842 47296 7858 47360
rect 7922 47296 7930 47360
rect 7610 47295 7930 47296
rect 14277 47360 14597 47361
rect 14277 47296 14285 47360
rect 14349 47296 14365 47360
rect 14429 47296 14445 47360
rect 14509 47296 14525 47360
rect 14589 47296 14597 47360
rect 19520 47336 20000 47366
rect 14277 47295 14597 47296
rect 2865 47290 2931 47293
rect 4705 47290 4771 47293
rect 2865 47288 4771 47290
rect 2865 47232 2870 47288
rect 2926 47232 4710 47288
rect 4766 47232 4771 47288
rect 2865 47230 4771 47232
rect 2865 47227 2931 47230
rect 4705 47227 4771 47230
rect 12341 47290 12407 47293
rect 12566 47290 12572 47292
rect 12341 47288 12572 47290
rect 12341 47232 12346 47288
rect 12402 47232 12572 47288
rect 12341 47230 12572 47232
rect 12341 47227 12407 47230
rect 12566 47228 12572 47230
rect 12636 47290 12642 47292
rect 14089 47290 14155 47293
rect 12636 47288 14155 47290
rect 12636 47232 14094 47288
rect 14150 47232 14155 47288
rect 12636 47230 14155 47232
rect 12636 47228 12642 47230
rect 14089 47227 14155 47230
rect 4981 47154 5047 47157
rect 11697 47154 11763 47157
rect 13629 47154 13695 47157
rect 15561 47154 15627 47157
rect 4981 47152 5090 47154
rect 4981 47096 4986 47152
rect 5042 47096 5090 47152
rect 4981 47091 5090 47096
rect 11697 47152 15627 47154
rect 11697 47096 11702 47152
rect 11758 47096 13634 47152
rect 13690 47096 15566 47152
rect 15622 47096 15627 47152
rect 11697 47094 15627 47096
rect 11697 47091 11763 47094
rect 13629 47091 13695 47094
rect 15561 47091 15627 47094
rect 16389 47154 16455 47157
rect 17033 47154 17099 47157
rect 16389 47152 17099 47154
rect 16389 47096 16394 47152
rect 16450 47096 17038 47152
rect 17094 47096 17099 47152
rect 16389 47094 17099 47096
rect 16389 47091 16455 47094
rect 17033 47091 17099 47094
rect 1577 47016 1643 47021
rect 1577 46960 1582 47016
rect 1638 46960 1643 47016
rect 1577 46955 1643 46960
rect 0 46746 480 46776
rect 1580 46746 1640 46955
rect 5030 46885 5090 47091
rect 6494 46956 6500 47020
rect 6564 47018 6570 47020
rect 11605 47018 11671 47021
rect 6564 47016 11671 47018
rect 6564 46960 11610 47016
rect 11666 46960 11671 47016
rect 6564 46958 11671 46960
rect 6564 46956 6570 46958
rect 11605 46955 11671 46958
rect 16297 47018 16363 47021
rect 16941 47018 17007 47021
rect 16297 47016 17007 47018
rect 16297 46960 16302 47016
rect 16358 46960 16946 47016
rect 17002 46960 17007 47016
rect 16297 46958 17007 46960
rect 16297 46955 16363 46958
rect 16941 46955 17007 46958
rect 5030 46880 5139 46885
rect 8385 46884 8451 46885
rect 5030 46824 5078 46880
rect 5134 46824 5139 46880
rect 5030 46822 5139 46824
rect 5073 46819 5139 46822
rect 8334 46820 8340 46884
rect 8404 46882 8451 46884
rect 13169 46882 13235 46885
rect 13537 46882 13603 46885
rect 8404 46880 8496 46882
rect 8446 46824 8496 46880
rect 8404 46822 8496 46824
rect 13169 46880 13603 46882
rect 13169 46824 13174 46880
rect 13230 46824 13542 46880
rect 13598 46824 13603 46880
rect 13169 46822 13603 46824
rect 8404 46820 8451 46822
rect 8385 46819 8451 46820
rect 13169 46819 13235 46822
rect 13537 46819 13603 46822
rect 4277 46816 4597 46817
rect 4277 46752 4285 46816
rect 4349 46752 4365 46816
rect 4429 46752 4445 46816
rect 4509 46752 4525 46816
rect 4589 46752 4597 46816
rect 4277 46751 4597 46752
rect 10944 46816 11264 46817
rect 10944 46752 10952 46816
rect 11016 46752 11032 46816
rect 11096 46752 11112 46816
rect 11176 46752 11192 46816
rect 11256 46752 11264 46816
rect 10944 46751 11264 46752
rect 17610 46816 17930 46817
rect 17610 46752 17618 46816
rect 17682 46752 17698 46816
rect 17762 46752 17778 46816
rect 17842 46752 17858 46816
rect 17922 46752 17930 46816
rect 17610 46751 17930 46752
rect 3233 46748 3299 46749
rect 0 46686 1640 46746
rect 0 46656 480 46686
rect 3182 46684 3188 46748
rect 3252 46746 3299 46748
rect 15326 46746 15332 46748
rect 3252 46744 3344 46746
rect 3294 46688 3344 46744
rect 3252 46686 3344 46688
rect 12436 46686 15332 46746
rect 3252 46684 3299 46686
rect 3233 46683 3299 46684
rect 4521 46610 4587 46613
rect 12436 46610 12496 46686
rect 15326 46684 15332 46686
rect 15396 46684 15402 46748
rect 19520 46746 20000 46776
rect 18094 46686 20000 46746
rect 4521 46608 12496 46610
rect 4521 46552 4526 46608
rect 4582 46552 12496 46608
rect 4521 46550 12496 46552
rect 13261 46610 13327 46613
rect 18094 46610 18154 46686
rect 19520 46656 20000 46686
rect 13261 46608 18154 46610
rect 13261 46552 13266 46608
rect 13322 46552 18154 46608
rect 13261 46550 18154 46552
rect 4521 46547 4587 46550
rect 13261 46547 13327 46550
rect 5625 46474 5691 46477
rect 7046 46474 7052 46476
rect 5625 46472 7052 46474
rect 5625 46416 5630 46472
rect 5686 46416 7052 46472
rect 5625 46414 7052 46416
rect 5625 46411 5691 46414
rect 7046 46412 7052 46414
rect 7116 46412 7122 46476
rect 13537 46474 13603 46477
rect 13537 46472 14842 46474
rect 13537 46416 13542 46472
rect 13598 46416 14842 46472
rect 13537 46414 14842 46416
rect 13537 46411 13603 46414
rect 13302 46338 13308 46340
rect 8572 46278 13308 46338
rect 7610 46272 7930 46273
rect 7610 46208 7618 46272
rect 7682 46208 7698 46272
rect 7762 46208 7778 46272
rect 7842 46208 7858 46272
rect 7922 46208 7930 46272
rect 7610 46207 7930 46208
rect 8572 46205 8632 46278
rect 13302 46276 13308 46278
rect 13372 46276 13378 46340
rect 14277 46272 14597 46273
rect 14277 46208 14285 46272
rect 14349 46208 14365 46272
rect 14429 46208 14445 46272
rect 14509 46208 14525 46272
rect 14589 46208 14597 46272
rect 14277 46207 14597 46208
rect 8569 46200 8635 46205
rect 8569 46144 8574 46200
rect 8630 46144 8635 46200
rect 8569 46139 8635 46144
rect 12198 46140 12204 46204
rect 12268 46202 12274 46204
rect 12566 46202 12572 46204
rect 12268 46142 12572 46202
rect 12268 46140 12274 46142
rect 12566 46140 12572 46142
rect 12636 46140 12642 46204
rect 3601 46066 3667 46069
rect 5022 46066 5028 46068
rect 3601 46064 5028 46066
rect 3601 46008 3606 46064
rect 3662 46008 5028 46064
rect 3601 46006 5028 46008
rect 3601 46003 3667 46006
rect 5022 46004 5028 46006
rect 5092 46004 5098 46068
rect 10685 46066 10751 46069
rect 13261 46066 13327 46069
rect 10685 46064 13327 46066
rect 10685 46008 10690 46064
rect 10746 46008 13266 46064
rect 13322 46008 13327 46064
rect 10685 46006 13327 46008
rect 14782 46066 14842 46414
rect 16982 46412 16988 46476
rect 17052 46474 17058 46476
rect 17217 46474 17283 46477
rect 17052 46472 17283 46474
rect 17052 46416 17222 46472
rect 17278 46416 17283 46472
rect 17052 46414 17283 46416
rect 17052 46412 17058 46414
rect 17217 46411 17283 46414
rect 19520 46066 20000 46096
rect 14782 46006 20000 46066
rect 10685 46003 10751 46006
rect 13261 46003 13327 46006
rect 19520 45976 20000 46006
rect 0 45930 480 45960
rect 1761 45930 1827 45933
rect 0 45928 1827 45930
rect 0 45872 1766 45928
rect 1822 45872 1827 45928
rect 0 45870 1827 45872
rect 0 45840 480 45870
rect 1761 45867 1827 45870
rect 2262 45868 2268 45932
rect 2332 45930 2338 45932
rect 2497 45930 2563 45933
rect 2332 45928 2563 45930
rect 2332 45872 2502 45928
rect 2558 45872 2563 45928
rect 2332 45870 2563 45872
rect 2332 45868 2338 45870
rect 2497 45867 2563 45870
rect 3233 45930 3299 45933
rect 4838 45930 4844 45932
rect 3233 45928 4844 45930
rect 3233 45872 3238 45928
rect 3294 45872 4844 45928
rect 3233 45870 4844 45872
rect 3233 45867 3299 45870
rect 4838 45868 4844 45870
rect 4908 45868 4914 45932
rect 10358 45868 10364 45932
rect 10428 45930 10434 45932
rect 15101 45930 15167 45933
rect 10428 45928 15167 45930
rect 10428 45872 15106 45928
rect 15162 45872 15167 45928
rect 10428 45870 15167 45872
rect 10428 45868 10434 45870
rect 15101 45867 15167 45870
rect 8702 45732 8708 45796
rect 8772 45794 8778 45796
rect 9806 45794 9812 45796
rect 8772 45734 9812 45794
rect 8772 45732 8778 45734
rect 9806 45732 9812 45734
rect 9876 45732 9882 45796
rect 11646 45732 11652 45796
rect 11716 45794 11722 45796
rect 12382 45794 12388 45796
rect 11716 45734 12388 45794
rect 11716 45732 11722 45734
rect 12382 45732 12388 45734
rect 12452 45732 12458 45796
rect 4277 45728 4597 45729
rect 4277 45664 4285 45728
rect 4349 45664 4365 45728
rect 4429 45664 4445 45728
rect 4509 45664 4525 45728
rect 4589 45664 4597 45728
rect 4277 45663 4597 45664
rect 10944 45728 11264 45729
rect 10944 45664 10952 45728
rect 11016 45664 11032 45728
rect 11096 45664 11112 45728
rect 11176 45664 11192 45728
rect 11256 45664 11264 45728
rect 10944 45663 11264 45664
rect 17610 45728 17930 45729
rect 17610 45664 17618 45728
rect 17682 45664 17698 45728
rect 17762 45664 17778 45728
rect 17842 45664 17858 45728
rect 17922 45664 17930 45728
rect 17610 45663 17930 45664
rect 7046 45596 7052 45660
rect 7116 45658 7122 45660
rect 7925 45658 7991 45661
rect 8937 45660 9003 45661
rect 8886 45658 8892 45660
rect 7116 45656 7991 45658
rect 7116 45600 7930 45656
rect 7986 45600 7991 45656
rect 7116 45598 7991 45600
rect 8846 45598 8892 45658
rect 8956 45656 9003 45660
rect 8998 45600 9003 45656
rect 7116 45596 7122 45598
rect 7925 45595 7991 45598
rect 8886 45596 8892 45598
rect 8956 45596 9003 45600
rect 8937 45595 9003 45596
rect 14825 45658 14891 45661
rect 15326 45658 15332 45660
rect 14825 45656 15332 45658
rect 14825 45600 14830 45656
rect 14886 45600 15332 45656
rect 14825 45598 15332 45600
rect 14825 45595 14891 45598
rect 15326 45596 15332 45598
rect 15396 45596 15402 45660
rect 6177 45524 6243 45525
rect 9857 45524 9923 45525
rect 6126 45460 6132 45524
rect 6196 45522 6243 45524
rect 6196 45520 6288 45522
rect 6238 45464 6288 45520
rect 6196 45462 6288 45464
rect 6196 45460 6243 45462
rect 9806 45460 9812 45524
rect 9876 45522 9923 45524
rect 10869 45522 10935 45525
rect 11513 45522 11579 45525
rect 11789 45522 11855 45525
rect 9876 45520 9968 45522
rect 9918 45464 9968 45520
rect 9876 45462 9968 45464
rect 10869 45520 11579 45522
rect 10869 45464 10874 45520
rect 10930 45464 11518 45520
rect 11574 45464 11579 45520
rect 10869 45462 11579 45464
rect 9876 45460 9923 45462
rect 6177 45459 6243 45460
rect 9857 45459 9923 45460
rect 10869 45459 10935 45462
rect 11513 45459 11579 45462
rect 11654 45520 11855 45522
rect 11654 45464 11794 45520
rect 11850 45464 11855 45520
rect 11654 45462 11855 45464
rect 10225 45386 10291 45389
rect 11654 45386 11714 45462
rect 11789 45459 11855 45462
rect 10225 45384 11714 45386
rect 10225 45328 10230 45384
rect 10286 45328 11714 45384
rect 10225 45326 11714 45328
rect 13537 45386 13603 45389
rect 19520 45386 20000 45416
rect 13537 45384 20000 45386
rect 13537 45328 13542 45384
rect 13598 45328 20000 45384
rect 13537 45326 20000 45328
rect 10225 45323 10291 45326
rect 13537 45323 13603 45326
rect 19520 45296 20000 45326
rect 9949 45250 10015 45253
rect 12198 45250 12204 45252
rect 9949 45248 12204 45250
rect 9949 45192 9954 45248
rect 10010 45192 12204 45248
rect 9949 45190 12204 45192
rect 9949 45187 10015 45190
rect 12198 45188 12204 45190
rect 12268 45188 12274 45252
rect 7610 45184 7930 45185
rect 0 45114 480 45144
rect 7610 45120 7618 45184
rect 7682 45120 7698 45184
rect 7762 45120 7778 45184
rect 7842 45120 7858 45184
rect 7922 45120 7930 45184
rect 7610 45119 7930 45120
rect 14277 45184 14597 45185
rect 14277 45120 14285 45184
rect 14349 45120 14365 45184
rect 14429 45120 14445 45184
rect 14509 45120 14525 45184
rect 14589 45120 14597 45184
rect 14277 45119 14597 45120
rect 2405 45114 2471 45117
rect 0 45112 2471 45114
rect 0 45056 2410 45112
rect 2466 45056 2471 45112
rect 0 45054 2471 45056
rect 0 45024 480 45054
rect 2405 45051 2471 45054
rect 4245 45114 4311 45117
rect 4654 45114 4660 45116
rect 4245 45112 4660 45114
rect 4245 45056 4250 45112
rect 4306 45056 4660 45112
rect 4245 45054 4660 45056
rect 4245 45051 4311 45054
rect 4654 45052 4660 45054
rect 4724 45052 4730 45116
rect 7005 45112 7071 45117
rect 7005 45056 7010 45112
rect 7066 45056 7071 45112
rect 7005 45051 7071 45056
rect 15694 45052 15700 45116
rect 15764 45114 15770 45116
rect 15929 45114 15995 45117
rect 15764 45112 15995 45114
rect 15764 45056 15934 45112
rect 15990 45056 15995 45112
rect 15764 45054 15995 45056
rect 15764 45052 15770 45054
rect 15929 45051 15995 45054
rect 7008 44978 7068 45051
rect 7557 44978 7623 44981
rect 7008 44976 7623 44978
rect 7008 44920 7562 44976
rect 7618 44920 7623 44976
rect 7008 44918 7623 44920
rect 7557 44915 7623 44918
rect 12065 44706 12131 44709
rect 14549 44706 14615 44709
rect 19520 44706 20000 44736
rect 12065 44704 14615 44706
rect 12065 44648 12070 44704
rect 12126 44648 14554 44704
rect 14610 44648 14615 44704
rect 12065 44646 14615 44648
rect 12065 44643 12131 44646
rect 14549 44643 14615 44646
rect 18094 44646 20000 44706
rect 4277 44640 4597 44641
rect 4277 44576 4285 44640
rect 4349 44576 4365 44640
rect 4429 44576 4445 44640
rect 4509 44576 4525 44640
rect 4589 44576 4597 44640
rect 4277 44575 4597 44576
rect 10944 44640 11264 44641
rect 10944 44576 10952 44640
rect 11016 44576 11032 44640
rect 11096 44576 11112 44640
rect 11176 44576 11192 44640
rect 11256 44576 11264 44640
rect 10944 44575 11264 44576
rect 17610 44640 17930 44641
rect 17610 44576 17618 44640
rect 17682 44576 17698 44640
rect 17762 44576 17778 44640
rect 17842 44576 17858 44640
rect 17922 44576 17930 44640
rect 17610 44575 17930 44576
rect 3969 44436 4035 44437
rect 3918 44372 3924 44436
rect 3988 44434 4035 44436
rect 5625 44434 5691 44437
rect 9254 44434 9260 44436
rect 3988 44432 4080 44434
rect 4030 44376 4080 44432
rect 3988 44374 4080 44376
rect 5625 44432 9260 44434
rect 5625 44376 5630 44432
rect 5686 44376 9260 44432
rect 5625 44374 9260 44376
rect 3988 44372 4035 44374
rect 3969 44371 4035 44372
rect 5625 44371 5691 44374
rect 9254 44372 9260 44374
rect 9324 44372 9330 44436
rect 10869 44434 10935 44437
rect 12065 44434 12131 44437
rect 10869 44432 12131 44434
rect 10869 44376 10874 44432
rect 10930 44376 12070 44432
rect 12126 44376 12131 44432
rect 10869 44374 12131 44376
rect 10869 44371 10935 44374
rect 12065 44371 12131 44374
rect 13537 44434 13603 44437
rect 18094 44434 18154 44646
rect 19520 44616 20000 44646
rect 13537 44432 18154 44434
rect 13537 44376 13542 44432
rect 13598 44376 18154 44432
rect 13537 44374 18154 44376
rect 13537 44371 13603 44374
rect 0 44298 480 44328
rect 1485 44298 1551 44301
rect 0 44296 1551 44298
rect 0 44240 1490 44296
rect 1546 44240 1551 44296
rect 0 44238 1551 44240
rect 0 44208 480 44238
rect 1485 44235 1551 44238
rect 9070 44236 9076 44300
rect 9140 44298 9146 44300
rect 9140 44238 13876 44298
rect 9140 44236 9146 44238
rect 9029 44162 9095 44165
rect 9438 44162 9444 44164
rect 9029 44160 9444 44162
rect 9029 44104 9034 44160
rect 9090 44104 9444 44160
rect 9029 44102 9444 44104
rect 9029 44099 9095 44102
rect 9438 44100 9444 44102
rect 9508 44100 9514 44164
rect 7610 44096 7930 44097
rect 7610 44032 7618 44096
rect 7682 44032 7698 44096
rect 7762 44032 7778 44096
rect 7842 44032 7858 44096
rect 7922 44032 7930 44096
rect 7610 44031 7930 44032
rect 13816 44029 13876 44238
rect 14277 44096 14597 44097
rect 14277 44032 14285 44096
rect 14349 44032 14365 44096
rect 14429 44032 14445 44096
rect 14509 44032 14525 44096
rect 14589 44032 14597 44096
rect 14277 44031 14597 44032
rect 2497 44026 2563 44029
rect 6913 44026 6979 44029
rect 2497 44024 6979 44026
rect 2497 43968 2502 44024
rect 2558 43968 6918 44024
rect 6974 43968 6979 44024
rect 2497 43966 6979 43968
rect 2497 43963 2563 43966
rect 6913 43963 6979 43966
rect 13813 44024 13879 44029
rect 13813 43968 13818 44024
rect 13874 43968 13879 44024
rect 13813 43963 13879 43968
rect 15653 44026 15719 44029
rect 19520 44026 20000 44056
rect 15653 44024 20000 44026
rect 15653 43968 15658 44024
rect 15714 43968 20000 44024
rect 15653 43966 20000 43968
rect 15653 43963 15719 43966
rect 19520 43936 20000 43966
rect 5257 43890 5323 43893
rect 5390 43890 5396 43892
rect 5257 43888 5396 43890
rect 5257 43832 5262 43888
rect 5318 43832 5396 43888
rect 5257 43830 5396 43832
rect 5257 43827 5323 43830
rect 5390 43828 5396 43830
rect 5460 43828 5466 43892
rect 9990 43828 9996 43892
rect 10060 43890 10066 43892
rect 10317 43890 10383 43893
rect 10060 43888 10383 43890
rect 10060 43832 10322 43888
rect 10378 43832 10383 43888
rect 10060 43830 10383 43832
rect 10060 43828 10066 43830
rect 10317 43827 10383 43830
rect 15009 43890 15075 43893
rect 15510 43890 15516 43892
rect 15009 43888 15516 43890
rect 15009 43832 15014 43888
rect 15070 43832 15516 43888
rect 15009 43830 15516 43832
rect 15009 43827 15075 43830
rect 15510 43828 15516 43830
rect 15580 43828 15586 43892
rect 7005 43754 7071 43757
rect 9857 43754 9923 43757
rect 7005 43752 9923 43754
rect 7005 43696 7010 43752
rect 7066 43696 9862 43752
rect 9918 43696 9923 43752
rect 7005 43694 9923 43696
rect 7005 43691 7071 43694
rect 9857 43691 9923 43694
rect 13670 43692 13676 43756
rect 13740 43754 13746 43756
rect 16389 43754 16455 43757
rect 13740 43752 16455 43754
rect 13740 43696 16394 43752
rect 16450 43696 16455 43752
rect 13740 43694 16455 43696
rect 13740 43692 13746 43694
rect 16389 43691 16455 43694
rect 4277 43552 4597 43553
rect 0 43482 480 43512
rect 4277 43488 4285 43552
rect 4349 43488 4365 43552
rect 4429 43488 4445 43552
rect 4509 43488 4525 43552
rect 4589 43488 4597 43552
rect 4277 43487 4597 43488
rect 10944 43552 11264 43553
rect 10944 43488 10952 43552
rect 11016 43488 11032 43552
rect 11096 43488 11112 43552
rect 11176 43488 11192 43552
rect 11256 43488 11264 43552
rect 10944 43487 11264 43488
rect 17610 43552 17930 43553
rect 17610 43488 17618 43552
rect 17682 43488 17698 43552
rect 17762 43488 17778 43552
rect 17842 43488 17858 43552
rect 17922 43488 17930 43552
rect 17610 43487 17930 43488
rect 1577 43482 1643 43485
rect 0 43480 1643 43482
rect 0 43424 1582 43480
rect 1638 43424 1643 43480
rect 0 43422 1643 43424
rect 0 43392 480 43422
rect 1577 43419 1643 43422
rect 15837 43482 15903 43485
rect 16430 43482 16436 43484
rect 15837 43480 16436 43482
rect 15837 43424 15842 43480
rect 15898 43424 16436 43480
rect 15837 43422 16436 43424
rect 15837 43419 15903 43422
rect 16430 43420 16436 43422
rect 16500 43420 16506 43484
rect 3233 43346 3299 43349
rect 8518 43346 8524 43348
rect 3233 43344 8524 43346
rect 3233 43288 3238 43344
rect 3294 43288 8524 43344
rect 3233 43286 8524 43288
rect 3233 43283 3299 43286
rect 8518 43284 8524 43286
rect 8588 43284 8594 43348
rect 10174 43284 10180 43348
rect 10244 43284 10250 43348
rect 12525 43346 12591 43349
rect 13813 43346 13879 43349
rect 12525 43344 13879 43346
rect 12525 43288 12530 43344
rect 12586 43288 13818 43344
rect 13874 43288 13879 43344
rect 12525 43286 13879 43288
rect 3969 43074 4035 43077
rect 3742 43072 4035 43074
rect 3742 43016 3974 43072
rect 4030 43016 4035 43072
rect 3742 43014 4035 43016
rect 3742 42805 3802 43014
rect 3969 43011 4035 43014
rect 6177 43074 6243 43077
rect 6310 43074 6316 43076
rect 6177 43072 6316 43074
rect 6177 43016 6182 43072
rect 6238 43016 6316 43072
rect 6177 43014 6316 43016
rect 6177 43011 6243 43014
rect 6310 43012 6316 43014
rect 6380 43012 6386 43076
rect 7610 43008 7930 43009
rect 7610 42944 7618 43008
rect 7682 42944 7698 43008
rect 7762 42944 7778 43008
rect 7842 42944 7858 43008
rect 7922 42944 7930 43008
rect 7610 42943 7930 42944
rect 3969 42938 4035 42941
rect 6862 42938 6868 42940
rect 3969 42936 6868 42938
rect 3969 42880 3974 42936
rect 4030 42880 6868 42936
rect 3969 42878 6868 42880
rect 3969 42875 4035 42878
rect 6862 42876 6868 42878
rect 6932 42876 6938 42940
rect 9070 42876 9076 42940
rect 9140 42938 9146 42940
rect 9990 42938 9996 42940
rect 9140 42878 9996 42938
rect 9140 42876 9146 42878
rect 9990 42876 9996 42878
rect 10060 42876 10066 42940
rect 10182 42805 10242 43284
rect 12525 43283 12591 43286
rect 13813 43283 13879 43286
rect 15101 43346 15167 43349
rect 19520 43346 20000 43376
rect 15101 43344 20000 43346
rect 15101 43288 15106 43344
rect 15162 43288 20000 43344
rect 15101 43286 20000 43288
rect 15101 43283 15167 43286
rect 19520 43256 20000 43286
rect 15101 43210 15167 43213
rect 15326 43210 15332 43212
rect 15101 43208 15332 43210
rect 15101 43152 15106 43208
rect 15162 43152 15332 43208
rect 15101 43150 15332 43152
rect 15101 43147 15167 43150
rect 15326 43148 15332 43150
rect 15396 43148 15402 43212
rect 14277 43008 14597 43009
rect 14277 42944 14285 43008
rect 14349 42944 14365 43008
rect 14429 42944 14445 43008
rect 14509 42944 14525 43008
rect 14589 42944 14597 43008
rect 14277 42943 14597 42944
rect 10409 42940 10475 42941
rect 10358 42938 10364 42940
rect 10318 42878 10364 42938
rect 10428 42936 10475 42940
rect 10470 42880 10475 42936
rect 10358 42876 10364 42878
rect 10428 42876 10475 42880
rect 10409 42875 10475 42876
rect 2446 42740 2452 42804
rect 2516 42802 2522 42804
rect 2865 42802 2931 42805
rect 2516 42800 2931 42802
rect 2516 42744 2870 42800
rect 2926 42744 2931 42800
rect 2516 42742 2931 42744
rect 3742 42800 3851 42805
rect 6177 42804 6243 42805
rect 3742 42744 3790 42800
rect 3846 42744 3851 42800
rect 3742 42742 3851 42744
rect 2516 42740 2522 42742
rect 2865 42739 2931 42742
rect 3785 42739 3851 42742
rect 6126 42740 6132 42804
rect 6196 42802 6243 42804
rect 8293 42804 8359 42805
rect 6196 42800 6288 42802
rect 6238 42744 6288 42800
rect 6196 42742 6288 42744
rect 8293 42800 8340 42804
rect 8404 42802 8410 42804
rect 8293 42744 8298 42800
rect 6196 42740 6243 42742
rect 6177 42739 6243 42740
rect 8293 42740 8340 42744
rect 8404 42742 8450 42802
rect 10182 42800 10291 42805
rect 10961 42802 11027 42805
rect 10182 42744 10230 42800
rect 10286 42744 10291 42800
rect 10182 42742 10291 42744
rect 8404 42740 8410 42742
rect 8293 42739 8359 42740
rect 10225 42739 10291 42742
rect 10366 42800 11027 42802
rect 10366 42744 10966 42800
rect 11022 42744 11027 42800
rect 10366 42742 11027 42744
rect 0 42666 480 42696
rect 1945 42666 2011 42669
rect 0 42664 2011 42666
rect 0 42608 1950 42664
rect 2006 42608 2011 42664
rect 0 42606 2011 42608
rect 0 42576 480 42606
rect 1945 42603 2011 42606
rect 7557 42666 7623 42669
rect 9581 42666 9647 42669
rect 7557 42664 9647 42666
rect 7557 42608 7562 42664
rect 7618 42608 9586 42664
rect 9642 42608 9647 42664
rect 7557 42606 9647 42608
rect 7557 42603 7623 42606
rect 9581 42603 9647 42606
rect 10225 42666 10291 42669
rect 10366 42666 10426 42742
rect 10961 42739 11027 42742
rect 16021 42804 16087 42805
rect 16021 42800 16068 42804
rect 16132 42802 16138 42804
rect 16389 42802 16455 42805
rect 16021 42744 16026 42800
rect 16021 42740 16068 42744
rect 16132 42742 16178 42802
rect 16389 42800 18154 42802
rect 16389 42744 16394 42800
rect 16450 42744 18154 42800
rect 16389 42742 18154 42744
rect 16132 42740 16138 42742
rect 16021 42739 16087 42740
rect 16389 42739 16455 42742
rect 10225 42664 10426 42666
rect 10225 42608 10230 42664
rect 10286 42608 10426 42664
rect 10225 42606 10426 42608
rect 10777 42666 10843 42669
rect 13169 42666 13235 42669
rect 10777 42664 13235 42666
rect 10777 42608 10782 42664
rect 10838 42608 13174 42664
rect 13230 42608 13235 42664
rect 10777 42606 13235 42608
rect 10225 42603 10291 42606
rect 10777 42603 10843 42606
rect 13169 42603 13235 42606
rect 4277 42464 4597 42465
rect 4277 42400 4285 42464
rect 4349 42400 4365 42464
rect 4429 42400 4445 42464
rect 4509 42400 4525 42464
rect 4589 42400 4597 42464
rect 4277 42399 4597 42400
rect 10944 42464 11264 42465
rect 10944 42400 10952 42464
rect 11016 42400 11032 42464
rect 11096 42400 11112 42464
rect 11176 42400 11192 42464
rect 11256 42400 11264 42464
rect 10944 42399 11264 42400
rect 17610 42464 17930 42465
rect 17610 42400 17618 42464
rect 17682 42400 17698 42464
rect 17762 42400 17778 42464
rect 17842 42400 17858 42464
rect 17922 42400 17930 42464
rect 17610 42399 17930 42400
rect 5165 42394 5231 42397
rect 5030 42392 5231 42394
rect 5030 42336 5170 42392
rect 5226 42336 5231 42392
rect 5030 42334 5231 42336
rect 0 41850 480 41880
rect 5030 41853 5090 42334
rect 5165 42331 5231 42334
rect 15929 42392 15995 42397
rect 15929 42336 15934 42392
rect 15990 42336 15995 42392
rect 15929 42331 15995 42336
rect 5165 42258 5231 42261
rect 6913 42258 6979 42261
rect 5165 42256 6979 42258
rect 5165 42200 5170 42256
rect 5226 42200 6918 42256
rect 6974 42200 6979 42256
rect 5165 42198 6979 42200
rect 5165 42195 5231 42198
rect 6913 42195 6979 42198
rect 7741 42258 7807 42261
rect 11605 42260 11671 42261
rect 8702 42258 8708 42260
rect 7741 42256 8708 42258
rect 7741 42200 7746 42256
rect 7802 42200 8708 42256
rect 7741 42198 8708 42200
rect 7741 42195 7807 42198
rect 8702 42196 8708 42198
rect 8772 42196 8778 42260
rect 11605 42256 11652 42260
rect 11716 42258 11722 42260
rect 12985 42258 13051 42261
rect 15285 42258 15351 42261
rect 15932 42258 15992 42331
rect 11605 42200 11610 42256
rect 11605 42196 11652 42200
rect 11716 42198 11762 42258
rect 12985 42256 14658 42258
rect 12985 42200 12990 42256
rect 13046 42200 14658 42256
rect 12985 42198 14658 42200
rect 11716 42196 11722 42198
rect 11605 42195 11671 42196
rect 12985 42195 13051 42198
rect 6678 42060 6684 42124
rect 6748 42122 6754 42124
rect 6913 42122 6979 42125
rect 6748 42120 6979 42122
rect 6748 42064 6918 42120
rect 6974 42064 6979 42120
rect 6748 42062 6979 42064
rect 14598 42122 14658 42198
rect 15285 42256 15992 42258
rect 15285 42200 15290 42256
rect 15346 42200 15992 42256
rect 15285 42198 15992 42200
rect 15285 42195 15351 42198
rect 17953 42122 18019 42125
rect 14598 42120 18019 42122
rect 14598 42064 17958 42120
rect 18014 42064 18019 42120
rect 14598 42062 18019 42064
rect 6748 42060 6754 42062
rect 6913 42059 6979 42062
rect 17953 42059 18019 42062
rect 5574 41924 5580 41988
rect 5644 41986 5650 41988
rect 5717 41986 5783 41989
rect 5644 41984 5783 41986
rect 5644 41928 5722 41984
rect 5778 41928 5783 41984
rect 5644 41926 5783 41928
rect 18094 41986 18154 42742
rect 18229 42666 18295 42669
rect 19520 42666 20000 42696
rect 18229 42664 20000 42666
rect 18229 42608 18234 42664
rect 18290 42608 20000 42664
rect 18229 42606 20000 42608
rect 18229 42603 18295 42606
rect 19520 42576 20000 42606
rect 19520 41986 20000 42016
rect 18094 41926 20000 41986
rect 5644 41924 5650 41926
rect 5717 41923 5783 41926
rect 7610 41920 7930 41921
rect 7610 41856 7618 41920
rect 7682 41856 7698 41920
rect 7762 41856 7778 41920
rect 7842 41856 7858 41920
rect 7922 41856 7930 41920
rect 7610 41855 7930 41856
rect 14277 41920 14597 41921
rect 14277 41856 14285 41920
rect 14349 41856 14365 41920
rect 14429 41856 14445 41920
rect 14509 41856 14525 41920
rect 14589 41856 14597 41920
rect 19520 41896 20000 41926
rect 14277 41855 14597 41856
rect 1485 41850 1551 41853
rect 0 41848 1551 41850
rect 0 41792 1490 41848
rect 1546 41792 1551 41848
rect 0 41790 1551 41792
rect 5030 41848 5139 41853
rect 5030 41792 5078 41848
rect 5134 41792 5139 41848
rect 5030 41790 5139 41792
rect 0 41760 480 41790
rect 1485 41787 1551 41790
rect 5073 41787 5139 41790
rect 16798 41788 16804 41852
rect 16868 41850 16874 41852
rect 17769 41850 17835 41853
rect 16868 41848 17835 41850
rect 16868 41792 17774 41848
rect 17830 41792 17835 41848
rect 16868 41790 17835 41792
rect 16868 41788 16874 41790
rect 17769 41787 17835 41790
rect 5993 41714 6059 41717
rect 8937 41714 9003 41717
rect 5993 41712 9003 41714
rect 5993 41656 5998 41712
rect 6054 41656 8942 41712
rect 8998 41656 9003 41712
rect 5993 41654 9003 41656
rect 5993 41651 6059 41654
rect 8937 41651 9003 41654
rect 15561 41714 15627 41717
rect 15745 41714 15811 41717
rect 15561 41712 15811 41714
rect 15561 41656 15566 41712
rect 15622 41656 15750 41712
rect 15806 41656 15811 41712
rect 15561 41654 15811 41656
rect 15561 41651 15627 41654
rect 15745 41651 15811 41654
rect 16757 41714 16823 41717
rect 16982 41714 16988 41716
rect 16757 41712 16988 41714
rect 16757 41656 16762 41712
rect 16818 41656 16988 41712
rect 16757 41654 16988 41656
rect 16757 41651 16823 41654
rect 16982 41652 16988 41654
rect 17052 41652 17058 41716
rect 2865 41578 2931 41581
rect 7097 41578 7163 41581
rect 2865 41576 7163 41578
rect 2865 41520 2870 41576
rect 2926 41520 7102 41576
rect 7158 41520 7163 41576
rect 2865 41518 7163 41520
rect 2865 41515 2931 41518
rect 1577 41440 1643 41445
rect 1577 41384 1582 41440
rect 1638 41384 1643 41440
rect 1577 41379 1643 41384
rect 0 41034 480 41064
rect 1580 41034 1640 41379
rect 4110 41170 4170 41518
rect 7097 41515 7163 41518
rect 9213 41578 9279 41581
rect 13169 41578 13235 41581
rect 9213 41576 13235 41578
rect 9213 41520 9218 41576
rect 9274 41520 13174 41576
rect 13230 41520 13235 41576
rect 9213 41518 13235 41520
rect 9213 41515 9279 41518
rect 13169 41515 13235 41518
rect 15326 41516 15332 41580
rect 15396 41578 15402 41580
rect 15469 41578 15535 41581
rect 15396 41576 15535 41578
rect 15396 41520 15474 41576
rect 15530 41520 15535 41576
rect 15396 41518 15535 41520
rect 15396 41516 15402 41518
rect 15469 41515 15535 41518
rect 16389 41580 16455 41581
rect 16389 41576 16436 41580
rect 16500 41578 16506 41580
rect 16389 41520 16394 41576
rect 16389 41516 16436 41520
rect 16500 41518 16546 41578
rect 16500 41516 16506 41518
rect 16389 41515 16455 41516
rect 5625 41442 5691 41445
rect 5758 41442 5764 41444
rect 5625 41440 5764 41442
rect 5625 41384 5630 41440
rect 5686 41384 5764 41440
rect 5625 41382 5764 41384
rect 5625 41379 5691 41382
rect 5758 41380 5764 41382
rect 5828 41380 5834 41444
rect 6269 41442 6335 41445
rect 6678 41442 6684 41444
rect 6269 41440 6684 41442
rect 6269 41384 6274 41440
rect 6330 41384 6684 41440
rect 6269 41382 6684 41384
rect 6269 41379 6335 41382
rect 6678 41380 6684 41382
rect 6748 41380 6754 41444
rect 9254 41380 9260 41444
rect 9324 41442 9330 41444
rect 9489 41442 9555 41445
rect 9324 41440 9555 41442
rect 9324 41384 9494 41440
rect 9550 41384 9555 41440
rect 9324 41382 9555 41384
rect 9324 41380 9330 41382
rect 9489 41379 9555 41382
rect 11513 41442 11579 41445
rect 13997 41442 14063 41445
rect 17033 41444 17099 41445
rect 16798 41442 16804 41444
rect 11513 41440 12312 41442
rect 11513 41384 11518 41440
rect 11574 41384 12312 41440
rect 11513 41382 12312 41384
rect 11513 41379 11579 41382
rect 4277 41376 4597 41377
rect 4277 41312 4285 41376
rect 4349 41312 4365 41376
rect 4429 41312 4445 41376
rect 4509 41312 4525 41376
rect 4589 41312 4597 41376
rect 4277 41311 4597 41312
rect 10944 41376 11264 41377
rect 10944 41312 10952 41376
rect 11016 41312 11032 41376
rect 11096 41312 11112 41376
rect 11176 41312 11192 41376
rect 11256 41312 11264 41376
rect 10944 41311 11264 41312
rect 6269 41306 6335 41309
rect 6678 41306 6684 41308
rect 6269 41304 6684 41306
rect 6269 41248 6274 41304
rect 6330 41248 6684 41304
rect 6269 41246 6684 41248
rect 6269 41243 6335 41246
rect 6678 41244 6684 41246
rect 6748 41244 6754 41308
rect 7005 41306 7071 41309
rect 8334 41306 8340 41308
rect 7005 41304 8340 41306
rect 7005 41248 7010 41304
rect 7066 41248 8340 41304
rect 7005 41246 8340 41248
rect 7005 41243 7071 41246
rect 8334 41244 8340 41246
rect 8404 41244 8410 41308
rect 12252 41173 12312 41382
rect 13997 41440 16804 41442
rect 13997 41384 14002 41440
rect 14058 41384 16804 41440
rect 13997 41382 16804 41384
rect 13997 41379 14063 41382
rect 16798 41380 16804 41382
rect 16868 41380 16874 41444
rect 16982 41380 16988 41444
rect 17052 41442 17099 41444
rect 17052 41440 17144 41442
rect 17094 41384 17144 41440
rect 17052 41382 17144 41384
rect 17052 41380 17099 41382
rect 17033 41379 17099 41380
rect 17610 41376 17930 41377
rect 17610 41312 17618 41376
rect 17682 41312 17698 41376
rect 17762 41312 17778 41376
rect 17842 41312 17858 41376
rect 17922 41312 17930 41376
rect 17610 41311 17930 41312
rect 14917 41306 14983 41309
rect 14917 41304 15210 41306
rect 14917 41248 14922 41304
rect 14978 41248 15210 41304
rect 14917 41246 15210 41248
rect 14917 41243 14983 41246
rect 4245 41170 4311 41173
rect 4110 41168 4311 41170
rect 4110 41112 4250 41168
rect 4306 41112 4311 41168
rect 4110 41110 4311 41112
rect 4245 41107 4311 41110
rect 5625 41170 5691 41173
rect 5758 41170 5764 41172
rect 5625 41168 5764 41170
rect 5625 41112 5630 41168
rect 5686 41112 5764 41168
rect 5625 41110 5764 41112
rect 5625 41107 5691 41110
rect 5758 41108 5764 41110
rect 5828 41108 5834 41172
rect 12249 41168 12315 41173
rect 12249 41112 12254 41168
rect 12310 41112 12315 41168
rect 12249 41107 12315 41112
rect 13670 41108 13676 41172
rect 13740 41170 13746 41172
rect 14774 41170 14780 41172
rect 13740 41110 14780 41170
rect 13740 41108 13746 41110
rect 14774 41108 14780 41110
rect 14844 41108 14850 41172
rect 15150 41170 15210 41246
rect 15326 41244 15332 41308
rect 15396 41306 15402 41308
rect 15561 41306 15627 41309
rect 15396 41304 15627 41306
rect 15396 41248 15566 41304
rect 15622 41248 15627 41304
rect 15396 41246 15627 41248
rect 15396 41244 15402 41246
rect 15561 41243 15627 41246
rect 16798 41244 16804 41308
rect 16868 41306 16874 41308
rect 17033 41306 17099 41309
rect 19520 41306 20000 41336
rect 16868 41304 17099 41306
rect 16868 41248 17038 41304
rect 17094 41248 17099 41304
rect 16868 41246 17099 41248
rect 16868 41244 16874 41246
rect 17033 41243 17099 41246
rect 18094 41246 20000 41306
rect 15878 41170 15884 41172
rect 15150 41110 15884 41170
rect 15878 41108 15884 41110
rect 15948 41108 15954 41172
rect 16297 41170 16363 41173
rect 18094 41170 18154 41246
rect 19520 41216 20000 41246
rect 16297 41168 18154 41170
rect 16297 41112 16302 41168
rect 16358 41112 18154 41168
rect 16297 41110 18154 41112
rect 16297 41107 16363 41110
rect 0 40974 1640 41034
rect 5625 41034 5691 41037
rect 7281 41034 7347 41037
rect 5625 41032 7347 41034
rect 5625 40976 5630 41032
rect 5686 40976 7286 41032
rect 7342 40976 7347 41032
rect 5625 40974 7347 40976
rect 0 40944 480 40974
rect 5625 40971 5691 40974
rect 7281 40971 7347 40974
rect 7465 41034 7531 41037
rect 13486 41034 13492 41036
rect 7465 41032 13492 41034
rect 7465 40976 7470 41032
rect 7526 40976 13492 41032
rect 7465 40974 13492 40976
rect 7465 40971 7531 40974
rect 13486 40972 13492 40974
rect 13556 41034 13562 41036
rect 14549 41034 14615 41037
rect 13556 41032 14615 41034
rect 13556 40976 14554 41032
rect 14610 40976 14615 41032
rect 13556 40974 14615 40976
rect 13556 40972 13562 40974
rect 14549 40971 14615 40974
rect 14774 40972 14780 41036
rect 14844 41034 14850 41036
rect 15142 41034 15148 41036
rect 14844 40974 15148 41034
rect 14844 40972 14850 40974
rect 15142 40972 15148 40974
rect 15212 40972 15218 41036
rect 5533 40900 5599 40901
rect 5533 40898 5580 40900
rect 5488 40896 5580 40898
rect 5488 40840 5538 40896
rect 5488 40838 5580 40840
rect 5533 40836 5580 40838
rect 5644 40836 5650 40900
rect 5533 40835 5599 40836
rect 7610 40832 7930 40833
rect 7610 40768 7618 40832
rect 7682 40768 7698 40832
rect 7762 40768 7778 40832
rect 7842 40768 7858 40832
rect 7922 40768 7930 40832
rect 7610 40767 7930 40768
rect 14277 40832 14597 40833
rect 14277 40768 14285 40832
rect 14349 40768 14365 40832
rect 14429 40768 14445 40832
rect 14509 40768 14525 40832
rect 14589 40768 14597 40832
rect 14277 40767 14597 40768
rect 15193 40762 15259 40765
rect 15510 40762 15516 40764
rect 15193 40760 15516 40762
rect 15193 40704 15198 40760
rect 15254 40704 15516 40760
rect 15193 40702 15516 40704
rect 15193 40699 15259 40702
rect 15510 40700 15516 40702
rect 15580 40700 15586 40764
rect 2681 40626 2747 40629
rect 8334 40626 8340 40628
rect 2681 40624 8340 40626
rect 2681 40568 2686 40624
rect 2742 40568 8340 40624
rect 2681 40566 8340 40568
rect 2681 40563 2747 40566
rect 8334 40564 8340 40566
rect 8404 40626 8410 40628
rect 10317 40626 10383 40629
rect 8404 40624 10383 40626
rect 8404 40568 10322 40624
rect 10378 40568 10383 40624
rect 8404 40566 10383 40568
rect 8404 40564 8410 40566
rect 10317 40563 10383 40566
rect 10869 40626 10935 40629
rect 13813 40626 13879 40629
rect 10869 40624 13879 40626
rect 10869 40568 10874 40624
rect 10930 40568 13818 40624
rect 13874 40568 13879 40624
rect 10869 40566 13879 40568
rect 10869 40563 10935 40566
rect 13813 40563 13879 40566
rect 16205 40626 16271 40629
rect 19520 40626 20000 40656
rect 16205 40624 20000 40626
rect 16205 40568 16210 40624
rect 16266 40568 20000 40624
rect 16205 40566 20000 40568
rect 16205 40563 16271 40566
rect 19520 40536 20000 40566
rect 6177 40490 6243 40493
rect 9029 40490 9095 40493
rect 12341 40490 12407 40493
rect 6177 40488 12407 40490
rect 6177 40432 6182 40488
rect 6238 40432 9034 40488
rect 9090 40432 12346 40488
rect 12402 40432 12407 40488
rect 6177 40430 12407 40432
rect 6177 40427 6243 40430
rect 9029 40427 9095 40430
rect 12341 40427 12407 40430
rect 0 40354 480 40384
rect 1577 40354 1643 40357
rect 0 40352 1643 40354
rect 0 40296 1582 40352
rect 1638 40296 1643 40352
rect 0 40294 1643 40296
rect 0 40264 480 40294
rect 1577 40291 1643 40294
rect 16430 40292 16436 40356
rect 16500 40354 16506 40356
rect 17217 40354 17283 40357
rect 16500 40352 17283 40354
rect 16500 40296 17222 40352
rect 17278 40296 17283 40352
rect 16500 40294 17283 40296
rect 16500 40292 16506 40294
rect 17217 40291 17283 40294
rect 4277 40288 4597 40289
rect 4277 40224 4285 40288
rect 4349 40224 4365 40288
rect 4429 40224 4445 40288
rect 4509 40224 4525 40288
rect 4589 40224 4597 40288
rect 4277 40223 4597 40224
rect 10944 40288 11264 40289
rect 10944 40224 10952 40288
rect 11016 40224 11032 40288
rect 11096 40224 11112 40288
rect 11176 40224 11192 40288
rect 11256 40224 11264 40288
rect 10944 40223 11264 40224
rect 17610 40288 17930 40289
rect 17610 40224 17618 40288
rect 17682 40224 17698 40288
rect 17762 40224 17778 40288
rect 17842 40224 17858 40288
rect 17922 40224 17930 40288
rect 17610 40223 17930 40224
rect 3693 40218 3759 40221
rect 3918 40218 3924 40220
rect 3693 40216 3924 40218
rect 3693 40160 3698 40216
rect 3754 40160 3924 40216
rect 3693 40158 3924 40160
rect 3693 40155 3759 40158
rect 3918 40156 3924 40158
rect 3988 40156 3994 40220
rect 17217 40084 17283 40085
rect 17166 40020 17172 40084
rect 17236 40082 17283 40084
rect 17236 40080 17328 40082
rect 17278 40024 17328 40080
rect 17236 40022 17328 40024
rect 17236 40020 17283 40022
rect 17217 40019 17283 40020
rect 4102 39884 4108 39948
rect 4172 39946 4178 39948
rect 4337 39946 4403 39949
rect 4172 39944 4403 39946
rect 4172 39888 4342 39944
rect 4398 39888 4403 39944
rect 4172 39886 4403 39888
rect 4172 39884 4178 39886
rect 4337 39883 4403 39886
rect 6177 39946 6243 39949
rect 11697 39948 11763 39949
rect 11462 39946 11468 39948
rect 6177 39944 11468 39946
rect 6177 39888 6182 39944
rect 6238 39888 11468 39944
rect 6177 39886 11468 39888
rect 6177 39883 6243 39886
rect 11462 39884 11468 39886
rect 11532 39884 11538 39948
rect 11646 39884 11652 39948
rect 11716 39946 11763 39948
rect 16481 39946 16547 39949
rect 19520 39946 20000 39976
rect 11716 39944 11808 39946
rect 11758 39888 11808 39944
rect 11716 39886 11808 39888
rect 16481 39944 20000 39946
rect 16481 39888 16486 39944
rect 16542 39888 20000 39944
rect 16481 39886 20000 39888
rect 11716 39884 11763 39886
rect 11697 39883 11763 39884
rect 16481 39883 16547 39886
rect 19520 39856 20000 39886
rect 6177 39810 6243 39813
rect 6310 39810 6316 39812
rect 6177 39808 6316 39810
rect 6177 39752 6182 39808
rect 6238 39752 6316 39808
rect 6177 39750 6316 39752
rect 6177 39747 6243 39750
rect 6310 39748 6316 39750
rect 6380 39748 6386 39812
rect 10869 39810 10935 39813
rect 13077 39810 13143 39813
rect 10869 39808 13143 39810
rect 10869 39752 10874 39808
rect 10930 39752 13082 39808
rect 13138 39752 13143 39808
rect 10869 39750 13143 39752
rect 10869 39747 10935 39750
rect 13077 39747 13143 39750
rect 7610 39744 7930 39745
rect 7610 39680 7618 39744
rect 7682 39680 7698 39744
rect 7762 39680 7778 39744
rect 7842 39680 7858 39744
rect 7922 39680 7930 39744
rect 7610 39679 7930 39680
rect 14277 39744 14597 39745
rect 14277 39680 14285 39744
rect 14349 39680 14365 39744
rect 14429 39680 14445 39744
rect 14509 39680 14525 39744
rect 14589 39680 14597 39744
rect 14277 39679 14597 39680
rect 8109 39674 8175 39677
rect 11697 39674 11763 39677
rect 8109 39672 11763 39674
rect 8109 39616 8114 39672
rect 8170 39616 11702 39672
rect 11758 39616 11763 39672
rect 8109 39614 11763 39616
rect 8109 39611 8175 39614
rect 11697 39611 11763 39614
rect 0 39538 480 39568
rect 2129 39538 2195 39541
rect 0 39536 2195 39538
rect 0 39480 2134 39536
rect 2190 39480 2195 39536
rect 0 39478 2195 39480
rect 0 39448 480 39478
rect 2129 39475 2195 39478
rect 5993 39538 6059 39541
rect 9397 39538 9463 39541
rect 5993 39536 9463 39538
rect 5993 39480 5998 39536
rect 6054 39480 9402 39536
rect 9458 39480 9463 39536
rect 5993 39478 9463 39480
rect 5993 39475 6059 39478
rect 9397 39475 9463 39478
rect 13486 39476 13492 39540
rect 13556 39538 13562 39540
rect 14641 39538 14707 39541
rect 13556 39536 14707 39538
rect 13556 39480 14646 39536
rect 14702 39480 14707 39536
rect 13556 39478 14707 39480
rect 13556 39476 13562 39478
rect 14641 39475 14707 39478
rect 15929 39538 15995 39541
rect 16062 39538 16068 39540
rect 15929 39536 16068 39538
rect 15929 39480 15934 39536
rect 15990 39480 16068 39536
rect 15929 39478 16068 39480
rect 15929 39475 15995 39478
rect 16062 39476 16068 39478
rect 16132 39476 16138 39540
rect 16297 39538 16363 39541
rect 18229 39538 18295 39541
rect 16297 39536 18295 39538
rect 16297 39480 16302 39536
rect 16358 39480 18234 39536
rect 18290 39480 18295 39536
rect 16297 39478 18295 39480
rect 16297 39475 16363 39478
rect 18229 39475 18295 39478
rect 2681 39402 2747 39405
rect 7557 39402 7623 39405
rect 11513 39402 11579 39405
rect 12566 39402 12572 39404
rect 2681 39400 12572 39402
rect 2681 39344 2686 39400
rect 2742 39344 7562 39400
rect 7618 39344 11518 39400
rect 11574 39344 12572 39400
rect 2681 39342 12572 39344
rect 2681 39339 2747 39342
rect 7557 39339 7623 39342
rect 11513 39339 11579 39342
rect 12566 39340 12572 39342
rect 12636 39340 12642 39404
rect 15101 39402 15167 39405
rect 15101 39400 18154 39402
rect 15101 39344 15106 39400
rect 15162 39344 18154 39400
rect 15101 39342 18154 39344
rect 15101 39339 15167 39342
rect 15510 39204 15516 39268
rect 15580 39266 15586 39268
rect 15653 39266 15719 39269
rect 15580 39264 15719 39266
rect 15580 39208 15658 39264
rect 15714 39208 15719 39264
rect 15580 39206 15719 39208
rect 18094 39266 18154 39342
rect 19520 39266 20000 39296
rect 18094 39206 20000 39266
rect 15580 39204 15586 39206
rect 15653 39203 15719 39206
rect 4277 39200 4597 39201
rect 4277 39136 4285 39200
rect 4349 39136 4365 39200
rect 4429 39136 4445 39200
rect 4509 39136 4525 39200
rect 4589 39136 4597 39200
rect 4277 39135 4597 39136
rect 10944 39200 11264 39201
rect 10944 39136 10952 39200
rect 11016 39136 11032 39200
rect 11096 39136 11112 39200
rect 11176 39136 11192 39200
rect 11256 39136 11264 39200
rect 10944 39135 11264 39136
rect 17610 39200 17930 39201
rect 17610 39136 17618 39200
rect 17682 39136 17698 39200
rect 17762 39136 17778 39200
rect 17842 39136 17858 39200
rect 17922 39136 17930 39200
rect 19520 39176 20000 39206
rect 17610 39135 17930 39136
rect 9990 39068 9996 39132
rect 10060 39130 10066 39132
rect 10317 39130 10383 39133
rect 10060 39128 10383 39130
rect 10060 39072 10322 39128
rect 10378 39072 10383 39128
rect 10060 39070 10383 39072
rect 10060 39068 10066 39070
rect 10317 39067 10383 39070
rect 7649 38994 7715 38997
rect 9213 38994 9279 38997
rect 12198 38994 12204 38996
rect 7649 38992 12204 38994
rect 7649 38936 7654 38992
rect 7710 38936 9218 38992
rect 9274 38936 12204 38992
rect 7649 38934 12204 38936
rect 7649 38931 7715 38934
rect 9213 38931 9279 38934
rect 12198 38932 12204 38934
rect 12268 38932 12274 38996
rect 11973 38858 12039 38861
rect 614 38856 12039 38858
rect 614 38800 11978 38856
rect 12034 38800 12039 38856
rect 614 38798 12039 38800
rect 0 38722 480 38752
rect 614 38722 674 38798
rect 11973 38795 12039 38798
rect 0 38662 674 38722
rect 9213 38722 9279 38725
rect 9673 38722 9739 38725
rect 9213 38720 9739 38722
rect 9213 38664 9218 38720
rect 9274 38664 9678 38720
rect 9734 38664 9739 38720
rect 9213 38662 9739 38664
rect 0 38632 480 38662
rect 9213 38659 9279 38662
rect 9673 38659 9739 38662
rect 9949 38722 10015 38725
rect 10501 38722 10567 38725
rect 11053 38722 11119 38725
rect 9949 38720 11119 38722
rect 9949 38664 9954 38720
rect 10010 38664 10506 38720
rect 10562 38664 11058 38720
rect 11114 38664 11119 38720
rect 9949 38662 11119 38664
rect 9949 38659 10015 38662
rect 10501 38659 10567 38662
rect 11053 38659 11119 38662
rect 11237 38722 11303 38725
rect 12750 38722 12756 38724
rect 11237 38720 12756 38722
rect 11237 38664 11242 38720
rect 11298 38664 12756 38720
rect 11237 38662 12756 38664
rect 11237 38659 11303 38662
rect 12750 38660 12756 38662
rect 12820 38660 12826 38724
rect 7610 38656 7930 38657
rect 7610 38592 7618 38656
rect 7682 38592 7698 38656
rect 7762 38592 7778 38656
rect 7842 38592 7858 38656
rect 7922 38592 7930 38656
rect 7610 38591 7930 38592
rect 14277 38656 14597 38657
rect 14277 38592 14285 38656
rect 14349 38592 14365 38656
rect 14429 38592 14445 38656
rect 14509 38592 14525 38656
rect 14589 38592 14597 38656
rect 14277 38591 14597 38592
rect 8293 38586 8359 38589
rect 13721 38586 13787 38589
rect 8293 38584 13787 38586
rect 8293 38528 8298 38584
rect 8354 38528 13726 38584
rect 13782 38528 13787 38584
rect 8293 38526 13787 38528
rect 8293 38523 8359 38526
rect 13721 38523 13787 38526
rect 15878 38524 15884 38588
rect 15948 38586 15954 38588
rect 19520 38586 20000 38616
rect 15948 38526 20000 38586
rect 15948 38524 15954 38526
rect 19520 38496 20000 38526
rect 2589 38450 2655 38453
rect 8293 38450 8359 38453
rect 2589 38448 8359 38450
rect 2589 38392 2594 38448
rect 2650 38392 8298 38448
rect 8354 38392 8359 38448
rect 2589 38390 8359 38392
rect 2589 38387 2655 38390
rect 8293 38387 8359 38390
rect 8702 38388 8708 38452
rect 8772 38450 8778 38452
rect 10501 38450 10567 38453
rect 8772 38448 10567 38450
rect 8772 38392 10506 38448
rect 10562 38392 10567 38448
rect 8772 38390 10567 38392
rect 8772 38388 8778 38390
rect 10501 38387 10567 38390
rect 3233 38314 3299 38317
rect 9029 38314 9095 38317
rect 12341 38314 12407 38317
rect 3233 38312 12407 38314
rect 3233 38256 3238 38312
rect 3294 38256 9034 38312
rect 9090 38256 12346 38312
rect 12402 38256 12407 38312
rect 3233 38254 12407 38256
rect 3233 38251 3299 38254
rect 9029 38251 9095 38254
rect 12341 38251 12407 38254
rect 14641 38314 14707 38317
rect 15142 38314 15148 38316
rect 14641 38312 15148 38314
rect 14641 38256 14646 38312
rect 14702 38256 15148 38312
rect 14641 38254 15148 38256
rect 14641 38251 14707 38254
rect 15142 38252 15148 38254
rect 15212 38252 15218 38316
rect 6862 38116 6868 38180
rect 6932 38178 6938 38180
rect 7281 38178 7347 38181
rect 6932 38176 7347 38178
rect 6932 38120 7286 38176
rect 7342 38120 7347 38176
rect 6932 38118 7347 38120
rect 6932 38116 6938 38118
rect 7281 38115 7347 38118
rect 11973 38178 12039 38181
rect 12709 38178 12775 38181
rect 13353 38178 13419 38181
rect 11973 38176 13419 38178
rect 11973 38120 11978 38176
rect 12034 38120 12714 38176
rect 12770 38120 13358 38176
rect 13414 38120 13419 38176
rect 11973 38118 13419 38120
rect 11973 38115 12039 38118
rect 12709 38115 12775 38118
rect 13353 38115 13419 38118
rect 4277 38112 4597 38113
rect 4277 38048 4285 38112
rect 4349 38048 4365 38112
rect 4429 38048 4445 38112
rect 4509 38048 4525 38112
rect 4589 38048 4597 38112
rect 4277 38047 4597 38048
rect 10944 38112 11264 38113
rect 10944 38048 10952 38112
rect 11016 38048 11032 38112
rect 11096 38048 11112 38112
rect 11176 38048 11192 38112
rect 11256 38048 11264 38112
rect 10944 38047 11264 38048
rect 17610 38112 17930 38113
rect 17610 38048 17618 38112
rect 17682 38048 17698 38112
rect 17762 38048 17778 38112
rect 17842 38048 17858 38112
rect 17922 38048 17930 38112
rect 17610 38047 17930 38048
rect 0 37906 480 37936
rect 3509 37906 3575 37909
rect 0 37904 3575 37906
rect 0 37848 3514 37904
rect 3570 37848 3575 37904
rect 0 37846 3575 37848
rect 0 37816 480 37846
rect 3509 37843 3575 37846
rect 9121 37906 9187 37909
rect 11237 37906 11303 37909
rect 9121 37904 11303 37906
rect 9121 37848 9126 37904
rect 9182 37848 11242 37904
rect 11298 37848 11303 37904
rect 9121 37846 11303 37848
rect 9121 37843 9187 37846
rect 11237 37843 11303 37846
rect 15101 37906 15167 37909
rect 19520 37906 20000 37936
rect 15101 37904 20000 37906
rect 15101 37848 15106 37904
rect 15162 37848 20000 37904
rect 15101 37846 20000 37848
rect 15101 37843 15167 37846
rect 19520 37816 20000 37846
rect 6729 37770 6795 37773
rect 9581 37770 9647 37773
rect 6729 37768 9647 37770
rect 6729 37712 6734 37768
rect 6790 37712 9586 37768
rect 9642 37712 9647 37768
rect 6729 37710 9647 37712
rect 6729 37707 6795 37710
rect 9581 37707 9647 37710
rect 7610 37568 7930 37569
rect 7610 37504 7618 37568
rect 7682 37504 7698 37568
rect 7762 37504 7778 37568
rect 7842 37504 7858 37568
rect 7922 37504 7930 37568
rect 7610 37503 7930 37504
rect 14277 37568 14597 37569
rect 14277 37504 14285 37568
rect 14349 37504 14365 37568
rect 14429 37504 14445 37568
rect 14509 37504 14525 37568
rect 14589 37504 14597 37568
rect 14277 37503 14597 37504
rect 15377 37500 15443 37501
rect 15326 37436 15332 37500
rect 15396 37498 15443 37500
rect 15396 37496 15488 37498
rect 15438 37440 15488 37496
rect 15396 37438 15488 37440
rect 15396 37436 15443 37438
rect 15334 37435 15443 37436
rect 5257 37362 5323 37365
rect 7373 37362 7439 37365
rect 5257 37360 7439 37362
rect 5257 37304 5262 37360
rect 5318 37304 7378 37360
rect 7434 37304 7439 37360
rect 5257 37302 7439 37304
rect 5257 37299 5323 37302
rect 7373 37299 7439 37302
rect 12893 37362 12959 37365
rect 15334 37362 15394 37435
rect 12893 37360 15394 37362
rect 12893 37304 12898 37360
rect 12954 37304 15394 37360
rect 12893 37302 15394 37304
rect 12893 37299 12959 37302
rect 14774 37226 14780 37228
rect 9676 37166 14780 37226
rect 0 37090 480 37120
rect 3785 37090 3851 37093
rect 0 37088 3851 37090
rect 0 37032 3790 37088
rect 3846 37032 3851 37088
rect 0 37030 3851 37032
rect 0 37000 480 37030
rect 3785 37027 3851 37030
rect 6729 37090 6795 37093
rect 7230 37090 7236 37092
rect 6729 37088 7236 37090
rect 6729 37032 6734 37088
rect 6790 37032 7236 37088
rect 6729 37030 7236 37032
rect 6729 37027 6795 37030
rect 7230 37028 7236 37030
rect 7300 37090 7306 37092
rect 7925 37090 7991 37093
rect 7300 37088 7991 37090
rect 7300 37032 7930 37088
rect 7986 37032 7991 37088
rect 7300 37030 7991 37032
rect 7300 37028 7306 37030
rect 7925 37027 7991 37030
rect 4277 37024 4597 37025
rect 4277 36960 4285 37024
rect 4349 36960 4365 37024
rect 4429 36960 4445 37024
rect 4509 36960 4525 37024
rect 4589 36960 4597 37024
rect 4277 36959 4597 36960
rect 3417 36818 3483 36821
rect 9676 36818 9736 37166
rect 14774 37164 14780 37166
rect 14844 37164 14850 37228
rect 15377 37226 15443 37229
rect 16798 37226 16804 37228
rect 15377 37224 16804 37226
rect 15377 37168 15382 37224
rect 15438 37168 16804 37224
rect 15377 37166 16804 37168
rect 15377 37163 15443 37166
rect 16798 37164 16804 37166
rect 16868 37164 16874 37228
rect 17493 37226 17559 37229
rect 19520 37226 20000 37256
rect 17493 37224 20000 37226
rect 17493 37168 17498 37224
rect 17554 37168 20000 37224
rect 17493 37166 20000 37168
rect 17493 37163 17559 37166
rect 19520 37136 20000 37166
rect 10944 37024 11264 37025
rect 10944 36960 10952 37024
rect 11016 36960 11032 37024
rect 11096 36960 11112 37024
rect 11176 36960 11192 37024
rect 11256 36960 11264 37024
rect 10944 36959 11264 36960
rect 17610 37024 17930 37025
rect 17610 36960 17618 37024
rect 17682 36960 17698 37024
rect 17762 36960 17778 37024
rect 17842 36960 17858 37024
rect 17922 36960 17930 37024
rect 17610 36959 17930 36960
rect 3417 36816 9736 36818
rect 3417 36760 3422 36816
rect 3478 36760 9736 36816
rect 3417 36758 9736 36760
rect 3417 36755 3483 36758
rect 9806 36756 9812 36820
rect 9876 36818 9882 36820
rect 10501 36818 10567 36821
rect 9876 36816 10567 36818
rect 9876 36760 10506 36816
rect 10562 36760 10567 36816
rect 9876 36758 10567 36760
rect 9876 36756 9882 36758
rect 10501 36755 10567 36758
rect 6269 36682 6335 36685
rect 6269 36680 6378 36682
rect 6269 36624 6274 36680
rect 6330 36624 6378 36680
rect 6269 36619 6378 36624
rect 5809 36412 5875 36413
rect 5758 36348 5764 36412
rect 5828 36410 5875 36412
rect 6318 36410 6378 36619
rect 17125 36546 17191 36549
rect 19520 36546 20000 36576
rect 17125 36544 20000 36546
rect 17125 36488 17130 36544
rect 17186 36488 20000 36544
rect 17125 36486 20000 36488
rect 17125 36483 17191 36486
rect 7610 36480 7930 36481
rect 7610 36416 7618 36480
rect 7682 36416 7698 36480
rect 7762 36416 7778 36480
rect 7842 36416 7858 36480
rect 7922 36416 7930 36480
rect 7610 36415 7930 36416
rect 14277 36480 14597 36481
rect 14277 36416 14285 36480
rect 14349 36416 14365 36480
rect 14429 36416 14445 36480
rect 14509 36416 14525 36480
rect 14589 36416 14597 36480
rect 19520 36456 20000 36486
rect 14277 36415 14597 36416
rect 6821 36410 6887 36413
rect 5828 36408 5920 36410
rect 5870 36352 5920 36408
rect 5828 36350 5920 36352
rect 6318 36408 6887 36410
rect 6318 36352 6826 36408
rect 6882 36352 6887 36408
rect 6318 36350 6887 36352
rect 5828 36348 5875 36350
rect 5809 36347 5875 36348
rect 6821 36347 6887 36350
rect 0 36274 480 36304
rect 1853 36274 1919 36277
rect 0 36272 1919 36274
rect 0 36216 1858 36272
rect 1914 36216 1919 36272
rect 0 36214 1919 36216
rect 0 36184 480 36214
rect 1853 36211 1919 36214
rect 5993 36274 6059 36277
rect 13077 36274 13143 36277
rect 5993 36272 13143 36274
rect 5993 36216 5998 36272
rect 6054 36216 13082 36272
rect 13138 36216 13143 36272
rect 5993 36214 13143 36216
rect 5993 36211 6059 36214
rect 13077 36211 13143 36214
rect 4277 35936 4597 35937
rect 4277 35872 4285 35936
rect 4349 35872 4365 35936
rect 4429 35872 4445 35936
rect 4509 35872 4525 35936
rect 4589 35872 4597 35936
rect 4277 35871 4597 35872
rect 10944 35936 11264 35937
rect 10944 35872 10952 35936
rect 11016 35872 11032 35936
rect 11096 35872 11112 35936
rect 11176 35872 11192 35936
rect 11256 35872 11264 35936
rect 10944 35871 11264 35872
rect 17610 35936 17930 35937
rect 17610 35872 17618 35936
rect 17682 35872 17698 35936
rect 17762 35872 17778 35936
rect 17842 35872 17858 35936
rect 17922 35872 17930 35936
rect 17610 35871 17930 35872
rect 18045 35866 18111 35869
rect 19520 35866 20000 35896
rect 18045 35864 20000 35866
rect 18045 35808 18050 35864
rect 18106 35808 20000 35864
rect 18045 35806 20000 35808
rect 18045 35803 18111 35806
rect 19520 35776 20000 35806
rect 15653 35732 15719 35733
rect 15653 35730 15700 35732
rect 15608 35728 15700 35730
rect 15608 35672 15658 35728
rect 15608 35670 15700 35672
rect 15653 35668 15700 35670
rect 15764 35668 15770 35732
rect 15653 35667 15719 35668
rect 0 35458 480 35488
rect 1485 35458 1551 35461
rect 0 35456 1551 35458
rect 0 35400 1490 35456
rect 1546 35400 1551 35456
rect 0 35398 1551 35400
rect 0 35368 480 35398
rect 1485 35395 1551 35398
rect 7610 35392 7930 35393
rect 7610 35328 7618 35392
rect 7682 35328 7698 35392
rect 7762 35328 7778 35392
rect 7842 35328 7858 35392
rect 7922 35328 7930 35392
rect 7610 35327 7930 35328
rect 14277 35392 14597 35393
rect 14277 35328 14285 35392
rect 14349 35328 14365 35392
rect 14429 35328 14445 35392
rect 14509 35328 14525 35392
rect 14589 35328 14597 35392
rect 14277 35327 14597 35328
rect 17493 35186 17559 35189
rect 19520 35186 20000 35216
rect 17493 35184 20000 35186
rect 17493 35128 17498 35184
rect 17554 35128 20000 35184
rect 17493 35126 20000 35128
rect 17493 35123 17559 35126
rect 19520 35096 20000 35126
rect 3969 35050 4035 35053
rect 13670 35050 13676 35052
rect 3969 35048 13676 35050
rect 3969 34992 3974 35048
rect 4030 34992 13676 35048
rect 3969 34990 13676 34992
rect 3969 34987 4035 34990
rect 13670 34988 13676 34990
rect 13740 34988 13746 35052
rect 4277 34848 4597 34849
rect 4277 34784 4285 34848
rect 4349 34784 4365 34848
rect 4429 34784 4445 34848
rect 4509 34784 4525 34848
rect 4589 34784 4597 34848
rect 4277 34783 4597 34784
rect 10944 34848 11264 34849
rect 10944 34784 10952 34848
rect 11016 34784 11032 34848
rect 11096 34784 11112 34848
rect 11176 34784 11192 34848
rect 11256 34784 11264 34848
rect 10944 34783 11264 34784
rect 17610 34848 17930 34849
rect 17610 34784 17618 34848
rect 17682 34784 17698 34848
rect 17762 34784 17778 34848
rect 17842 34784 17858 34848
rect 17922 34784 17930 34848
rect 17610 34783 17930 34784
rect 0 34642 480 34672
rect 2313 34642 2379 34645
rect 0 34640 2379 34642
rect 0 34584 2318 34640
rect 2374 34584 2379 34640
rect 0 34582 2379 34584
rect 0 34552 480 34582
rect 2313 34579 2379 34582
rect 7925 34642 7991 34645
rect 8937 34642 9003 34645
rect 7925 34640 9003 34642
rect 7925 34584 7930 34640
rect 7986 34584 8942 34640
rect 8998 34584 9003 34640
rect 7925 34582 9003 34584
rect 7925 34579 7991 34582
rect 8937 34579 9003 34582
rect 7465 34506 7531 34509
rect 9581 34506 9647 34509
rect 7465 34504 9647 34506
rect 7465 34448 7470 34504
rect 7526 34448 9586 34504
rect 9642 34448 9647 34504
rect 7465 34446 9647 34448
rect 7465 34443 7531 34446
rect 9581 34443 9647 34446
rect 10777 34506 10843 34509
rect 14089 34506 14155 34509
rect 10777 34504 14155 34506
rect 10777 34448 10782 34504
rect 10838 34448 14094 34504
rect 14150 34448 14155 34504
rect 10777 34446 14155 34448
rect 10777 34443 10843 34446
rect 14089 34443 14155 34446
rect 15561 34506 15627 34509
rect 16430 34506 16436 34508
rect 15561 34504 16436 34506
rect 15561 34448 15566 34504
rect 15622 34448 16436 34504
rect 15561 34446 16436 34448
rect 15561 34443 15627 34446
rect 16430 34444 16436 34446
rect 16500 34444 16506 34508
rect 17125 34506 17191 34509
rect 19520 34506 20000 34536
rect 17125 34504 20000 34506
rect 17125 34448 17130 34504
rect 17186 34448 20000 34504
rect 17125 34446 20000 34448
rect 17125 34443 17191 34446
rect 19520 34416 20000 34446
rect 7610 34304 7930 34305
rect 7610 34240 7618 34304
rect 7682 34240 7698 34304
rect 7762 34240 7778 34304
rect 7842 34240 7858 34304
rect 7922 34240 7930 34304
rect 7610 34239 7930 34240
rect 14277 34304 14597 34305
rect 14277 34240 14285 34304
rect 14349 34240 14365 34304
rect 14429 34240 14445 34304
rect 14509 34240 14525 34304
rect 14589 34240 14597 34304
rect 14277 34239 14597 34240
rect 6729 34098 6795 34101
rect 9121 34098 9187 34101
rect 6729 34096 9187 34098
rect 6729 34040 6734 34096
rect 6790 34040 9126 34096
rect 9182 34040 9187 34096
rect 6729 34038 9187 34040
rect 6729 34035 6795 34038
rect 9121 34035 9187 34038
rect 10358 34036 10364 34100
rect 10428 34098 10434 34100
rect 11421 34098 11487 34101
rect 10428 34096 11487 34098
rect 10428 34040 11426 34096
rect 11482 34040 11487 34096
rect 10428 34038 11487 34040
rect 10428 34036 10434 34038
rect 11421 34035 11487 34038
rect 14825 34098 14891 34101
rect 15142 34098 15148 34100
rect 14825 34096 15148 34098
rect 14825 34040 14830 34096
rect 14886 34040 15148 34096
rect 14825 34038 15148 34040
rect 14825 34035 14891 34038
rect 15142 34036 15148 34038
rect 15212 34036 15218 34100
rect 4889 33962 4955 33965
rect 13629 33962 13695 33965
rect 4889 33960 13695 33962
rect 4889 33904 4894 33960
rect 4950 33904 13634 33960
rect 13690 33904 13695 33960
rect 4889 33902 13695 33904
rect 4889 33899 4955 33902
rect 13629 33899 13695 33902
rect 17125 33962 17191 33965
rect 17125 33960 18338 33962
rect 17125 33904 17130 33960
rect 17186 33904 18338 33960
rect 17125 33902 18338 33904
rect 17125 33899 17191 33902
rect 0 33826 480 33856
rect 1577 33826 1643 33829
rect 0 33824 1643 33826
rect 0 33768 1582 33824
rect 1638 33768 1643 33824
rect 0 33766 1643 33768
rect 0 33736 480 33766
rect 1577 33763 1643 33766
rect 6821 33826 6887 33829
rect 8293 33826 8359 33829
rect 6821 33824 8359 33826
rect 6821 33768 6826 33824
rect 6882 33768 8298 33824
rect 8354 33768 8359 33824
rect 6821 33766 8359 33768
rect 18278 33826 18338 33902
rect 19520 33826 20000 33856
rect 18278 33766 20000 33826
rect 6821 33763 6887 33766
rect 8293 33763 8359 33766
rect 4277 33760 4597 33761
rect 4277 33696 4285 33760
rect 4349 33696 4365 33760
rect 4429 33696 4445 33760
rect 4509 33696 4525 33760
rect 4589 33696 4597 33760
rect 4277 33695 4597 33696
rect 10944 33760 11264 33761
rect 10944 33696 10952 33760
rect 11016 33696 11032 33760
rect 11096 33696 11112 33760
rect 11176 33696 11192 33760
rect 11256 33696 11264 33760
rect 10944 33695 11264 33696
rect 17610 33760 17930 33761
rect 17610 33696 17618 33760
rect 17682 33696 17698 33760
rect 17762 33696 17778 33760
rect 17842 33696 17858 33760
rect 17922 33696 17930 33760
rect 19520 33736 20000 33766
rect 17610 33695 17930 33696
rect 6821 33692 6887 33693
rect 6821 33688 6868 33692
rect 6932 33690 6938 33692
rect 6821 33632 6826 33688
rect 6821 33628 6868 33632
rect 6932 33630 6978 33690
rect 6932 33628 6938 33630
rect 6821 33627 6887 33628
rect 1393 33554 1459 33557
rect 6177 33554 6243 33557
rect 1393 33552 6243 33554
rect 1393 33496 1398 33552
rect 1454 33496 6182 33552
rect 6238 33496 6243 33552
rect 1393 33494 6243 33496
rect 1393 33491 1459 33494
rect 6177 33491 6243 33494
rect 12801 33554 12867 33557
rect 15561 33554 15627 33557
rect 17033 33556 17099 33557
rect 12801 33552 15627 33554
rect 12801 33496 12806 33552
rect 12862 33496 15566 33552
rect 15622 33496 15627 33552
rect 12801 33494 15627 33496
rect 12801 33491 12867 33494
rect 15561 33491 15627 33494
rect 16982 33492 16988 33556
rect 17052 33554 17099 33556
rect 17052 33552 17144 33554
rect 17094 33496 17144 33552
rect 17052 33494 17144 33496
rect 17052 33492 17099 33494
rect 17033 33491 17099 33492
rect 5717 33418 5783 33421
rect 16614 33418 16620 33420
rect 5717 33416 16620 33418
rect 5717 33360 5722 33416
rect 5778 33360 16620 33416
rect 5717 33358 16620 33360
rect 5717 33355 5783 33358
rect 16614 33356 16620 33358
rect 16684 33356 16690 33420
rect 10501 33282 10567 33285
rect 12617 33282 12683 33285
rect 10501 33280 12683 33282
rect 10501 33224 10506 33280
rect 10562 33224 12622 33280
rect 12678 33224 12683 33280
rect 10501 33222 12683 33224
rect 10501 33219 10567 33222
rect 12617 33219 12683 33222
rect 7610 33216 7930 33217
rect 0 33146 480 33176
rect 7610 33152 7618 33216
rect 7682 33152 7698 33216
rect 7762 33152 7778 33216
rect 7842 33152 7858 33216
rect 7922 33152 7930 33216
rect 7610 33151 7930 33152
rect 14277 33216 14597 33217
rect 14277 33152 14285 33216
rect 14349 33152 14365 33216
rect 14429 33152 14445 33216
rect 14509 33152 14525 33216
rect 14589 33152 14597 33216
rect 14277 33151 14597 33152
rect 0 33086 1410 33146
rect 0 33056 480 33086
rect 1350 33010 1410 33086
rect 2630 33084 2636 33148
rect 2700 33146 2706 33148
rect 2865 33146 2931 33149
rect 2700 33144 2931 33146
rect 2700 33088 2870 33144
rect 2926 33088 2931 33144
rect 2700 33086 2931 33088
rect 2700 33084 2706 33086
rect 2865 33083 2931 33086
rect 6361 33146 6427 33149
rect 11513 33146 11579 33149
rect 11646 33146 11652 33148
rect 6361 33144 6746 33146
rect 6361 33088 6366 33144
rect 6422 33088 6746 33144
rect 6361 33086 6746 33088
rect 6361 33083 6427 33086
rect 3785 33010 3851 33013
rect 1350 33008 3851 33010
rect 1350 32952 3790 33008
rect 3846 32952 3851 33008
rect 1350 32950 3851 32952
rect 6686 33010 6746 33086
rect 11513 33144 11652 33146
rect 11513 33088 11518 33144
rect 11574 33088 11652 33144
rect 11513 33086 11652 33088
rect 11513 33083 11579 33086
rect 11646 33084 11652 33086
rect 11716 33084 11722 33148
rect 17125 33146 17191 33149
rect 19520 33146 20000 33176
rect 17125 33144 20000 33146
rect 17125 33088 17130 33144
rect 17186 33088 20000 33144
rect 17125 33086 20000 33088
rect 17125 33083 17191 33086
rect 19520 33056 20000 33086
rect 6821 33010 6887 33013
rect 6686 33008 6887 33010
rect 6686 32952 6826 33008
rect 6882 32952 6887 33008
rect 6686 32950 6887 32952
rect 3785 32947 3851 32950
rect 6821 32947 6887 32950
rect 9857 33010 9923 33013
rect 10225 33010 10291 33013
rect 17401 33012 17467 33013
rect 9857 33008 10291 33010
rect 9857 32952 9862 33008
rect 9918 32952 10230 33008
rect 10286 32952 10291 33008
rect 9857 32950 10291 32952
rect 9857 32947 9923 32950
rect 10225 32947 10291 32950
rect 17350 32948 17356 33012
rect 17420 33010 17467 33012
rect 17420 33008 17512 33010
rect 17462 32952 17512 33008
rect 17420 32950 17512 32952
rect 17420 32948 17467 32950
rect 17401 32947 17467 32948
rect 8150 32812 8156 32876
rect 8220 32874 8226 32876
rect 9305 32874 9371 32877
rect 8220 32872 9371 32874
rect 8220 32816 9310 32872
rect 9366 32816 9371 32872
rect 8220 32814 9371 32816
rect 8220 32812 8226 32814
rect 9305 32811 9371 32814
rect 10041 32874 10107 32877
rect 15101 32874 15167 32877
rect 10041 32872 15167 32874
rect 10041 32816 10046 32872
rect 10102 32816 15106 32872
rect 15162 32816 15167 32872
rect 10041 32814 15167 32816
rect 10041 32811 10107 32814
rect 15101 32811 15167 32814
rect 17125 32876 17191 32877
rect 17125 32872 17172 32876
rect 17236 32874 17242 32876
rect 17125 32816 17130 32872
rect 17125 32812 17172 32816
rect 17236 32814 17282 32874
rect 17236 32812 17242 32814
rect 17125 32811 17191 32812
rect 7373 32738 7439 32741
rect 8293 32738 8359 32741
rect 7373 32736 8359 32738
rect 7373 32680 7378 32736
rect 7434 32680 8298 32736
rect 8354 32680 8359 32736
rect 7373 32678 8359 32680
rect 7373 32675 7439 32678
rect 8293 32675 8359 32678
rect 4277 32672 4597 32673
rect 4277 32608 4285 32672
rect 4349 32608 4365 32672
rect 4429 32608 4445 32672
rect 4509 32608 4525 32672
rect 4589 32608 4597 32672
rect 4277 32607 4597 32608
rect 10944 32672 11264 32673
rect 10944 32608 10952 32672
rect 11016 32608 11032 32672
rect 11096 32608 11112 32672
rect 11176 32608 11192 32672
rect 11256 32608 11264 32672
rect 10944 32607 11264 32608
rect 17610 32672 17930 32673
rect 17610 32608 17618 32672
rect 17682 32608 17698 32672
rect 17762 32608 17778 32672
rect 17842 32608 17858 32672
rect 17922 32608 17930 32672
rect 17610 32607 17930 32608
rect 7414 32540 7420 32604
rect 7484 32602 7490 32604
rect 8017 32602 8083 32605
rect 7484 32600 8083 32602
rect 7484 32544 8022 32600
rect 8078 32544 8083 32600
rect 7484 32542 8083 32544
rect 7484 32540 7490 32542
rect 8017 32539 8083 32542
rect 17493 32466 17559 32469
rect 19520 32466 20000 32496
rect 17493 32464 20000 32466
rect 17493 32408 17498 32464
rect 17554 32408 20000 32464
rect 17493 32406 20000 32408
rect 17493 32403 17559 32406
rect 19520 32376 20000 32406
rect 0 32330 480 32360
rect 1853 32330 1919 32333
rect 0 32328 1919 32330
rect 0 32272 1858 32328
rect 1914 32272 1919 32328
rect 0 32270 1919 32272
rect 0 32240 480 32270
rect 1853 32267 1919 32270
rect 6821 32330 6887 32333
rect 10225 32330 10291 32333
rect 14958 32330 14964 32332
rect 6821 32328 10291 32330
rect 6821 32272 6826 32328
rect 6882 32272 10230 32328
rect 10286 32272 10291 32328
rect 6821 32270 10291 32272
rect 6821 32267 6887 32270
rect 10225 32267 10291 32270
rect 10688 32270 14964 32330
rect 10225 32194 10291 32197
rect 10688 32194 10748 32270
rect 14958 32268 14964 32270
rect 15028 32268 15034 32332
rect 10225 32192 10748 32194
rect 10225 32136 10230 32192
rect 10286 32136 10748 32192
rect 10225 32134 10748 32136
rect 10225 32131 10291 32134
rect 7610 32128 7930 32129
rect 7610 32064 7618 32128
rect 7682 32064 7698 32128
rect 7762 32064 7778 32128
rect 7842 32064 7858 32128
rect 7922 32064 7930 32128
rect 7610 32063 7930 32064
rect 14277 32128 14597 32129
rect 14277 32064 14285 32128
rect 14349 32064 14365 32128
rect 14429 32064 14445 32128
rect 14509 32064 14525 32128
rect 14589 32064 14597 32128
rect 14277 32063 14597 32064
rect 1577 32056 1643 32061
rect 1577 32000 1582 32056
rect 1638 32000 1643 32056
rect 1577 31995 1643 32000
rect 1580 31922 1640 31995
rect 1945 31922 2011 31925
rect 1580 31920 2011 31922
rect 1580 31864 1950 31920
rect 2006 31864 2011 31920
rect 1580 31862 2011 31864
rect 1945 31859 2011 31862
rect 5809 31922 5875 31925
rect 10685 31922 10751 31925
rect 5809 31920 10751 31922
rect 5809 31864 5814 31920
rect 5870 31864 10690 31920
rect 10746 31864 10751 31920
rect 5809 31862 10751 31864
rect 5809 31859 5875 31862
rect 10685 31859 10751 31862
rect 11973 31922 12039 31925
rect 13854 31922 13860 31924
rect 11973 31920 13860 31922
rect 11973 31864 11978 31920
rect 12034 31864 13860 31920
rect 11973 31862 13860 31864
rect 11973 31859 12039 31862
rect 13854 31860 13860 31862
rect 13924 31860 13930 31924
rect 1761 31786 1827 31789
rect 1718 31784 1827 31786
rect 1718 31728 1766 31784
rect 1822 31728 1827 31784
rect 1718 31723 1827 31728
rect 6361 31786 6427 31789
rect 6821 31786 6887 31789
rect 6361 31784 6887 31786
rect 6361 31728 6366 31784
rect 6422 31728 6826 31784
rect 6882 31728 6887 31784
rect 6361 31726 6887 31728
rect 6361 31723 6427 31726
rect 6821 31723 6887 31726
rect 7046 31724 7052 31788
rect 7116 31786 7122 31788
rect 8753 31786 8819 31789
rect 11329 31786 11395 31789
rect 7116 31784 11395 31786
rect 7116 31728 8758 31784
rect 8814 31728 11334 31784
rect 11390 31728 11395 31784
rect 7116 31726 11395 31728
rect 7116 31724 7122 31726
rect 8753 31723 8819 31726
rect 11329 31723 11395 31726
rect 11881 31786 11947 31789
rect 13169 31786 13235 31789
rect 11881 31784 13235 31786
rect 11881 31728 11886 31784
rect 11942 31728 13174 31784
rect 13230 31728 13235 31784
rect 11881 31726 13235 31728
rect 11881 31723 11947 31726
rect 13169 31723 13235 31726
rect 17769 31786 17835 31789
rect 19520 31786 20000 31816
rect 17769 31784 20000 31786
rect 17769 31728 17774 31784
rect 17830 31728 20000 31784
rect 17769 31726 20000 31728
rect 17769 31723 17835 31726
rect 0 31514 480 31544
rect 1718 31514 1778 31723
rect 19520 31696 20000 31726
rect 4277 31584 4597 31585
rect 4277 31520 4285 31584
rect 4349 31520 4365 31584
rect 4429 31520 4445 31584
rect 4509 31520 4525 31584
rect 4589 31520 4597 31584
rect 4277 31519 4597 31520
rect 10944 31584 11264 31585
rect 10944 31520 10952 31584
rect 11016 31520 11032 31584
rect 11096 31520 11112 31584
rect 11176 31520 11192 31584
rect 11256 31520 11264 31584
rect 10944 31519 11264 31520
rect 17610 31584 17930 31585
rect 17610 31520 17618 31584
rect 17682 31520 17698 31584
rect 17762 31520 17778 31584
rect 17842 31520 17858 31584
rect 17922 31520 17930 31584
rect 17610 31519 17930 31520
rect 0 31454 1778 31514
rect 0 31424 480 31454
rect 10777 31380 10843 31381
rect 10726 31316 10732 31380
rect 10796 31378 10843 31380
rect 10796 31376 10888 31378
rect 10838 31320 10888 31376
rect 10796 31318 10888 31320
rect 10796 31316 10843 31318
rect 10777 31315 10843 31316
rect 9489 31242 9555 31245
rect 11513 31242 11579 31245
rect 9489 31240 11579 31242
rect 9489 31184 9494 31240
rect 9550 31184 11518 31240
rect 11574 31184 11579 31240
rect 9489 31182 11579 31184
rect 9489 31179 9555 31182
rect 11513 31179 11579 31182
rect 13813 31242 13879 31245
rect 15285 31242 15351 31245
rect 13813 31240 15351 31242
rect 13813 31184 13818 31240
rect 13874 31184 15290 31240
rect 15346 31184 15351 31240
rect 13813 31182 15351 31184
rect 13813 31179 13879 31182
rect 15285 31179 15351 31182
rect 17769 31106 17835 31109
rect 19520 31106 20000 31136
rect 17769 31104 20000 31106
rect 17769 31048 17774 31104
rect 17830 31048 20000 31104
rect 17769 31046 20000 31048
rect 17769 31043 17835 31046
rect 7610 31040 7930 31041
rect 7610 30976 7618 31040
rect 7682 30976 7698 31040
rect 7762 30976 7778 31040
rect 7842 30976 7858 31040
rect 7922 30976 7930 31040
rect 7610 30975 7930 30976
rect 14277 31040 14597 31041
rect 14277 30976 14285 31040
rect 14349 30976 14365 31040
rect 14429 30976 14445 31040
rect 14509 30976 14525 31040
rect 14589 30976 14597 31040
rect 19520 31016 20000 31046
rect 14277 30975 14597 30976
rect 4061 30834 4127 30837
rect 10225 30834 10291 30837
rect 4061 30832 10291 30834
rect 4061 30776 4066 30832
rect 4122 30776 10230 30832
rect 10286 30776 10291 30832
rect 4061 30774 10291 30776
rect 4061 30771 4127 30774
rect 10225 30771 10291 30774
rect 10593 30834 10659 30837
rect 11329 30834 11395 30837
rect 10593 30832 11395 30834
rect 10593 30776 10598 30832
rect 10654 30776 11334 30832
rect 11390 30776 11395 30832
rect 10593 30774 11395 30776
rect 10593 30771 10659 30774
rect 11329 30771 11395 30774
rect 0 30698 480 30728
rect 1577 30698 1643 30701
rect 0 30696 1643 30698
rect 0 30640 1582 30696
rect 1638 30640 1643 30696
rect 0 30638 1643 30640
rect 0 30608 480 30638
rect 1577 30635 1643 30638
rect 3693 30698 3759 30701
rect 14038 30698 14044 30700
rect 3693 30696 14044 30698
rect 3693 30640 3698 30696
rect 3754 30640 14044 30696
rect 3693 30638 14044 30640
rect 3693 30635 3759 30638
rect 14038 30636 14044 30638
rect 14108 30636 14114 30700
rect 4981 30562 5047 30565
rect 7649 30562 7715 30565
rect 10685 30562 10751 30565
rect 4981 30560 10751 30562
rect 4981 30504 4986 30560
rect 5042 30504 7654 30560
rect 7710 30504 10690 30560
rect 10746 30504 10751 30560
rect 4981 30502 10751 30504
rect 4981 30499 5047 30502
rect 7649 30499 7715 30502
rect 10685 30499 10751 30502
rect 4277 30496 4597 30497
rect 4277 30432 4285 30496
rect 4349 30432 4365 30496
rect 4429 30432 4445 30496
rect 4509 30432 4525 30496
rect 4589 30432 4597 30496
rect 4277 30431 4597 30432
rect 10944 30496 11264 30497
rect 10944 30432 10952 30496
rect 11016 30432 11032 30496
rect 11096 30432 11112 30496
rect 11176 30432 11192 30496
rect 11256 30432 11264 30496
rect 10944 30431 11264 30432
rect 17610 30496 17930 30497
rect 17610 30432 17618 30496
rect 17682 30432 17698 30496
rect 17762 30432 17778 30496
rect 17842 30432 17858 30496
rect 17922 30432 17930 30496
rect 17610 30431 17930 30432
rect 19520 30426 20000 30456
rect 18094 30366 20000 30426
rect 10501 30290 10567 30293
rect 11881 30290 11947 30293
rect 10501 30288 11947 30290
rect 10501 30232 10506 30288
rect 10562 30232 11886 30288
rect 11942 30232 11947 30288
rect 10501 30230 11947 30232
rect 10501 30227 10567 30230
rect 11881 30227 11947 30230
rect 14181 30290 14247 30293
rect 14825 30290 14891 30293
rect 15837 30290 15903 30293
rect 14181 30288 15903 30290
rect 14181 30232 14186 30288
rect 14242 30232 14830 30288
rect 14886 30232 15842 30288
rect 15898 30232 15903 30288
rect 14181 30230 15903 30232
rect 14181 30227 14247 30230
rect 14825 30227 14891 30230
rect 15837 30227 15903 30230
rect 17861 30290 17927 30293
rect 18094 30290 18154 30366
rect 19520 30336 20000 30366
rect 17861 30288 18154 30290
rect 17861 30232 17866 30288
rect 17922 30232 18154 30288
rect 17861 30230 18154 30232
rect 17861 30227 17927 30230
rect 2129 30018 2195 30021
rect 4521 30018 4587 30021
rect 2129 30016 4587 30018
rect 2129 29960 2134 30016
rect 2190 29960 4526 30016
rect 4582 29960 4587 30016
rect 2129 29958 4587 29960
rect 2129 29955 2195 29958
rect 4521 29955 4587 29958
rect 7610 29952 7930 29953
rect 0 29882 480 29912
rect 7610 29888 7618 29952
rect 7682 29888 7698 29952
rect 7762 29888 7778 29952
rect 7842 29888 7858 29952
rect 7922 29888 7930 29952
rect 7610 29887 7930 29888
rect 14277 29952 14597 29953
rect 14277 29888 14285 29952
rect 14349 29888 14365 29952
rect 14429 29888 14445 29952
rect 14509 29888 14525 29952
rect 14589 29888 14597 29952
rect 14277 29887 14597 29888
rect 1669 29882 1735 29885
rect 0 29880 1735 29882
rect 0 29824 1674 29880
rect 1730 29824 1735 29880
rect 0 29822 1735 29824
rect 0 29792 480 29822
rect 1669 29819 1735 29822
rect 10961 29746 11027 29749
rect 12014 29746 12020 29748
rect 10961 29744 12020 29746
rect 10961 29688 10966 29744
rect 11022 29688 12020 29744
rect 10961 29686 12020 29688
rect 10961 29683 11027 29686
rect 12014 29684 12020 29686
rect 12084 29684 12090 29748
rect 17217 29746 17283 29749
rect 19520 29746 20000 29776
rect 17217 29744 20000 29746
rect 17217 29688 17222 29744
rect 17278 29688 20000 29744
rect 17217 29686 20000 29688
rect 17217 29683 17283 29686
rect 19520 29656 20000 29686
rect 4277 29408 4597 29409
rect 4277 29344 4285 29408
rect 4349 29344 4365 29408
rect 4429 29344 4445 29408
rect 4509 29344 4525 29408
rect 4589 29344 4597 29408
rect 4277 29343 4597 29344
rect 10944 29408 11264 29409
rect 10944 29344 10952 29408
rect 11016 29344 11032 29408
rect 11096 29344 11112 29408
rect 11176 29344 11192 29408
rect 11256 29344 11264 29408
rect 10944 29343 11264 29344
rect 17610 29408 17930 29409
rect 17610 29344 17618 29408
rect 17682 29344 17698 29408
rect 17762 29344 17778 29408
rect 17842 29344 17858 29408
rect 17922 29344 17930 29408
rect 17610 29343 17930 29344
rect 5441 29202 5507 29205
rect 7189 29202 7255 29205
rect 8334 29202 8340 29204
rect 5441 29200 8340 29202
rect 5441 29144 5446 29200
rect 5502 29144 7194 29200
rect 7250 29144 8340 29200
rect 5441 29142 8340 29144
rect 5441 29139 5507 29142
rect 7189 29139 7255 29142
rect 8334 29140 8340 29142
rect 8404 29140 8410 29204
rect 0 29066 480 29096
rect 2129 29066 2195 29069
rect 0 29064 2195 29066
rect 0 29008 2134 29064
rect 2190 29008 2195 29064
rect 0 29006 2195 29008
rect 0 28976 480 29006
rect 2129 29003 2195 29006
rect 8109 29066 8175 29069
rect 17769 29066 17835 29069
rect 19520 29066 20000 29096
rect 8109 29064 8218 29066
rect 8109 29008 8114 29064
rect 8170 29008 8218 29064
rect 8109 29003 8218 29008
rect 17769 29064 20000 29066
rect 17769 29008 17774 29064
rect 17830 29008 20000 29064
rect 17769 29006 20000 29008
rect 17769 29003 17835 29006
rect 7610 28864 7930 28865
rect 7610 28800 7618 28864
rect 7682 28800 7698 28864
rect 7762 28800 7778 28864
rect 7842 28800 7858 28864
rect 7922 28800 7930 28864
rect 7610 28799 7930 28800
rect 8158 28661 8218 29003
rect 19520 28976 20000 29006
rect 11513 28932 11579 28933
rect 11462 28930 11468 28932
rect 11422 28870 11468 28930
rect 11532 28928 11579 28932
rect 11574 28872 11579 28928
rect 11462 28868 11468 28870
rect 11532 28868 11579 28872
rect 11513 28867 11579 28868
rect 14277 28864 14597 28865
rect 14277 28800 14285 28864
rect 14349 28800 14365 28864
rect 14429 28800 14445 28864
rect 14509 28800 14525 28864
rect 14589 28800 14597 28864
rect 14277 28799 14597 28800
rect 8109 28656 8218 28661
rect 8109 28600 8114 28656
rect 8170 28600 8218 28656
rect 8109 28598 8218 28600
rect 8109 28595 8175 28598
rect 1945 28522 2011 28525
rect 12157 28522 12223 28525
rect 1945 28520 12223 28522
rect 1945 28464 1950 28520
rect 2006 28464 12162 28520
rect 12218 28464 12223 28520
rect 1945 28462 12223 28464
rect 1945 28459 2011 28462
rect 12157 28459 12223 28462
rect 19520 28386 20000 28416
rect 18646 28326 20000 28386
rect 4277 28320 4597 28321
rect 0 28250 480 28280
rect 4277 28256 4285 28320
rect 4349 28256 4365 28320
rect 4429 28256 4445 28320
rect 4509 28256 4525 28320
rect 4589 28256 4597 28320
rect 4277 28255 4597 28256
rect 10944 28320 11264 28321
rect 10944 28256 10952 28320
rect 11016 28256 11032 28320
rect 11096 28256 11112 28320
rect 11176 28256 11192 28320
rect 11256 28256 11264 28320
rect 10944 28255 11264 28256
rect 17610 28320 17930 28321
rect 17610 28256 17618 28320
rect 17682 28256 17698 28320
rect 17762 28256 17778 28320
rect 17842 28256 17858 28320
rect 17922 28256 17930 28320
rect 17610 28255 17930 28256
rect 1577 28250 1643 28253
rect 0 28248 1643 28250
rect 0 28192 1582 28248
rect 1638 28192 1643 28248
rect 0 28190 1643 28192
rect 0 28160 480 28190
rect 1577 28187 1643 28190
rect 1669 28114 1735 28117
rect 11973 28114 12039 28117
rect 1669 28112 12039 28114
rect 1669 28056 1674 28112
rect 1730 28056 11978 28112
rect 12034 28056 12039 28112
rect 1669 28054 12039 28056
rect 1669 28051 1735 28054
rect 11973 28051 12039 28054
rect 17769 28114 17835 28117
rect 18646 28114 18706 28326
rect 19520 28296 20000 28326
rect 17769 28112 18706 28114
rect 17769 28056 17774 28112
rect 17830 28056 18706 28112
rect 17769 28054 18706 28056
rect 17769 28051 17835 28054
rect 11513 27978 11579 27981
rect 16297 27978 16363 27981
rect 11513 27976 16363 27978
rect 11513 27920 11518 27976
rect 11574 27920 16302 27976
rect 16358 27920 16363 27976
rect 11513 27918 16363 27920
rect 11513 27915 11579 27918
rect 16297 27915 16363 27918
rect 7610 27776 7930 27777
rect 7610 27712 7618 27776
rect 7682 27712 7698 27776
rect 7762 27712 7778 27776
rect 7842 27712 7858 27776
rect 7922 27712 7930 27776
rect 7610 27711 7930 27712
rect 14277 27776 14597 27777
rect 14277 27712 14285 27776
rect 14349 27712 14365 27776
rect 14429 27712 14445 27776
rect 14509 27712 14525 27776
rect 14589 27712 14597 27776
rect 14277 27711 14597 27712
rect 17493 27706 17559 27709
rect 19520 27706 20000 27736
rect 17493 27704 20000 27706
rect 17493 27648 17498 27704
rect 17554 27648 20000 27704
rect 17493 27646 20000 27648
rect 17493 27643 17559 27646
rect 19520 27616 20000 27646
rect 0 27434 480 27464
rect 4061 27434 4127 27437
rect 0 27432 4127 27434
rect 0 27376 4066 27432
rect 4122 27376 4127 27432
rect 0 27374 4127 27376
rect 0 27344 480 27374
rect 4061 27371 4127 27374
rect 4277 27232 4597 27233
rect 4277 27168 4285 27232
rect 4349 27168 4365 27232
rect 4429 27168 4445 27232
rect 4509 27168 4525 27232
rect 4589 27168 4597 27232
rect 4277 27167 4597 27168
rect 10944 27232 11264 27233
rect 10944 27168 10952 27232
rect 11016 27168 11032 27232
rect 11096 27168 11112 27232
rect 11176 27168 11192 27232
rect 11256 27168 11264 27232
rect 10944 27167 11264 27168
rect 17610 27232 17930 27233
rect 17610 27168 17618 27232
rect 17682 27168 17698 27232
rect 17762 27168 17778 27232
rect 17842 27168 17858 27232
rect 17922 27168 17930 27232
rect 17610 27167 17930 27168
rect 10501 27026 10567 27029
rect 13537 27026 13603 27029
rect 10501 27024 13603 27026
rect 10501 26968 10506 27024
rect 10562 26968 13542 27024
rect 13598 26968 13603 27024
rect 10501 26966 13603 26968
rect 10501 26963 10567 26966
rect 13537 26963 13603 26966
rect 17585 27026 17651 27029
rect 19520 27026 20000 27056
rect 17585 27024 20000 27026
rect 17585 26968 17590 27024
rect 17646 26968 20000 27024
rect 17585 26966 20000 26968
rect 17585 26963 17651 26966
rect 19520 26936 20000 26966
rect 0 26754 480 26784
rect 1577 26754 1643 26757
rect 0 26752 1643 26754
rect 0 26696 1582 26752
rect 1638 26696 1643 26752
rect 0 26694 1643 26696
rect 0 26664 480 26694
rect 1577 26691 1643 26694
rect 7610 26688 7930 26689
rect 7610 26624 7618 26688
rect 7682 26624 7698 26688
rect 7762 26624 7778 26688
rect 7842 26624 7858 26688
rect 7922 26624 7930 26688
rect 7610 26623 7930 26624
rect 14277 26688 14597 26689
rect 14277 26624 14285 26688
rect 14349 26624 14365 26688
rect 14429 26624 14445 26688
rect 14509 26624 14525 26688
rect 14589 26624 14597 26688
rect 14277 26623 14597 26624
rect 5165 26618 5231 26621
rect 5390 26618 5396 26620
rect 5165 26616 5396 26618
rect 5165 26560 5170 26616
rect 5226 26560 5396 26616
rect 5165 26558 5396 26560
rect 5165 26555 5231 26558
rect 5390 26556 5396 26558
rect 5460 26556 5466 26620
rect 9305 26482 9371 26485
rect 9622 26482 9628 26484
rect 9305 26480 9628 26482
rect 9305 26424 9310 26480
rect 9366 26424 9628 26480
rect 9305 26422 9628 26424
rect 9305 26419 9371 26422
rect 9622 26420 9628 26422
rect 9692 26420 9698 26484
rect 3417 26346 3483 26349
rect 11145 26346 11211 26349
rect 3417 26344 11211 26346
rect 3417 26288 3422 26344
rect 3478 26288 11150 26344
rect 11206 26288 11211 26344
rect 3417 26286 11211 26288
rect 3417 26283 3483 26286
rect 11145 26283 11211 26286
rect 19520 26210 20000 26240
rect 18094 26150 20000 26210
rect 4277 26144 4597 26145
rect 4277 26080 4285 26144
rect 4349 26080 4365 26144
rect 4429 26080 4445 26144
rect 4509 26080 4525 26144
rect 4589 26080 4597 26144
rect 4277 26079 4597 26080
rect 10944 26144 11264 26145
rect 10944 26080 10952 26144
rect 11016 26080 11032 26144
rect 11096 26080 11112 26144
rect 11176 26080 11192 26144
rect 11256 26080 11264 26144
rect 10944 26079 11264 26080
rect 17610 26144 17930 26145
rect 17610 26080 17618 26144
rect 17682 26080 17698 26144
rect 17762 26080 17778 26144
rect 17842 26080 17858 26144
rect 17922 26080 17930 26144
rect 17610 26079 17930 26080
rect 0 25938 480 25968
rect 2773 25938 2839 25941
rect 0 25936 2839 25938
rect 0 25880 2778 25936
rect 2834 25880 2839 25936
rect 0 25878 2839 25880
rect 0 25848 480 25878
rect 2773 25875 2839 25878
rect 15561 25938 15627 25941
rect 17033 25938 17099 25941
rect 15561 25936 17099 25938
rect 15561 25880 15566 25936
rect 15622 25880 17038 25936
rect 17094 25880 17099 25936
rect 15561 25878 17099 25880
rect 15561 25875 15627 25878
rect 17033 25875 17099 25878
rect 17585 25938 17651 25941
rect 18094 25938 18154 26150
rect 19520 26120 20000 26150
rect 17585 25936 18154 25938
rect 17585 25880 17590 25936
rect 17646 25880 18154 25936
rect 17585 25878 18154 25880
rect 17585 25875 17651 25878
rect 3233 25802 3299 25805
rect 12065 25802 12131 25805
rect 3233 25800 12131 25802
rect 3233 25744 3238 25800
rect 3294 25744 12070 25800
rect 12126 25744 12131 25800
rect 3233 25742 12131 25744
rect 3233 25739 3299 25742
rect 12065 25739 12131 25742
rect 9489 25666 9555 25669
rect 12157 25666 12223 25669
rect 9489 25664 12223 25666
rect 9489 25608 9494 25664
rect 9550 25608 12162 25664
rect 12218 25608 12223 25664
rect 9489 25606 12223 25608
rect 9489 25603 9555 25606
rect 12157 25603 12223 25606
rect 7610 25600 7930 25601
rect 7610 25536 7618 25600
rect 7682 25536 7698 25600
rect 7762 25536 7778 25600
rect 7842 25536 7858 25600
rect 7922 25536 7930 25600
rect 7610 25535 7930 25536
rect 14277 25600 14597 25601
rect 14277 25536 14285 25600
rect 14349 25536 14365 25600
rect 14429 25536 14445 25600
rect 14509 25536 14525 25600
rect 14589 25536 14597 25600
rect 14277 25535 14597 25536
rect 16389 25530 16455 25533
rect 19520 25530 20000 25560
rect 16389 25528 20000 25530
rect 16389 25472 16394 25528
rect 16450 25472 20000 25528
rect 16389 25470 20000 25472
rect 16389 25467 16455 25470
rect 19520 25440 20000 25470
rect 3141 25258 3207 25261
rect 4153 25258 4219 25261
rect 9029 25258 9095 25261
rect 11973 25258 12039 25261
rect 3141 25256 12039 25258
rect 3141 25200 3146 25256
rect 3202 25200 4158 25256
rect 4214 25200 9034 25256
rect 9090 25200 11978 25256
rect 12034 25200 12039 25256
rect 3141 25198 12039 25200
rect 3141 25195 3207 25198
rect 4153 25195 4219 25198
rect 9029 25195 9095 25198
rect 11973 25195 12039 25198
rect 0 25122 480 25152
rect 0 25062 1824 25122
rect 0 25032 480 25062
rect 1764 24853 1824 25062
rect 4277 25056 4597 25057
rect 4277 24992 4285 25056
rect 4349 24992 4365 25056
rect 4429 24992 4445 25056
rect 4509 24992 4525 25056
rect 4589 24992 4597 25056
rect 4277 24991 4597 24992
rect 10944 25056 11264 25057
rect 10944 24992 10952 25056
rect 11016 24992 11032 25056
rect 11096 24992 11112 25056
rect 11176 24992 11192 25056
rect 11256 24992 11264 25056
rect 10944 24991 11264 24992
rect 17610 25056 17930 25057
rect 17610 24992 17618 25056
rect 17682 24992 17698 25056
rect 17762 24992 17778 25056
rect 17842 24992 17858 25056
rect 17922 24992 17930 25056
rect 17610 24991 17930 24992
rect 11421 24986 11487 24989
rect 13445 24986 13511 24989
rect 15653 24986 15719 24989
rect 11421 24984 15719 24986
rect 11421 24928 11426 24984
rect 11482 24928 13450 24984
rect 13506 24928 15658 24984
rect 15714 24928 15719 24984
rect 11421 24926 15719 24928
rect 11421 24923 11487 24926
rect 13445 24923 13511 24926
rect 15653 24923 15719 24926
rect 16113 24986 16179 24989
rect 16665 24986 16731 24989
rect 16113 24984 16731 24986
rect 16113 24928 16118 24984
rect 16174 24928 16670 24984
rect 16726 24928 16731 24984
rect 16113 24926 16731 24928
rect 16113 24923 16179 24926
rect 16665 24923 16731 24926
rect 1761 24848 1827 24853
rect 1761 24792 1766 24848
rect 1822 24792 1827 24848
rect 1761 24787 1827 24792
rect 13997 24850 14063 24853
rect 15653 24850 15719 24853
rect 13997 24848 15719 24850
rect 13997 24792 14002 24848
rect 14058 24792 15658 24848
rect 15714 24792 15719 24848
rect 13997 24790 15719 24792
rect 13997 24787 14063 24790
rect 15653 24787 15719 24790
rect 17585 24850 17651 24853
rect 19520 24850 20000 24880
rect 17585 24848 20000 24850
rect 17585 24792 17590 24848
rect 17646 24792 20000 24848
rect 17585 24790 20000 24792
rect 17585 24787 17651 24790
rect 19520 24760 20000 24790
rect 7610 24512 7930 24513
rect 7610 24448 7618 24512
rect 7682 24448 7698 24512
rect 7762 24448 7778 24512
rect 7842 24448 7858 24512
rect 7922 24448 7930 24512
rect 7610 24447 7930 24448
rect 14277 24512 14597 24513
rect 14277 24448 14285 24512
rect 14349 24448 14365 24512
rect 14429 24448 14445 24512
rect 14509 24448 14525 24512
rect 14589 24448 14597 24512
rect 14277 24447 14597 24448
rect 5165 24442 5231 24445
rect 7005 24442 7071 24445
rect 5165 24440 7071 24442
rect 5165 24384 5170 24440
rect 5226 24384 7010 24440
rect 7066 24384 7071 24440
rect 5165 24382 7071 24384
rect 5165 24379 5231 24382
rect 7005 24379 7071 24382
rect 0 24306 480 24336
rect 2129 24306 2195 24309
rect 0 24304 2195 24306
rect 0 24248 2134 24304
rect 2190 24248 2195 24304
rect 0 24246 2195 24248
rect 0 24216 480 24246
rect 2129 24243 2195 24246
rect 10041 24306 10107 24309
rect 10542 24306 10548 24308
rect 10041 24304 10548 24306
rect 10041 24248 10046 24304
rect 10102 24248 10548 24304
rect 10041 24246 10548 24248
rect 10041 24243 10107 24246
rect 10542 24244 10548 24246
rect 10612 24244 10618 24308
rect 16389 24170 16455 24173
rect 19520 24170 20000 24200
rect 16389 24168 20000 24170
rect 16389 24112 16394 24168
rect 16450 24112 20000 24168
rect 16389 24110 20000 24112
rect 16389 24107 16455 24110
rect 19520 24080 20000 24110
rect 6637 24034 6703 24037
rect 7465 24034 7531 24037
rect 9765 24034 9831 24037
rect 6637 24032 9831 24034
rect 6637 23976 6642 24032
rect 6698 23976 7470 24032
rect 7526 23976 9770 24032
rect 9826 23976 9831 24032
rect 6637 23974 9831 23976
rect 6637 23971 6703 23974
rect 7465 23971 7531 23974
rect 9765 23971 9831 23974
rect 4277 23968 4597 23969
rect 4277 23904 4285 23968
rect 4349 23904 4365 23968
rect 4429 23904 4445 23968
rect 4509 23904 4525 23968
rect 4589 23904 4597 23968
rect 4277 23903 4597 23904
rect 10944 23968 11264 23969
rect 10944 23904 10952 23968
rect 11016 23904 11032 23968
rect 11096 23904 11112 23968
rect 11176 23904 11192 23968
rect 11256 23904 11264 23968
rect 10944 23903 11264 23904
rect 17610 23968 17930 23969
rect 17610 23904 17618 23968
rect 17682 23904 17698 23968
rect 17762 23904 17778 23968
rect 17842 23904 17858 23968
rect 17922 23904 17930 23968
rect 17610 23903 17930 23904
rect 11973 23762 12039 23765
rect 14641 23762 14707 23765
rect 11973 23760 14707 23762
rect 11973 23704 11978 23760
rect 12034 23704 14646 23760
rect 14702 23704 14707 23760
rect 11973 23702 14707 23704
rect 11973 23699 12039 23702
rect 14641 23699 14707 23702
rect 12893 23626 12959 23629
rect 15009 23626 15075 23629
rect 12893 23624 15075 23626
rect 12893 23568 12898 23624
rect 12954 23568 15014 23624
rect 15070 23568 15075 23624
rect 12893 23566 15075 23568
rect 12893 23563 12959 23566
rect 15009 23563 15075 23566
rect 0 23490 480 23520
rect 3325 23490 3391 23493
rect 0 23488 3391 23490
rect 0 23432 3330 23488
rect 3386 23432 3391 23488
rect 0 23430 3391 23432
rect 0 23400 480 23430
rect 3325 23427 3391 23430
rect 5073 23490 5139 23493
rect 5901 23490 5967 23493
rect 5073 23488 5967 23490
rect 5073 23432 5078 23488
rect 5134 23432 5906 23488
rect 5962 23432 5967 23488
rect 5073 23430 5967 23432
rect 5073 23427 5139 23430
rect 5901 23427 5967 23430
rect 17125 23490 17191 23493
rect 19520 23490 20000 23520
rect 17125 23488 20000 23490
rect 17125 23432 17130 23488
rect 17186 23432 20000 23488
rect 17125 23430 20000 23432
rect 17125 23427 17191 23430
rect 7610 23424 7930 23425
rect 7610 23360 7618 23424
rect 7682 23360 7698 23424
rect 7762 23360 7778 23424
rect 7842 23360 7858 23424
rect 7922 23360 7930 23424
rect 7610 23359 7930 23360
rect 14277 23424 14597 23425
rect 14277 23360 14285 23424
rect 14349 23360 14365 23424
rect 14429 23360 14445 23424
rect 14509 23360 14525 23424
rect 14589 23360 14597 23424
rect 19520 23400 20000 23430
rect 14277 23359 14597 23360
rect 4061 23218 4127 23221
rect 12893 23218 12959 23221
rect 4061 23216 12959 23218
rect 4061 23160 4066 23216
rect 4122 23160 12898 23216
rect 12954 23160 12959 23216
rect 4061 23158 12959 23160
rect 4061 23155 4127 23158
rect 12893 23155 12959 23158
rect 3141 23082 3207 23085
rect 13261 23082 13327 23085
rect 3141 23080 13327 23082
rect 3141 23024 3146 23080
rect 3202 23024 13266 23080
rect 13322 23024 13327 23080
rect 3141 23022 13327 23024
rect 3141 23019 3207 23022
rect 13261 23019 13327 23022
rect 4705 22946 4771 22949
rect 5165 22946 5231 22949
rect 10225 22946 10291 22949
rect 4705 22944 10291 22946
rect 4705 22888 4710 22944
rect 4766 22888 5170 22944
rect 5226 22888 10230 22944
rect 10286 22888 10291 22944
rect 4705 22886 10291 22888
rect 4705 22883 4771 22886
rect 5165 22883 5231 22886
rect 10225 22883 10291 22886
rect 4277 22880 4597 22881
rect 4277 22816 4285 22880
rect 4349 22816 4365 22880
rect 4429 22816 4445 22880
rect 4509 22816 4525 22880
rect 4589 22816 4597 22880
rect 4277 22815 4597 22816
rect 10944 22880 11264 22881
rect 10944 22816 10952 22880
rect 11016 22816 11032 22880
rect 11096 22816 11112 22880
rect 11176 22816 11192 22880
rect 11256 22816 11264 22880
rect 10944 22815 11264 22816
rect 17610 22880 17930 22881
rect 17610 22816 17618 22880
rect 17682 22816 17698 22880
rect 17762 22816 17778 22880
rect 17842 22816 17858 22880
rect 17922 22816 17930 22880
rect 17610 22815 17930 22816
rect 13813 22810 13879 22813
rect 16113 22810 16179 22813
rect 19520 22810 20000 22840
rect 13813 22808 16179 22810
rect 13813 22752 13818 22808
rect 13874 22752 16118 22808
rect 16174 22752 16179 22808
rect 13813 22750 16179 22752
rect 13813 22747 13879 22750
rect 16113 22747 16179 22750
rect 18094 22750 20000 22810
rect 0 22674 480 22704
rect 1669 22674 1735 22677
rect 11421 22676 11487 22677
rect 11421 22674 11468 22676
rect 0 22672 1735 22674
rect 0 22616 1674 22672
rect 1730 22616 1735 22672
rect 0 22614 1735 22616
rect 11376 22672 11468 22674
rect 11376 22616 11426 22672
rect 11376 22614 11468 22616
rect 0 22584 480 22614
rect 1669 22611 1735 22614
rect 11421 22612 11468 22614
rect 11532 22612 11538 22676
rect 16021 22674 16087 22677
rect 18094 22674 18154 22750
rect 19520 22720 20000 22750
rect 16021 22672 18154 22674
rect 16021 22616 16026 22672
rect 16082 22616 18154 22672
rect 16021 22614 18154 22616
rect 11421 22611 11487 22612
rect 16021 22611 16087 22614
rect 13629 22538 13695 22541
rect 15193 22538 15259 22541
rect 13629 22536 15259 22538
rect 13629 22480 13634 22536
rect 13690 22480 15198 22536
rect 15254 22480 15259 22536
rect 13629 22478 15259 22480
rect 13629 22475 13695 22478
rect 15193 22475 15259 22478
rect 7610 22336 7930 22337
rect 7610 22272 7618 22336
rect 7682 22272 7698 22336
rect 7762 22272 7778 22336
rect 7842 22272 7858 22336
rect 7922 22272 7930 22336
rect 7610 22271 7930 22272
rect 14277 22336 14597 22337
rect 14277 22272 14285 22336
rect 14349 22272 14365 22336
rect 14429 22272 14445 22336
rect 14509 22272 14525 22336
rect 14589 22272 14597 22336
rect 14277 22271 14597 22272
rect 8109 22266 8175 22269
rect 9857 22266 9923 22269
rect 8109 22264 9923 22266
rect 8109 22208 8114 22264
rect 8170 22208 9862 22264
rect 9918 22208 9923 22264
rect 8109 22206 9923 22208
rect 8109 22203 8175 22206
rect 9857 22203 9923 22206
rect 9673 22130 9739 22133
rect 10501 22130 10567 22133
rect 9673 22128 10567 22130
rect 9673 22072 9678 22128
rect 9734 22072 10506 22128
rect 10562 22072 10567 22128
rect 9673 22070 10567 22072
rect 9673 22067 9739 22070
rect 10501 22067 10567 22070
rect 14365 22130 14431 22133
rect 19520 22130 20000 22160
rect 14365 22128 20000 22130
rect 14365 22072 14370 22128
rect 14426 22072 20000 22128
rect 14365 22070 20000 22072
rect 14365 22067 14431 22070
rect 19520 22040 20000 22070
rect 0 21858 480 21888
rect 1485 21858 1551 21861
rect 0 21856 1551 21858
rect 0 21800 1490 21856
rect 1546 21800 1551 21856
rect 0 21798 1551 21800
rect 0 21768 480 21798
rect 1485 21795 1551 21798
rect 4277 21792 4597 21793
rect 4277 21728 4285 21792
rect 4349 21728 4365 21792
rect 4429 21728 4445 21792
rect 4509 21728 4525 21792
rect 4589 21728 4597 21792
rect 4277 21727 4597 21728
rect 10944 21792 11264 21793
rect 10944 21728 10952 21792
rect 11016 21728 11032 21792
rect 11096 21728 11112 21792
rect 11176 21728 11192 21792
rect 11256 21728 11264 21792
rect 10944 21727 11264 21728
rect 17610 21792 17930 21793
rect 17610 21728 17618 21792
rect 17682 21728 17698 21792
rect 17762 21728 17778 21792
rect 17842 21728 17858 21792
rect 17922 21728 17930 21792
rect 17610 21727 17930 21728
rect 3417 21586 3483 21589
rect 12525 21586 12591 21589
rect 3417 21584 12591 21586
rect 3417 21528 3422 21584
rect 3478 21528 12530 21584
rect 12586 21528 12591 21584
rect 3417 21526 12591 21528
rect 3417 21523 3483 21526
rect 12525 21523 12591 21526
rect 15193 21450 15259 21453
rect 19520 21450 20000 21480
rect 15193 21448 20000 21450
rect 15193 21392 15198 21448
rect 15254 21392 20000 21448
rect 15193 21390 20000 21392
rect 15193 21387 15259 21390
rect 19520 21360 20000 21390
rect 15101 21314 15167 21317
rect 15929 21314 15995 21317
rect 16573 21314 16639 21317
rect 15101 21312 16639 21314
rect 15101 21256 15106 21312
rect 15162 21256 15934 21312
rect 15990 21256 16578 21312
rect 16634 21256 16639 21312
rect 15101 21254 16639 21256
rect 15101 21251 15167 21254
rect 15929 21251 15995 21254
rect 16573 21251 16639 21254
rect 7610 21248 7930 21249
rect 7610 21184 7618 21248
rect 7682 21184 7698 21248
rect 7762 21184 7778 21248
rect 7842 21184 7858 21248
rect 7922 21184 7930 21248
rect 7610 21183 7930 21184
rect 14277 21248 14597 21249
rect 14277 21184 14285 21248
rect 14349 21184 14365 21248
rect 14429 21184 14445 21248
rect 14509 21184 14525 21248
rect 14589 21184 14597 21248
rect 14277 21183 14597 21184
rect 0 21042 480 21072
rect 3417 21042 3483 21045
rect 0 21040 3483 21042
rect 0 20984 3422 21040
rect 3478 20984 3483 21040
rect 0 20982 3483 20984
rect 0 20952 480 20982
rect 3417 20979 3483 20982
rect 15469 20906 15535 20909
rect 15469 20904 18154 20906
rect 15469 20848 15474 20904
rect 15530 20848 18154 20904
rect 15469 20846 18154 20848
rect 15469 20843 15535 20846
rect 18094 20770 18154 20846
rect 19520 20770 20000 20800
rect 18094 20710 20000 20770
rect 4277 20704 4597 20705
rect 4277 20640 4285 20704
rect 4349 20640 4365 20704
rect 4429 20640 4445 20704
rect 4509 20640 4525 20704
rect 4589 20640 4597 20704
rect 4277 20639 4597 20640
rect 10944 20704 11264 20705
rect 10944 20640 10952 20704
rect 11016 20640 11032 20704
rect 11096 20640 11112 20704
rect 11176 20640 11192 20704
rect 11256 20640 11264 20704
rect 10944 20639 11264 20640
rect 17610 20704 17930 20705
rect 17610 20640 17618 20704
rect 17682 20640 17698 20704
rect 17762 20640 17778 20704
rect 17842 20640 17858 20704
rect 17922 20640 17930 20704
rect 19520 20680 20000 20710
rect 17610 20639 17930 20640
rect 3325 20498 3391 20501
rect 9397 20498 9463 20501
rect 3325 20496 9463 20498
rect 3325 20440 3330 20496
rect 3386 20440 9402 20496
rect 9458 20440 9463 20496
rect 3325 20438 9463 20440
rect 3325 20435 3391 20438
rect 9397 20435 9463 20438
rect 0 20362 480 20392
rect 3509 20362 3575 20365
rect 0 20360 3575 20362
rect 0 20304 3514 20360
rect 3570 20304 3575 20360
rect 0 20302 3575 20304
rect 0 20272 480 20302
rect 3509 20299 3575 20302
rect 7610 20160 7930 20161
rect 7610 20096 7618 20160
rect 7682 20096 7698 20160
rect 7762 20096 7778 20160
rect 7842 20096 7858 20160
rect 7922 20096 7930 20160
rect 7610 20095 7930 20096
rect 14277 20160 14597 20161
rect 14277 20096 14285 20160
rect 14349 20096 14365 20160
rect 14429 20096 14445 20160
rect 14509 20096 14525 20160
rect 14589 20096 14597 20160
rect 14277 20095 14597 20096
rect 15377 20090 15443 20093
rect 19520 20090 20000 20120
rect 15377 20088 20000 20090
rect 15377 20032 15382 20088
rect 15438 20032 20000 20088
rect 15377 20030 20000 20032
rect 15377 20027 15443 20030
rect 19520 20000 20000 20030
rect 13813 19954 13879 19957
rect 15929 19954 15995 19957
rect 13813 19952 15995 19954
rect 13813 19896 13818 19952
rect 13874 19896 15934 19952
rect 15990 19896 15995 19952
rect 13813 19894 15995 19896
rect 13813 19891 13879 19894
rect 15929 19891 15995 19894
rect 2957 19818 3023 19821
rect 14733 19818 14799 19821
rect 2957 19816 14799 19818
rect 2957 19760 2962 19816
rect 3018 19760 14738 19816
rect 14794 19760 14799 19816
rect 2957 19758 14799 19760
rect 2957 19755 3023 19758
rect 14733 19755 14799 19758
rect 4277 19616 4597 19617
rect 0 19546 480 19576
rect 4277 19552 4285 19616
rect 4349 19552 4365 19616
rect 4429 19552 4445 19616
rect 4509 19552 4525 19616
rect 4589 19552 4597 19616
rect 4277 19551 4597 19552
rect 10944 19616 11264 19617
rect 10944 19552 10952 19616
rect 11016 19552 11032 19616
rect 11096 19552 11112 19616
rect 11176 19552 11192 19616
rect 11256 19552 11264 19616
rect 10944 19551 11264 19552
rect 17610 19616 17930 19617
rect 17610 19552 17618 19616
rect 17682 19552 17698 19616
rect 17762 19552 17778 19616
rect 17842 19552 17858 19616
rect 17922 19552 17930 19616
rect 17610 19551 17930 19552
rect 1761 19546 1827 19549
rect 0 19544 1827 19546
rect 0 19488 1766 19544
rect 1822 19488 1827 19544
rect 0 19486 1827 19488
rect 0 19456 480 19486
rect 1761 19483 1827 19486
rect 8477 19546 8543 19549
rect 9765 19546 9831 19549
rect 8477 19544 9831 19546
rect 8477 19488 8482 19544
rect 8538 19488 9770 19544
rect 9826 19488 9831 19544
rect 8477 19486 9831 19488
rect 8477 19483 8543 19486
rect 9765 19483 9831 19486
rect 4705 19410 4771 19413
rect 12157 19410 12223 19413
rect 4705 19408 12223 19410
rect 4705 19352 4710 19408
rect 4766 19352 12162 19408
rect 12218 19352 12223 19408
rect 4705 19350 12223 19352
rect 4705 19347 4771 19350
rect 12157 19347 12223 19350
rect 12617 19410 12683 19413
rect 19520 19410 20000 19440
rect 12617 19408 20000 19410
rect 12617 19352 12622 19408
rect 12678 19352 20000 19408
rect 12617 19350 20000 19352
rect 12617 19347 12683 19350
rect 19520 19320 20000 19350
rect 4061 19274 4127 19277
rect 14181 19274 14247 19277
rect 4061 19272 14247 19274
rect 4061 19216 4066 19272
rect 4122 19216 14186 19272
rect 14242 19216 14247 19272
rect 4061 19214 14247 19216
rect 4061 19211 4127 19214
rect 14181 19211 14247 19214
rect 11789 19138 11855 19141
rect 13537 19138 13603 19141
rect 11789 19136 13603 19138
rect 11789 19080 11794 19136
rect 11850 19080 13542 19136
rect 13598 19080 13603 19136
rect 11789 19078 13603 19080
rect 11789 19075 11855 19078
rect 13537 19075 13603 19078
rect 7610 19072 7930 19073
rect 7610 19008 7618 19072
rect 7682 19008 7698 19072
rect 7762 19008 7778 19072
rect 7842 19008 7858 19072
rect 7922 19008 7930 19072
rect 7610 19007 7930 19008
rect 14277 19072 14597 19073
rect 14277 19008 14285 19072
rect 14349 19008 14365 19072
rect 14429 19008 14445 19072
rect 14509 19008 14525 19072
rect 14589 19008 14597 19072
rect 14277 19007 14597 19008
rect 3785 18866 3851 18869
rect 10777 18866 10843 18869
rect 11237 18866 11303 18869
rect 3785 18864 11303 18866
rect 3785 18808 3790 18864
rect 3846 18808 10782 18864
rect 10838 18808 11242 18864
rect 11298 18808 11303 18864
rect 3785 18806 11303 18808
rect 3785 18803 3851 18806
rect 10777 18803 10843 18806
rect 11237 18803 11303 18806
rect 0 18730 480 18760
rect 1393 18730 1459 18733
rect 0 18728 1459 18730
rect 0 18672 1398 18728
rect 1454 18672 1459 18728
rect 0 18670 1459 18672
rect 0 18640 480 18670
rect 1393 18667 1459 18670
rect 15193 18730 15259 18733
rect 19520 18730 20000 18760
rect 15193 18728 20000 18730
rect 15193 18672 15198 18728
rect 15254 18672 20000 18728
rect 15193 18670 20000 18672
rect 15193 18667 15259 18670
rect 19520 18640 20000 18670
rect 4277 18528 4597 18529
rect 4277 18464 4285 18528
rect 4349 18464 4365 18528
rect 4429 18464 4445 18528
rect 4509 18464 4525 18528
rect 4589 18464 4597 18528
rect 4277 18463 4597 18464
rect 10944 18528 11264 18529
rect 10944 18464 10952 18528
rect 11016 18464 11032 18528
rect 11096 18464 11112 18528
rect 11176 18464 11192 18528
rect 11256 18464 11264 18528
rect 10944 18463 11264 18464
rect 17610 18528 17930 18529
rect 17610 18464 17618 18528
rect 17682 18464 17698 18528
rect 17762 18464 17778 18528
rect 17842 18464 17858 18528
rect 17922 18464 17930 18528
rect 17610 18463 17930 18464
rect 12065 18458 12131 18461
rect 14641 18458 14707 18461
rect 15009 18458 15075 18461
rect 16849 18458 16915 18461
rect 12065 18456 16915 18458
rect 12065 18400 12070 18456
rect 12126 18400 14646 18456
rect 14702 18400 15014 18456
rect 15070 18400 16854 18456
rect 16910 18400 16915 18456
rect 12065 18398 16915 18400
rect 12065 18395 12131 18398
rect 14641 18395 14707 18398
rect 15009 18395 15075 18398
rect 16849 18395 16915 18398
rect 13629 18322 13695 18325
rect 15193 18322 15259 18325
rect 13629 18320 15259 18322
rect 13629 18264 13634 18320
rect 13690 18264 15198 18320
rect 15254 18264 15259 18320
rect 13629 18262 15259 18264
rect 13629 18259 13695 18262
rect 15193 18259 15259 18262
rect 15101 18050 15167 18053
rect 19520 18050 20000 18080
rect 15101 18048 20000 18050
rect 15101 17992 15106 18048
rect 15162 17992 20000 18048
rect 15101 17990 20000 17992
rect 15101 17987 15167 17990
rect 7610 17984 7930 17985
rect 0 17914 480 17944
rect 7610 17920 7618 17984
rect 7682 17920 7698 17984
rect 7762 17920 7778 17984
rect 7842 17920 7858 17984
rect 7922 17920 7930 17984
rect 7610 17919 7930 17920
rect 14277 17984 14597 17985
rect 14277 17920 14285 17984
rect 14349 17920 14365 17984
rect 14429 17920 14445 17984
rect 14509 17920 14525 17984
rect 14589 17920 14597 17984
rect 19520 17960 20000 17990
rect 14277 17919 14597 17920
rect 3785 17914 3851 17917
rect 0 17912 3851 17914
rect 0 17856 3790 17912
rect 3846 17856 3851 17912
rect 0 17854 3851 17856
rect 0 17824 480 17854
rect 3785 17851 3851 17854
rect 3509 17778 3575 17781
rect 9397 17778 9463 17781
rect 3509 17776 9463 17778
rect 3509 17720 3514 17776
rect 3570 17720 9402 17776
rect 9458 17720 9463 17776
rect 3509 17718 9463 17720
rect 3509 17715 3575 17718
rect 9397 17715 9463 17718
rect 3141 17642 3207 17645
rect 11789 17642 11855 17645
rect 3141 17640 11855 17642
rect 3141 17584 3146 17640
rect 3202 17584 11794 17640
rect 11850 17584 11855 17640
rect 3141 17582 11855 17584
rect 3141 17579 3207 17582
rect 11789 17579 11855 17582
rect 15193 17642 15259 17645
rect 15193 17640 18154 17642
rect 15193 17584 15198 17640
rect 15254 17584 18154 17640
rect 15193 17582 18154 17584
rect 15193 17579 15259 17582
rect 4277 17440 4597 17441
rect 4277 17376 4285 17440
rect 4349 17376 4365 17440
rect 4429 17376 4445 17440
rect 4509 17376 4525 17440
rect 4589 17376 4597 17440
rect 4277 17375 4597 17376
rect 10944 17440 11264 17441
rect 10944 17376 10952 17440
rect 11016 17376 11032 17440
rect 11096 17376 11112 17440
rect 11176 17376 11192 17440
rect 11256 17376 11264 17440
rect 10944 17375 11264 17376
rect 17610 17440 17930 17441
rect 17610 17376 17618 17440
rect 17682 17376 17698 17440
rect 17762 17376 17778 17440
rect 17842 17376 17858 17440
rect 17922 17376 17930 17440
rect 17610 17375 17930 17376
rect 18094 17370 18154 17582
rect 19520 17370 20000 17400
rect 18094 17310 20000 17370
rect 19520 17280 20000 17310
rect 1669 17236 1735 17237
rect 1669 17234 1716 17236
rect 1624 17232 1716 17234
rect 1624 17176 1674 17232
rect 1624 17174 1716 17176
rect 1669 17172 1716 17174
rect 1780 17172 1786 17236
rect 1669 17171 1735 17172
rect 0 17098 480 17128
rect 2773 17098 2839 17101
rect 0 17096 2839 17098
rect 0 17040 2778 17096
rect 2834 17040 2839 17096
rect 0 17038 2839 17040
rect 0 17008 480 17038
rect 2773 17035 2839 17038
rect 8017 16962 8083 16965
rect 9765 16962 9831 16965
rect 8017 16960 9831 16962
rect 8017 16904 8022 16960
rect 8078 16904 9770 16960
rect 9826 16904 9831 16960
rect 8017 16902 9831 16904
rect 8017 16899 8083 16902
rect 9765 16899 9831 16902
rect 7610 16896 7930 16897
rect 7610 16832 7618 16896
rect 7682 16832 7698 16896
rect 7762 16832 7778 16896
rect 7842 16832 7858 16896
rect 7922 16832 7930 16896
rect 7610 16831 7930 16832
rect 14277 16896 14597 16897
rect 14277 16832 14285 16896
rect 14349 16832 14365 16896
rect 14429 16832 14445 16896
rect 14509 16832 14525 16896
rect 14589 16832 14597 16896
rect 14277 16831 14597 16832
rect 6913 16690 6979 16693
rect 9673 16690 9739 16693
rect 6913 16688 9739 16690
rect 6913 16632 6918 16688
rect 6974 16632 9678 16688
rect 9734 16632 9739 16688
rect 6913 16630 9739 16632
rect 6913 16627 6979 16630
rect 9673 16627 9739 16630
rect 11329 16690 11395 16693
rect 19520 16690 20000 16720
rect 11329 16688 20000 16690
rect 11329 16632 11334 16688
rect 11390 16632 20000 16688
rect 11329 16630 20000 16632
rect 11329 16627 11395 16630
rect 19520 16600 20000 16630
rect 4277 16352 4597 16353
rect 0 16282 480 16312
rect 4277 16288 4285 16352
rect 4349 16288 4365 16352
rect 4429 16288 4445 16352
rect 4509 16288 4525 16352
rect 4589 16288 4597 16352
rect 4277 16287 4597 16288
rect 10944 16352 11264 16353
rect 10944 16288 10952 16352
rect 11016 16288 11032 16352
rect 11096 16288 11112 16352
rect 11176 16288 11192 16352
rect 11256 16288 11264 16352
rect 10944 16287 11264 16288
rect 17610 16352 17930 16353
rect 17610 16288 17618 16352
rect 17682 16288 17698 16352
rect 17762 16288 17778 16352
rect 17842 16288 17858 16352
rect 17922 16288 17930 16352
rect 17610 16287 17930 16288
rect 2589 16282 2655 16285
rect 0 16280 2655 16282
rect 0 16224 2594 16280
rect 2650 16224 2655 16280
rect 0 16222 2655 16224
rect 0 16192 480 16222
rect 2589 16219 2655 16222
rect 5901 16146 5967 16149
rect 12525 16146 12591 16149
rect 5901 16144 12591 16146
rect 5901 16088 5906 16144
rect 5962 16088 12530 16144
rect 12586 16088 12591 16144
rect 5901 16086 12591 16088
rect 5901 16083 5967 16086
rect 12525 16083 12591 16086
rect 3141 16010 3207 16013
rect 15561 16010 15627 16013
rect 19520 16010 20000 16040
rect 3141 16008 15394 16010
rect 3141 15952 3146 16008
rect 3202 15952 15394 16008
rect 3141 15950 15394 15952
rect 3141 15947 3207 15950
rect 15334 15874 15394 15950
rect 15561 16008 20000 16010
rect 15561 15952 15566 16008
rect 15622 15952 20000 16008
rect 15561 15950 20000 15952
rect 15561 15947 15627 15950
rect 19520 15920 20000 15950
rect 16941 15874 17007 15877
rect 15334 15872 17007 15874
rect 15334 15816 16946 15872
rect 17002 15816 17007 15872
rect 15334 15814 17007 15816
rect 16941 15811 17007 15814
rect 7610 15808 7930 15809
rect 7610 15744 7618 15808
rect 7682 15744 7698 15808
rect 7762 15744 7778 15808
rect 7842 15744 7858 15808
rect 7922 15744 7930 15808
rect 7610 15743 7930 15744
rect 14277 15808 14597 15809
rect 14277 15744 14285 15808
rect 14349 15744 14365 15808
rect 14429 15744 14445 15808
rect 14509 15744 14525 15808
rect 14589 15744 14597 15808
rect 14277 15743 14597 15744
rect 0 15466 480 15496
rect 1209 15466 1275 15469
rect 0 15464 1275 15466
rect 0 15408 1214 15464
rect 1270 15408 1275 15464
rect 0 15406 1275 15408
rect 0 15376 480 15406
rect 1209 15403 1275 15406
rect 16389 15466 16455 15469
rect 16389 15464 18154 15466
rect 16389 15408 16394 15464
rect 16450 15408 18154 15464
rect 16389 15406 18154 15408
rect 16389 15403 16455 15406
rect 14273 15330 14339 15333
rect 16021 15330 16087 15333
rect 14273 15328 16087 15330
rect 14273 15272 14278 15328
rect 14334 15272 16026 15328
rect 16082 15272 16087 15328
rect 14273 15270 16087 15272
rect 18094 15330 18154 15406
rect 19520 15330 20000 15360
rect 18094 15270 20000 15330
rect 14273 15267 14339 15270
rect 16021 15267 16087 15270
rect 4277 15264 4597 15265
rect 4277 15200 4285 15264
rect 4349 15200 4365 15264
rect 4429 15200 4445 15264
rect 4509 15200 4525 15264
rect 4589 15200 4597 15264
rect 4277 15199 4597 15200
rect 10944 15264 11264 15265
rect 10944 15200 10952 15264
rect 11016 15200 11032 15264
rect 11096 15200 11112 15264
rect 11176 15200 11192 15264
rect 11256 15200 11264 15264
rect 10944 15199 11264 15200
rect 17610 15264 17930 15265
rect 17610 15200 17618 15264
rect 17682 15200 17698 15264
rect 17762 15200 17778 15264
rect 17842 15200 17858 15264
rect 17922 15200 17930 15264
rect 19520 15240 20000 15270
rect 17610 15199 17930 15200
rect 5073 14922 5139 14925
rect 15377 14922 15443 14925
rect 5073 14920 15443 14922
rect 5073 14864 5078 14920
rect 5134 14864 15382 14920
rect 15438 14864 15443 14920
rect 5073 14862 15443 14864
rect 5073 14859 5139 14862
rect 15377 14859 15443 14862
rect 7610 14720 7930 14721
rect 0 14650 480 14680
rect 7610 14656 7618 14720
rect 7682 14656 7698 14720
rect 7762 14656 7778 14720
rect 7842 14656 7858 14720
rect 7922 14656 7930 14720
rect 7610 14655 7930 14656
rect 14277 14720 14597 14721
rect 14277 14656 14285 14720
rect 14349 14656 14365 14720
rect 14429 14656 14445 14720
rect 14509 14656 14525 14720
rect 14589 14656 14597 14720
rect 14277 14655 14597 14656
rect 3233 14650 3299 14653
rect 0 14648 3299 14650
rect 0 14592 3238 14648
rect 3294 14592 3299 14648
rect 0 14590 3299 14592
rect 0 14560 480 14590
rect 3233 14587 3299 14590
rect 16205 14650 16271 14653
rect 19520 14650 20000 14680
rect 16205 14648 20000 14650
rect 16205 14592 16210 14648
rect 16266 14592 20000 14648
rect 16205 14590 20000 14592
rect 16205 14587 16271 14590
rect 19520 14560 20000 14590
rect 7281 14514 7347 14517
rect 9857 14514 9923 14517
rect 7281 14512 9923 14514
rect 7281 14456 7286 14512
rect 7342 14456 9862 14512
rect 9918 14456 9923 14512
rect 7281 14454 9923 14456
rect 7281 14451 7347 14454
rect 9857 14451 9923 14454
rect 3969 14378 4035 14381
rect 16849 14378 16915 14381
rect 3969 14376 16915 14378
rect 3969 14320 3974 14376
rect 4030 14320 16854 14376
rect 16910 14320 16915 14376
rect 3969 14318 16915 14320
rect 3969 14315 4035 14318
rect 16849 14315 16915 14318
rect 4277 14176 4597 14177
rect 4277 14112 4285 14176
rect 4349 14112 4365 14176
rect 4429 14112 4445 14176
rect 4509 14112 4525 14176
rect 4589 14112 4597 14176
rect 4277 14111 4597 14112
rect 10944 14176 11264 14177
rect 10944 14112 10952 14176
rect 11016 14112 11032 14176
rect 11096 14112 11112 14176
rect 11176 14112 11192 14176
rect 11256 14112 11264 14176
rect 10944 14111 11264 14112
rect 17610 14176 17930 14177
rect 17610 14112 17618 14176
rect 17682 14112 17698 14176
rect 17762 14112 17778 14176
rect 17842 14112 17858 14176
rect 17922 14112 17930 14176
rect 17610 14111 17930 14112
rect 8293 13970 8359 13973
rect 13813 13970 13879 13973
rect 8293 13968 13879 13970
rect 8293 13912 8298 13968
rect 8354 13912 13818 13968
rect 13874 13912 13879 13968
rect 8293 13910 13879 13912
rect 8293 13907 8359 13910
rect 13813 13907 13879 13910
rect 15561 13970 15627 13973
rect 19520 13970 20000 14000
rect 15561 13968 20000 13970
rect 15561 13912 15566 13968
rect 15622 13912 20000 13968
rect 15561 13910 20000 13912
rect 15561 13907 15627 13910
rect 19520 13880 20000 13910
rect 0 13834 480 13864
rect 3785 13834 3851 13837
rect 0 13832 3851 13834
rect 0 13776 3790 13832
rect 3846 13776 3851 13832
rect 0 13774 3851 13776
rect 0 13744 480 13774
rect 3785 13771 3851 13774
rect 12341 13834 12407 13837
rect 15193 13834 15259 13837
rect 12341 13832 15259 13834
rect 12341 13776 12346 13832
rect 12402 13776 15198 13832
rect 15254 13776 15259 13832
rect 12341 13774 15259 13776
rect 12341 13771 12407 13774
rect 15193 13771 15259 13774
rect 7610 13632 7930 13633
rect 7610 13568 7618 13632
rect 7682 13568 7698 13632
rect 7762 13568 7778 13632
rect 7842 13568 7858 13632
rect 7922 13568 7930 13632
rect 7610 13567 7930 13568
rect 14277 13632 14597 13633
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 13567 14597 13568
rect 9489 13426 9555 13429
rect 15653 13426 15719 13429
rect 9489 13424 15719 13426
rect 9489 13368 9494 13424
rect 9550 13368 15658 13424
rect 15714 13368 15719 13424
rect 9489 13366 15719 13368
rect 9489 13363 9555 13366
rect 15653 13363 15719 13366
rect 4613 13290 4679 13293
rect 10317 13290 10383 13293
rect 4613 13288 10383 13290
rect 4613 13232 4618 13288
rect 4674 13232 10322 13288
rect 10378 13232 10383 13288
rect 4613 13230 10383 13232
rect 4613 13227 4679 13230
rect 10317 13227 10383 13230
rect 16757 13290 16823 13293
rect 19520 13290 20000 13320
rect 16757 13288 20000 13290
rect 16757 13232 16762 13288
rect 16818 13232 20000 13288
rect 16757 13230 20000 13232
rect 16757 13227 16823 13230
rect 19520 13200 20000 13230
rect 0 13154 480 13184
rect 1577 13154 1643 13157
rect 0 13152 1643 13154
rect 0 13096 1582 13152
rect 1638 13096 1643 13152
rect 0 13094 1643 13096
rect 0 13064 480 13094
rect 1577 13091 1643 13094
rect 5625 13154 5691 13157
rect 9765 13154 9831 13157
rect 5625 13152 9831 13154
rect 5625 13096 5630 13152
rect 5686 13096 9770 13152
rect 9826 13096 9831 13152
rect 5625 13094 9831 13096
rect 5625 13091 5691 13094
rect 9765 13091 9831 13094
rect 4277 13088 4597 13089
rect 4277 13024 4285 13088
rect 4349 13024 4365 13088
rect 4429 13024 4445 13088
rect 4509 13024 4525 13088
rect 4589 13024 4597 13088
rect 4277 13023 4597 13024
rect 10944 13088 11264 13089
rect 10944 13024 10952 13088
rect 11016 13024 11032 13088
rect 11096 13024 11112 13088
rect 11176 13024 11192 13088
rect 11256 13024 11264 13088
rect 10944 13023 11264 13024
rect 17610 13088 17930 13089
rect 17610 13024 17618 13088
rect 17682 13024 17698 13088
rect 17762 13024 17778 13088
rect 17842 13024 17858 13088
rect 17922 13024 17930 13088
rect 17610 13023 17930 13024
rect 9489 13018 9555 13021
rect 10225 13018 10291 13021
rect 9489 13016 10291 13018
rect 9489 12960 9494 13016
rect 9550 12960 10230 13016
rect 10286 12960 10291 13016
rect 9489 12958 10291 12960
rect 9489 12955 9555 12958
rect 10225 12955 10291 12958
rect 3049 12882 3115 12885
rect 16113 12882 16179 12885
rect 3049 12880 16179 12882
rect 3049 12824 3054 12880
rect 3110 12824 16118 12880
rect 16174 12824 16179 12880
rect 3049 12822 16179 12824
rect 3049 12819 3115 12822
rect 16113 12819 16179 12822
rect 2957 12746 3023 12749
rect 8293 12746 8359 12749
rect 2957 12744 8359 12746
rect 2957 12688 2962 12744
rect 3018 12688 8298 12744
rect 8354 12688 8359 12744
rect 2957 12686 8359 12688
rect 2957 12683 3023 12686
rect 8293 12683 8359 12686
rect 13721 12746 13787 12749
rect 13721 12744 15210 12746
rect 13721 12688 13726 12744
rect 13782 12688 15210 12744
rect 13721 12686 15210 12688
rect 13721 12683 13787 12686
rect 7610 12544 7930 12545
rect 7610 12480 7618 12544
rect 7682 12480 7698 12544
rect 7762 12480 7778 12544
rect 7842 12480 7858 12544
rect 7922 12480 7930 12544
rect 7610 12479 7930 12480
rect 14277 12544 14597 12545
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 12479 14597 12480
rect 0 12338 480 12368
rect 3785 12338 3851 12341
rect 0 12336 3851 12338
rect 0 12280 3790 12336
rect 3846 12280 3851 12336
rect 0 12278 3851 12280
rect 0 12248 480 12278
rect 3785 12275 3851 12278
rect 12249 12338 12315 12341
rect 14181 12338 14247 12341
rect 12249 12336 14247 12338
rect 12249 12280 12254 12336
rect 12310 12280 14186 12336
rect 14242 12280 14247 12336
rect 12249 12278 14247 12280
rect 12249 12275 12315 12278
rect 14181 12275 14247 12278
rect 15150 12202 15210 12686
rect 16389 12610 16455 12613
rect 19520 12610 20000 12640
rect 16389 12608 20000 12610
rect 16389 12552 16394 12608
rect 16450 12552 20000 12608
rect 16389 12550 20000 12552
rect 16389 12547 16455 12550
rect 19520 12520 20000 12550
rect 15150 12142 18154 12202
rect 4277 12000 4597 12001
rect 4277 11936 4285 12000
rect 4349 11936 4365 12000
rect 4429 11936 4445 12000
rect 4509 11936 4525 12000
rect 4589 11936 4597 12000
rect 4277 11935 4597 11936
rect 10944 12000 11264 12001
rect 10944 11936 10952 12000
rect 11016 11936 11032 12000
rect 11096 11936 11112 12000
rect 11176 11936 11192 12000
rect 11256 11936 11264 12000
rect 10944 11935 11264 11936
rect 17610 12000 17930 12001
rect 17610 11936 17618 12000
rect 17682 11936 17698 12000
rect 17762 11936 17778 12000
rect 17842 11936 17858 12000
rect 17922 11936 17930 12000
rect 17610 11935 17930 11936
rect 14181 11930 14247 11933
rect 16757 11930 16823 11933
rect 13494 11928 16823 11930
rect 13494 11872 14186 11928
rect 14242 11872 16762 11928
rect 16818 11872 16823 11928
rect 13494 11870 16823 11872
rect 18094 11930 18154 12142
rect 19520 11930 20000 11960
rect 18094 11870 20000 11930
rect 5809 11794 5875 11797
rect 13494 11794 13554 11870
rect 14181 11867 14247 11870
rect 16757 11867 16823 11870
rect 19520 11840 20000 11870
rect 5809 11792 13554 11794
rect 5809 11736 5814 11792
rect 5870 11736 13554 11792
rect 5809 11734 13554 11736
rect 13629 11794 13695 11797
rect 15377 11794 15443 11797
rect 13629 11792 15443 11794
rect 13629 11736 13634 11792
rect 13690 11736 15382 11792
rect 15438 11736 15443 11792
rect 13629 11734 15443 11736
rect 5809 11731 5875 11734
rect 13629 11731 13695 11734
rect 15377 11731 15443 11734
rect 9581 11658 9647 11661
rect 614 11656 9647 11658
rect 614 11600 9586 11656
rect 9642 11600 9647 11656
rect 614 11598 9647 11600
rect 0 11522 480 11552
rect 614 11522 674 11598
rect 9581 11595 9647 11598
rect 12249 11658 12315 11661
rect 14273 11658 14339 11661
rect 12249 11656 14339 11658
rect 12249 11600 12254 11656
rect 12310 11600 14278 11656
rect 14334 11600 14339 11656
rect 12249 11598 14339 11600
rect 12249 11595 12315 11598
rect 14273 11595 14339 11598
rect 0 11462 674 11522
rect 0 11432 480 11462
rect 7610 11456 7930 11457
rect 7610 11392 7618 11456
rect 7682 11392 7698 11456
rect 7762 11392 7778 11456
rect 7842 11392 7858 11456
rect 7922 11392 7930 11456
rect 7610 11391 7930 11392
rect 14277 11456 14597 11457
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 11391 14597 11392
rect 8109 11386 8175 11389
rect 11053 11386 11119 11389
rect 8109 11384 11119 11386
rect 8109 11328 8114 11384
rect 8170 11328 11058 11384
rect 11114 11328 11119 11384
rect 8109 11326 11119 11328
rect 8109 11323 8175 11326
rect 11053 11323 11119 11326
rect 15193 11250 15259 11253
rect 19520 11250 20000 11280
rect 15193 11248 20000 11250
rect 15193 11192 15198 11248
rect 15254 11192 20000 11248
rect 15193 11190 20000 11192
rect 15193 11187 15259 11190
rect 19520 11160 20000 11190
rect 3969 11114 4035 11117
rect 7465 11114 7531 11117
rect 3969 11112 7531 11114
rect 3969 11056 3974 11112
rect 4030 11056 7470 11112
rect 7526 11056 7531 11112
rect 3969 11054 7531 11056
rect 3969 11051 4035 11054
rect 7465 11051 7531 11054
rect 4277 10912 4597 10913
rect 4277 10848 4285 10912
rect 4349 10848 4365 10912
rect 4429 10848 4445 10912
rect 4509 10848 4525 10912
rect 4589 10848 4597 10912
rect 4277 10847 4597 10848
rect 10944 10912 11264 10913
rect 10944 10848 10952 10912
rect 11016 10848 11032 10912
rect 11096 10848 11112 10912
rect 11176 10848 11192 10912
rect 11256 10848 11264 10912
rect 10944 10847 11264 10848
rect 17610 10912 17930 10913
rect 17610 10848 17618 10912
rect 17682 10848 17698 10912
rect 17762 10848 17778 10912
rect 17842 10848 17858 10912
rect 17922 10848 17930 10912
rect 17610 10847 17930 10848
rect 0 10706 480 10736
rect 8753 10706 8819 10709
rect 11605 10706 11671 10709
rect 11789 10706 11855 10709
rect 0 10646 674 10706
rect 0 10616 480 10646
rect 614 10570 674 10646
rect 8753 10704 11855 10706
rect 8753 10648 8758 10704
rect 8814 10648 11610 10704
rect 11666 10648 11794 10704
rect 11850 10648 11855 10704
rect 8753 10646 11855 10648
rect 8753 10643 8819 10646
rect 11605 10643 11671 10646
rect 11789 10643 11855 10646
rect 9397 10570 9463 10573
rect 614 10568 9463 10570
rect 614 10512 9402 10568
rect 9458 10512 9463 10568
rect 614 10510 9463 10512
rect 9397 10507 9463 10510
rect 12249 10570 12315 10573
rect 13813 10570 13879 10573
rect 12249 10568 13879 10570
rect 12249 10512 12254 10568
rect 12310 10512 13818 10568
rect 13874 10512 13879 10568
rect 12249 10510 13879 10512
rect 12249 10507 12315 10510
rect 13813 10507 13879 10510
rect 15009 10570 15075 10573
rect 19520 10570 20000 10600
rect 15009 10568 20000 10570
rect 15009 10512 15014 10568
rect 15070 10512 20000 10568
rect 15009 10510 20000 10512
rect 15009 10507 15075 10510
rect 19520 10480 20000 10510
rect 8477 10434 8543 10437
rect 10777 10434 10843 10437
rect 12985 10434 13051 10437
rect 8477 10432 13051 10434
rect 8477 10376 8482 10432
rect 8538 10376 10782 10432
rect 10838 10376 12990 10432
rect 13046 10376 13051 10432
rect 8477 10374 13051 10376
rect 8477 10371 8543 10374
rect 10777 10371 10843 10374
rect 12985 10371 13051 10374
rect 7610 10368 7930 10369
rect 7610 10304 7618 10368
rect 7682 10304 7698 10368
rect 7762 10304 7778 10368
rect 7842 10304 7858 10368
rect 7922 10304 7930 10368
rect 7610 10303 7930 10304
rect 14277 10368 14597 10369
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 10303 14597 10304
rect 8109 10298 8175 10301
rect 10133 10298 10199 10301
rect 8109 10296 10199 10298
rect 8109 10240 8114 10296
rect 8170 10240 10138 10296
rect 10194 10240 10199 10296
rect 8109 10238 10199 10240
rect 8109 10235 8175 10238
rect 10133 10235 10199 10238
rect 3141 10162 3207 10165
rect 17309 10162 17375 10165
rect 3141 10160 17375 10162
rect 3141 10104 3146 10160
rect 3202 10104 17314 10160
rect 17370 10104 17375 10160
rect 3141 10102 17375 10104
rect 3141 10099 3207 10102
rect 17309 10099 17375 10102
rect 15377 10026 15443 10029
rect 15377 10024 18154 10026
rect 15377 9968 15382 10024
rect 15438 9968 18154 10024
rect 15377 9966 18154 9968
rect 15377 9963 15443 9966
rect 0 9890 480 9920
rect 3969 9890 4035 9893
rect 0 9888 4035 9890
rect 0 9832 3974 9888
rect 4030 9832 4035 9888
rect 0 9830 4035 9832
rect 18094 9890 18154 9966
rect 19520 9890 20000 9920
rect 18094 9830 20000 9890
rect 0 9800 480 9830
rect 3969 9827 4035 9830
rect 4277 9824 4597 9825
rect 4277 9760 4285 9824
rect 4349 9760 4365 9824
rect 4429 9760 4445 9824
rect 4509 9760 4525 9824
rect 4589 9760 4597 9824
rect 4277 9759 4597 9760
rect 10944 9824 11264 9825
rect 10944 9760 10952 9824
rect 11016 9760 11032 9824
rect 11096 9760 11112 9824
rect 11176 9760 11192 9824
rect 11256 9760 11264 9824
rect 10944 9759 11264 9760
rect 17610 9824 17930 9825
rect 17610 9760 17618 9824
rect 17682 9760 17698 9824
rect 17762 9760 17778 9824
rect 17842 9760 17858 9824
rect 17922 9760 17930 9824
rect 19520 9800 20000 9830
rect 17610 9759 17930 9760
rect 11145 9618 11211 9621
rect 13997 9618 14063 9621
rect 15193 9618 15259 9621
rect 11145 9616 15259 9618
rect 11145 9560 11150 9616
rect 11206 9560 14002 9616
rect 14058 9560 15198 9616
rect 15254 9560 15259 9616
rect 11145 9558 15259 9560
rect 11145 9555 11211 9558
rect 13997 9555 14063 9558
rect 15193 9555 15259 9558
rect 7833 9482 7899 9485
rect 13169 9482 13235 9485
rect 14181 9482 14247 9485
rect 7833 9480 14247 9482
rect 7833 9424 7838 9480
rect 7894 9424 13174 9480
rect 13230 9424 14186 9480
rect 14242 9424 14247 9480
rect 7833 9422 14247 9424
rect 7833 9419 7899 9422
rect 13169 9419 13235 9422
rect 14181 9419 14247 9422
rect 8569 9346 8635 9349
rect 11513 9346 11579 9349
rect 8569 9344 11579 9346
rect 8569 9288 8574 9344
rect 8630 9288 11518 9344
rect 11574 9288 11579 9344
rect 8569 9286 11579 9288
rect 8569 9283 8635 9286
rect 11513 9283 11579 9286
rect 11697 9346 11763 9349
rect 12433 9346 12499 9349
rect 11697 9344 12499 9346
rect 11697 9288 11702 9344
rect 11758 9288 12438 9344
rect 12494 9288 12499 9344
rect 11697 9286 12499 9288
rect 11697 9283 11763 9286
rect 12433 9283 12499 9286
rect 7610 9280 7930 9281
rect 7610 9216 7618 9280
rect 7682 9216 7698 9280
rect 7762 9216 7778 9280
rect 7842 9216 7858 9280
rect 7922 9216 7930 9280
rect 7610 9215 7930 9216
rect 14277 9280 14597 9281
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 9215 14597 9216
rect 15561 9210 15627 9213
rect 19520 9210 20000 9240
rect 15561 9208 20000 9210
rect 15561 9152 15566 9208
rect 15622 9152 20000 9208
rect 15561 9150 20000 9152
rect 15561 9147 15627 9150
rect 19520 9120 20000 9150
rect 0 9074 480 9104
rect 9765 9074 9831 9077
rect 0 9072 9831 9074
rect 0 9016 9770 9072
rect 9826 9016 9831 9072
rect 0 9014 9831 9016
rect 0 8984 480 9014
rect 9765 9011 9831 9014
rect 10593 8938 10659 8941
rect 12985 8938 13051 8941
rect 10593 8936 13051 8938
rect 10593 8880 10598 8936
rect 10654 8880 12990 8936
rect 13046 8880 13051 8936
rect 10593 8878 13051 8880
rect 10593 8875 10659 8878
rect 12985 8875 13051 8878
rect 4277 8736 4597 8737
rect 4277 8672 4285 8736
rect 4349 8672 4365 8736
rect 4429 8672 4445 8736
rect 4509 8672 4525 8736
rect 4589 8672 4597 8736
rect 4277 8671 4597 8672
rect 10944 8736 11264 8737
rect 10944 8672 10952 8736
rect 11016 8672 11032 8736
rect 11096 8672 11112 8736
rect 11176 8672 11192 8736
rect 11256 8672 11264 8736
rect 10944 8671 11264 8672
rect 17610 8736 17930 8737
rect 17610 8672 17618 8736
rect 17682 8672 17698 8736
rect 17762 8672 17778 8736
rect 17842 8672 17858 8736
rect 17922 8672 17930 8736
rect 17610 8671 17930 8672
rect 10501 8530 10567 8533
rect 11973 8530 12039 8533
rect 19520 8530 20000 8560
rect 10501 8528 12039 8530
rect 10501 8472 10506 8528
rect 10562 8472 11978 8528
rect 12034 8472 12039 8528
rect 10501 8470 12039 8472
rect 10501 8467 10567 8470
rect 11973 8467 12039 8470
rect 15886 8470 20000 8530
rect 10869 8394 10935 8397
rect 14181 8394 14247 8397
rect 15653 8394 15719 8397
rect 10869 8392 15719 8394
rect 10869 8336 10874 8392
rect 10930 8336 14186 8392
rect 14242 8336 15658 8392
rect 15714 8336 15719 8392
rect 10869 8334 15719 8336
rect 10869 8331 10935 8334
rect 14181 8331 14247 8334
rect 15653 8331 15719 8334
rect 0 8258 480 8288
rect 0 8198 7482 8258
rect 0 8168 480 8198
rect 7422 7986 7482 8198
rect 7610 8192 7930 8193
rect 7610 8128 7618 8192
rect 7682 8128 7698 8192
rect 7762 8128 7778 8192
rect 7842 8128 7858 8192
rect 7922 8128 7930 8192
rect 7610 8127 7930 8128
rect 14277 8192 14597 8193
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 8127 14597 8128
rect 10133 7986 10199 7989
rect 7422 7984 10199 7986
rect 7422 7928 10138 7984
rect 10194 7928 10199 7984
rect 7422 7926 10199 7928
rect 10133 7923 10199 7926
rect 11605 7986 11671 7989
rect 15886 7986 15946 8470
rect 19520 8440 20000 8470
rect 11605 7984 15946 7986
rect 11605 7928 11610 7984
rect 11666 7928 15946 7984
rect 11605 7926 15946 7928
rect 11605 7923 11671 7926
rect 8937 7850 9003 7853
rect 11881 7850 11947 7853
rect 15653 7850 15719 7853
rect 8937 7848 15719 7850
rect 8937 7792 8942 7848
rect 8998 7792 11886 7848
rect 11942 7792 15658 7848
rect 15714 7792 15719 7848
rect 8937 7790 15719 7792
rect 8937 7787 9003 7790
rect 11881 7787 11947 7790
rect 15653 7787 15719 7790
rect 16021 7850 16087 7853
rect 19520 7850 20000 7880
rect 16021 7848 20000 7850
rect 16021 7792 16026 7848
rect 16082 7792 20000 7848
rect 16021 7790 20000 7792
rect 16021 7787 16087 7790
rect 19520 7760 20000 7790
rect 4277 7648 4597 7649
rect 4277 7584 4285 7648
rect 4349 7584 4365 7648
rect 4429 7584 4445 7648
rect 4509 7584 4525 7648
rect 4589 7584 4597 7648
rect 4277 7583 4597 7584
rect 10944 7648 11264 7649
rect 10944 7584 10952 7648
rect 11016 7584 11032 7648
rect 11096 7584 11112 7648
rect 11176 7584 11192 7648
rect 11256 7584 11264 7648
rect 10944 7583 11264 7584
rect 17610 7648 17930 7649
rect 17610 7584 17618 7648
rect 17682 7584 17698 7648
rect 17762 7584 17778 7648
rect 17842 7584 17858 7648
rect 17922 7584 17930 7648
rect 17610 7583 17930 7584
rect 0 7442 480 7472
rect 8753 7442 8819 7445
rect 0 7440 8819 7442
rect 0 7384 8758 7440
rect 8814 7384 8819 7440
rect 0 7382 8819 7384
rect 0 7352 480 7382
rect 8753 7379 8819 7382
rect 5717 7306 5783 7309
rect 9673 7306 9739 7309
rect 5717 7304 9739 7306
rect 5717 7248 5722 7304
rect 5778 7248 9678 7304
rect 9734 7248 9739 7304
rect 5717 7246 9739 7248
rect 5717 7243 5783 7246
rect 9673 7243 9739 7246
rect 4061 7170 4127 7173
rect 5533 7170 5599 7173
rect 4061 7168 5599 7170
rect 4061 7112 4066 7168
rect 4122 7112 5538 7168
rect 5594 7112 5599 7168
rect 4061 7110 5599 7112
rect 4061 7107 4127 7110
rect 5533 7107 5599 7110
rect 15193 7170 15259 7173
rect 19520 7170 20000 7200
rect 15193 7168 20000 7170
rect 15193 7112 15198 7168
rect 15254 7112 20000 7168
rect 15193 7110 20000 7112
rect 15193 7107 15259 7110
rect 7610 7104 7930 7105
rect 7610 7040 7618 7104
rect 7682 7040 7698 7104
rect 7762 7040 7778 7104
rect 7842 7040 7858 7104
rect 7922 7040 7930 7104
rect 7610 7039 7930 7040
rect 14277 7104 14597 7105
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 19520 7080 20000 7110
rect 14277 7039 14597 7040
rect 0 6762 480 6792
rect 3417 6762 3483 6765
rect 0 6760 3483 6762
rect 0 6704 3422 6760
rect 3478 6704 3483 6760
rect 0 6702 3483 6704
rect 0 6672 480 6702
rect 3417 6699 3483 6702
rect 7281 6762 7347 6765
rect 15929 6762 15995 6765
rect 17401 6762 17467 6765
rect 7281 6760 17467 6762
rect 7281 6704 7286 6760
rect 7342 6704 15934 6760
rect 15990 6704 17406 6760
rect 17462 6704 17467 6760
rect 7281 6702 17467 6704
rect 7281 6699 7347 6702
rect 15929 6699 15995 6702
rect 17401 6699 17467 6702
rect 4277 6560 4597 6561
rect 4277 6496 4285 6560
rect 4349 6496 4365 6560
rect 4429 6496 4445 6560
rect 4509 6496 4525 6560
rect 4589 6496 4597 6560
rect 4277 6495 4597 6496
rect 10944 6560 11264 6561
rect 10944 6496 10952 6560
rect 11016 6496 11032 6560
rect 11096 6496 11112 6560
rect 11176 6496 11192 6560
rect 11256 6496 11264 6560
rect 10944 6495 11264 6496
rect 17610 6560 17930 6561
rect 17610 6496 17618 6560
rect 17682 6496 17698 6560
rect 17762 6496 17778 6560
rect 17842 6496 17858 6560
rect 17922 6496 17930 6560
rect 17610 6495 17930 6496
rect 19520 6490 20000 6520
rect 18094 6430 20000 6490
rect 13629 6354 13695 6357
rect 18094 6354 18154 6430
rect 19520 6400 20000 6430
rect 13629 6352 18154 6354
rect 13629 6296 13634 6352
rect 13690 6296 18154 6352
rect 13629 6294 18154 6296
rect 13629 6291 13695 6294
rect 11789 6218 11855 6221
rect 11789 6216 15946 6218
rect 11789 6160 11794 6216
rect 11850 6160 15946 6216
rect 11789 6158 15946 6160
rect 11789 6155 11855 6158
rect 7610 6016 7930 6017
rect 0 5946 480 5976
rect 7610 5952 7618 6016
rect 7682 5952 7698 6016
rect 7762 5952 7778 6016
rect 7842 5952 7858 6016
rect 7922 5952 7930 6016
rect 7610 5951 7930 5952
rect 14277 6016 14597 6017
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 5951 14597 5952
rect 4061 5946 4127 5949
rect 0 5944 4127 5946
rect 0 5888 4066 5944
rect 4122 5888 4127 5944
rect 0 5886 4127 5888
rect 0 5856 480 5886
rect 4061 5883 4127 5886
rect 3785 5810 3851 5813
rect 14089 5810 14155 5813
rect 14641 5810 14707 5813
rect 3785 5808 14707 5810
rect 3785 5752 3790 5808
rect 3846 5752 14094 5808
rect 14150 5752 14646 5808
rect 14702 5752 14707 5808
rect 3785 5750 14707 5752
rect 15886 5810 15946 6158
rect 16297 6082 16363 6085
rect 16665 6082 16731 6085
rect 16297 6080 16731 6082
rect 16297 6024 16302 6080
rect 16358 6024 16670 6080
rect 16726 6024 16731 6080
rect 16297 6022 16731 6024
rect 16297 6019 16363 6022
rect 16665 6019 16731 6022
rect 19520 5810 20000 5840
rect 15886 5750 20000 5810
rect 3785 5747 3851 5750
rect 14089 5747 14155 5750
rect 14641 5747 14707 5750
rect 19520 5720 20000 5750
rect 11421 5674 11487 5677
rect 16021 5674 16087 5677
rect 11421 5672 16087 5674
rect 11421 5616 11426 5672
rect 11482 5616 16026 5672
rect 16082 5616 16087 5672
rect 11421 5614 16087 5616
rect 11421 5611 11487 5614
rect 16021 5611 16087 5614
rect 4277 5472 4597 5473
rect 4277 5408 4285 5472
rect 4349 5408 4365 5472
rect 4429 5408 4445 5472
rect 4509 5408 4525 5472
rect 4589 5408 4597 5472
rect 4277 5407 4597 5408
rect 10944 5472 11264 5473
rect 10944 5408 10952 5472
rect 11016 5408 11032 5472
rect 11096 5408 11112 5472
rect 11176 5408 11192 5472
rect 11256 5408 11264 5472
rect 10944 5407 11264 5408
rect 17610 5472 17930 5473
rect 17610 5408 17618 5472
rect 17682 5408 17698 5472
rect 17762 5408 17778 5472
rect 17842 5408 17858 5472
rect 17922 5408 17930 5472
rect 17610 5407 17930 5408
rect 0 5130 480 5160
rect 2129 5130 2195 5133
rect 0 5128 2195 5130
rect 0 5072 2134 5128
rect 2190 5072 2195 5128
rect 0 5070 2195 5072
rect 0 5040 480 5070
rect 2129 5067 2195 5070
rect 16113 5130 16179 5133
rect 19520 5130 20000 5160
rect 16113 5128 20000 5130
rect 16113 5072 16118 5128
rect 16174 5072 20000 5128
rect 16113 5070 20000 5072
rect 16113 5067 16179 5070
rect 19520 5040 20000 5070
rect 7610 4928 7930 4929
rect 7610 4864 7618 4928
rect 7682 4864 7698 4928
rect 7762 4864 7778 4928
rect 7842 4864 7858 4928
rect 7922 4864 7930 4928
rect 7610 4863 7930 4864
rect 14277 4928 14597 4929
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 4863 14597 4864
rect 4061 4722 4127 4725
rect 9857 4722 9923 4725
rect 10041 4722 10107 4725
rect 14641 4722 14707 4725
rect 4061 4720 9923 4722
rect 4061 4664 4066 4720
rect 4122 4664 9862 4720
rect 9918 4664 9923 4720
rect 4061 4662 9923 4664
rect 4061 4659 4127 4662
rect 9857 4659 9923 4662
rect 9998 4720 14707 4722
rect 9998 4664 10046 4720
rect 10102 4664 14646 4720
rect 14702 4664 14707 4720
rect 9998 4662 14707 4664
rect 9998 4659 10107 4662
rect 14641 4659 14707 4662
rect 3049 4586 3115 4589
rect 9998 4586 10058 4659
rect 3049 4584 10058 4586
rect 3049 4528 3054 4584
rect 3110 4528 10058 4584
rect 3049 4526 10058 4528
rect 17033 4586 17099 4589
rect 17033 4584 18154 4586
rect 17033 4528 17038 4584
rect 17094 4528 18154 4584
rect 17033 4526 18154 4528
rect 3049 4523 3115 4526
rect 17033 4523 17099 4526
rect 18094 4450 18154 4526
rect 19520 4450 20000 4480
rect 18094 4390 20000 4450
rect 4277 4384 4597 4385
rect 0 4314 480 4344
rect 4277 4320 4285 4384
rect 4349 4320 4365 4384
rect 4429 4320 4445 4384
rect 4509 4320 4525 4384
rect 4589 4320 4597 4384
rect 4277 4319 4597 4320
rect 10944 4384 11264 4385
rect 10944 4320 10952 4384
rect 11016 4320 11032 4384
rect 11096 4320 11112 4384
rect 11176 4320 11192 4384
rect 11256 4320 11264 4384
rect 10944 4319 11264 4320
rect 17610 4384 17930 4385
rect 17610 4320 17618 4384
rect 17682 4320 17698 4384
rect 17762 4320 17778 4384
rect 17842 4320 17858 4384
rect 17922 4320 17930 4384
rect 19520 4360 20000 4390
rect 17610 4319 17930 4320
rect 1669 4314 1735 4317
rect 0 4312 1735 4314
rect 0 4256 1674 4312
rect 1730 4256 1735 4312
rect 0 4254 1735 4256
rect 0 4224 480 4254
rect 1669 4251 1735 4254
rect 7610 3840 7930 3841
rect 7610 3776 7618 3840
rect 7682 3776 7698 3840
rect 7762 3776 7778 3840
rect 7842 3776 7858 3840
rect 7922 3776 7930 3840
rect 7610 3775 7930 3776
rect 14277 3840 14597 3841
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 3775 14597 3776
rect 16389 3770 16455 3773
rect 19520 3770 20000 3800
rect 16389 3768 20000 3770
rect 16389 3712 16394 3768
rect 16450 3712 20000 3768
rect 16389 3710 20000 3712
rect 16389 3707 16455 3710
rect 19520 3680 20000 3710
rect 0 3498 480 3528
rect 4061 3498 4127 3501
rect 0 3496 4127 3498
rect 0 3440 4066 3496
rect 4122 3440 4127 3496
rect 0 3438 4127 3440
rect 0 3408 480 3438
rect 4061 3435 4127 3438
rect 4277 3296 4597 3297
rect 4277 3232 4285 3296
rect 4349 3232 4365 3296
rect 4429 3232 4445 3296
rect 4509 3232 4525 3296
rect 4589 3232 4597 3296
rect 4277 3231 4597 3232
rect 10944 3296 11264 3297
rect 10944 3232 10952 3296
rect 11016 3232 11032 3296
rect 11096 3232 11112 3296
rect 11176 3232 11192 3296
rect 11256 3232 11264 3296
rect 10944 3231 11264 3232
rect 17610 3296 17930 3297
rect 17610 3232 17618 3296
rect 17682 3232 17698 3296
rect 17762 3232 17778 3296
rect 17842 3232 17858 3296
rect 17922 3232 17930 3296
rect 17610 3231 17930 3232
rect 15561 3090 15627 3093
rect 19520 3090 20000 3120
rect 15561 3088 20000 3090
rect 15561 3032 15566 3088
rect 15622 3032 20000 3088
rect 15561 3030 20000 3032
rect 15561 3027 15627 3030
rect 19520 3000 20000 3030
rect 7610 2752 7930 2753
rect 0 2682 480 2712
rect 7610 2688 7618 2752
rect 7682 2688 7698 2752
rect 7762 2688 7778 2752
rect 7842 2688 7858 2752
rect 7922 2688 7930 2752
rect 7610 2687 7930 2688
rect 14277 2752 14597 2753
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2687 14597 2688
rect 7281 2682 7347 2685
rect 0 2680 7347 2682
rect 0 2624 7286 2680
rect 7342 2624 7347 2680
rect 0 2622 7347 2624
rect 0 2592 480 2622
rect 7281 2619 7347 2622
rect 3417 2546 3483 2549
rect 10041 2546 10107 2549
rect 3417 2544 10107 2546
rect 3417 2488 3422 2544
rect 3478 2488 10046 2544
rect 10102 2488 10107 2544
rect 3417 2486 10107 2488
rect 3417 2483 3483 2486
rect 10041 2483 10107 2486
rect 16481 2410 16547 2413
rect 19520 2410 20000 2440
rect 16481 2408 20000 2410
rect 16481 2352 16486 2408
rect 16542 2352 20000 2408
rect 16481 2350 20000 2352
rect 16481 2347 16547 2350
rect 19520 2320 20000 2350
rect 4277 2208 4597 2209
rect 4277 2144 4285 2208
rect 4349 2144 4365 2208
rect 4429 2144 4445 2208
rect 4509 2144 4525 2208
rect 4589 2144 4597 2208
rect 4277 2143 4597 2144
rect 10944 2208 11264 2209
rect 10944 2144 10952 2208
rect 11016 2144 11032 2208
rect 11096 2144 11112 2208
rect 11176 2144 11192 2208
rect 11256 2144 11264 2208
rect 10944 2143 11264 2144
rect 17610 2208 17930 2209
rect 17610 2144 17618 2208
rect 17682 2144 17698 2208
rect 17762 2144 17778 2208
rect 17842 2144 17858 2208
rect 17922 2144 17930 2208
rect 17610 2143 17930 2144
rect 0 1866 480 1896
rect 3417 1866 3483 1869
rect 0 1864 3483 1866
rect 0 1808 3422 1864
rect 3478 1808 3483 1864
rect 0 1806 3483 1808
rect 0 1776 480 1806
rect 3417 1803 3483 1806
rect 16297 1730 16363 1733
rect 19520 1730 20000 1760
rect 16297 1728 20000 1730
rect 16297 1672 16302 1728
rect 16358 1672 20000 1728
rect 16297 1670 20000 1672
rect 16297 1667 16363 1670
rect 19520 1640 20000 1670
rect 9489 1458 9555 1461
rect 3374 1456 9555 1458
rect 3374 1400 9494 1456
rect 9550 1400 9555 1456
rect 3374 1398 9555 1400
rect 0 1050 480 1080
rect 3374 1050 3434 1398
rect 9489 1395 9555 1398
rect 0 990 3434 1050
rect 15193 1050 15259 1053
rect 19520 1050 20000 1080
rect 15193 1048 20000 1050
rect 15193 992 15198 1048
rect 15254 992 20000 1048
rect 15193 990 20000 992
rect 0 960 480 990
rect 15193 987 15259 990
rect 19520 960 20000 990
rect 0 370 480 400
rect 9305 370 9371 373
rect 0 368 9371 370
rect 0 312 9310 368
rect 9366 312 9371 368
rect 0 310 9371 312
rect 0 280 480 310
rect 9305 307 9371 310
rect 11329 370 11395 373
rect 19520 370 20000 400
rect 11329 368 20000 370
rect 11329 312 11334 368
rect 11390 312 20000 368
rect 11329 310 20000 312
rect 11329 307 11395 310
rect 19520 280 20000 310
<< via3 >>
rect 5396 79596 5460 79660
rect 7618 77820 7682 77824
rect 7618 77764 7622 77820
rect 7622 77764 7678 77820
rect 7678 77764 7682 77820
rect 7618 77760 7682 77764
rect 7698 77820 7762 77824
rect 7698 77764 7702 77820
rect 7702 77764 7758 77820
rect 7758 77764 7762 77820
rect 7698 77760 7762 77764
rect 7778 77820 7842 77824
rect 7778 77764 7782 77820
rect 7782 77764 7838 77820
rect 7838 77764 7842 77820
rect 7778 77760 7842 77764
rect 7858 77820 7922 77824
rect 7858 77764 7862 77820
rect 7862 77764 7918 77820
rect 7918 77764 7922 77820
rect 7858 77760 7922 77764
rect 14285 77820 14349 77824
rect 14285 77764 14289 77820
rect 14289 77764 14345 77820
rect 14345 77764 14349 77820
rect 14285 77760 14349 77764
rect 14365 77820 14429 77824
rect 14365 77764 14369 77820
rect 14369 77764 14425 77820
rect 14425 77764 14429 77820
rect 14365 77760 14429 77764
rect 14445 77820 14509 77824
rect 14445 77764 14449 77820
rect 14449 77764 14505 77820
rect 14505 77764 14509 77820
rect 14445 77760 14509 77764
rect 14525 77820 14589 77824
rect 14525 77764 14529 77820
rect 14529 77764 14585 77820
rect 14585 77764 14589 77820
rect 14525 77760 14589 77764
rect 14964 77420 15028 77484
rect 4285 77276 4349 77280
rect 4285 77220 4289 77276
rect 4289 77220 4345 77276
rect 4345 77220 4349 77276
rect 4285 77216 4349 77220
rect 4365 77276 4429 77280
rect 4365 77220 4369 77276
rect 4369 77220 4425 77276
rect 4425 77220 4429 77276
rect 4365 77216 4429 77220
rect 4445 77276 4509 77280
rect 4445 77220 4449 77276
rect 4449 77220 4505 77276
rect 4505 77220 4509 77276
rect 4445 77216 4509 77220
rect 4525 77276 4589 77280
rect 4525 77220 4529 77276
rect 4529 77220 4585 77276
rect 4585 77220 4589 77276
rect 4525 77216 4589 77220
rect 10952 77276 11016 77280
rect 10952 77220 10956 77276
rect 10956 77220 11012 77276
rect 11012 77220 11016 77276
rect 10952 77216 11016 77220
rect 11032 77276 11096 77280
rect 11032 77220 11036 77276
rect 11036 77220 11092 77276
rect 11092 77220 11096 77276
rect 11032 77216 11096 77220
rect 11112 77276 11176 77280
rect 11112 77220 11116 77276
rect 11116 77220 11172 77276
rect 11172 77220 11176 77276
rect 11112 77216 11176 77220
rect 11192 77276 11256 77280
rect 11192 77220 11196 77276
rect 11196 77220 11252 77276
rect 11252 77220 11256 77276
rect 11192 77216 11256 77220
rect 17618 77276 17682 77280
rect 17618 77220 17622 77276
rect 17622 77220 17678 77276
rect 17678 77220 17682 77276
rect 17618 77216 17682 77220
rect 17698 77276 17762 77280
rect 17698 77220 17702 77276
rect 17702 77220 17758 77276
rect 17758 77220 17762 77276
rect 17698 77216 17762 77220
rect 17778 77276 17842 77280
rect 17778 77220 17782 77276
rect 17782 77220 17838 77276
rect 17838 77220 17842 77276
rect 17778 77216 17842 77220
rect 17858 77276 17922 77280
rect 17858 77220 17862 77276
rect 17862 77220 17918 77276
rect 17918 77220 17922 77276
rect 17858 77216 17922 77220
rect 7618 76732 7682 76736
rect 7618 76676 7622 76732
rect 7622 76676 7678 76732
rect 7678 76676 7682 76732
rect 7618 76672 7682 76676
rect 7698 76732 7762 76736
rect 7698 76676 7702 76732
rect 7702 76676 7758 76732
rect 7758 76676 7762 76732
rect 7698 76672 7762 76676
rect 7778 76732 7842 76736
rect 7778 76676 7782 76732
rect 7782 76676 7838 76732
rect 7838 76676 7842 76732
rect 7778 76672 7842 76676
rect 7858 76732 7922 76736
rect 7858 76676 7862 76732
rect 7862 76676 7918 76732
rect 7918 76676 7922 76732
rect 7858 76672 7922 76676
rect 14285 76732 14349 76736
rect 14285 76676 14289 76732
rect 14289 76676 14345 76732
rect 14345 76676 14349 76732
rect 14285 76672 14349 76676
rect 14365 76732 14429 76736
rect 14365 76676 14369 76732
rect 14369 76676 14425 76732
rect 14425 76676 14429 76732
rect 14365 76672 14429 76676
rect 14445 76732 14509 76736
rect 14445 76676 14449 76732
rect 14449 76676 14505 76732
rect 14505 76676 14509 76732
rect 14445 76672 14509 76676
rect 14525 76732 14589 76736
rect 14525 76676 14529 76732
rect 14529 76676 14585 76732
rect 14585 76676 14589 76732
rect 14525 76672 14589 76676
rect 5212 76332 5276 76396
rect 4285 76188 4349 76192
rect 4285 76132 4289 76188
rect 4289 76132 4345 76188
rect 4345 76132 4349 76188
rect 4285 76128 4349 76132
rect 4365 76188 4429 76192
rect 4365 76132 4369 76188
rect 4369 76132 4425 76188
rect 4425 76132 4429 76188
rect 4365 76128 4429 76132
rect 4445 76188 4509 76192
rect 4445 76132 4449 76188
rect 4449 76132 4505 76188
rect 4505 76132 4509 76188
rect 4445 76128 4509 76132
rect 4525 76188 4589 76192
rect 4525 76132 4529 76188
rect 4529 76132 4585 76188
rect 4585 76132 4589 76188
rect 4525 76128 4589 76132
rect 10952 76188 11016 76192
rect 10952 76132 10956 76188
rect 10956 76132 11012 76188
rect 11012 76132 11016 76188
rect 10952 76128 11016 76132
rect 11032 76188 11096 76192
rect 11032 76132 11036 76188
rect 11036 76132 11092 76188
rect 11092 76132 11096 76188
rect 11032 76128 11096 76132
rect 11112 76188 11176 76192
rect 11112 76132 11116 76188
rect 11116 76132 11172 76188
rect 11172 76132 11176 76188
rect 11112 76128 11176 76132
rect 11192 76188 11256 76192
rect 11192 76132 11196 76188
rect 11196 76132 11252 76188
rect 11252 76132 11256 76188
rect 11192 76128 11256 76132
rect 17618 76188 17682 76192
rect 17618 76132 17622 76188
rect 17622 76132 17678 76188
rect 17678 76132 17682 76188
rect 17618 76128 17682 76132
rect 17698 76188 17762 76192
rect 17698 76132 17702 76188
rect 17702 76132 17758 76188
rect 17758 76132 17762 76188
rect 17698 76128 17762 76132
rect 17778 76188 17842 76192
rect 17778 76132 17782 76188
rect 17782 76132 17838 76188
rect 17838 76132 17842 76188
rect 17778 76128 17842 76132
rect 17858 76188 17922 76192
rect 17858 76132 17862 76188
rect 17862 76132 17918 76188
rect 17918 76132 17922 76188
rect 17858 76128 17922 76132
rect 4844 75924 4908 75988
rect 7618 75644 7682 75648
rect 7618 75588 7622 75644
rect 7622 75588 7678 75644
rect 7678 75588 7682 75644
rect 7618 75584 7682 75588
rect 7698 75644 7762 75648
rect 7698 75588 7702 75644
rect 7702 75588 7758 75644
rect 7758 75588 7762 75644
rect 7698 75584 7762 75588
rect 7778 75644 7842 75648
rect 7778 75588 7782 75644
rect 7782 75588 7838 75644
rect 7838 75588 7842 75644
rect 7778 75584 7842 75588
rect 7858 75644 7922 75648
rect 7858 75588 7862 75644
rect 7862 75588 7918 75644
rect 7918 75588 7922 75644
rect 7858 75584 7922 75588
rect 14285 75644 14349 75648
rect 14285 75588 14289 75644
rect 14289 75588 14345 75644
rect 14345 75588 14349 75644
rect 14285 75584 14349 75588
rect 14365 75644 14429 75648
rect 14365 75588 14369 75644
rect 14369 75588 14425 75644
rect 14425 75588 14429 75644
rect 14365 75584 14429 75588
rect 14445 75644 14509 75648
rect 14445 75588 14449 75644
rect 14449 75588 14505 75644
rect 14505 75588 14509 75644
rect 14445 75584 14509 75588
rect 14525 75644 14589 75648
rect 14525 75588 14529 75644
rect 14529 75588 14585 75644
rect 14585 75588 14589 75644
rect 14525 75584 14589 75588
rect 5028 75380 5092 75444
rect 4285 75100 4349 75104
rect 4285 75044 4289 75100
rect 4289 75044 4345 75100
rect 4345 75044 4349 75100
rect 4285 75040 4349 75044
rect 4365 75100 4429 75104
rect 4365 75044 4369 75100
rect 4369 75044 4425 75100
rect 4425 75044 4429 75100
rect 4365 75040 4429 75044
rect 4445 75100 4509 75104
rect 4445 75044 4449 75100
rect 4449 75044 4505 75100
rect 4505 75044 4509 75100
rect 4445 75040 4509 75044
rect 4525 75100 4589 75104
rect 4525 75044 4529 75100
rect 4529 75044 4585 75100
rect 4585 75044 4589 75100
rect 4525 75040 4589 75044
rect 10952 75100 11016 75104
rect 10952 75044 10956 75100
rect 10956 75044 11012 75100
rect 11012 75044 11016 75100
rect 10952 75040 11016 75044
rect 11032 75100 11096 75104
rect 11032 75044 11036 75100
rect 11036 75044 11092 75100
rect 11092 75044 11096 75100
rect 11032 75040 11096 75044
rect 11112 75100 11176 75104
rect 11112 75044 11116 75100
rect 11116 75044 11172 75100
rect 11172 75044 11176 75100
rect 11112 75040 11176 75044
rect 11192 75100 11256 75104
rect 11192 75044 11196 75100
rect 11196 75044 11252 75100
rect 11252 75044 11256 75100
rect 11192 75040 11256 75044
rect 17618 75100 17682 75104
rect 17618 75044 17622 75100
rect 17622 75044 17678 75100
rect 17678 75044 17682 75100
rect 17618 75040 17682 75044
rect 17698 75100 17762 75104
rect 17698 75044 17702 75100
rect 17702 75044 17758 75100
rect 17758 75044 17762 75100
rect 17698 75040 17762 75044
rect 17778 75100 17842 75104
rect 17778 75044 17782 75100
rect 17782 75044 17838 75100
rect 17838 75044 17842 75100
rect 17778 75040 17842 75044
rect 17858 75100 17922 75104
rect 17858 75044 17862 75100
rect 17862 75044 17918 75100
rect 17918 75044 17922 75100
rect 17858 75040 17922 75044
rect 2452 74700 2516 74764
rect 7618 74556 7682 74560
rect 7618 74500 7622 74556
rect 7622 74500 7678 74556
rect 7678 74500 7682 74556
rect 7618 74496 7682 74500
rect 7698 74556 7762 74560
rect 7698 74500 7702 74556
rect 7702 74500 7758 74556
rect 7758 74500 7762 74556
rect 7698 74496 7762 74500
rect 7778 74556 7842 74560
rect 7778 74500 7782 74556
rect 7782 74500 7838 74556
rect 7838 74500 7842 74556
rect 7778 74496 7842 74500
rect 7858 74556 7922 74560
rect 7858 74500 7862 74556
rect 7862 74500 7918 74556
rect 7918 74500 7922 74556
rect 7858 74496 7922 74500
rect 14285 74556 14349 74560
rect 14285 74500 14289 74556
rect 14289 74500 14345 74556
rect 14345 74500 14349 74556
rect 14285 74496 14349 74500
rect 14365 74556 14429 74560
rect 14365 74500 14369 74556
rect 14369 74500 14425 74556
rect 14425 74500 14429 74556
rect 14365 74496 14429 74500
rect 14445 74556 14509 74560
rect 14445 74500 14449 74556
rect 14449 74500 14505 74556
rect 14505 74500 14509 74556
rect 14445 74496 14509 74500
rect 14525 74556 14589 74560
rect 14525 74500 14529 74556
rect 14529 74500 14585 74556
rect 14585 74500 14589 74556
rect 14525 74496 14589 74500
rect 4285 74012 4349 74016
rect 4285 73956 4289 74012
rect 4289 73956 4345 74012
rect 4345 73956 4349 74012
rect 4285 73952 4349 73956
rect 4365 74012 4429 74016
rect 4365 73956 4369 74012
rect 4369 73956 4425 74012
rect 4425 73956 4429 74012
rect 4365 73952 4429 73956
rect 4445 74012 4509 74016
rect 4445 73956 4449 74012
rect 4449 73956 4505 74012
rect 4505 73956 4509 74012
rect 4445 73952 4509 73956
rect 4525 74012 4589 74016
rect 4525 73956 4529 74012
rect 4529 73956 4585 74012
rect 4585 73956 4589 74012
rect 4525 73952 4589 73956
rect 10952 74012 11016 74016
rect 10952 73956 10956 74012
rect 10956 73956 11012 74012
rect 11012 73956 11016 74012
rect 10952 73952 11016 73956
rect 11032 74012 11096 74016
rect 11032 73956 11036 74012
rect 11036 73956 11092 74012
rect 11092 73956 11096 74012
rect 11032 73952 11096 73956
rect 11112 74012 11176 74016
rect 11112 73956 11116 74012
rect 11116 73956 11172 74012
rect 11172 73956 11176 74012
rect 11112 73952 11176 73956
rect 11192 74012 11256 74016
rect 11192 73956 11196 74012
rect 11196 73956 11252 74012
rect 11252 73956 11256 74012
rect 11192 73952 11256 73956
rect 17618 74012 17682 74016
rect 17618 73956 17622 74012
rect 17622 73956 17678 74012
rect 17678 73956 17682 74012
rect 17618 73952 17682 73956
rect 17698 74012 17762 74016
rect 17698 73956 17702 74012
rect 17702 73956 17758 74012
rect 17758 73956 17762 74012
rect 17698 73952 17762 73956
rect 17778 74012 17842 74016
rect 17778 73956 17782 74012
rect 17782 73956 17838 74012
rect 17838 73956 17842 74012
rect 17778 73952 17842 73956
rect 17858 74012 17922 74016
rect 17858 73956 17862 74012
rect 17862 73956 17918 74012
rect 17918 73956 17922 74012
rect 17858 73952 17922 73956
rect 7236 73748 7300 73812
rect 7618 73468 7682 73472
rect 7618 73412 7622 73468
rect 7622 73412 7678 73468
rect 7678 73412 7682 73468
rect 7618 73408 7682 73412
rect 7698 73468 7762 73472
rect 7698 73412 7702 73468
rect 7702 73412 7758 73468
rect 7758 73412 7762 73468
rect 7698 73408 7762 73412
rect 7778 73468 7842 73472
rect 7778 73412 7782 73468
rect 7782 73412 7838 73468
rect 7838 73412 7842 73468
rect 7778 73408 7842 73412
rect 7858 73468 7922 73472
rect 7858 73412 7862 73468
rect 7862 73412 7918 73468
rect 7918 73412 7922 73468
rect 7858 73408 7922 73412
rect 14285 73468 14349 73472
rect 14285 73412 14289 73468
rect 14289 73412 14345 73468
rect 14345 73412 14349 73468
rect 14285 73408 14349 73412
rect 14365 73468 14429 73472
rect 14365 73412 14369 73468
rect 14369 73412 14425 73468
rect 14425 73412 14429 73468
rect 14365 73408 14429 73412
rect 14445 73468 14509 73472
rect 14445 73412 14449 73468
rect 14449 73412 14505 73468
rect 14505 73412 14509 73468
rect 14445 73408 14509 73412
rect 14525 73468 14589 73472
rect 14525 73412 14529 73468
rect 14529 73412 14585 73468
rect 14585 73412 14589 73468
rect 14525 73408 14589 73412
rect 10732 73264 10796 73268
rect 10732 73208 10746 73264
rect 10746 73208 10796 73264
rect 10732 73204 10796 73208
rect 4285 72924 4349 72928
rect 4285 72868 4289 72924
rect 4289 72868 4345 72924
rect 4345 72868 4349 72924
rect 4285 72864 4349 72868
rect 4365 72924 4429 72928
rect 4365 72868 4369 72924
rect 4369 72868 4425 72924
rect 4425 72868 4429 72924
rect 4365 72864 4429 72868
rect 4445 72924 4509 72928
rect 4445 72868 4449 72924
rect 4449 72868 4505 72924
rect 4505 72868 4509 72924
rect 4445 72864 4509 72868
rect 4525 72924 4589 72928
rect 4525 72868 4529 72924
rect 4529 72868 4585 72924
rect 4585 72868 4589 72924
rect 4525 72864 4589 72868
rect 10952 72924 11016 72928
rect 10952 72868 10956 72924
rect 10956 72868 11012 72924
rect 11012 72868 11016 72924
rect 10952 72864 11016 72868
rect 11032 72924 11096 72928
rect 11032 72868 11036 72924
rect 11036 72868 11092 72924
rect 11092 72868 11096 72924
rect 11032 72864 11096 72868
rect 11112 72924 11176 72928
rect 11112 72868 11116 72924
rect 11116 72868 11172 72924
rect 11172 72868 11176 72924
rect 11112 72864 11176 72868
rect 11192 72924 11256 72928
rect 11192 72868 11196 72924
rect 11196 72868 11252 72924
rect 11252 72868 11256 72924
rect 11192 72864 11256 72868
rect 17618 72924 17682 72928
rect 17618 72868 17622 72924
rect 17622 72868 17678 72924
rect 17678 72868 17682 72924
rect 17618 72864 17682 72868
rect 17698 72924 17762 72928
rect 17698 72868 17702 72924
rect 17702 72868 17758 72924
rect 17758 72868 17762 72924
rect 17698 72864 17762 72868
rect 17778 72924 17842 72928
rect 17778 72868 17782 72924
rect 17782 72868 17838 72924
rect 17838 72868 17842 72924
rect 17778 72864 17842 72868
rect 17858 72924 17922 72928
rect 17858 72868 17862 72924
rect 17862 72868 17918 72924
rect 17918 72868 17922 72924
rect 17858 72864 17922 72868
rect 7618 72380 7682 72384
rect 7618 72324 7622 72380
rect 7622 72324 7678 72380
rect 7678 72324 7682 72380
rect 7618 72320 7682 72324
rect 7698 72380 7762 72384
rect 7698 72324 7702 72380
rect 7702 72324 7758 72380
rect 7758 72324 7762 72380
rect 7698 72320 7762 72324
rect 7778 72380 7842 72384
rect 7778 72324 7782 72380
rect 7782 72324 7838 72380
rect 7838 72324 7842 72380
rect 7778 72320 7842 72324
rect 7858 72380 7922 72384
rect 7858 72324 7862 72380
rect 7862 72324 7918 72380
rect 7918 72324 7922 72380
rect 7858 72320 7922 72324
rect 14285 72380 14349 72384
rect 14285 72324 14289 72380
rect 14289 72324 14345 72380
rect 14345 72324 14349 72380
rect 14285 72320 14349 72324
rect 14365 72380 14429 72384
rect 14365 72324 14369 72380
rect 14369 72324 14425 72380
rect 14425 72324 14429 72380
rect 14365 72320 14429 72324
rect 14445 72380 14509 72384
rect 14445 72324 14449 72380
rect 14449 72324 14505 72380
rect 14505 72324 14509 72380
rect 14445 72320 14509 72324
rect 14525 72380 14589 72384
rect 14525 72324 14529 72380
rect 14529 72324 14585 72380
rect 14585 72324 14589 72380
rect 14525 72320 14589 72324
rect 4285 71836 4349 71840
rect 4285 71780 4289 71836
rect 4289 71780 4345 71836
rect 4345 71780 4349 71836
rect 4285 71776 4349 71780
rect 4365 71836 4429 71840
rect 4365 71780 4369 71836
rect 4369 71780 4425 71836
rect 4425 71780 4429 71836
rect 4365 71776 4429 71780
rect 4445 71836 4509 71840
rect 4445 71780 4449 71836
rect 4449 71780 4505 71836
rect 4505 71780 4509 71836
rect 4445 71776 4509 71780
rect 4525 71836 4589 71840
rect 4525 71780 4529 71836
rect 4529 71780 4585 71836
rect 4585 71780 4589 71836
rect 4525 71776 4589 71780
rect 10952 71836 11016 71840
rect 10952 71780 10956 71836
rect 10956 71780 11012 71836
rect 11012 71780 11016 71836
rect 10952 71776 11016 71780
rect 11032 71836 11096 71840
rect 11032 71780 11036 71836
rect 11036 71780 11092 71836
rect 11092 71780 11096 71836
rect 11032 71776 11096 71780
rect 11112 71836 11176 71840
rect 11112 71780 11116 71836
rect 11116 71780 11172 71836
rect 11172 71780 11176 71836
rect 11112 71776 11176 71780
rect 11192 71836 11256 71840
rect 11192 71780 11196 71836
rect 11196 71780 11252 71836
rect 11252 71780 11256 71836
rect 11192 71776 11256 71780
rect 17618 71836 17682 71840
rect 17618 71780 17622 71836
rect 17622 71780 17678 71836
rect 17678 71780 17682 71836
rect 17618 71776 17682 71780
rect 17698 71836 17762 71840
rect 17698 71780 17702 71836
rect 17702 71780 17758 71836
rect 17758 71780 17762 71836
rect 17698 71776 17762 71780
rect 17778 71836 17842 71840
rect 17778 71780 17782 71836
rect 17782 71780 17838 71836
rect 17838 71780 17842 71836
rect 17778 71776 17842 71780
rect 17858 71836 17922 71840
rect 17858 71780 17862 71836
rect 17862 71780 17918 71836
rect 17918 71780 17922 71836
rect 17858 71776 17922 71780
rect 4108 71436 4172 71500
rect 16620 71300 16684 71364
rect 7618 71292 7682 71296
rect 7618 71236 7622 71292
rect 7622 71236 7678 71292
rect 7678 71236 7682 71292
rect 7618 71232 7682 71236
rect 7698 71292 7762 71296
rect 7698 71236 7702 71292
rect 7702 71236 7758 71292
rect 7758 71236 7762 71292
rect 7698 71232 7762 71236
rect 7778 71292 7842 71296
rect 7778 71236 7782 71292
rect 7782 71236 7838 71292
rect 7838 71236 7842 71292
rect 7778 71232 7842 71236
rect 7858 71292 7922 71296
rect 7858 71236 7862 71292
rect 7862 71236 7918 71292
rect 7918 71236 7922 71292
rect 7858 71232 7922 71236
rect 14285 71292 14349 71296
rect 14285 71236 14289 71292
rect 14289 71236 14345 71292
rect 14345 71236 14349 71292
rect 14285 71232 14349 71236
rect 14365 71292 14429 71296
rect 14365 71236 14369 71292
rect 14369 71236 14425 71292
rect 14425 71236 14429 71292
rect 14365 71232 14429 71236
rect 14445 71292 14509 71296
rect 14445 71236 14449 71292
rect 14449 71236 14505 71292
rect 14505 71236 14509 71292
rect 14445 71232 14509 71236
rect 14525 71292 14589 71296
rect 14525 71236 14529 71292
rect 14529 71236 14585 71292
rect 14585 71236 14589 71292
rect 14525 71232 14589 71236
rect 4285 70748 4349 70752
rect 4285 70692 4289 70748
rect 4289 70692 4345 70748
rect 4345 70692 4349 70748
rect 4285 70688 4349 70692
rect 4365 70748 4429 70752
rect 4365 70692 4369 70748
rect 4369 70692 4425 70748
rect 4425 70692 4429 70748
rect 4365 70688 4429 70692
rect 4445 70748 4509 70752
rect 4445 70692 4449 70748
rect 4449 70692 4505 70748
rect 4505 70692 4509 70748
rect 4445 70688 4509 70692
rect 4525 70748 4589 70752
rect 4525 70692 4529 70748
rect 4529 70692 4585 70748
rect 4585 70692 4589 70748
rect 4525 70688 4589 70692
rect 10952 70748 11016 70752
rect 10952 70692 10956 70748
rect 10956 70692 11012 70748
rect 11012 70692 11016 70748
rect 10952 70688 11016 70692
rect 11032 70748 11096 70752
rect 11032 70692 11036 70748
rect 11036 70692 11092 70748
rect 11092 70692 11096 70748
rect 11032 70688 11096 70692
rect 11112 70748 11176 70752
rect 11112 70692 11116 70748
rect 11116 70692 11172 70748
rect 11172 70692 11176 70748
rect 11112 70688 11176 70692
rect 11192 70748 11256 70752
rect 11192 70692 11196 70748
rect 11196 70692 11252 70748
rect 11252 70692 11256 70748
rect 11192 70688 11256 70692
rect 17618 70748 17682 70752
rect 17618 70692 17622 70748
rect 17622 70692 17678 70748
rect 17678 70692 17682 70748
rect 17618 70688 17682 70692
rect 17698 70748 17762 70752
rect 17698 70692 17702 70748
rect 17702 70692 17758 70748
rect 17758 70692 17762 70748
rect 17698 70688 17762 70692
rect 17778 70748 17842 70752
rect 17778 70692 17782 70748
rect 17782 70692 17838 70748
rect 17838 70692 17842 70748
rect 17778 70688 17842 70692
rect 17858 70748 17922 70752
rect 17858 70692 17862 70748
rect 17862 70692 17918 70748
rect 17918 70692 17922 70748
rect 17858 70688 17922 70692
rect 9628 70680 9692 70684
rect 9628 70624 9642 70680
rect 9642 70624 9692 70680
rect 9628 70620 9692 70624
rect 4660 70484 4724 70548
rect 8156 70348 8220 70412
rect 7618 70204 7682 70208
rect 7618 70148 7622 70204
rect 7622 70148 7678 70204
rect 7678 70148 7682 70204
rect 7618 70144 7682 70148
rect 7698 70204 7762 70208
rect 7698 70148 7702 70204
rect 7702 70148 7758 70204
rect 7758 70148 7762 70204
rect 7698 70144 7762 70148
rect 7778 70204 7842 70208
rect 7778 70148 7782 70204
rect 7782 70148 7838 70204
rect 7838 70148 7842 70204
rect 7778 70144 7842 70148
rect 7858 70204 7922 70208
rect 7858 70148 7862 70204
rect 7862 70148 7918 70204
rect 7918 70148 7922 70204
rect 7858 70144 7922 70148
rect 14285 70204 14349 70208
rect 14285 70148 14289 70204
rect 14289 70148 14345 70204
rect 14345 70148 14349 70204
rect 14285 70144 14349 70148
rect 14365 70204 14429 70208
rect 14365 70148 14369 70204
rect 14369 70148 14425 70204
rect 14425 70148 14429 70204
rect 14365 70144 14429 70148
rect 14445 70204 14509 70208
rect 14445 70148 14449 70204
rect 14449 70148 14505 70204
rect 14505 70148 14509 70204
rect 14445 70144 14509 70148
rect 14525 70204 14589 70208
rect 14525 70148 14529 70204
rect 14529 70148 14585 70204
rect 14585 70148 14589 70204
rect 14525 70144 14589 70148
rect 6868 69668 6932 69732
rect 4285 69660 4349 69664
rect 4285 69604 4289 69660
rect 4289 69604 4345 69660
rect 4345 69604 4349 69660
rect 4285 69600 4349 69604
rect 4365 69660 4429 69664
rect 4365 69604 4369 69660
rect 4369 69604 4425 69660
rect 4425 69604 4429 69660
rect 4365 69600 4429 69604
rect 4445 69660 4509 69664
rect 4445 69604 4449 69660
rect 4449 69604 4505 69660
rect 4505 69604 4509 69660
rect 4445 69600 4509 69604
rect 4525 69660 4589 69664
rect 4525 69604 4529 69660
rect 4529 69604 4585 69660
rect 4585 69604 4589 69660
rect 4525 69600 4589 69604
rect 10952 69660 11016 69664
rect 10952 69604 10956 69660
rect 10956 69604 11012 69660
rect 11012 69604 11016 69660
rect 10952 69600 11016 69604
rect 11032 69660 11096 69664
rect 11032 69604 11036 69660
rect 11036 69604 11092 69660
rect 11092 69604 11096 69660
rect 11032 69600 11096 69604
rect 11112 69660 11176 69664
rect 11112 69604 11116 69660
rect 11116 69604 11172 69660
rect 11172 69604 11176 69660
rect 11112 69600 11176 69604
rect 11192 69660 11256 69664
rect 11192 69604 11196 69660
rect 11196 69604 11252 69660
rect 11252 69604 11256 69660
rect 11192 69600 11256 69604
rect 17618 69660 17682 69664
rect 17618 69604 17622 69660
rect 17622 69604 17678 69660
rect 17678 69604 17682 69660
rect 17618 69600 17682 69604
rect 17698 69660 17762 69664
rect 17698 69604 17702 69660
rect 17702 69604 17758 69660
rect 17758 69604 17762 69660
rect 17698 69600 17762 69604
rect 17778 69660 17842 69664
rect 17778 69604 17782 69660
rect 17782 69604 17838 69660
rect 17838 69604 17842 69660
rect 17778 69600 17842 69604
rect 17858 69660 17922 69664
rect 17858 69604 17862 69660
rect 17862 69604 17918 69660
rect 17918 69604 17922 69660
rect 17858 69600 17922 69604
rect 7618 69116 7682 69120
rect 7618 69060 7622 69116
rect 7622 69060 7678 69116
rect 7678 69060 7682 69116
rect 7618 69056 7682 69060
rect 7698 69116 7762 69120
rect 7698 69060 7702 69116
rect 7702 69060 7758 69116
rect 7758 69060 7762 69116
rect 7698 69056 7762 69060
rect 7778 69116 7842 69120
rect 7778 69060 7782 69116
rect 7782 69060 7838 69116
rect 7838 69060 7842 69116
rect 7778 69056 7842 69060
rect 7858 69116 7922 69120
rect 7858 69060 7862 69116
rect 7862 69060 7918 69116
rect 7918 69060 7922 69116
rect 7858 69056 7922 69060
rect 14285 69116 14349 69120
rect 14285 69060 14289 69116
rect 14289 69060 14345 69116
rect 14345 69060 14349 69116
rect 14285 69056 14349 69060
rect 14365 69116 14429 69120
rect 14365 69060 14369 69116
rect 14369 69060 14425 69116
rect 14425 69060 14429 69116
rect 14365 69056 14429 69060
rect 14445 69116 14509 69120
rect 14445 69060 14449 69116
rect 14449 69060 14505 69116
rect 14505 69060 14509 69116
rect 14445 69056 14509 69060
rect 14525 69116 14589 69120
rect 14525 69060 14529 69116
rect 14529 69060 14585 69116
rect 14585 69060 14589 69116
rect 14525 69056 14589 69060
rect 12020 69048 12084 69052
rect 12020 68992 12034 69048
rect 12034 68992 12084 69048
rect 12020 68988 12084 68992
rect 2636 68716 2700 68780
rect 4285 68572 4349 68576
rect 4285 68516 4289 68572
rect 4289 68516 4345 68572
rect 4345 68516 4349 68572
rect 4285 68512 4349 68516
rect 4365 68572 4429 68576
rect 4365 68516 4369 68572
rect 4369 68516 4425 68572
rect 4425 68516 4429 68572
rect 4365 68512 4429 68516
rect 4445 68572 4509 68576
rect 4445 68516 4449 68572
rect 4449 68516 4505 68572
rect 4505 68516 4509 68572
rect 4445 68512 4509 68516
rect 4525 68572 4589 68576
rect 4525 68516 4529 68572
rect 4529 68516 4585 68572
rect 4585 68516 4589 68572
rect 4525 68512 4589 68516
rect 10952 68572 11016 68576
rect 10952 68516 10956 68572
rect 10956 68516 11012 68572
rect 11012 68516 11016 68572
rect 10952 68512 11016 68516
rect 11032 68572 11096 68576
rect 11032 68516 11036 68572
rect 11036 68516 11092 68572
rect 11092 68516 11096 68572
rect 11032 68512 11096 68516
rect 11112 68572 11176 68576
rect 11112 68516 11116 68572
rect 11116 68516 11172 68572
rect 11172 68516 11176 68572
rect 11112 68512 11176 68516
rect 11192 68572 11256 68576
rect 11192 68516 11196 68572
rect 11196 68516 11252 68572
rect 11252 68516 11256 68572
rect 11192 68512 11256 68516
rect 17618 68572 17682 68576
rect 17618 68516 17622 68572
rect 17622 68516 17678 68572
rect 17678 68516 17682 68572
rect 17618 68512 17682 68516
rect 17698 68572 17762 68576
rect 17698 68516 17702 68572
rect 17702 68516 17758 68572
rect 17758 68516 17762 68572
rect 17698 68512 17762 68516
rect 17778 68572 17842 68576
rect 17778 68516 17782 68572
rect 17782 68516 17838 68572
rect 17838 68516 17842 68572
rect 17778 68512 17842 68516
rect 17858 68572 17922 68576
rect 17858 68516 17862 68572
rect 17862 68516 17918 68572
rect 17918 68516 17922 68572
rect 17858 68512 17922 68516
rect 14044 68308 14108 68372
rect 13860 68096 13924 68100
rect 13860 68040 13910 68096
rect 13910 68040 13924 68096
rect 13860 68036 13924 68040
rect 7618 68028 7682 68032
rect 7618 67972 7622 68028
rect 7622 67972 7678 68028
rect 7678 67972 7682 68028
rect 7618 67968 7682 67972
rect 7698 68028 7762 68032
rect 7698 67972 7702 68028
rect 7702 67972 7758 68028
rect 7758 67972 7762 68028
rect 7698 67968 7762 67972
rect 7778 68028 7842 68032
rect 7778 67972 7782 68028
rect 7782 67972 7838 68028
rect 7838 67972 7842 68028
rect 7778 67968 7842 67972
rect 7858 68028 7922 68032
rect 7858 67972 7862 68028
rect 7862 67972 7918 68028
rect 7918 67972 7922 68028
rect 7858 67968 7922 67972
rect 14285 68028 14349 68032
rect 14285 67972 14289 68028
rect 14289 67972 14345 68028
rect 14345 67972 14349 68028
rect 14285 67968 14349 67972
rect 14365 68028 14429 68032
rect 14365 67972 14369 68028
rect 14369 67972 14425 68028
rect 14425 67972 14429 68028
rect 14365 67968 14429 67972
rect 14445 68028 14509 68032
rect 14445 67972 14449 68028
rect 14449 67972 14505 68028
rect 14505 67972 14509 68028
rect 14445 67968 14509 67972
rect 14525 68028 14589 68032
rect 14525 67972 14529 68028
rect 14529 67972 14585 68028
rect 14585 67972 14589 68028
rect 14525 67968 14589 67972
rect 4285 67484 4349 67488
rect 4285 67428 4289 67484
rect 4289 67428 4345 67484
rect 4345 67428 4349 67484
rect 4285 67424 4349 67428
rect 4365 67484 4429 67488
rect 4365 67428 4369 67484
rect 4369 67428 4425 67484
rect 4425 67428 4429 67484
rect 4365 67424 4429 67428
rect 4445 67484 4509 67488
rect 4445 67428 4449 67484
rect 4449 67428 4505 67484
rect 4505 67428 4509 67484
rect 4445 67424 4509 67428
rect 4525 67484 4589 67488
rect 4525 67428 4529 67484
rect 4529 67428 4585 67484
rect 4585 67428 4589 67484
rect 4525 67424 4589 67428
rect 10952 67484 11016 67488
rect 10952 67428 10956 67484
rect 10956 67428 11012 67484
rect 11012 67428 11016 67484
rect 10952 67424 11016 67428
rect 11032 67484 11096 67488
rect 11032 67428 11036 67484
rect 11036 67428 11092 67484
rect 11092 67428 11096 67484
rect 11032 67424 11096 67428
rect 11112 67484 11176 67488
rect 11112 67428 11116 67484
rect 11116 67428 11172 67484
rect 11172 67428 11176 67484
rect 11112 67424 11176 67428
rect 11192 67484 11256 67488
rect 11192 67428 11196 67484
rect 11196 67428 11252 67484
rect 11252 67428 11256 67484
rect 11192 67424 11256 67428
rect 17618 67484 17682 67488
rect 17618 67428 17622 67484
rect 17622 67428 17678 67484
rect 17678 67428 17682 67484
rect 17618 67424 17682 67428
rect 17698 67484 17762 67488
rect 17698 67428 17702 67484
rect 17702 67428 17758 67484
rect 17758 67428 17762 67484
rect 17698 67424 17762 67428
rect 17778 67484 17842 67488
rect 17778 67428 17782 67484
rect 17782 67428 17838 67484
rect 17838 67428 17842 67484
rect 17778 67424 17842 67428
rect 17858 67484 17922 67488
rect 17858 67428 17862 67484
rect 17862 67428 17918 67484
rect 17918 67428 17922 67484
rect 17858 67424 17922 67428
rect 7618 66940 7682 66944
rect 7618 66884 7622 66940
rect 7622 66884 7678 66940
rect 7678 66884 7682 66940
rect 7618 66880 7682 66884
rect 7698 66940 7762 66944
rect 7698 66884 7702 66940
rect 7702 66884 7758 66940
rect 7758 66884 7762 66940
rect 7698 66880 7762 66884
rect 7778 66940 7842 66944
rect 7778 66884 7782 66940
rect 7782 66884 7838 66940
rect 7838 66884 7842 66940
rect 7778 66880 7842 66884
rect 7858 66940 7922 66944
rect 7858 66884 7862 66940
rect 7862 66884 7918 66940
rect 7918 66884 7922 66940
rect 7858 66880 7922 66884
rect 14285 66940 14349 66944
rect 14285 66884 14289 66940
rect 14289 66884 14345 66940
rect 14345 66884 14349 66940
rect 14285 66880 14349 66884
rect 14365 66940 14429 66944
rect 14365 66884 14369 66940
rect 14369 66884 14425 66940
rect 14425 66884 14429 66940
rect 14365 66880 14429 66884
rect 14445 66940 14509 66944
rect 14445 66884 14449 66940
rect 14449 66884 14505 66940
rect 14505 66884 14509 66940
rect 14445 66880 14509 66884
rect 14525 66940 14589 66944
rect 14525 66884 14529 66940
rect 14529 66884 14585 66940
rect 14585 66884 14589 66940
rect 14525 66880 14589 66884
rect 4285 66396 4349 66400
rect 4285 66340 4289 66396
rect 4289 66340 4345 66396
rect 4345 66340 4349 66396
rect 4285 66336 4349 66340
rect 4365 66396 4429 66400
rect 4365 66340 4369 66396
rect 4369 66340 4425 66396
rect 4425 66340 4429 66396
rect 4365 66336 4429 66340
rect 4445 66396 4509 66400
rect 4445 66340 4449 66396
rect 4449 66340 4505 66396
rect 4505 66340 4509 66396
rect 4445 66336 4509 66340
rect 4525 66396 4589 66400
rect 4525 66340 4529 66396
rect 4529 66340 4585 66396
rect 4585 66340 4589 66396
rect 4525 66336 4589 66340
rect 10952 66396 11016 66400
rect 10952 66340 10956 66396
rect 10956 66340 11012 66396
rect 11012 66340 11016 66396
rect 10952 66336 11016 66340
rect 11032 66396 11096 66400
rect 11032 66340 11036 66396
rect 11036 66340 11092 66396
rect 11092 66340 11096 66396
rect 11032 66336 11096 66340
rect 11112 66396 11176 66400
rect 11112 66340 11116 66396
rect 11116 66340 11172 66396
rect 11172 66340 11176 66396
rect 11112 66336 11176 66340
rect 11192 66396 11256 66400
rect 11192 66340 11196 66396
rect 11196 66340 11252 66396
rect 11252 66340 11256 66396
rect 11192 66336 11256 66340
rect 17618 66396 17682 66400
rect 17618 66340 17622 66396
rect 17622 66340 17678 66396
rect 17678 66340 17682 66396
rect 17618 66336 17682 66340
rect 17698 66396 17762 66400
rect 17698 66340 17702 66396
rect 17702 66340 17758 66396
rect 17758 66340 17762 66396
rect 17698 66336 17762 66340
rect 17778 66396 17842 66400
rect 17778 66340 17782 66396
rect 17782 66340 17838 66396
rect 17838 66340 17842 66396
rect 17778 66336 17842 66340
rect 17858 66396 17922 66400
rect 17858 66340 17862 66396
rect 17862 66340 17918 66396
rect 17918 66340 17922 66396
rect 17858 66336 17922 66340
rect 10364 65860 10428 65924
rect 14780 65920 14844 65924
rect 14780 65864 14794 65920
rect 14794 65864 14844 65920
rect 14780 65860 14844 65864
rect 7618 65852 7682 65856
rect 7618 65796 7622 65852
rect 7622 65796 7678 65852
rect 7678 65796 7682 65852
rect 7618 65792 7682 65796
rect 7698 65852 7762 65856
rect 7698 65796 7702 65852
rect 7702 65796 7758 65852
rect 7758 65796 7762 65852
rect 7698 65792 7762 65796
rect 7778 65852 7842 65856
rect 7778 65796 7782 65852
rect 7782 65796 7838 65852
rect 7838 65796 7842 65852
rect 7778 65792 7842 65796
rect 7858 65852 7922 65856
rect 7858 65796 7862 65852
rect 7862 65796 7918 65852
rect 7918 65796 7922 65852
rect 7858 65792 7922 65796
rect 14285 65852 14349 65856
rect 14285 65796 14289 65852
rect 14289 65796 14345 65852
rect 14345 65796 14349 65852
rect 14285 65792 14349 65796
rect 14365 65852 14429 65856
rect 14365 65796 14369 65852
rect 14369 65796 14425 65852
rect 14425 65796 14429 65852
rect 14365 65792 14429 65796
rect 14445 65852 14509 65856
rect 14445 65796 14449 65852
rect 14449 65796 14505 65852
rect 14505 65796 14509 65852
rect 14445 65792 14509 65796
rect 14525 65852 14589 65856
rect 14525 65796 14529 65852
rect 14529 65796 14585 65852
rect 14585 65796 14589 65852
rect 14525 65792 14589 65796
rect 11468 65724 11532 65788
rect 4285 65308 4349 65312
rect 4285 65252 4289 65308
rect 4289 65252 4345 65308
rect 4345 65252 4349 65308
rect 4285 65248 4349 65252
rect 4365 65308 4429 65312
rect 4365 65252 4369 65308
rect 4369 65252 4425 65308
rect 4425 65252 4429 65308
rect 4365 65248 4429 65252
rect 4445 65308 4509 65312
rect 4445 65252 4449 65308
rect 4449 65252 4505 65308
rect 4505 65252 4509 65308
rect 4445 65248 4509 65252
rect 4525 65308 4589 65312
rect 4525 65252 4529 65308
rect 4529 65252 4585 65308
rect 4585 65252 4589 65308
rect 4525 65248 4589 65252
rect 10952 65308 11016 65312
rect 10952 65252 10956 65308
rect 10956 65252 11012 65308
rect 11012 65252 11016 65308
rect 10952 65248 11016 65252
rect 11032 65308 11096 65312
rect 11032 65252 11036 65308
rect 11036 65252 11092 65308
rect 11092 65252 11096 65308
rect 11032 65248 11096 65252
rect 11112 65308 11176 65312
rect 11112 65252 11116 65308
rect 11116 65252 11172 65308
rect 11172 65252 11176 65308
rect 11112 65248 11176 65252
rect 11192 65308 11256 65312
rect 11192 65252 11196 65308
rect 11196 65252 11252 65308
rect 11252 65252 11256 65308
rect 11192 65248 11256 65252
rect 17618 65308 17682 65312
rect 17618 65252 17622 65308
rect 17622 65252 17678 65308
rect 17678 65252 17682 65308
rect 17618 65248 17682 65252
rect 17698 65308 17762 65312
rect 17698 65252 17702 65308
rect 17702 65252 17758 65308
rect 17758 65252 17762 65308
rect 17698 65248 17762 65252
rect 17778 65308 17842 65312
rect 17778 65252 17782 65308
rect 17782 65252 17838 65308
rect 17838 65252 17842 65308
rect 17778 65248 17842 65252
rect 17858 65308 17922 65312
rect 17858 65252 17862 65308
rect 17862 65252 17918 65308
rect 17918 65252 17922 65308
rect 17858 65248 17922 65252
rect 10548 65180 10612 65244
rect 7618 64764 7682 64768
rect 7618 64708 7622 64764
rect 7622 64708 7678 64764
rect 7678 64708 7682 64764
rect 7618 64704 7682 64708
rect 7698 64764 7762 64768
rect 7698 64708 7702 64764
rect 7702 64708 7758 64764
rect 7758 64708 7762 64764
rect 7698 64704 7762 64708
rect 7778 64764 7842 64768
rect 7778 64708 7782 64764
rect 7782 64708 7838 64764
rect 7838 64708 7842 64764
rect 7778 64704 7842 64708
rect 7858 64764 7922 64768
rect 7858 64708 7862 64764
rect 7862 64708 7918 64764
rect 7918 64708 7922 64764
rect 7858 64704 7922 64708
rect 14285 64764 14349 64768
rect 14285 64708 14289 64764
rect 14289 64708 14345 64764
rect 14345 64708 14349 64764
rect 14285 64704 14349 64708
rect 14365 64764 14429 64768
rect 14365 64708 14369 64764
rect 14369 64708 14425 64764
rect 14425 64708 14429 64764
rect 14365 64704 14429 64708
rect 14445 64764 14509 64768
rect 14445 64708 14449 64764
rect 14449 64708 14505 64764
rect 14505 64708 14509 64764
rect 14445 64704 14509 64708
rect 14525 64764 14589 64768
rect 14525 64708 14529 64764
rect 14529 64708 14585 64764
rect 14585 64708 14589 64764
rect 14525 64704 14589 64708
rect 7420 64500 7484 64564
rect 4285 64220 4349 64224
rect 4285 64164 4289 64220
rect 4289 64164 4345 64220
rect 4345 64164 4349 64220
rect 4285 64160 4349 64164
rect 4365 64220 4429 64224
rect 4365 64164 4369 64220
rect 4369 64164 4425 64220
rect 4425 64164 4429 64220
rect 4365 64160 4429 64164
rect 4445 64220 4509 64224
rect 4445 64164 4449 64220
rect 4449 64164 4505 64220
rect 4505 64164 4509 64220
rect 4445 64160 4509 64164
rect 4525 64220 4589 64224
rect 4525 64164 4529 64220
rect 4529 64164 4585 64220
rect 4585 64164 4589 64220
rect 4525 64160 4589 64164
rect 10952 64220 11016 64224
rect 10952 64164 10956 64220
rect 10956 64164 11012 64220
rect 11012 64164 11016 64220
rect 10952 64160 11016 64164
rect 11032 64220 11096 64224
rect 11032 64164 11036 64220
rect 11036 64164 11092 64220
rect 11092 64164 11096 64220
rect 11032 64160 11096 64164
rect 11112 64220 11176 64224
rect 11112 64164 11116 64220
rect 11116 64164 11172 64220
rect 11172 64164 11176 64220
rect 11112 64160 11176 64164
rect 11192 64220 11256 64224
rect 11192 64164 11196 64220
rect 11196 64164 11252 64220
rect 11252 64164 11256 64220
rect 11192 64160 11256 64164
rect 17618 64220 17682 64224
rect 17618 64164 17622 64220
rect 17622 64164 17678 64220
rect 17678 64164 17682 64220
rect 17618 64160 17682 64164
rect 17698 64220 17762 64224
rect 17698 64164 17702 64220
rect 17702 64164 17758 64220
rect 17758 64164 17762 64220
rect 17698 64160 17762 64164
rect 17778 64220 17842 64224
rect 17778 64164 17782 64220
rect 17782 64164 17838 64220
rect 17838 64164 17842 64220
rect 17778 64160 17842 64164
rect 17858 64220 17922 64224
rect 17858 64164 17862 64220
rect 17862 64164 17918 64220
rect 17918 64164 17922 64220
rect 17858 64160 17922 64164
rect 9812 63956 9876 64020
rect 7052 63548 7116 63612
rect 7618 63676 7682 63680
rect 7618 63620 7622 63676
rect 7622 63620 7678 63676
rect 7678 63620 7682 63676
rect 7618 63616 7682 63620
rect 7698 63676 7762 63680
rect 7698 63620 7702 63676
rect 7702 63620 7758 63676
rect 7758 63620 7762 63676
rect 7698 63616 7762 63620
rect 7778 63676 7842 63680
rect 7778 63620 7782 63676
rect 7782 63620 7838 63676
rect 7838 63620 7842 63676
rect 7778 63616 7842 63620
rect 7858 63676 7922 63680
rect 7858 63620 7862 63676
rect 7862 63620 7918 63676
rect 7918 63620 7922 63676
rect 7858 63616 7922 63620
rect 14285 63676 14349 63680
rect 14285 63620 14289 63676
rect 14289 63620 14345 63676
rect 14345 63620 14349 63676
rect 14285 63616 14349 63620
rect 14365 63676 14429 63680
rect 14365 63620 14369 63676
rect 14369 63620 14425 63676
rect 14425 63620 14429 63676
rect 14365 63616 14429 63620
rect 14445 63676 14509 63680
rect 14445 63620 14449 63676
rect 14449 63620 14505 63676
rect 14505 63620 14509 63676
rect 14445 63616 14509 63620
rect 14525 63676 14589 63680
rect 14525 63620 14529 63676
rect 14529 63620 14585 63676
rect 14585 63620 14589 63676
rect 14525 63616 14589 63620
rect 4285 63132 4349 63136
rect 4285 63076 4289 63132
rect 4289 63076 4345 63132
rect 4345 63076 4349 63132
rect 4285 63072 4349 63076
rect 4365 63132 4429 63136
rect 4365 63076 4369 63132
rect 4369 63076 4425 63132
rect 4425 63076 4429 63132
rect 4365 63072 4429 63076
rect 4445 63132 4509 63136
rect 4445 63076 4449 63132
rect 4449 63076 4505 63132
rect 4505 63076 4509 63132
rect 4445 63072 4509 63076
rect 4525 63132 4589 63136
rect 4525 63076 4529 63132
rect 4529 63076 4585 63132
rect 4585 63076 4589 63132
rect 4525 63072 4589 63076
rect 10952 63132 11016 63136
rect 10952 63076 10956 63132
rect 10956 63076 11012 63132
rect 11012 63076 11016 63132
rect 10952 63072 11016 63076
rect 11032 63132 11096 63136
rect 11032 63076 11036 63132
rect 11036 63076 11092 63132
rect 11092 63076 11096 63132
rect 11032 63072 11096 63076
rect 11112 63132 11176 63136
rect 11112 63076 11116 63132
rect 11116 63076 11172 63132
rect 11172 63076 11176 63132
rect 11112 63072 11176 63076
rect 11192 63132 11256 63136
rect 11192 63076 11196 63132
rect 11196 63076 11252 63132
rect 11252 63076 11256 63132
rect 11192 63072 11256 63076
rect 17618 63132 17682 63136
rect 17618 63076 17622 63132
rect 17622 63076 17678 63132
rect 17678 63076 17682 63132
rect 17618 63072 17682 63076
rect 17698 63132 17762 63136
rect 17698 63076 17702 63132
rect 17702 63076 17758 63132
rect 17758 63076 17762 63132
rect 17698 63072 17762 63076
rect 17778 63132 17842 63136
rect 17778 63076 17782 63132
rect 17782 63076 17838 63132
rect 17838 63076 17842 63132
rect 17778 63072 17842 63076
rect 17858 63132 17922 63136
rect 17858 63076 17862 63132
rect 17862 63076 17918 63132
rect 17918 63076 17922 63132
rect 17858 63072 17922 63076
rect 7236 63004 7300 63068
rect 8340 63004 8404 63068
rect 3372 62868 3436 62932
rect 7618 62588 7682 62592
rect 7618 62532 7622 62588
rect 7622 62532 7678 62588
rect 7678 62532 7682 62588
rect 7618 62528 7682 62532
rect 7698 62588 7762 62592
rect 7698 62532 7702 62588
rect 7702 62532 7758 62588
rect 7758 62532 7762 62588
rect 7698 62528 7762 62532
rect 7778 62588 7842 62592
rect 7778 62532 7782 62588
rect 7782 62532 7838 62588
rect 7838 62532 7842 62588
rect 7778 62528 7842 62532
rect 7858 62588 7922 62592
rect 7858 62532 7862 62588
rect 7862 62532 7918 62588
rect 7918 62532 7922 62588
rect 7858 62528 7922 62532
rect 14285 62588 14349 62592
rect 14285 62532 14289 62588
rect 14289 62532 14345 62588
rect 14345 62532 14349 62588
rect 14285 62528 14349 62532
rect 14365 62588 14429 62592
rect 14365 62532 14369 62588
rect 14369 62532 14425 62588
rect 14425 62532 14429 62588
rect 14365 62528 14429 62532
rect 14445 62588 14509 62592
rect 14445 62532 14449 62588
rect 14449 62532 14505 62588
rect 14505 62532 14509 62588
rect 14445 62528 14509 62532
rect 14525 62588 14589 62592
rect 14525 62532 14529 62588
rect 14529 62532 14585 62588
rect 14585 62532 14589 62588
rect 14525 62528 14589 62532
rect 12020 62324 12084 62388
rect 9996 62188 10060 62252
rect 12204 62188 12268 62252
rect 10180 62052 10244 62116
rect 4285 62044 4349 62048
rect 4285 61988 4289 62044
rect 4289 61988 4345 62044
rect 4345 61988 4349 62044
rect 4285 61984 4349 61988
rect 4365 62044 4429 62048
rect 4365 61988 4369 62044
rect 4369 61988 4425 62044
rect 4425 61988 4429 62044
rect 4365 61984 4429 61988
rect 4445 62044 4509 62048
rect 4445 61988 4449 62044
rect 4449 61988 4505 62044
rect 4505 61988 4509 62044
rect 4445 61984 4509 61988
rect 4525 62044 4589 62048
rect 4525 61988 4529 62044
rect 4529 61988 4585 62044
rect 4585 61988 4589 62044
rect 4525 61984 4589 61988
rect 10952 62044 11016 62048
rect 10952 61988 10956 62044
rect 10956 61988 11012 62044
rect 11012 61988 11016 62044
rect 10952 61984 11016 61988
rect 11032 62044 11096 62048
rect 11032 61988 11036 62044
rect 11036 61988 11092 62044
rect 11092 61988 11096 62044
rect 11032 61984 11096 61988
rect 11112 62044 11176 62048
rect 11112 61988 11116 62044
rect 11116 61988 11172 62044
rect 11172 61988 11176 62044
rect 11112 61984 11176 61988
rect 11192 62044 11256 62048
rect 11192 61988 11196 62044
rect 11196 61988 11252 62044
rect 11252 61988 11256 62044
rect 11192 61984 11256 61988
rect 17618 62044 17682 62048
rect 17618 61988 17622 62044
rect 17622 61988 17678 62044
rect 17678 61988 17682 62044
rect 17618 61984 17682 61988
rect 17698 62044 17762 62048
rect 17698 61988 17702 62044
rect 17702 61988 17758 62044
rect 17758 61988 17762 62044
rect 17698 61984 17762 61988
rect 17778 62044 17842 62048
rect 17778 61988 17782 62044
rect 17782 61988 17838 62044
rect 17838 61988 17842 62044
rect 17778 61984 17842 61988
rect 17858 62044 17922 62048
rect 17858 61988 17862 62044
rect 17862 61988 17918 62044
rect 17918 61988 17922 62044
rect 17858 61984 17922 61988
rect 7618 61500 7682 61504
rect 7618 61444 7622 61500
rect 7622 61444 7678 61500
rect 7678 61444 7682 61500
rect 7618 61440 7682 61444
rect 7698 61500 7762 61504
rect 7698 61444 7702 61500
rect 7702 61444 7758 61500
rect 7758 61444 7762 61500
rect 7698 61440 7762 61444
rect 7778 61500 7842 61504
rect 7778 61444 7782 61500
rect 7782 61444 7838 61500
rect 7838 61444 7842 61500
rect 7778 61440 7842 61444
rect 7858 61500 7922 61504
rect 7858 61444 7862 61500
rect 7862 61444 7918 61500
rect 7918 61444 7922 61500
rect 7858 61440 7922 61444
rect 14285 61500 14349 61504
rect 14285 61444 14289 61500
rect 14289 61444 14345 61500
rect 14345 61444 14349 61500
rect 14285 61440 14349 61444
rect 14365 61500 14429 61504
rect 14365 61444 14369 61500
rect 14369 61444 14425 61500
rect 14425 61444 14429 61500
rect 14365 61440 14429 61444
rect 14445 61500 14509 61504
rect 14445 61444 14449 61500
rect 14449 61444 14505 61500
rect 14505 61444 14509 61500
rect 14445 61440 14509 61444
rect 14525 61500 14589 61504
rect 14525 61444 14529 61500
rect 14529 61444 14585 61500
rect 14585 61444 14589 61500
rect 14525 61440 14589 61444
rect 10548 61236 10612 61300
rect 14780 61236 14844 61300
rect 15332 61236 15396 61300
rect 10548 61100 10612 61164
rect 14044 60964 14108 61028
rect 4285 60956 4349 60960
rect 4285 60900 4289 60956
rect 4289 60900 4345 60956
rect 4345 60900 4349 60956
rect 4285 60896 4349 60900
rect 4365 60956 4429 60960
rect 4365 60900 4369 60956
rect 4369 60900 4425 60956
rect 4425 60900 4429 60956
rect 4365 60896 4429 60900
rect 4445 60956 4509 60960
rect 4445 60900 4449 60956
rect 4449 60900 4505 60956
rect 4505 60900 4509 60956
rect 4445 60896 4509 60900
rect 4525 60956 4589 60960
rect 4525 60900 4529 60956
rect 4529 60900 4585 60956
rect 4585 60900 4589 60956
rect 4525 60896 4589 60900
rect 10952 60956 11016 60960
rect 10952 60900 10956 60956
rect 10956 60900 11012 60956
rect 11012 60900 11016 60956
rect 10952 60896 11016 60900
rect 11032 60956 11096 60960
rect 11032 60900 11036 60956
rect 11036 60900 11092 60956
rect 11092 60900 11096 60956
rect 11032 60896 11096 60900
rect 11112 60956 11176 60960
rect 11112 60900 11116 60956
rect 11116 60900 11172 60956
rect 11172 60900 11176 60956
rect 11112 60896 11176 60900
rect 11192 60956 11256 60960
rect 11192 60900 11196 60956
rect 11196 60900 11252 60956
rect 11252 60900 11256 60956
rect 11192 60896 11256 60900
rect 17618 60956 17682 60960
rect 17618 60900 17622 60956
rect 17622 60900 17678 60956
rect 17678 60900 17682 60956
rect 17618 60896 17682 60900
rect 17698 60956 17762 60960
rect 17698 60900 17702 60956
rect 17702 60900 17758 60956
rect 17758 60900 17762 60956
rect 17698 60896 17762 60900
rect 17778 60956 17842 60960
rect 17778 60900 17782 60956
rect 17782 60900 17838 60956
rect 17838 60900 17842 60956
rect 17778 60896 17842 60900
rect 17858 60956 17922 60960
rect 17858 60900 17862 60956
rect 17862 60900 17918 60956
rect 17918 60900 17922 60956
rect 17858 60896 17922 60900
rect 3372 60616 3436 60620
rect 3372 60560 3386 60616
rect 3386 60560 3436 60616
rect 3372 60556 3436 60560
rect 9812 60692 9876 60756
rect 14044 60752 14108 60756
rect 14044 60696 14094 60752
rect 14094 60696 14108 60752
rect 14044 60692 14108 60696
rect 14780 60752 14844 60756
rect 14780 60696 14794 60752
rect 14794 60696 14844 60752
rect 14780 60692 14844 60696
rect 7618 60412 7682 60416
rect 7618 60356 7622 60412
rect 7622 60356 7678 60412
rect 7678 60356 7682 60412
rect 7618 60352 7682 60356
rect 7698 60412 7762 60416
rect 7698 60356 7702 60412
rect 7702 60356 7758 60412
rect 7758 60356 7762 60412
rect 7698 60352 7762 60356
rect 7778 60412 7842 60416
rect 7778 60356 7782 60412
rect 7782 60356 7838 60412
rect 7838 60356 7842 60412
rect 7778 60352 7842 60356
rect 7858 60412 7922 60416
rect 7858 60356 7862 60412
rect 7862 60356 7918 60412
rect 7918 60356 7922 60412
rect 7858 60352 7922 60356
rect 14285 60412 14349 60416
rect 14285 60356 14289 60412
rect 14289 60356 14345 60412
rect 14345 60356 14349 60412
rect 14285 60352 14349 60356
rect 14365 60412 14429 60416
rect 14365 60356 14369 60412
rect 14369 60356 14425 60412
rect 14425 60356 14429 60412
rect 14365 60352 14429 60356
rect 14445 60412 14509 60416
rect 14445 60356 14449 60412
rect 14449 60356 14505 60412
rect 14505 60356 14509 60412
rect 14445 60352 14509 60356
rect 14525 60412 14589 60416
rect 14525 60356 14529 60412
rect 14529 60356 14585 60412
rect 14585 60356 14589 60412
rect 14525 60352 14589 60356
rect 9260 60012 9324 60076
rect 4285 59868 4349 59872
rect 4285 59812 4289 59868
rect 4289 59812 4345 59868
rect 4345 59812 4349 59868
rect 4285 59808 4349 59812
rect 4365 59868 4429 59872
rect 4365 59812 4369 59868
rect 4369 59812 4425 59868
rect 4425 59812 4429 59868
rect 4365 59808 4429 59812
rect 4445 59868 4509 59872
rect 4445 59812 4449 59868
rect 4449 59812 4505 59868
rect 4505 59812 4509 59868
rect 4445 59808 4509 59812
rect 4525 59868 4589 59872
rect 4525 59812 4529 59868
rect 4529 59812 4585 59868
rect 4585 59812 4589 59868
rect 4525 59808 4589 59812
rect 10952 59868 11016 59872
rect 10952 59812 10956 59868
rect 10956 59812 11012 59868
rect 11012 59812 11016 59868
rect 10952 59808 11016 59812
rect 11032 59868 11096 59872
rect 11032 59812 11036 59868
rect 11036 59812 11092 59868
rect 11092 59812 11096 59868
rect 11032 59808 11096 59812
rect 11112 59868 11176 59872
rect 11112 59812 11116 59868
rect 11116 59812 11172 59868
rect 11172 59812 11176 59868
rect 11112 59808 11176 59812
rect 11192 59868 11256 59872
rect 11192 59812 11196 59868
rect 11196 59812 11252 59868
rect 11252 59812 11256 59868
rect 11192 59808 11256 59812
rect 17618 59868 17682 59872
rect 17618 59812 17622 59868
rect 17622 59812 17678 59868
rect 17678 59812 17682 59868
rect 17618 59808 17682 59812
rect 17698 59868 17762 59872
rect 17698 59812 17702 59868
rect 17702 59812 17758 59868
rect 17758 59812 17762 59868
rect 17698 59808 17762 59812
rect 17778 59868 17842 59872
rect 17778 59812 17782 59868
rect 17782 59812 17838 59868
rect 17838 59812 17842 59868
rect 17778 59808 17842 59812
rect 17858 59868 17922 59872
rect 17858 59812 17862 59868
rect 17862 59812 17918 59868
rect 17918 59812 17922 59868
rect 17858 59808 17922 59812
rect 3372 59392 3436 59396
rect 3372 59336 3422 59392
rect 3422 59336 3436 59392
rect 3372 59332 3436 59336
rect 7618 59324 7682 59328
rect 7618 59268 7622 59324
rect 7622 59268 7678 59324
rect 7678 59268 7682 59324
rect 7618 59264 7682 59268
rect 7698 59324 7762 59328
rect 7698 59268 7702 59324
rect 7702 59268 7758 59324
rect 7758 59268 7762 59324
rect 7698 59264 7762 59268
rect 7778 59324 7842 59328
rect 7778 59268 7782 59324
rect 7782 59268 7838 59324
rect 7838 59268 7842 59324
rect 7778 59264 7842 59268
rect 7858 59324 7922 59328
rect 7858 59268 7862 59324
rect 7862 59268 7918 59324
rect 7918 59268 7922 59324
rect 7858 59264 7922 59268
rect 7236 58924 7300 58988
rect 4285 58780 4349 58784
rect 4285 58724 4289 58780
rect 4289 58724 4345 58780
rect 4345 58724 4349 58780
rect 4285 58720 4349 58724
rect 4365 58780 4429 58784
rect 4365 58724 4369 58780
rect 4369 58724 4425 58780
rect 4425 58724 4429 58780
rect 4365 58720 4429 58724
rect 4445 58780 4509 58784
rect 4445 58724 4449 58780
rect 4449 58724 4505 58780
rect 4505 58724 4509 58780
rect 4445 58720 4509 58724
rect 4525 58780 4589 58784
rect 4525 58724 4529 58780
rect 4529 58724 4585 58780
rect 4585 58724 4589 58780
rect 4525 58720 4589 58724
rect 3556 58652 3620 58716
rect 14285 59324 14349 59328
rect 14285 59268 14289 59324
rect 14289 59268 14345 59324
rect 14345 59268 14349 59324
rect 14285 59264 14349 59268
rect 14365 59324 14429 59328
rect 14365 59268 14369 59324
rect 14369 59268 14425 59324
rect 14425 59268 14429 59324
rect 14365 59264 14429 59268
rect 14445 59324 14509 59328
rect 14445 59268 14449 59324
rect 14449 59268 14505 59324
rect 14505 59268 14509 59324
rect 14445 59264 14509 59268
rect 14525 59324 14589 59328
rect 14525 59268 14529 59324
rect 14529 59268 14585 59324
rect 14585 59268 14589 59324
rect 14525 59264 14589 59268
rect 10952 58780 11016 58784
rect 10952 58724 10956 58780
rect 10956 58724 11012 58780
rect 11012 58724 11016 58780
rect 10952 58720 11016 58724
rect 11032 58780 11096 58784
rect 11032 58724 11036 58780
rect 11036 58724 11092 58780
rect 11092 58724 11096 58780
rect 11032 58720 11096 58724
rect 11112 58780 11176 58784
rect 11112 58724 11116 58780
rect 11116 58724 11172 58780
rect 11172 58724 11176 58780
rect 11112 58720 11176 58724
rect 11192 58780 11256 58784
rect 11192 58724 11196 58780
rect 11196 58724 11252 58780
rect 11252 58724 11256 58780
rect 11192 58720 11256 58724
rect 17618 58780 17682 58784
rect 17618 58724 17622 58780
rect 17622 58724 17678 58780
rect 17678 58724 17682 58780
rect 17618 58720 17682 58724
rect 17698 58780 17762 58784
rect 17698 58724 17702 58780
rect 17702 58724 17758 58780
rect 17758 58724 17762 58780
rect 17698 58720 17762 58724
rect 17778 58780 17842 58784
rect 17778 58724 17782 58780
rect 17782 58724 17838 58780
rect 17838 58724 17842 58780
rect 17778 58720 17842 58724
rect 17858 58780 17922 58784
rect 17858 58724 17862 58780
rect 17862 58724 17918 58780
rect 17918 58724 17922 58780
rect 17858 58720 17922 58724
rect 7618 58236 7682 58240
rect 7618 58180 7622 58236
rect 7622 58180 7678 58236
rect 7678 58180 7682 58236
rect 7618 58176 7682 58180
rect 7698 58236 7762 58240
rect 7698 58180 7702 58236
rect 7702 58180 7758 58236
rect 7758 58180 7762 58236
rect 7698 58176 7762 58180
rect 7778 58236 7842 58240
rect 7778 58180 7782 58236
rect 7782 58180 7838 58236
rect 7838 58180 7842 58236
rect 7778 58176 7842 58180
rect 7858 58236 7922 58240
rect 7858 58180 7862 58236
rect 7862 58180 7918 58236
rect 7918 58180 7922 58236
rect 7858 58176 7922 58180
rect 14285 58236 14349 58240
rect 14285 58180 14289 58236
rect 14289 58180 14345 58236
rect 14345 58180 14349 58236
rect 14285 58176 14349 58180
rect 14365 58236 14429 58240
rect 14365 58180 14369 58236
rect 14369 58180 14425 58236
rect 14425 58180 14429 58236
rect 14365 58176 14429 58180
rect 14445 58236 14509 58240
rect 14445 58180 14449 58236
rect 14449 58180 14505 58236
rect 14505 58180 14509 58236
rect 14445 58176 14509 58180
rect 14525 58236 14589 58240
rect 14525 58180 14529 58236
rect 14529 58180 14585 58236
rect 14585 58180 14589 58236
rect 14525 58176 14589 58180
rect 11836 57700 11900 57764
rect 4285 57692 4349 57696
rect 4285 57636 4289 57692
rect 4289 57636 4345 57692
rect 4345 57636 4349 57692
rect 4285 57632 4349 57636
rect 4365 57692 4429 57696
rect 4365 57636 4369 57692
rect 4369 57636 4425 57692
rect 4425 57636 4429 57692
rect 4365 57632 4429 57636
rect 4445 57692 4509 57696
rect 4445 57636 4449 57692
rect 4449 57636 4505 57692
rect 4505 57636 4509 57692
rect 4445 57632 4509 57636
rect 4525 57692 4589 57696
rect 4525 57636 4529 57692
rect 4529 57636 4585 57692
rect 4585 57636 4589 57692
rect 4525 57632 4589 57636
rect 10952 57692 11016 57696
rect 10952 57636 10956 57692
rect 10956 57636 11012 57692
rect 11012 57636 11016 57692
rect 10952 57632 11016 57636
rect 11032 57692 11096 57696
rect 11032 57636 11036 57692
rect 11036 57636 11092 57692
rect 11092 57636 11096 57692
rect 11032 57632 11096 57636
rect 11112 57692 11176 57696
rect 11112 57636 11116 57692
rect 11116 57636 11172 57692
rect 11172 57636 11176 57692
rect 11112 57632 11176 57636
rect 11192 57692 11256 57696
rect 11192 57636 11196 57692
rect 11196 57636 11252 57692
rect 11252 57636 11256 57692
rect 11192 57632 11256 57636
rect 17618 57692 17682 57696
rect 17618 57636 17622 57692
rect 17622 57636 17678 57692
rect 17678 57636 17682 57692
rect 17618 57632 17682 57636
rect 17698 57692 17762 57696
rect 17698 57636 17702 57692
rect 17702 57636 17758 57692
rect 17758 57636 17762 57692
rect 17698 57632 17762 57636
rect 17778 57692 17842 57696
rect 17778 57636 17782 57692
rect 17782 57636 17838 57692
rect 17838 57636 17842 57692
rect 17778 57632 17842 57636
rect 17858 57692 17922 57696
rect 17858 57636 17862 57692
rect 17862 57636 17918 57692
rect 17918 57636 17922 57692
rect 17858 57632 17922 57636
rect 10364 57428 10428 57492
rect 9444 57292 9508 57356
rect 7618 57148 7682 57152
rect 7618 57092 7622 57148
rect 7622 57092 7678 57148
rect 7678 57092 7682 57148
rect 7618 57088 7682 57092
rect 7698 57148 7762 57152
rect 7698 57092 7702 57148
rect 7702 57092 7758 57148
rect 7758 57092 7762 57148
rect 7698 57088 7762 57092
rect 7778 57148 7842 57152
rect 7778 57092 7782 57148
rect 7782 57092 7838 57148
rect 7838 57092 7842 57148
rect 7778 57088 7842 57092
rect 7858 57148 7922 57152
rect 7858 57092 7862 57148
rect 7862 57092 7918 57148
rect 7918 57092 7922 57148
rect 7858 57088 7922 57092
rect 14285 57148 14349 57152
rect 14285 57092 14289 57148
rect 14289 57092 14345 57148
rect 14345 57092 14349 57148
rect 14285 57088 14349 57092
rect 14365 57148 14429 57152
rect 14365 57092 14369 57148
rect 14369 57092 14425 57148
rect 14425 57092 14429 57148
rect 14365 57088 14429 57092
rect 14445 57148 14509 57152
rect 14445 57092 14449 57148
rect 14449 57092 14505 57148
rect 14505 57092 14509 57148
rect 14445 57088 14509 57092
rect 14525 57148 14589 57152
rect 14525 57092 14529 57148
rect 14529 57092 14585 57148
rect 14585 57092 14589 57148
rect 14525 57088 14589 57092
rect 12572 56612 12636 56676
rect 4285 56604 4349 56608
rect 4285 56548 4289 56604
rect 4289 56548 4345 56604
rect 4345 56548 4349 56604
rect 4285 56544 4349 56548
rect 4365 56604 4429 56608
rect 4365 56548 4369 56604
rect 4369 56548 4425 56604
rect 4425 56548 4429 56604
rect 4365 56544 4429 56548
rect 4445 56604 4509 56608
rect 4445 56548 4449 56604
rect 4449 56548 4505 56604
rect 4505 56548 4509 56604
rect 4445 56544 4509 56548
rect 4525 56604 4589 56608
rect 4525 56548 4529 56604
rect 4529 56548 4585 56604
rect 4585 56548 4589 56604
rect 4525 56544 4589 56548
rect 10952 56604 11016 56608
rect 10952 56548 10956 56604
rect 10956 56548 11012 56604
rect 11012 56548 11016 56604
rect 10952 56544 11016 56548
rect 11032 56604 11096 56608
rect 11032 56548 11036 56604
rect 11036 56548 11092 56604
rect 11092 56548 11096 56604
rect 11032 56544 11096 56548
rect 11112 56604 11176 56608
rect 11112 56548 11116 56604
rect 11116 56548 11172 56604
rect 11172 56548 11176 56604
rect 11112 56544 11176 56548
rect 11192 56604 11256 56608
rect 11192 56548 11196 56604
rect 11196 56548 11252 56604
rect 11252 56548 11256 56604
rect 11192 56544 11256 56548
rect 17618 56604 17682 56608
rect 17618 56548 17622 56604
rect 17622 56548 17678 56604
rect 17678 56548 17682 56604
rect 17618 56544 17682 56548
rect 17698 56604 17762 56608
rect 17698 56548 17702 56604
rect 17702 56548 17758 56604
rect 17758 56548 17762 56604
rect 17698 56544 17762 56548
rect 17778 56604 17842 56608
rect 17778 56548 17782 56604
rect 17782 56548 17838 56604
rect 17838 56548 17842 56604
rect 17778 56544 17842 56548
rect 17858 56604 17922 56608
rect 17858 56548 17862 56604
rect 17862 56548 17918 56604
rect 17918 56548 17922 56604
rect 17858 56544 17922 56548
rect 12388 56476 12452 56540
rect 9076 56340 9140 56404
rect 10364 56400 10428 56404
rect 10364 56344 10414 56400
rect 10414 56344 10428 56400
rect 10364 56340 10428 56344
rect 8892 56204 8956 56268
rect 5580 56068 5644 56132
rect 7618 56060 7682 56064
rect 7618 56004 7622 56060
rect 7622 56004 7678 56060
rect 7678 56004 7682 56060
rect 7618 56000 7682 56004
rect 7698 56060 7762 56064
rect 7698 56004 7702 56060
rect 7702 56004 7758 56060
rect 7758 56004 7762 56060
rect 7698 56000 7762 56004
rect 7778 56060 7842 56064
rect 7778 56004 7782 56060
rect 7782 56004 7838 56060
rect 7838 56004 7842 56060
rect 7778 56000 7842 56004
rect 7858 56060 7922 56064
rect 7858 56004 7862 56060
rect 7862 56004 7918 56060
rect 7918 56004 7922 56060
rect 7858 56000 7922 56004
rect 14285 56060 14349 56064
rect 14285 56004 14289 56060
rect 14289 56004 14345 56060
rect 14345 56004 14349 56060
rect 14285 56000 14349 56004
rect 14365 56060 14429 56064
rect 14365 56004 14369 56060
rect 14369 56004 14425 56060
rect 14425 56004 14429 56060
rect 14365 56000 14429 56004
rect 14445 56060 14509 56064
rect 14445 56004 14449 56060
rect 14449 56004 14505 56060
rect 14505 56004 14509 56060
rect 14445 56000 14509 56004
rect 14525 56060 14589 56064
rect 14525 56004 14529 56060
rect 14529 56004 14585 56060
rect 14585 56004 14589 56060
rect 14525 56000 14589 56004
rect 3188 55932 3252 55996
rect 8524 55796 8588 55860
rect 3740 55660 3804 55724
rect 5212 55660 5276 55724
rect 5948 55660 6012 55724
rect 4285 55516 4349 55520
rect 4285 55460 4289 55516
rect 4289 55460 4345 55516
rect 4345 55460 4349 55516
rect 4285 55456 4349 55460
rect 4365 55516 4429 55520
rect 4365 55460 4369 55516
rect 4369 55460 4425 55516
rect 4425 55460 4429 55516
rect 4365 55456 4429 55460
rect 4445 55516 4509 55520
rect 4445 55460 4449 55516
rect 4449 55460 4505 55516
rect 4505 55460 4509 55516
rect 4445 55456 4509 55460
rect 4525 55516 4589 55520
rect 4525 55460 4529 55516
rect 4529 55460 4585 55516
rect 4585 55460 4589 55516
rect 4525 55456 4589 55460
rect 10952 55516 11016 55520
rect 10952 55460 10956 55516
rect 10956 55460 11012 55516
rect 11012 55460 11016 55516
rect 10952 55456 11016 55460
rect 11032 55516 11096 55520
rect 11032 55460 11036 55516
rect 11036 55460 11092 55516
rect 11092 55460 11096 55516
rect 11032 55456 11096 55460
rect 11112 55516 11176 55520
rect 11112 55460 11116 55516
rect 11116 55460 11172 55516
rect 11172 55460 11176 55516
rect 11112 55456 11176 55460
rect 11192 55516 11256 55520
rect 11192 55460 11196 55516
rect 11196 55460 11252 55516
rect 11252 55460 11256 55516
rect 11192 55456 11256 55460
rect 17618 55516 17682 55520
rect 17618 55460 17622 55516
rect 17622 55460 17678 55516
rect 17678 55460 17682 55516
rect 17618 55456 17682 55460
rect 17698 55516 17762 55520
rect 17698 55460 17702 55516
rect 17702 55460 17758 55516
rect 17758 55460 17762 55516
rect 17698 55456 17762 55460
rect 17778 55516 17842 55520
rect 17778 55460 17782 55516
rect 17782 55460 17838 55516
rect 17838 55460 17842 55516
rect 17778 55456 17842 55460
rect 17858 55516 17922 55520
rect 17858 55460 17862 55516
rect 17862 55460 17918 55516
rect 17918 55460 17922 55516
rect 17858 55456 17922 55460
rect 3924 55388 3988 55452
rect 8708 55388 8772 55452
rect 11652 55252 11716 55316
rect 8892 55116 8956 55180
rect 12020 55116 12084 55180
rect 12572 55116 12636 55180
rect 3004 54980 3068 55044
rect 6132 54980 6196 55044
rect 9260 54980 9324 55044
rect 7618 54972 7682 54976
rect 7618 54916 7622 54972
rect 7622 54916 7678 54972
rect 7678 54916 7682 54972
rect 7618 54912 7682 54916
rect 7698 54972 7762 54976
rect 7698 54916 7702 54972
rect 7702 54916 7758 54972
rect 7758 54916 7762 54972
rect 7698 54912 7762 54916
rect 7778 54972 7842 54976
rect 7778 54916 7782 54972
rect 7782 54916 7838 54972
rect 7838 54916 7842 54972
rect 7778 54912 7842 54916
rect 7858 54972 7922 54976
rect 7858 54916 7862 54972
rect 7862 54916 7918 54972
rect 7918 54916 7922 54972
rect 7858 54912 7922 54916
rect 14285 54972 14349 54976
rect 14285 54916 14289 54972
rect 14289 54916 14345 54972
rect 14345 54916 14349 54972
rect 14285 54912 14349 54916
rect 14365 54972 14429 54976
rect 14365 54916 14369 54972
rect 14369 54916 14425 54972
rect 14425 54916 14429 54972
rect 14365 54912 14429 54916
rect 14445 54972 14509 54976
rect 14445 54916 14449 54972
rect 14449 54916 14505 54972
rect 14505 54916 14509 54972
rect 14445 54912 14509 54916
rect 14525 54972 14589 54976
rect 14525 54916 14529 54972
rect 14529 54916 14585 54972
rect 14585 54916 14589 54972
rect 14525 54912 14589 54916
rect 9812 54844 9876 54908
rect 12388 54844 12452 54908
rect 4285 54428 4349 54432
rect 4285 54372 4289 54428
rect 4289 54372 4345 54428
rect 4345 54372 4349 54428
rect 4285 54368 4349 54372
rect 4365 54428 4429 54432
rect 4365 54372 4369 54428
rect 4369 54372 4425 54428
rect 4425 54372 4429 54428
rect 4365 54368 4429 54372
rect 4445 54428 4509 54432
rect 4445 54372 4449 54428
rect 4449 54372 4505 54428
rect 4505 54372 4509 54428
rect 4445 54368 4509 54372
rect 4525 54428 4589 54432
rect 4525 54372 4529 54428
rect 4529 54372 4585 54428
rect 4585 54372 4589 54428
rect 4525 54368 4589 54372
rect 5764 54028 5828 54092
rect 10952 54428 11016 54432
rect 10952 54372 10956 54428
rect 10956 54372 11012 54428
rect 11012 54372 11016 54428
rect 10952 54368 11016 54372
rect 11032 54428 11096 54432
rect 11032 54372 11036 54428
rect 11036 54372 11092 54428
rect 11092 54372 11096 54428
rect 11032 54368 11096 54372
rect 11112 54428 11176 54432
rect 11112 54372 11116 54428
rect 11116 54372 11172 54428
rect 11172 54372 11176 54428
rect 11112 54368 11176 54372
rect 11192 54428 11256 54432
rect 11192 54372 11196 54428
rect 11196 54372 11252 54428
rect 11252 54372 11256 54428
rect 11192 54368 11256 54372
rect 17618 54428 17682 54432
rect 17618 54372 17622 54428
rect 17622 54372 17678 54428
rect 17678 54372 17682 54428
rect 17618 54368 17682 54372
rect 17698 54428 17762 54432
rect 17698 54372 17702 54428
rect 17702 54372 17758 54428
rect 17758 54372 17762 54428
rect 17698 54368 17762 54372
rect 17778 54428 17842 54432
rect 17778 54372 17782 54428
rect 17782 54372 17838 54428
rect 17838 54372 17842 54428
rect 17778 54368 17842 54372
rect 17858 54428 17922 54432
rect 17858 54372 17862 54428
rect 17862 54372 17918 54428
rect 17918 54372 17922 54428
rect 17858 54368 17922 54372
rect 6684 54360 6748 54364
rect 6684 54304 6734 54360
rect 6734 54304 6748 54360
rect 6684 54300 6748 54304
rect 11836 54164 11900 54228
rect 12388 54224 12452 54228
rect 12388 54168 12402 54224
rect 12402 54168 12452 54224
rect 12388 54164 12452 54168
rect 7236 54028 7300 54092
rect 6500 53892 6564 53956
rect 7236 53892 7300 53956
rect 7618 53884 7682 53888
rect 7618 53828 7622 53884
rect 7622 53828 7678 53884
rect 7678 53828 7682 53884
rect 7618 53824 7682 53828
rect 7698 53884 7762 53888
rect 7698 53828 7702 53884
rect 7702 53828 7758 53884
rect 7758 53828 7762 53884
rect 7698 53824 7762 53828
rect 7778 53884 7842 53888
rect 7778 53828 7782 53884
rect 7782 53828 7838 53884
rect 7838 53828 7842 53884
rect 7778 53824 7842 53828
rect 7858 53884 7922 53888
rect 7858 53828 7862 53884
rect 7862 53828 7918 53884
rect 7918 53828 7922 53884
rect 7858 53824 7922 53828
rect 11836 53892 11900 53956
rect 14285 53884 14349 53888
rect 14285 53828 14289 53884
rect 14289 53828 14345 53884
rect 14345 53828 14349 53884
rect 14285 53824 14349 53828
rect 14365 53884 14429 53888
rect 14365 53828 14369 53884
rect 14369 53828 14425 53884
rect 14425 53828 14429 53884
rect 14365 53824 14429 53828
rect 14445 53884 14509 53888
rect 14445 53828 14449 53884
rect 14449 53828 14505 53884
rect 14505 53828 14509 53884
rect 14445 53824 14509 53828
rect 14525 53884 14589 53888
rect 14525 53828 14529 53884
rect 14529 53828 14585 53884
rect 14585 53828 14589 53884
rect 14525 53824 14589 53828
rect 13124 53756 13188 53820
rect 9444 53620 9508 53684
rect 4285 53340 4349 53344
rect 4285 53284 4289 53340
rect 4289 53284 4345 53340
rect 4345 53284 4349 53340
rect 4285 53280 4349 53284
rect 4365 53340 4429 53344
rect 4365 53284 4369 53340
rect 4369 53284 4425 53340
rect 4425 53284 4429 53340
rect 4365 53280 4429 53284
rect 4445 53340 4509 53344
rect 4445 53284 4449 53340
rect 4449 53284 4505 53340
rect 4505 53284 4509 53340
rect 4445 53280 4509 53284
rect 4525 53340 4589 53344
rect 4525 53284 4529 53340
rect 4529 53284 4585 53340
rect 4585 53284 4589 53340
rect 4525 53280 4589 53284
rect 10952 53340 11016 53344
rect 10952 53284 10956 53340
rect 10956 53284 11012 53340
rect 11012 53284 11016 53340
rect 10952 53280 11016 53284
rect 11032 53340 11096 53344
rect 11032 53284 11036 53340
rect 11036 53284 11092 53340
rect 11092 53284 11096 53340
rect 11032 53280 11096 53284
rect 11112 53340 11176 53344
rect 11112 53284 11116 53340
rect 11116 53284 11172 53340
rect 11172 53284 11176 53340
rect 11112 53280 11176 53284
rect 11192 53340 11256 53344
rect 11192 53284 11196 53340
rect 11196 53284 11252 53340
rect 11252 53284 11256 53340
rect 11192 53280 11256 53284
rect 17172 53348 17236 53412
rect 17618 53340 17682 53344
rect 17618 53284 17622 53340
rect 17622 53284 17678 53340
rect 17678 53284 17682 53340
rect 17618 53280 17682 53284
rect 17698 53340 17762 53344
rect 17698 53284 17702 53340
rect 17702 53284 17758 53340
rect 17758 53284 17762 53340
rect 17698 53280 17762 53284
rect 17778 53340 17842 53344
rect 17778 53284 17782 53340
rect 17782 53284 17838 53340
rect 17838 53284 17842 53340
rect 17778 53280 17842 53284
rect 17858 53340 17922 53344
rect 17858 53284 17862 53340
rect 17862 53284 17918 53340
rect 17918 53284 17922 53340
rect 17858 53280 17922 53284
rect 5948 53076 6012 53140
rect 6316 52940 6380 53004
rect 10364 52804 10428 52868
rect 14964 52804 15028 52868
rect 15332 52804 15396 52868
rect 7618 52796 7682 52800
rect 7618 52740 7622 52796
rect 7622 52740 7678 52796
rect 7678 52740 7682 52796
rect 7618 52736 7682 52740
rect 7698 52796 7762 52800
rect 7698 52740 7702 52796
rect 7702 52740 7758 52796
rect 7758 52740 7762 52796
rect 7698 52736 7762 52740
rect 7778 52796 7842 52800
rect 7778 52740 7782 52796
rect 7782 52740 7838 52796
rect 7838 52740 7842 52796
rect 7778 52736 7842 52740
rect 7858 52796 7922 52800
rect 7858 52740 7862 52796
rect 7862 52740 7918 52796
rect 7918 52740 7922 52796
rect 7858 52736 7922 52740
rect 14285 52796 14349 52800
rect 14285 52740 14289 52796
rect 14289 52740 14345 52796
rect 14345 52740 14349 52796
rect 14285 52736 14349 52740
rect 14365 52796 14429 52800
rect 14365 52740 14369 52796
rect 14369 52740 14425 52796
rect 14425 52740 14429 52796
rect 14365 52736 14429 52740
rect 14445 52796 14509 52800
rect 14445 52740 14449 52796
rect 14449 52740 14505 52796
rect 14505 52740 14509 52796
rect 14445 52736 14509 52740
rect 14525 52796 14589 52800
rect 14525 52740 14529 52796
rect 14529 52740 14585 52796
rect 14585 52740 14589 52796
rect 14525 52736 14589 52740
rect 8524 52668 8588 52732
rect 12572 52668 12636 52732
rect 13492 52668 13556 52732
rect 10364 52532 10428 52596
rect 13308 52396 13372 52460
rect 17356 52260 17420 52324
rect 4285 52252 4349 52256
rect 4285 52196 4289 52252
rect 4289 52196 4345 52252
rect 4345 52196 4349 52252
rect 4285 52192 4349 52196
rect 4365 52252 4429 52256
rect 4365 52196 4369 52252
rect 4369 52196 4425 52252
rect 4425 52196 4429 52252
rect 4365 52192 4429 52196
rect 4445 52252 4509 52256
rect 4445 52196 4449 52252
rect 4449 52196 4505 52252
rect 4505 52196 4509 52252
rect 4445 52192 4509 52196
rect 4525 52252 4589 52256
rect 4525 52196 4529 52252
rect 4529 52196 4585 52252
rect 4585 52196 4589 52252
rect 4525 52192 4589 52196
rect 10952 52252 11016 52256
rect 10952 52196 10956 52252
rect 10956 52196 11012 52252
rect 11012 52196 11016 52252
rect 10952 52192 11016 52196
rect 11032 52252 11096 52256
rect 11032 52196 11036 52252
rect 11036 52196 11092 52252
rect 11092 52196 11096 52252
rect 11032 52192 11096 52196
rect 11112 52252 11176 52256
rect 11112 52196 11116 52252
rect 11116 52196 11172 52252
rect 11172 52196 11176 52252
rect 11112 52192 11176 52196
rect 11192 52252 11256 52256
rect 11192 52196 11196 52252
rect 11196 52196 11252 52252
rect 11252 52196 11256 52252
rect 11192 52192 11256 52196
rect 17618 52252 17682 52256
rect 17618 52196 17622 52252
rect 17622 52196 17678 52252
rect 17678 52196 17682 52252
rect 17618 52192 17682 52196
rect 17698 52252 17762 52256
rect 17698 52196 17702 52252
rect 17702 52196 17758 52252
rect 17758 52196 17762 52252
rect 17698 52192 17762 52196
rect 17778 52252 17842 52256
rect 17778 52196 17782 52252
rect 17782 52196 17838 52252
rect 17838 52196 17842 52252
rect 17778 52192 17842 52196
rect 17858 52252 17922 52256
rect 17858 52196 17862 52252
rect 17862 52196 17918 52252
rect 17918 52196 17922 52252
rect 17858 52192 17922 52196
rect 5580 52124 5644 52188
rect 10548 51716 10612 51780
rect 7618 51708 7682 51712
rect 7618 51652 7622 51708
rect 7622 51652 7678 51708
rect 7678 51652 7682 51708
rect 7618 51648 7682 51652
rect 7698 51708 7762 51712
rect 7698 51652 7702 51708
rect 7702 51652 7758 51708
rect 7758 51652 7762 51708
rect 7698 51648 7762 51652
rect 7778 51708 7842 51712
rect 7778 51652 7782 51708
rect 7782 51652 7838 51708
rect 7838 51652 7842 51708
rect 7778 51648 7842 51652
rect 7858 51708 7922 51712
rect 7858 51652 7862 51708
rect 7862 51652 7918 51708
rect 7918 51652 7922 51708
rect 7858 51648 7922 51652
rect 14285 51708 14349 51712
rect 14285 51652 14289 51708
rect 14289 51652 14345 51708
rect 14345 51652 14349 51708
rect 14285 51648 14349 51652
rect 14365 51708 14429 51712
rect 14365 51652 14369 51708
rect 14369 51652 14425 51708
rect 14425 51652 14429 51708
rect 14365 51648 14429 51652
rect 14445 51708 14509 51712
rect 14445 51652 14449 51708
rect 14449 51652 14505 51708
rect 14505 51652 14509 51708
rect 14445 51648 14509 51652
rect 14525 51708 14589 51712
rect 14525 51652 14529 51708
rect 14529 51652 14585 51708
rect 14585 51652 14589 51708
rect 14525 51648 14589 51652
rect 3556 51580 3620 51644
rect 6684 51580 6748 51644
rect 3372 51444 3436 51508
rect 3004 51308 3068 51372
rect 3924 51308 3988 51372
rect 5948 51444 6012 51508
rect 12756 51444 12820 51508
rect 5212 51172 5276 51236
rect 4285 51164 4349 51168
rect 4285 51108 4289 51164
rect 4289 51108 4345 51164
rect 4345 51108 4349 51164
rect 4285 51104 4349 51108
rect 4365 51164 4429 51168
rect 4365 51108 4369 51164
rect 4369 51108 4425 51164
rect 4425 51108 4429 51164
rect 4365 51104 4429 51108
rect 4445 51164 4509 51168
rect 4445 51108 4449 51164
rect 4449 51108 4505 51164
rect 4505 51108 4509 51164
rect 4445 51104 4509 51108
rect 4525 51164 4589 51168
rect 4525 51108 4529 51164
rect 4529 51108 4585 51164
rect 4585 51108 4589 51164
rect 4525 51104 4589 51108
rect 6684 51308 6748 51372
rect 7052 51308 7116 51372
rect 8340 51308 8404 51372
rect 5948 51172 6012 51236
rect 7052 51172 7116 51236
rect 7420 51172 7484 51236
rect 8708 51172 8772 51236
rect 9260 51172 9324 51236
rect 10952 51164 11016 51168
rect 10952 51108 10956 51164
rect 10956 51108 11012 51164
rect 11012 51108 11016 51164
rect 10952 51104 11016 51108
rect 11032 51164 11096 51168
rect 11032 51108 11036 51164
rect 11036 51108 11092 51164
rect 11092 51108 11096 51164
rect 11032 51104 11096 51108
rect 11112 51164 11176 51168
rect 11112 51108 11116 51164
rect 11116 51108 11172 51164
rect 11172 51108 11176 51164
rect 11112 51104 11176 51108
rect 11192 51164 11256 51168
rect 11192 51108 11196 51164
rect 11196 51108 11252 51164
rect 11252 51108 11256 51164
rect 11192 51104 11256 51108
rect 7420 51036 7484 51100
rect 5764 50960 5828 50964
rect 5764 50904 5778 50960
rect 5778 50904 5828 50960
rect 5764 50900 5828 50904
rect 9076 51036 9140 51100
rect 9444 50900 9508 50964
rect 10548 50900 10612 50964
rect 12940 51036 13004 51100
rect 5948 50764 6012 50828
rect 6868 50764 6932 50828
rect 1716 50628 1780 50692
rect 6684 50492 6748 50556
rect 11652 50764 11716 50828
rect 9076 50628 9140 50692
rect 9444 50628 9508 50692
rect 14780 51036 14844 51100
rect 15148 51036 15212 51100
rect 17618 51164 17682 51168
rect 17618 51108 17622 51164
rect 17622 51108 17678 51164
rect 17678 51108 17682 51164
rect 17618 51104 17682 51108
rect 17698 51164 17762 51168
rect 17698 51108 17702 51164
rect 17702 51108 17758 51164
rect 17758 51108 17762 51164
rect 17698 51104 17762 51108
rect 17778 51164 17842 51168
rect 17778 51108 17782 51164
rect 17782 51108 17838 51164
rect 17838 51108 17842 51164
rect 17778 51104 17842 51108
rect 17858 51164 17922 51168
rect 17858 51108 17862 51164
rect 17862 51108 17918 51164
rect 17918 51108 17922 51164
rect 17858 51104 17922 51108
rect 13492 50960 13556 50964
rect 13492 50904 13506 50960
rect 13506 50904 13556 50960
rect 13492 50900 13556 50904
rect 13676 50960 13740 50964
rect 13676 50904 13726 50960
rect 13726 50904 13740 50960
rect 13676 50900 13740 50904
rect 14780 50960 14844 50964
rect 14780 50904 14830 50960
rect 14830 50904 14844 50960
rect 14780 50900 14844 50904
rect 13492 50628 13556 50692
rect 7618 50620 7682 50624
rect 7618 50564 7622 50620
rect 7622 50564 7678 50620
rect 7678 50564 7682 50620
rect 7618 50560 7682 50564
rect 7698 50620 7762 50624
rect 7698 50564 7702 50620
rect 7702 50564 7758 50620
rect 7758 50564 7762 50620
rect 7698 50560 7762 50564
rect 7778 50620 7842 50624
rect 7778 50564 7782 50620
rect 7782 50564 7838 50620
rect 7838 50564 7842 50620
rect 7778 50560 7842 50564
rect 7858 50620 7922 50624
rect 7858 50564 7862 50620
rect 7862 50564 7918 50620
rect 7918 50564 7922 50620
rect 7858 50560 7922 50564
rect 14285 50620 14349 50624
rect 14285 50564 14289 50620
rect 14289 50564 14345 50620
rect 14345 50564 14349 50620
rect 14285 50560 14349 50564
rect 14365 50620 14429 50624
rect 14365 50564 14369 50620
rect 14369 50564 14425 50620
rect 14425 50564 14429 50620
rect 14365 50560 14429 50564
rect 14445 50620 14509 50624
rect 14445 50564 14449 50620
rect 14449 50564 14505 50620
rect 14505 50564 14509 50620
rect 14445 50560 14509 50564
rect 14525 50620 14589 50624
rect 14525 50564 14529 50620
rect 14529 50564 14585 50620
rect 14585 50564 14589 50620
rect 14525 50560 14589 50564
rect 11468 50492 11532 50556
rect 6132 50356 6196 50420
rect 6132 50084 6196 50148
rect 8340 50084 8404 50148
rect 13308 50220 13372 50284
rect 13308 50084 13372 50148
rect 4285 50076 4349 50080
rect 4285 50020 4289 50076
rect 4289 50020 4345 50076
rect 4345 50020 4349 50076
rect 4285 50016 4349 50020
rect 4365 50076 4429 50080
rect 4365 50020 4369 50076
rect 4369 50020 4425 50076
rect 4425 50020 4429 50076
rect 4365 50016 4429 50020
rect 4445 50076 4509 50080
rect 4445 50020 4449 50076
rect 4449 50020 4505 50076
rect 4505 50020 4509 50076
rect 4445 50016 4509 50020
rect 4525 50076 4589 50080
rect 4525 50020 4529 50076
rect 4529 50020 4585 50076
rect 4585 50020 4589 50076
rect 4525 50016 4589 50020
rect 10952 50076 11016 50080
rect 10952 50020 10956 50076
rect 10956 50020 11012 50076
rect 11012 50020 11016 50076
rect 10952 50016 11016 50020
rect 11032 50076 11096 50080
rect 11032 50020 11036 50076
rect 11036 50020 11092 50076
rect 11092 50020 11096 50076
rect 11032 50016 11096 50020
rect 11112 50076 11176 50080
rect 11112 50020 11116 50076
rect 11116 50020 11172 50076
rect 11172 50020 11176 50076
rect 11112 50016 11176 50020
rect 11192 50076 11256 50080
rect 11192 50020 11196 50076
rect 11196 50020 11252 50076
rect 11252 50020 11256 50076
rect 11192 50016 11256 50020
rect 17618 50076 17682 50080
rect 17618 50020 17622 50076
rect 17622 50020 17678 50076
rect 17678 50020 17682 50076
rect 17618 50016 17682 50020
rect 17698 50076 17762 50080
rect 17698 50020 17702 50076
rect 17702 50020 17758 50076
rect 17758 50020 17762 50076
rect 17698 50016 17762 50020
rect 17778 50076 17842 50080
rect 17778 50020 17782 50076
rect 17782 50020 17838 50076
rect 17838 50020 17842 50076
rect 17778 50016 17842 50020
rect 17858 50076 17922 50080
rect 17858 50020 17862 50076
rect 17862 50020 17918 50076
rect 17918 50020 17922 50076
rect 17858 50016 17922 50020
rect 2268 49948 2332 50012
rect 6868 49812 6932 49876
rect 9260 49872 9324 49876
rect 9260 49816 9274 49872
rect 9274 49816 9324 49872
rect 9260 49812 9324 49816
rect 6868 49540 6932 49604
rect 7618 49532 7682 49536
rect 7618 49476 7622 49532
rect 7622 49476 7678 49532
rect 7678 49476 7682 49532
rect 7618 49472 7682 49476
rect 7698 49532 7762 49536
rect 7698 49476 7702 49532
rect 7702 49476 7758 49532
rect 7758 49476 7762 49532
rect 7698 49472 7762 49476
rect 7778 49532 7842 49536
rect 7778 49476 7782 49532
rect 7782 49476 7838 49532
rect 7838 49476 7842 49532
rect 7778 49472 7842 49476
rect 7858 49532 7922 49536
rect 7858 49476 7862 49532
rect 7862 49476 7918 49532
rect 7918 49476 7922 49532
rect 7858 49472 7922 49476
rect 9260 49404 9324 49468
rect 9628 50008 9692 50012
rect 9628 49952 9678 50008
rect 9678 49952 9692 50008
rect 9628 49948 9692 49952
rect 9628 49812 9692 49876
rect 10548 49812 10612 49876
rect 10548 49736 10612 49740
rect 10548 49680 10562 49736
rect 10562 49680 10612 49736
rect 10548 49676 10612 49680
rect 14285 49532 14349 49536
rect 14285 49476 14289 49532
rect 14289 49476 14345 49532
rect 14345 49476 14349 49532
rect 14285 49472 14349 49476
rect 14365 49532 14429 49536
rect 14365 49476 14369 49532
rect 14369 49476 14425 49532
rect 14425 49476 14429 49532
rect 14365 49472 14429 49476
rect 14445 49532 14509 49536
rect 14445 49476 14449 49532
rect 14449 49476 14505 49532
rect 14505 49476 14509 49532
rect 14445 49472 14509 49476
rect 14525 49532 14589 49536
rect 14525 49476 14529 49532
rect 14529 49476 14585 49532
rect 14585 49476 14589 49532
rect 14525 49472 14589 49476
rect 12572 49268 12636 49332
rect 5396 49132 5460 49196
rect 8892 49132 8956 49196
rect 13124 49132 13188 49196
rect 13492 49132 13556 49196
rect 4285 48988 4349 48992
rect 4285 48932 4289 48988
rect 4289 48932 4345 48988
rect 4345 48932 4349 48988
rect 4285 48928 4349 48932
rect 4365 48988 4429 48992
rect 4365 48932 4369 48988
rect 4369 48932 4425 48988
rect 4425 48932 4429 48988
rect 4365 48928 4429 48932
rect 4445 48988 4509 48992
rect 4445 48932 4449 48988
rect 4449 48932 4505 48988
rect 4505 48932 4509 48988
rect 4445 48928 4509 48932
rect 4525 48988 4589 48992
rect 4525 48932 4529 48988
rect 4529 48932 4585 48988
rect 4585 48932 4589 48988
rect 4525 48928 4589 48932
rect 10952 48988 11016 48992
rect 10952 48932 10956 48988
rect 10956 48932 11012 48988
rect 11012 48932 11016 48988
rect 10952 48928 11016 48932
rect 11032 48988 11096 48992
rect 11032 48932 11036 48988
rect 11036 48932 11092 48988
rect 11092 48932 11096 48988
rect 11032 48928 11096 48932
rect 11112 48988 11176 48992
rect 11112 48932 11116 48988
rect 11116 48932 11172 48988
rect 11172 48932 11176 48988
rect 11112 48928 11176 48932
rect 11192 48988 11256 48992
rect 11192 48932 11196 48988
rect 11196 48932 11252 48988
rect 11252 48932 11256 48988
rect 11192 48928 11256 48932
rect 17618 48988 17682 48992
rect 17618 48932 17622 48988
rect 17622 48932 17678 48988
rect 17678 48932 17682 48988
rect 17618 48928 17682 48932
rect 17698 48988 17762 48992
rect 17698 48932 17702 48988
rect 17702 48932 17758 48988
rect 17758 48932 17762 48988
rect 17698 48928 17762 48932
rect 17778 48988 17842 48992
rect 17778 48932 17782 48988
rect 17782 48932 17838 48988
rect 17838 48932 17842 48988
rect 17778 48928 17842 48932
rect 17858 48988 17922 48992
rect 17858 48932 17862 48988
rect 17862 48932 17918 48988
rect 17918 48932 17922 48988
rect 17858 48928 17922 48932
rect 5396 48860 5460 48924
rect 12756 48724 12820 48788
rect 7618 48444 7682 48448
rect 7618 48388 7622 48444
rect 7622 48388 7678 48444
rect 7678 48388 7682 48444
rect 7618 48384 7682 48388
rect 7698 48444 7762 48448
rect 7698 48388 7702 48444
rect 7702 48388 7758 48444
rect 7758 48388 7762 48444
rect 7698 48384 7762 48388
rect 7778 48444 7842 48448
rect 7778 48388 7782 48444
rect 7782 48388 7838 48444
rect 7838 48388 7842 48444
rect 7778 48384 7842 48388
rect 7858 48444 7922 48448
rect 7858 48388 7862 48444
rect 7862 48388 7918 48444
rect 7918 48388 7922 48444
rect 7858 48384 7922 48388
rect 14285 48444 14349 48448
rect 14285 48388 14289 48444
rect 14289 48388 14345 48444
rect 14345 48388 14349 48444
rect 14285 48384 14349 48388
rect 14365 48444 14429 48448
rect 14365 48388 14369 48444
rect 14369 48388 14425 48444
rect 14425 48388 14429 48444
rect 14365 48384 14429 48388
rect 14445 48444 14509 48448
rect 14445 48388 14449 48444
rect 14449 48388 14505 48444
rect 14505 48388 14509 48444
rect 14445 48384 14509 48388
rect 14525 48444 14589 48448
rect 14525 48388 14529 48444
rect 14529 48388 14585 48444
rect 14585 48388 14589 48444
rect 14525 48384 14589 48388
rect 5764 48316 5828 48380
rect 8708 48316 8772 48380
rect 3740 48180 3804 48244
rect 12940 48316 13004 48380
rect 4285 47900 4349 47904
rect 4285 47844 4289 47900
rect 4289 47844 4345 47900
rect 4345 47844 4349 47900
rect 4285 47840 4349 47844
rect 4365 47900 4429 47904
rect 4365 47844 4369 47900
rect 4369 47844 4425 47900
rect 4425 47844 4429 47900
rect 4365 47840 4429 47844
rect 4445 47900 4509 47904
rect 4445 47844 4449 47900
rect 4449 47844 4505 47900
rect 4505 47844 4509 47900
rect 4445 47840 4509 47844
rect 4525 47900 4589 47904
rect 4525 47844 4529 47900
rect 4529 47844 4585 47900
rect 4585 47844 4589 47900
rect 4525 47840 4589 47844
rect 10952 47900 11016 47904
rect 10952 47844 10956 47900
rect 10956 47844 11012 47900
rect 11012 47844 11016 47900
rect 10952 47840 11016 47844
rect 11032 47900 11096 47904
rect 11032 47844 11036 47900
rect 11036 47844 11092 47900
rect 11092 47844 11096 47900
rect 11032 47840 11096 47844
rect 11112 47900 11176 47904
rect 11112 47844 11116 47900
rect 11116 47844 11172 47900
rect 11172 47844 11176 47900
rect 11112 47840 11176 47844
rect 11192 47900 11256 47904
rect 11192 47844 11196 47900
rect 11196 47844 11252 47900
rect 11252 47844 11256 47900
rect 11192 47840 11256 47844
rect 17618 47900 17682 47904
rect 17618 47844 17622 47900
rect 17622 47844 17678 47900
rect 17678 47844 17682 47900
rect 17618 47840 17682 47844
rect 17698 47900 17762 47904
rect 17698 47844 17702 47900
rect 17702 47844 17758 47900
rect 17758 47844 17762 47900
rect 17698 47840 17762 47844
rect 17778 47900 17842 47904
rect 17778 47844 17782 47900
rect 17782 47844 17838 47900
rect 17838 47844 17842 47900
rect 17778 47840 17842 47844
rect 17858 47900 17922 47904
rect 17858 47844 17862 47900
rect 17862 47844 17918 47900
rect 17918 47844 17922 47900
rect 17858 47840 17922 47844
rect 6684 47772 6748 47836
rect 6316 47636 6380 47700
rect 12388 47636 12452 47700
rect 3924 47500 3988 47564
rect 12756 47364 12820 47428
rect 7618 47356 7682 47360
rect 7618 47300 7622 47356
rect 7622 47300 7678 47356
rect 7678 47300 7682 47356
rect 7618 47296 7682 47300
rect 7698 47356 7762 47360
rect 7698 47300 7702 47356
rect 7702 47300 7758 47356
rect 7758 47300 7762 47356
rect 7698 47296 7762 47300
rect 7778 47356 7842 47360
rect 7778 47300 7782 47356
rect 7782 47300 7838 47356
rect 7838 47300 7842 47356
rect 7778 47296 7842 47300
rect 7858 47356 7922 47360
rect 7858 47300 7862 47356
rect 7862 47300 7918 47356
rect 7918 47300 7922 47356
rect 7858 47296 7922 47300
rect 14285 47356 14349 47360
rect 14285 47300 14289 47356
rect 14289 47300 14345 47356
rect 14345 47300 14349 47356
rect 14285 47296 14349 47300
rect 14365 47356 14429 47360
rect 14365 47300 14369 47356
rect 14369 47300 14425 47356
rect 14425 47300 14429 47356
rect 14365 47296 14429 47300
rect 14445 47356 14509 47360
rect 14445 47300 14449 47356
rect 14449 47300 14505 47356
rect 14505 47300 14509 47356
rect 14445 47296 14509 47300
rect 14525 47356 14589 47360
rect 14525 47300 14529 47356
rect 14529 47300 14585 47356
rect 14585 47300 14589 47356
rect 14525 47296 14589 47300
rect 12572 47228 12636 47292
rect 6500 46956 6564 47020
rect 8340 46880 8404 46884
rect 8340 46824 8390 46880
rect 8390 46824 8404 46880
rect 8340 46820 8404 46824
rect 4285 46812 4349 46816
rect 4285 46756 4289 46812
rect 4289 46756 4345 46812
rect 4345 46756 4349 46812
rect 4285 46752 4349 46756
rect 4365 46812 4429 46816
rect 4365 46756 4369 46812
rect 4369 46756 4425 46812
rect 4425 46756 4429 46812
rect 4365 46752 4429 46756
rect 4445 46812 4509 46816
rect 4445 46756 4449 46812
rect 4449 46756 4505 46812
rect 4505 46756 4509 46812
rect 4445 46752 4509 46756
rect 4525 46812 4589 46816
rect 4525 46756 4529 46812
rect 4529 46756 4585 46812
rect 4585 46756 4589 46812
rect 4525 46752 4589 46756
rect 10952 46812 11016 46816
rect 10952 46756 10956 46812
rect 10956 46756 11012 46812
rect 11012 46756 11016 46812
rect 10952 46752 11016 46756
rect 11032 46812 11096 46816
rect 11032 46756 11036 46812
rect 11036 46756 11092 46812
rect 11092 46756 11096 46812
rect 11032 46752 11096 46756
rect 11112 46812 11176 46816
rect 11112 46756 11116 46812
rect 11116 46756 11172 46812
rect 11172 46756 11176 46812
rect 11112 46752 11176 46756
rect 11192 46812 11256 46816
rect 11192 46756 11196 46812
rect 11196 46756 11252 46812
rect 11252 46756 11256 46812
rect 11192 46752 11256 46756
rect 17618 46812 17682 46816
rect 17618 46756 17622 46812
rect 17622 46756 17678 46812
rect 17678 46756 17682 46812
rect 17618 46752 17682 46756
rect 17698 46812 17762 46816
rect 17698 46756 17702 46812
rect 17702 46756 17758 46812
rect 17758 46756 17762 46812
rect 17698 46752 17762 46756
rect 17778 46812 17842 46816
rect 17778 46756 17782 46812
rect 17782 46756 17838 46812
rect 17838 46756 17842 46812
rect 17778 46752 17842 46756
rect 17858 46812 17922 46816
rect 17858 46756 17862 46812
rect 17862 46756 17918 46812
rect 17918 46756 17922 46812
rect 17858 46752 17922 46756
rect 3188 46744 3252 46748
rect 3188 46688 3238 46744
rect 3238 46688 3252 46744
rect 3188 46684 3252 46688
rect 15332 46684 15396 46748
rect 7052 46412 7116 46476
rect 7618 46268 7682 46272
rect 7618 46212 7622 46268
rect 7622 46212 7678 46268
rect 7678 46212 7682 46268
rect 7618 46208 7682 46212
rect 7698 46268 7762 46272
rect 7698 46212 7702 46268
rect 7702 46212 7758 46268
rect 7758 46212 7762 46268
rect 7698 46208 7762 46212
rect 7778 46268 7842 46272
rect 7778 46212 7782 46268
rect 7782 46212 7838 46268
rect 7838 46212 7842 46268
rect 7778 46208 7842 46212
rect 7858 46268 7922 46272
rect 7858 46212 7862 46268
rect 7862 46212 7918 46268
rect 7918 46212 7922 46268
rect 7858 46208 7922 46212
rect 13308 46276 13372 46340
rect 14285 46268 14349 46272
rect 14285 46212 14289 46268
rect 14289 46212 14345 46268
rect 14345 46212 14349 46268
rect 14285 46208 14349 46212
rect 14365 46268 14429 46272
rect 14365 46212 14369 46268
rect 14369 46212 14425 46268
rect 14425 46212 14429 46268
rect 14365 46208 14429 46212
rect 14445 46268 14509 46272
rect 14445 46212 14449 46268
rect 14449 46212 14505 46268
rect 14505 46212 14509 46268
rect 14445 46208 14509 46212
rect 14525 46268 14589 46272
rect 14525 46212 14529 46268
rect 14529 46212 14585 46268
rect 14585 46212 14589 46268
rect 14525 46208 14589 46212
rect 12204 46140 12268 46204
rect 12572 46140 12636 46204
rect 5028 46004 5092 46068
rect 16988 46412 17052 46476
rect 2268 45868 2332 45932
rect 4844 45868 4908 45932
rect 10364 45868 10428 45932
rect 8708 45732 8772 45796
rect 9812 45732 9876 45796
rect 11652 45732 11716 45796
rect 12388 45732 12452 45796
rect 4285 45724 4349 45728
rect 4285 45668 4289 45724
rect 4289 45668 4345 45724
rect 4345 45668 4349 45724
rect 4285 45664 4349 45668
rect 4365 45724 4429 45728
rect 4365 45668 4369 45724
rect 4369 45668 4425 45724
rect 4425 45668 4429 45724
rect 4365 45664 4429 45668
rect 4445 45724 4509 45728
rect 4445 45668 4449 45724
rect 4449 45668 4505 45724
rect 4505 45668 4509 45724
rect 4445 45664 4509 45668
rect 4525 45724 4589 45728
rect 4525 45668 4529 45724
rect 4529 45668 4585 45724
rect 4585 45668 4589 45724
rect 4525 45664 4589 45668
rect 10952 45724 11016 45728
rect 10952 45668 10956 45724
rect 10956 45668 11012 45724
rect 11012 45668 11016 45724
rect 10952 45664 11016 45668
rect 11032 45724 11096 45728
rect 11032 45668 11036 45724
rect 11036 45668 11092 45724
rect 11092 45668 11096 45724
rect 11032 45664 11096 45668
rect 11112 45724 11176 45728
rect 11112 45668 11116 45724
rect 11116 45668 11172 45724
rect 11172 45668 11176 45724
rect 11112 45664 11176 45668
rect 11192 45724 11256 45728
rect 11192 45668 11196 45724
rect 11196 45668 11252 45724
rect 11252 45668 11256 45724
rect 11192 45664 11256 45668
rect 17618 45724 17682 45728
rect 17618 45668 17622 45724
rect 17622 45668 17678 45724
rect 17678 45668 17682 45724
rect 17618 45664 17682 45668
rect 17698 45724 17762 45728
rect 17698 45668 17702 45724
rect 17702 45668 17758 45724
rect 17758 45668 17762 45724
rect 17698 45664 17762 45668
rect 17778 45724 17842 45728
rect 17778 45668 17782 45724
rect 17782 45668 17838 45724
rect 17838 45668 17842 45724
rect 17778 45664 17842 45668
rect 17858 45724 17922 45728
rect 17858 45668 17862 45724
rect 17862 45668 17918 45724
rect 17918 45668 17922 45724
rect 17858 45664 17922 45668
rect 7052 45596 7116 45660
rect 8892 45656 8956 45660
rect 8892 45600 8942 45656
rect 8942 45600 8956 45656
rect 8892 45596 8956 45600
rect 15332 45596 15396 45660
rect 6132 45520 6196 45524
rect 6132 45464 6182 45520
rect 6182 45464 6196 45520
rect 6132 45460 6196 45464
rect 9812 45520 9876 45524
rect 9812 45464 9862 45520
rect 9862 45464 9876 45520
rect 9812 45460 9876 45464
rect 12204 45188 12268 45252
rect 7618 45180 7682 45184
rect 7618 45124 7622 45180
rect 7622 45124 7678 45180
rect 7678 45124 7682 45180
rect 7618 45120 7682 45124
rect 7698 45180 7762 45184
rect 7698 45124 7702 45180
rect 7702 45124 7758 45180
rect 7758 45124 7762 45180
rect 7698 45120 7762 45124
rect 7778 45180 7842 45184
rect 7778 45124 7782 45180
rect 7782 45124 7838 45180
rect 7838 45124 7842 45180
rect 7778 45120 7842 45124
rect 7858 45180 7922 45184
rect 7858 45124 7862 45180
rect 7862 45124 7918 45180
rect 7918 45124 7922 45180
rect 7858 45120 7922 45124
rect 14285 45180 14349 45184
rect 14285 45124 14289 45180
rect 14289 45124 14345 45180
rect 14345 45124 14349 45180
rect 14285 45120 14349 45124
rect 14365 45180 14429 45184
rect 14365 45124 14369 45180
rect 14369 45124 14425 45180
rect 14425 45124 14429 45180
rect 14365 45120 14429 45124
rect 14445 45180 14509 45184
rect 14445 45124 14449 45180
rect 14449 45124 14505 45180
rect 14505 45124 14509 45180
rect 14445 45120 14509 45124
rect 14525 45180 14589 45184
rect 14525 45124 14529 45180
rect 14529 45124 14585 45180
rect 14585 45124 14589 45180
rect 14525 45120 14589 45124
rect 4660 45052 4724 45116
rect 15700 45052 15764 45116
rect 4285 44636 4349 44640
rect 4285 44580 4289 44636
rect 4289 44580 4345 44636
rect 4345 44580 4349 44636
rect 4285 44576 4349 44580
rect 4365 44636 4429 44640
rect 4365 44580 4369 44636
rect 4369 44580 4425 44636
rect 4425 44580 4429 44636
rect 4365 44576 4429 44580
rect 4445 44636 4509 44640
rect 4445 44580 4449 44636
rect 4449 44580 4505 44636
rect 4505 44580 4509 44636
rect 4445 44576 4509 44580
rect 4525 44636 4589 44640
rect 4525 44580 4529 44636
rect 4529 44580 4585 44636
rect 4585 44580 4589 44636
rect 4525 44576 4589 44580
rect 10952 44636 11016 44640
rect 10952 44580 10956 44636
rect 10956 44580 11012 44636
rect 11012 44580 11016 44636
rect 10952 44576 11016 44580
rect 11032 44636 11096 44640
rect 11032 44580 11036 44636
rect 11036 44580 11092 44636
rect 11092 44580 11096 44636
rect 11032 44576 11096 44580
rect 11112 44636 11176 44640
rect 11112 44580 11116 44636
rect 11116 44580 11172 44636
rect 11172 44580 11176 44636
rect 11112 44576 11176 44580
rect 11192 44636 11256 44640
rect 11192 44580 11196 44636
rect 11196 44580 11252 44636
rect 11252 44580 11256 44636
rect 11192 44576 11256 44580
rect 17618 44636 17682 44640
rect 17618 44580 17622 44636
rect 17622 44580 17678 44636
rect 17678 44580 17682 44636
rect 17618 44576 17682 44580
rect 17698 44636 17762 44640
rect 17698 44580 17702 44636
rect 17702 44580 17758 44636
rect 17758 44580 17762 44636
rect 17698 44576 17762 44580
rect 17778 44636 17842 44640
rect 17778 44580 17782 44636
rect 17782 44580 17838 44636
rect 17838 44580 17842 44636
rect 17778 44576 17842 44580
rect 17858 44636 17922 44640
rect 17858 44580 17862 44636
rect 17862 44580 17918 44636
rect 17918 44580 17922 44636
rect 17858 44576 17922 44580
rect 3924 44432 3988 44436
rect 3924 44376 3974 44432
rect 3974 44376 3988 44432
rect 3924 44372 3988 44376
rect 9260 44372 9324 44436
rect 9076 44236 9140 44300
rect 9444 44100 9508 44164
rect 7618 44092 7682 44096
rect 7618 44036 7622 44092
rect 7622 44036 7678 44092
rect 7678 44036 7682 44092
rect 7618 44032 7682 44036
rect 7698 44092 7762 44096
rect 7698 44036 7702 44092
rect 7702 44036 7758 44092
rect 7758 44036 7762 44092
rect 7698 44032 7762 44036
rect 7778 44092 7842 44096
rect 7778 44036 7782 44092
rect 7782 44036 7838 44092
rect 7838 44036 7842 44092
rect 7778 44032 7842 44036
rect 7858 44092 7922 44096
rect 7858 44036 7862 44092
rect 7862 44036 7918 44092
rect 7918 44036 7922 44092
rect 7858 44032 7922 44036
rect 14285 44092 14349 44096
rect 14285 44036 14289 44092
rect 14289 44036 14345 44092
rect 14345 44036 14349 44092
rect 14285 44032 14349 44036
rect 14365 44092 14429 44096
rect 14365 44036 14369 44092
rect 14369 44036 14425 44092
rect 14425 44036 14429 44092
rect 14365 44032 14429 44036
rect 14445 44092 14509 44096
rect 14445 44036 14449 44092
rect 14449 44036 14505 44092
rect 14505 44036 14509 44092
rect 14445 44032 14509 44036
rect 14525 44092 14589 44096
rect 14525 44036 14529 44092
rect 14529 44036 14585 44092
rect 14585 44036 14589 44092
rect 14525 44032 14589 44036
rect 5396 43828 5460 43892
rect 9996 43828 10060 43892
rect 15516 43828 15580 43892
rect 13676 43692 13740 43756
rect 4285 43548 4349 43552
rect 4285 43492 4289 43548
rect 4289 43492 4345 43548
rect 4345 43492 4349 43548
rect 4285 43488 4349 43492
rect 4365 43548 4429 43552
rect 4365 43492 4369 43548
rect 4369 43492 4425 43548
rect 4425 43492 4429 43548
rect 4365 43488 4429 43492
rect 4445 43548 4509 43552
rect 4445 43492 4449 43548
rect 4449 43492 4505 43548
rect 4505 43492 4509 43548
rect 4445 43488 4509 43492
rect 4525 43548 4589 43552
rect 4525 43492 4529 43548
rect 4529 43492 4585 43548
rect 4585 43492 4589 43548
rect 4525 43488 4589 43492
rect 10952 43548 11016 43552
rect 10952 43492 10956 43548
rect 10956 43492 11012 43548
rect 11012 43492 11016 43548
rect 10952 43488 11016 43492
rect 11032 43548 11096 43552
rect 11032 43492 11036 43548
rect 11036 43492 11092 43548
rect 11092 43492 11096 43548
rect 11032 43488 11096 43492
rect 11112 43548 11176 43552
rect 11112 43492 11116 43548
rect 11116 43492 11172 43548
rect 11172 43492 11176 43548
rect 11112 43488 11176 43492
rect 11192 43548 11256 43552
rect 11192 43492 11196 43548
rect 11196 43492 11252 43548
rect 11252 43492 11256 43548
rect 11192 43488 11256 43492
rect 17618 43548 17682 43552
rect 17618 43492 17622 43548
rect 17622 43492 17678 43548
rect 17678 43492 17682 43548
rect 17618 43488 17682 43492
rect 17698 43548 17762 43552
rect 17698 43492 17702 43548
rect 17702 43492 17758 43548
rect 17758 43492 17762 43548
rect 17698 43488 17762 43492
rect 17778 43548 17842 43552
rect 17778 43492 17782 43548
rect 17782 43492 17838 43548
rect 17838 43492 17842 43548
rect 17778 43488 17842 43492
rect 17858 43548 17922 43552
rect 17858 43492 17862 43548
rect 17862 43492 17918 43548
rect 17918 43492 17922 43548
rect 17858 43488 17922 43492
rect 16436 43420 16500 43484
rect 8524 43284 8588 43348
rect 10180 43284 10244 43348
rect 6316 43012 6380 43076
rect 7618 43004 7682 43008
rect 7618 42948 7622 43004
rect 7622 42948 7678 43004
rect 7678 42948 7682 43004
rect 7618 42944 7682 42948
rect 7698 43004 7762 43008
rect 7698 42948 7702 43004
rect 7702 42948 7758 43004
rect 7758 42948 7762 43004
rect 7698 42944 7762 42948
rect 7778 43004 7842 43008
rect 7778 42948 7782 43004
rect 7782 42948 7838 43004
rect 7838 42948 7842 43004
rect 7778 42944 7842 42948
rect 7858 43004 7922 43008
rect 7858 42948 7862 43004
rect 7862 42948 7918 43004
rect 7918 42948 7922 43004
rect 7858 42944 7922 42948
rect 6868 42876 6932 42940
rect 9076 42876 9140 42940
rect 9996 42876 10060 42940
rect 15332 43148 15396 43212
rect 14285 43004 14349 43008
rect 14285 42948 14289 43004
rect 14289 42948 14345 43004
rect 14345 42948 14349 43004
rect 14285 42944 14349 42948
rect 14365 43004 14429 43008
rect 14365 42948 14369 43004
rect 14369 42948 14425 43004
rect 14425 42948 14429 43004
rect 14365 42944 14429 42948
rect 14445 43004 14509 43008
rect 14445 42948 14449 43004
rect 14449 42948 14505 43004
rect 14505 42948 14509 43004
rect 14445 42944 14509 42948
rect 14525 43004 14589 43008
rect 14525 42948 14529 43004
rect 14529 42948 14585 43004
rect 14585 42948 14589 43004
rect 14525 42944 14589 42948
rect 10364 42936 10428 42940
rect 10364 42880 10414 42936
rect 10414 42880 10428 42936
rect 10364 42876 10428 42880
rect 2452 42740 2516 42804
rect 6132 42800 6196 42804
rect 6132 42744 6182 42800
rect 6182 42744 6196 42800
rect 6132 42740 6196 42744
rect 8340 42800 8404 42804
rect 8340 42744 8354 42800
rect 8354 42744 8404 42800
rect 8340 42740 8404 42744
rect 16068 42800 16132 42804
rect 16068 42744 16082 42800
rect 16082 42744 16132 42800
rect 16068 42740 16132 42744
rect 4285 42460 4349 42464
rect 4285 42404 4289 42460
rect 4289 42404 4345 42460
rect 4345 42404 4349 42460
rect 4285 42400 4349 42404
rect 4365 42460 4429 42464
rect 4365 42404 4369 42460
rect 4369 42404 4425 42460
rect 4425 42404 4429 42460
rect 4365 42400 4429 42404
rect 4445 42460 4509 42464
rect 4445 42404 4449 42460
rect 4449 42404 4505 42460
rect 4505 42404 4509 42460
rect 4445 42400 4509 42404
rect 4525 42460 4589 42464
rect 4525 42404 4529 42460
rect 4529 42404 4585 42460
rect 4585 42404 4589 42460
rect 4525 42400 4589 42404
rect 10952 42460 11016 42464
rect 10952 42404 10956 42460
rect 10956 42404 11012 42460
rect 11012 42404 11016 42460
rect 10952 42400 11016 42404
rect 11032 42460 11096 42464
rect 11032 42404 11036 42460
rect 11036 42404 11092 42460
rect 11092 42404 11096 42460
rect 11032 42400 11096 42404
rect 11112 42460 11176 42464
rect 11112 42404 11116 42460
rect 11116 42404 11172 42460
rect 11172 42404 11176 42460
rect 11112 42400 11176 42404
rect 11192 42460 11256 42464
rect 11192 42404 11196 42460
rect 11196 42404 11252 42460
rect 11252 42404 11256 42460
rect 11192 42400 11256 42404
rect 17618 42460 17682 42464
rect 17618 42404 17622 42460
rect 17622 42404 17678 42460
rect 17678 42404 17682 42460
rect 17618 42400 17682 42404
rect 17698 42460 17762 42464
rect 17698 42404 17702 42460
rect 17702 42404 17758 42460
rect 17758 42404 17762 42460
rect 17698 42400 17762 42404
rect 17778 42460 17842 42464
rect 17778 42404 17782 42460
rect 17782 42404 17838 42460
rect 17838 42404 17842 42460
rect 17778 42400 17842 42404
rect 17858 42460 17922 42464
rect 17858 42404 17862 42460
rect 17862 42404 17918 42460
rect 17918 42404 17922 42460
rect 17858 42400 17922 42404
rect 8708 42196 8772 42260
rect 11652 42256 11716 42260
rect 11652 42200 11666 42256
rect 11666 42200 11716 42256
rect 11652 42196 11716 42200
rect 6684 42060 6748 42124
rect 5580 41924 5644 41988
rect 7618 41916 7682 41920
rect 7618 41860 7622 41916
rect 7622 41860 7678 41916
rect 7678 41860 7682 41916
rect 7618 41856 7682 41860
rect 7698 41916 7762 41920
rect 7698 41860 7702 41916
rect 7702 41860 7758 41916
rect 7758 41860 7762 41916
rect 7698 41856 7762 41860
rect 7778 41916 7842 41920
rect 7778 41860 7782 41916
rect 7782 41860 7838 41916
rect 7838 41860 7842 41916
rect 7778 41856 7842 41860
rect 7858 41916 7922 41920
rect 7858 41860 7862 41916
rect 7862 41860 7918 41916
rect 7918 41860 7922 41916
rect 7858 41856 7922 41860
rect 14285 41916 14349 41920
rect 14285 41860 14289 41916
rect 14289 41860 14345 41916
rect 14345 41860 14349 41916
rect 14285 41856 14349 41860
rect 14365 41916 14429 41920
rect 14365 41860 14369 41916
rect 14369 41860 14425 41916
rect 14425 41860 14429 41916
rect 14365 41856 14429 41860
rect 14445 41916 14509 41920
rect 14445 41860 14449 41916
rect 14449 41860 14505 41916
rect 14505 41860 14509 41916
rect 14445 41856 14509 41860
rect 14525 41916 14589 41920
rect 14525 41860 14529 41916
rect 14529 41860 14585 41916
rect 14585 41860 14589 41916
rect 14525 41856 14589 41860
rect 16804 41788 16868 41852
rect 16988 41652 17052 41716
rect 15332 41516 15396 41580
rect 16436 41576 16500 41580
rect 16436 41520 16450 41576
rect 16450 41520 16500 41576
rect 16436 41516 16500 41520
rect 5764 41380 5828 41444
rect 6684 41380 6748 41444
rect 9260 41380 9324 41444
rect 4285 41372 4349 41376
rect 4285 41316 4289 41372
rect 4289 41316 4345 41372
rect 4345 41316 4349 41372
rect 4285 41312 4349 41316
rect 4365 41372 4429 41376
rect 4365 41316 4369 41372
rect 4369 41316 4425 41372
rect 4425 41316 4429 41372
rect 4365 41312 4429 41316
rect 4445 41372 4509 41376
rect 4445 41316 4449 41372
rect 4449 41316 4505 41372
rect 4505 41316 4509 41372
rect 4445 41312 4509 41316
rect 4525 41372 4589 41376
rect 4525 41316 4529 41372
rect 4529 41316 4585 41372
rect 4585 41316 4589 41372
rect 4525 41312 4589 41316
rect 10952 41372 11016 41376
rect 10952 41316 10956 41372
rect 10956 41316 11012 41372
rect 11012 41316 11016 41372
rect 10952 41312 11016 41316
rect 11032 41372 11096 41376
rect 11032 41316 11036 41372
rect 11036 41316 11092 41372
rect 11092 41316 11096 41372
rect 11032 41312 11096 41316
rect 11112 41372 11176 41376
rect 11112 41316 11116 41372
rect 11116 41316 11172 41372
rect 11172 41316 11176 41372
rect 11112 41312 11176 41316
rect 11192 41372 11256 41376
rect 11192 41316 11196 41372
rect 11196 41316 11252 41372
rect 11252 41316 11256 41372
rect 11192 41312 11256 41316
rect 6684 41244 6748 41308
rect 8340 41244 8404 41308
rect 16804 41380 16868 41444
rect 16988 41440 17052 41444
rect 16988 41384 17038 41440
rect 17038 41384 17052 41440
rect 16988 41380 17052 41384
rect 17618 41372 17682 41376
rect 17618 41316 17622 41372
rect 17622 41316 17678 41372
rect 17678 41316 17682 41372
rect 17618 41312 17682 41316
rect 17698 41372 17762 41376
rect 17698 41316 17702 41372
rect 17702 41316 17758 41372
rect 17758 41316 17762 41372
rect 17698 41312 17762 41316
rect 17778 41372 17842 41376
rect 17778 41316 17782 41372
rect 17782 41316 17838 41372
rect 17838 41316 17842 41372
rect 17778 41312 17842 41316
rect 17858 41372 17922 41376
rect 17858 41316 17862 41372
rect 17862 41316 17918 41372
rect 17918 41316 17922 41372
rect 17858 41312 17922 41316
rect 5764 41108 5828 41172
rect 13676 41108 13740 41172
rect 14780 41108 14844 41172
rect 15332 41244 15396 41308
rect 16804 41244 16868 41308
rect 15884 41108 15948 41172
rect 13492 40972 13556 41036
rect 14780 40972 14844 41036
rect 15148 40972 15212 41036
rect 5580 40896 5644 40900
rect 5580 40840 5594 40896
rect 5594 40840 5644 40896
rect 5580 40836 5644 40840
rect 7618 40828 7682 40832
rect 7618 40772 7622 40828
rect 7622 40772 7678 40828
rect 7678 40772 7682 40828
rect 7618 40768 7682 40772
rect 7698 40828 7762 40832
rect 7698 40772 7702 40828
rect 7702 40772 7758 40828
rect 7758 40772 7762 40828
rect 7698 40768 7762 40772
rect 7778 40828 7842 40832
rect 7778 40772 7782 40828
rect 7782 40772 7838 40828
rect 7838 40772 7842 40828
rect 7778 40768 7842 40772
rect 7858 40828 7922 40832
rect 7858 40772 7862 40828
rect 7862 40772 7918 40828
rect 7918 40772 7922 40828
rect 7858 40768 7922 40772
rect 14285 40828 14349 40832
rect 14285 40772 14289 40828
rect 14289 40772 14345 40828
rect 14345 40772 14349 40828
rect 14285 40768 14349 40772
rect 14365 40828 14429 40832
rect 14365 40772 14369 40828
rect 14369 40772 14425 40828
rect 14425 40772 14429 40828
rect 14365 40768 14429 40772
rect 14445 40828 14509 40832
rect 14445 40772 14449 40828
rect 14449 40772 14505 40828
rect 14505 40772 14509 40828
rect 14445 40768 14509 40772
rect 14525 40828 14589 40832
rect 14525 40772 14529 40828
rect 14529 40772 14585 40828
rect 14585 40772 14589 40828
rect 14525 40768 14589 40772
rect 15516 40700 15580 40764
rect 8340 40564 8404 40628
rect 16436 40292 16500 40356
rect 4285 40284 4349 40288
rect 4285 40228 4289 40284
rect 4289 40228 4345 40284
rect 4345 40228 4349 40284
rect 4285 40224 4349 40228
rect 4365 40284 4429 40288
rect 4365 40228 4369 40284
rect 4369 40228 4425 40284
rect 4425 40228 4429 40284
rect 4365 40224 4429 40228
rect 4445 40284 4509 40288
rect 4445 40228 4449 40284
rect 4449 40228 4505 40284
rect 4505 40228 4509 40284
rect 4445 40224 4509 40228
rect 4525 40284 4589 40288
rect 4525 40228 4529 40284
rect 4529 40228 4585 40284
rect 4585 40228 4589 40284
rect 4525 40224 4589 40228
rect 10952 40284 11016 40288
rect 10952 40228 10956 40284
rect 10956 40228 11012 40284
rect 11012 40228 11016 40284
rect 10952 40224 11016 40228
rect 11032 40284 11096 40288
rect 11032 40228 11036 40284
rect 11036 40228 11092 40284
rect 11092 40228 11096 40284
rect 11032 40224 11096 40228
rect 11112 40284 11176 40288
rect 11112 40228 11116 40284
rect 11116 40228 11172 40284
rect 11172 40228 11176 40284
rect 11112 40224 11176 40228
rect 11192 40284 11256 40288
rect 11192 40228 11196 40284
rect 11196 40228 11252 40284
rect 11252 40228 11256 40284
rect 11192 40224 11256 40228
rect 17618 40284 17682 40288
rect 17618 40228 17622 40284
rect 17622 40228 17678 40284
rect 17678 40228 17682 40284
rect 17618 40224 17682 40228
rect 17698 40284 17762 40288
rect 17698 40228 17702 40284
rect 17702 40228 17758 40284
rect 17758 40228 17762 40284
rect 17698 40224 17762 40228
rect 17778 40284 17842 40288
rect 17778 40228 17782 40284
rect 17782 40228 17838 40284
rect 17838 40228 17842 40284
rect 17778 40224 17842 40228
rect 17858 40284 17922 40288
rect 17858 40228 17862 40284
rect 17862 40228 17918 40284
rect 17918 40228 17922 40284
rect 17858 40224 17922 40228
rect 3924 40156 3988 40220
rect 17172 40080 17236 40084
rect 17172 40024 17222 40080
rect 17222 40024 17236 40080
rect 17172 40020 17236 40024
rect 4108 39884 4172 39948
rect 11468 39884 11532 39948
rect 11652 39944 11716 39948
rect 11652 39888 11702 39944
rect 11702 39888 11716 39944
rect 11652 39884 11716 39888
rect 6316 39748 6380 39812
rect 7618 39740 7682 39744
rect 7618 39684 7622 39740
rect 7622 39684 7678 39740
rect 7678 39684 7682 39740
rect 7618 39680 7682 39684
rect 7698 39740 7762 39744
rect 7698 39684 7702 39740
rect 7702 39684 7758 39740
rect 7758 39684 7762 39740
rect 7698 39680 7762 39684
rect 7778 39740 7842 39744
rect 7778 39684 7782 39740
rect 7782 39684 7838 39740
rect 7838 39684 7842 39740
rect 7778 39680 7842 39684
rect 7858 39740 7922 39744
rect 7858 39684 7862 39740
rect 7862 39684 7918 39740
rect 7918 39684 7922 39740
rect 7858 39680 7922 39684
rect 14285 39740 14349 39744
rect 14285 39684 14289 39740
rect 14289 39684 14345 39740
rect 14345 39684 14349 39740
rect 14285 39680 14349 39684
rect 14365 39740 14429 39744
rect 14365 39684 14369 39740
rect 14369 39684 14425 39740
rect 14425 39684 14429 39740
rect 14365 39680 14429 39684
rect 14445 39740 14509 39744
rect 14445 39684 14449 39740
rect 14449 39684 14505 39740
rect 14505 39684 14509 39740
rect 14445 39680 14509 39684
rect 14525 39740 14589 39744
rect 14525 39684 14529 39740
rect 14529 39684 14585 39740
rect 14585 39684 14589 39740
rect 14525 39680 14589 39684
rect 13492 39476 13556 39540
rect 16068 39476 16132 39540
rect 12572 39340 12636 39404
rect 15516 39204 15580 39268
rect 4285 39196 4349 39200
rect 4285 39140 4289 39196
rect 4289 39140 4345 39196
rect 4345 39140 4349 39196
rect 4285 39136 4349 39140
rect 4365 39196 4429 39200
rect 4365 39140 4369 39196
rect 4369 39140 4425 39196
rect 4425 39140 4429 39196
rect 4365 39136 4429 39140
rect 4445 39196 4509 39200
rect 4445 39140 4449 39196
rect 4449 39140 4505 39196
rect 4505 39140 4509 39196
rect 4445 39136 4509 39140
rect 4525 39196 4589 39200
rect 4525 39140 4529 39196
rect 4529 39140 4585 39196
rect 4585 39140 4589 39196
rect 4525 39136 4589 39140
rect 10952 39196 11016 39200
rect 10952 39140 10956 39196
rect 10956 39140 11012 39196
rect 11012 39140 11016 39196
rect 10952 39136 11016 39140
rect 11032 39196 11096 39200
rect 11032 39140 11036 39196
rect 11036 39140 11092 39196
rect 11092 39140 11096 39196
rect 11032 39136 11096 39140
rect 11112 39196 11176 39200
rect 11112 39140 11116 39196
rect 11116 39140 11172 39196
rect 11172 39140 11176 39196
rect 11112 39136 11176 39140
rect 11192 39196 11256 39200
rect 11192 39140 11196 39196
rect 11196 39140 11252 39196
rect 11252 39140 11256 39196
rect 11192 39136 11256 39140
rect 17618 39196 17682 39200
rect 17618 39140 17622 39196
rect 17622 39140 17678 39196
rect 17678 39140 17682 39196
rect 17618 39136 17682 39140
rect 17698 39196 17762 39200
rect 17698 39140 17702 39196
rect 17702 39140 17758 39196
rect 17758 39140 17762 39196
rect 17698 39136 17762 39140
rect 17778 39196 17842 39200
rect 17778 39140 17782 39196
rect 17782 39140 17838 39196
rect 17838 39140 17842 39196
rect 17778 39136 17842 39140
rect 17858 39196 17922 39200
rect 17858 39140 17862 39196
rect 17862 39140 17918 39196
rect 17918 39140 17922 39196
rect 17858 39136 17922 39140
rect 9996 39068 10060 39132
rect 12204 38932 12268 38996
rect 12756 38660 12820 38724
rect 7618 38652 7682 38656
rect 7618 38596 7622 38652
rect 7622 38596 7678 38652
rect 7678 38596 7682 38652
rect 7618 38592 7682 38596
rect 7698 38652 7762 38656
rect 7698 38596 7702 38652
rect 7702 38596 7758 38652
rect 7758 38596 7762 38652
rect 7698 38592 7762 38596
rect 7778 38652 7842 38656
rect 7778 38596 7782 38652
rect 7782 38596 7838 38652
rect 7838 38596 7842 38652
rect 7778 38592 7842 38596
rect 7858 38652 7922 38656
rect 7858 38596 7862 38652
rect 7862 38596 7918 38652
rect 7918 38596 7922 38652
rect 7858 38592 7922 38596
rect 14285 38652 14349 38656
rect 14285 38596 14289 38652
rect 14289 38596 14345 38652
rect 14345 38596 14349 38652
rect 14285 38592 14349 38596
rect 14365 38652 14429 38656
rect 14365 38596 14369 38652
rect 14369 38596 14425 38652
rect 14425 38596 14429 38652
rect 14365 38592 14429 38596
rect 14445 38652 14509 38656
rect 14445 38596 14449 38652
rect 14449 38596 14505 38652
rect 14505 38596 14509 38652
rect 14445 38592 14509 38596
rect 14525 38652 14589 38656
rect 14525 38596 14529 38652
rect 14529 38596 14585 38652
rect 14585 38596 14589 38652
rect 14525 38592 14589 38596
rect 15884 38524 15948 38588
rect 8708 38388 8772 38452
rect 15148 38252 15212 38316
rect 6868 38116 6932 38180
rect 4285 38108 4349 38112
rect 4285 38052 4289 38108
rect 4289 38052 4345 38108
rect 4345 38052 4349 38108
rect 4285 38048 4349 38052
rect 4365 38108 4429 38112
rect 4365 38052 4369 38108
rect 4369 38052 4425 38108
rect 4425 38052 4429 38108
rect 4365 38048 4429 38052
rect 4445 38108 4509 38112
rect 4445 38052 4449 38108
rect 4449 38052 4505 38108
rect 4505 38052 4509 38108
rect 4445 38048 4509 38052
rect 4525 38108 4589 38112
rect 4525 38052 4529 38108
rect 4529 38052 4585 38108
rect 4585 38052 4589 38108
rect 4525 38048 4589 38052
rect 10952 38108 11016 38112
rect 10952 38052 10956 38108
rect 10956 38052 11012 38108
rect 11012 38052 11016 38108
rect 10952 38048 11016 38052
rect 11032 38108 11096 38112
rect 11032 38052 11036 38108
rect 11036 38052 11092 38108
rect 11092 38052 11096 38108
rect 11032 38048 11096 38052
rect 11112 38108 11176 38112
rect 11112 38052 11116 38108
rect 11116 38052 11172 38108
rect 11172 38052 11176 38108
rect 11112 38048 11176 38052
rect 11192 38108 11256 38112
rect 11192 38052 11196 38108
rect 11196 38052 11252 38108
rect 11252 38052 11256 38108
rect 11192 38048 11256 38052
rect 17618 38108 17682 38112
rect 17618 38052 17622 38108
rect 17622 38052 17678 38108
rect 17678 38052 17682 38108
rect 17618 38048 17682 38052
rect 17698 38108 17762 38112
rect 17698 38052 17702 38108
rect 17702 38052 17758 38108
rect 17758 38052 17762 38108
rect 17698 38048 17762 38052
rect 17778 38108 17842 38112
rect 17778 38052 17782 38108
rect 17782 38052 17838 38108
rect 17838 38052 17842 38108
rect 17778 38048 17842 38052
rect 17858 38108 17922 38112
rect 17858 38052 17862 38108
rect 17862 38052 17918 38108
rect 17918 38052 17922 38108
rect 17858 38048 17922 38052
rect 7618 37564 7682 37568
rect 7618 37508 7622 37564
rect 7622 37508 7678 37564
rect 7678 37508 7682 37564
rect 7618 37504 7682 37508
rect 7698 37564 7762 37568
rect 7698 37508 7702 37564
rect 7702 37508 7758 37564
rect 7758 37508 7762 37564
rect 7698 37504 7762 37508
rect 7778 37564 7842 37568
rect 7778 37508 7782 37564
rect 7782 37508 7838 37564
rect 7838 37508 7842 37564
rect 7778 37504 7842 37508
rect 7858 37564 7922 37568
rect 7858 37508 7862 37564
rect 7862 37508 7918 37564
rect 7918 37508 7922 37564
rect 7858 37504 7922 37508
rect 14285 37564 14349 37568
rect 14285 37508 14289 37564
rect 14289 37508 14345 37564
rect 14345 37508 14349 37564
rect 14285 37504 14349 37508
rect 14365 37564 14429 37568
rect 14365 37508 14369 37564
rect 14369 37508 14425 37564
rect 14425 37508 14429 37564
rect 14365 37504 14429 37508
rect 14445 37564 14509 37568
rect 14445 37508 14449 37564
rect 14449 37508 14505 37564
rect 14505 37508 14509 37564
rect 14445 37504 14509 37508
rect 14525 37564 14589 37568
rect 14525 37508 14529 37564
rect 14529 37508 14585 37564
rect 14585 37508 14589 37564
rect 14525 37504 14589 37508
rect 15332 37496 15396 37500
rect 15332 37440 15382 37496
rect 15382 37440 15396 37496
rect 15332 37436 15396 37440
rect 7236 37028 7300 37092
rect 4285 37020 4349 37024
rect 4285 36964 4289 37020
rect 4289 36964 4345 37020
rect 4345 36964 4349 37020
rect 4285 36960 4349 36964
rect 4365 37020 4429 37024
rect 4365 36964 4369 37020
rect 4369 36964 4425 37020
rect 4425 36964 4429 37020
rect 4365 36960 4429 36964
rect 4445 37020 4509 37024
rect 4445 36964 4449 37020
rect 4449 36964 4505 37020
rect 4505 36964 4509 37020
rect 4445 36960 4509 36964
rect 4525 37020 4589 37024
rect 4525 36964 4529 37020
rect 4529 36964 4585 37020
rect 4585 36964 4589 37020
rect 4525 36960 4589 36964
rect 14780 37164 14844 37228
rect 16804 37164 16868 37228
rect 10952 37020 11016 37024
rect 10952 36964 10956 37020
rect 10956 36964 11012 37020
rect 11012 36964 11016 37020
rect 10952 36960 11016 36964
rect 11032 37020 11096 37024
rect 11032 36964 11036 37020
rect 11036 36964 11092 37020
rect 11092 36964 11096 37020
rect 11032 36960 11096 36964
rect 11112 37020 11176 37024
rect 11112 36964 11116 37020
rect 11116 36964 11172 37020
rect 11172 36964 11176 37020
rect 11112 36960 11176 36964
rect 11192 37020 11256 37024
rect 11192 36964 11196 37020
rect 11196 36964 11252 37020
rect 11252 36964 11256 37020
rect 11192 36960 11256 36964
rect 17618 37020 17682 37024
rect 17618 36964 17622 37020
rect 17622 36964 17678 37020
rect 17678 36964 17682 37020
rect 17618 36960 17682 36964
rect 17698 37020 17762 37024
rect 17698 36964 17702 37020
rect 17702 36964 17758 37020
rect 17758 36964 17762 37020
rect 17698 36960 17762 36964
rect 17778 37020 17842 37024
rect 17778 36964 17782 37020
rect 17782 36964 17838 37020
rect 17838 36964 17842 37020
rect 17778 36960 17842 36964
rect 17858 37020 17922 37024
rect 17858 36964 17862 37020
rect 17862 36964 17918 37020
rect 17918 36964 17922 37020
rect 17858 36960 17922 36964
rect 9812 36756 9876 36820
rect 5764 36408 5828 36412
rect 7618 36476 7682 36480
rect 7618 36420 7622 36476
rect 7622 36420 7678 36476
rect 7678 36420 7682 36476
rect 7618 36416 7682 36420
rect 7698 36476 7762 36480
rect 7698 36420 7702 36476
rect 7702 36420 7758 36476
rect 7758 36420 7762 36476
rect 7698 36416 7762 36420
rect 7778 36476 7842 36480
rect 7778 36420 7782 36476
rect 7782 36420 7838 36476
rect 7838 36420 7842 36476
rect 7778 36416 7842 36420
rect 7858 36476 7922 36480
rect 7858 36420 7862 36476
rect 7862 36420 7918 36476
rect 7918 36420 7922 36476
rect 7858 36416 7922 36420
rect 14285 36476 14349 36480
rect 14285 36420 14289 36476
rect 14289 36420 14345 36476
rect 14345 36420 14349 36476
rect 14285 36416 14349 36420
rect 14365 36476 14429 36480
rect 14365 36420 14369 36476
rect 14369 36420 14425 36476
rect 14425 36420 14429 36476
rect 14365 36416 14429 36420
rect 14445 36476 14509 36480
rect 14445 36420 14449 36476
rect 14449 36420 14505 36476
rect 14505 36420 14509 36476
rect 14445 36416 14509 36420
rect 14525 36476 14589 36480
rect 14525 36420 14529 36476
rect 14529 36420 14585 36476
rect 14585 36420 14589 36476
rect 14525 36416 14589 36420
rect 5764 36352 5814 36408
rect 5814 36352 5828 36408
rect 5764 36348 5828 36352
rect 4285 35932 4349 35936
rect 4285 35876 4289 35932
rect 4289 35876 4345 35932
rect 4345 35876 4349 35932
rect 4285 35872 4349 35876
rect 4365 35932 4429 35936
rect 4365 35876 4369 35932
rect 4369 35876 4425 35932
rect 4425 35876 4429 35932
rect 4365 35872 4429 35876
rect 4445 35932 4509 35936
rect 4445 35876 4449 35932
rect 4449 35876 4505 35932
rect 4505 35876 4509 35932
rect 4445 35872 4509 35876
rect 4525 35932 4589 35936
rect 4525 35876 4529 35932
rect 4529 35876 4585 35932
rect 4585 35876 4589 35932
rect 4525 35872 4589 35876
rect 10952 35932 11016 35936
rect 10952 35876 10956 35932
rect 10956 35876 11012 35932
rect 11012 35876 11016 35932
rect 10952 35872 11016 35876
rect 11032 35932 11096 35936
rect 11032 35876 11036 35932
rect 11036 35876 11092 35932
rect 11092 35876 11096 35932
rect 11032 35872 11096 35876
rect 11112 35932 11176 35936
rect 11112 35876 11116 35932
rect 11116 35876 11172 35932
rect 11172 35876 11176 35932
rect 11112 35872 11176 35876
rect 11192 35932 11256 35936
rect 11192 35876 11196 35932
rect 11196 35876 11252 35932
rect 11252 35876 11256 35932
rect 11192 35872 11256 35876
rect 17618 35932 17682 35936
rect 17618 35876 17622 35932
rect 17622 35876 17678 35932
rect 17678 35876 17682 35932
rect 17618 35872 17682 35876
rect 17698 35932 17762 35936
rect 17698 35876 17702 35932
rect 17702 35876 17758 35932
rect 17758 35876 17762 35932
rect 17698 35872 17762 35876
rect 17778 35932 17842 35936
rect 17778 35876 17782 35932
rect 17782 35876 17838 35932
rect 17838 35876 17842 35932
rect 17778 35872 17842 35876
rect 17858 35932 17922 35936
rect 17858 35876 17862 35932
rect 17862 35876 17918 35932
rect 17918 35876 17922 35932
rect 17858 35872 17922 35876
rect 15700 35728 15764 35732
rect 15700 35672 15714 35728
rect 15714 35672 15764 35728
rect 15700 35668 15764 35672
rect 7618 35388 7682 35392
rect 7618 35332 7622 35388
rect 7622 35332 7678 35388
rect 7678 35332 7682 35388
rect 7618 35328 7682 35332
rect 7698 35388 7762 35392
rect 7698 35332 7702 35388
rect 7702 35332 7758 35388
rect 7758 35332 7762 35388
rect 7698 35328 7762 35332
rect 7778 35388 7842 35392
rect 7778 35332 7782 35388
rect 7782 35332 7838 35388
rect 7838 35332 7842 35388
rect 7778 35328 7842 35332
rect 7858 35388 7922 35392
rect 7858 35332 7862 35388
rect 7862 35332 7918 35388
rect 7918 35332 7922 35388
rect 7858 35328 7922 35332
rect 14285 35388 14349 35392
rect 14285 35332 14289 35388
rect 14289 35332 14345 35388
rect 14345 35332 14349 35388
rect 14285 35328 14349 35332
rect 14365 35388 14429 35392
rect 14365 35332 14369 35388
rect 14369 35332 14425 35388
rect 14425 35332 14429 35388
rect 14365 35328 14429 35332
rect 14445 35388 14509 35392
rect 14445 35332 14449 35388
rect 14449 35332 14505 35388
rect 14505 35332 14509 35388
rect 14445 35328 14509 35332
rect 14525 35388 14589 35392
rect 14525 35332 14529 35388
rect 14529 35332 14585 35388
rect 14585 35332 14589 35388
rect 14525 35328 14589 35332
rect 13676 34988 13740 35052
rect 4285 34844 4349 34848
rect 4285 34788 4289 34844
rect 4289 34788 4345 34844
rect 4345 34788 4349 34844
rect 4285 34784 4349 34788
rect 4365 34844 4429 34848
rect 4365 34788 4369 34844
rect 4369 34788 4425 34844
rect 4425 34788 4429 34844
rect 4365 34784 4429 34788
rect 4445 34844 4509 34848
rect 4445 34788 4449 34844
rect 4449 34788 4505 34844
rect 4505 34788 4509 34844
rect 4445 34784 4509 34788
rect 4525 34844 4589 34848
rect 4525 34788 4529 34844
rect 4529 34788 4585 34844
rect 4585 34788 4589 34844
rect 4525 34784 4589 34788
rect 10952 34844 11016 34848
rect 10952 34788 10956 34844
rect 10956 34788 11012 34844
rect 11012 34788 11016 34844
rect 10952 34784 11016 34788
rect 11032 34844 11096 34848
rect 11032 34788 11036 34844
rect 11036 34788 11092 34844
rect 11092 34788 11096 34844
rect 11032 34784 11096 34788
rect 11112 34844 11176 34848
rect 11112 34788 11116 34844
rect 11116 34788 11172 34844
rect 11172 34788 11176 34844
rect 11112 34784 11176 34788
rect 11192 34844 11256 34848
rect 11192 34788 11196 34844
rect 11196 34788 11252 34844
rect 11252 34788 11256 34844
rect 11192 34784 11256 34788
rect 17618 34844 17682 34848
rect 17618 34788 17622 34844
rect 17622 34788 17678 34844
rect 17678 34788 17682 34844
rect 17618 34784 17682 34788
rect 17698 34844 17762 34848
rect 17698 34788 17702 34844
rect 17702 34788 17758 34844
rect 17758 34788 17762 34844
rect 17698 34784 17762 34788
rect 17778 34844 17842 34848
rect 17778 34788 17782 34844
rect 17782 34788 17838 34844
rect 17838 34788 17842 34844
rect 17778 34784 17842 34788
rect 17858 34844 17922 34848
rect 17858 34788 17862 34844
rect 17862 34788 17918 34844
rect 17918 34788 17922 34844
rect 17858 34784 17922 34788
rect 16436 34444 16500 34508
rect 7618 34300 7682 34304
rect 7618 34244 7622 34300
rect 7622 34244 7678 34300
rect 7678 34244 7682 34300
rect 7618 34240 7682 34244
rect 7698 34300 7762 34304
rect 7698 34244 7702 34300
rect 7702 34244 7758 34300
rect 7758 34244 7762 34300
rect 7698 34240 7762 34244
rect 7778 34300 7842 34304
rect 7778 34244 7782 34300
rect 7782 34244 7838 34300
rect 7838 34244 7842 34300
rect 7778 34240 7842 34244
rect 7858 34300 7922 34304
rect 7858 34244 7862 34300
rect 7862 34244 7918 34300
rect 7918 34244 7922 34300
rect 7858 34240 7922 34244
rect 14285 34300 14349 34304
rect 14285 34244 14289 34300
rect 14289 34244 14345 34300
rect 14345 34244 14349 34300
rect 14285 34240 14349 34244
rect 14365 34300 14429 34304
rect 14365 34244 14369 34300
rect 14369 34244 14425 34300
rect 14425 34244 14429 34300
rect 14365 34240 14429 34244
rect 14445 34300 14509 34304
rect 14445 34244 14449 34300
rect 14449 34244 14505 34300
rect 14505 34244 14509 34300
rect 14445 34240 14509 34244
rect 14525 34300 14589 34304
rect 14525 34244 14529 34300
rect 14529 34244 14585 34300
rect 14585 34244 14589 34300
rect 14525 34240 14589 34244
rect 10364 34036 10428 34100
rect 15148 34036 15212 34100
rect 4285 33756 4349 33760
rect 4285 33700 4289 33756
rect 4289 33700 4345 33756
rect 4345 33700 4349 33756
rect 4285 33696 4349 33700
rect 4365 33756 4429 33760
rect 4365 33700 4369 33756
rect 4369 33700 4425 33756
rect 4425 33700 4429 33756
rect 4365 33696 4429 33700
rect 4445 33756 4509 33760
rect 4445 33700 4449 33756
rect 4449 33700 4505 33756
rect 4505 33700 4509 33756
rect 4445 33696 4509 33700
rect 4525 33756 4589 33760
rect 4525 33700 4529 33756
rect 4529 33700 4585 33756
rect 4585 33700 4589 33756
rect 4525 33696 4589 33700
rect 10952 33756 11016 33760
rect 10952 33700 10956 33756
rect 10956 33700 11012 33756
rect 11012 33700 11016 33756
rect 10952 33696 11016 33700
rect 11032 33756 11096 33760
rect 11032 33700 11036 33756
rect 11036 33700 11092 33756
rect 11092 33700 11096 33756
rect 11032 33696 11096 33700
rect 11112 33756 11176 33760
rect 11112 33700 11116 33756
rect 11116 33700 11172 33756
rect 11172 33700 11176 33756
rect 11112 33696 11176 33700
rect 11192 33756 11256 33760
rect 11192 33700 11196 33756
rect 11196 33700 11252 33756
rect 11252 33700 11256 33756
rect 11192 33696 11256 33700
rect 17618 33756 17682 33760
rect 17618 33700 17622 33756
rect 17622 33700 17678 33756
rect 17678 33700 17682 33756
rect 17618 33696 17682 33700
rect 17698 33756 17762 33760
rect 17698 33700 17702 33756
rect 17702 33700 17758 33756
rect 17758 33700 17762 33756
rect 17698 33696 17762 33700
rect 17778 33756 17842 33760
rect 17778 33700 17782 33756
rect 17782 33700 17838 33756
rect 17838 33700 17842 33756
rect 17778 33696 17842 33700
rect 17858 33756 17922 33760
rect 17858 33700 17862 33756
rect 17862 33700 17918 33756
rect 17918 33700 17922 33756
rect 17858 33696 17922 33700
rect 6868 33688 6932 33692
rect 6868 33632 6882 33688
rect 6882 33632 6932 33688
rect 6868 33628 6932 33632
rect 16988 33552 17052 33556
rect 16988 33496 17038 33552
rect 17038 33496 17052 33552
rect 16988 33492 17052 33496
rect 16620 33356 16684 33420
rect 7618 33212 7682 33216
rect 7618 33156 7622 33212
rect 7622 33156 7678 33212
rect 7678 33156 7682 33212
rect 7618 33152 7682 33156
rect 7698 33212 7762 33216
rect 7698 33156 7702 33212
rect 7702 33156 7758 33212
rect 7758 33156 7762 33212
rect 7698 33152 7762 33156
rect 7778 33212 7842 33216
rect 7778 33156 7782 33212
rect 7782 33156 7838 33212
rect 7838 33156 7842 33212
rect 7778 33152 7842 33156
rect 7858 33212 7922 33216
rect 7858 33156 7862 33212
rect 7862 33156 7918 33212
rect 7918 33156 7922 33212
rect 7858 33152 7922 33156
rect 14285 33212 14349 33216
rect 14285 33156 14289 33212
rect 14289 33156 14345 33212
rect 14345 33156 14349 33212
rect 14285 33152 14349 33156
rect 14365 33212 14429 33216
rect 14365 33156 14369 33212
rect 14369 33156 14425 33212
rect 14425 33156 14429 33212
rect 14365 33152 14429 33156
rect 14445 33212 14509 33216
rect 14445 33156 14449 33212
rect 14449 33156 14505 33212
rect 14505 33156 14509 33212
rect 14445 33152 14509 33156
rect 14525 33212 14589 33216
rect 14525 33156 14529 33212
rect 14529 33156 14585 33212
rect 14585 33156 14589 33212
rect 14525 33152 14589 33156
rect 2636 33084 2700 33148
rect 11652 33084 11716 33148
rect 17356 33008 17420 33012
rect 17356 32952 17406 33008
rect 17406 32952 17420 33008
rect 17356 32948 17420 32952
rect 8156 32812 8220 32876
rect 17172 32872 17236 32876
rect 17172 32816 17186 32872
rect 17186 32816 17236 32872
rect 17172 32812 17236 32816
rect 4285 32668 4349 32672
rect 4285 32612 4289 32668
rect 4289 32612 4345 32668
rect 4345 32612 4349 32668
rect 4285 32608 4349 32612
rect 4365 32668 4429 32672
rect 4365 32612 4369 32668
rect 4369 32612 4425 32668
rect 4425 32612 4429 32668
rect 4365 32608 4429 32612
rect 4445 32668 4509 32672
rect 4445 32612 4449 32668
rect 4449 32612 4505 32668
rect 4505 32612 4509 32668
rect 4445 32608 4509 32612
rect 4525 32668 4589 32672
rect 4525 32612 4529 32668
rect 4529 32612 4585 32668
rect 4585 32612 4589 32668
rect 4525 32608 4589 32612
rect 10952 32668 11016 32672
rect 10952 32612 10956 32668
rect 10956 32612 11012 32668
rect 11012 32612 11016 32668
rect 10952 32608 11016 32612
rect 11032 32668 11096 32672
rect 11032 32612 11036 32668
rect 11036 32612 11092 32668
rect 11092 32612 11096 32668
rect 11032 32608 11096 32612
rect 11112 32668 11176 32672
rect 11112 32612 11116 32668
rect 11116 32612 11172 32668
rect 11172 32612 11176 32668
rect 11112 32608 11176 32612
rect 11192 32668 11256 32672
rect 11192 32612 11196 32668
rect 11196 32612 11252 32668
rect 11252 32612 11256 32668
rect 11192 32608 11256 32612
rect 17618 32668 17682 32672
rect 17618 32612 17622 32668
rect 17622 32612 17678 32668
rect 17678 32612 17682 32668
rect 17618 32608 17682 32612
rect 17698 32668 17762 32672
rect 17698 32612 17702 32668
rect 17702 32612 17758 32668
rect 17758 32612 17762 32668
rect 17698 32608 17762 32612
rect 17778 32668 17842 32672
rect 17778 32612 17782 32668
rect 17782 32612 17838 32668
rect 17838 32612 17842 32668
rect 17778 32608 17842 32612
rect 17858 32668 17922 32672
rect 17858 32612 17862 32668
rect 17862 32612 17918 32668
rect 17918 32612 17922 32668
rect 17858 32608 17922 32612
rect 7420 32540 7484 32604
rect 14964 32268 15028 32332
rect 7618 32124 7682 32128
rect 7618 32068 7622 32124
rect 7622 32068 7678 32124
rect 7678 32068 7682 32124
rect 7618 32064 7682 32068
rect 7698 32124 7762 32128
rect 7698 32068 7702 32124
rect 7702 32068 7758 32124
rect 7758 32068 7762 32124
rect 7698 32064 7762 32068
rect 7778 32124 7842 32128
rect 7778 32068 7782 32124
rect 7782 32068 7838 32124
rect 7838 32068 7842 32124
rect 7778 32064 7842 32068
rect 7858 32124 7922 32128
rect 7858 32068 7862 32124
rect 7862 32068 7918 32124
rect 7918 32068 7922 32124
rect 7858 32064 7922 32068
rect 14285 32124 14349 32128
rect 14285 32068 14289 32124
rect 14289 32068 14345 32124
rect 14345 32068 14349 32124
rect 14285 32064 14349 32068
rect 14365 32124 14429 32128
rect 14365 32068 14369 32124
rect 14369 32068 14425 32124
rect 14425 32068 14429 32124
rect 14365 32064 14429 32068
rect 14445 32124 14509 32128
rect 14445 32068 14449 32124
rect 14449 32068 14505 32124
rect 14505 32068 14509 32124
rect 14445 32064 14509 32068
rect 14525 32124 14589 32128
rect 14525 32068 14529 32124
rect 14529 32068 14585 32124
rect 14585 32068 14589 32124
rect 14525 32064 14589 32068
rect 13860 31860 13924 31924
rect 7052 31724 7116 31788
rect 4285 31580 4349 31584
rect 4285 31524 4289 31580
rect 4289 31524 4345 31580
rect 4345 31524 4349 31580
rect 4285 31520 4349 31524
rect 4365 31580 4429 31584
rect 4365 31524 4369 31580
rect 4369 31524 4425 31580
rect 4425 31524 4429 31580
rect 4365 31520 4429 31524
rect 4445 31580 4509 31584
rect 4445 31524 4449 31580
rect 4449 31524 4505 31580
rect 4505 31524 4509 31580
rect 4445 31520 4509 31524
rect 4525 31580 4589 31584
rect 4525 31524 4529 31580
rect 4529 31524 4585 31580
rect 4585 31524 4589 31580
rect 4525 31520 4589 31524
rect 10952 31580 11016 31584
rect 10952 31524 10956 31580
rect 10956 31524 11012 31580
rect 11012 31524 11016 31580
rect 10952 31520 11016 31524
rect 11032 31580 11096 31584
rect 11032 31524 11036 31580
rect 11036 31524 11092 31580
rect 11092 31524 11096 31580
rect 11032 31520 11096 31524
rect 11112 31580 11176 31584
rect 11112 31524 11116 31580
rect 11116 31524 11172 31580
rect 11172 31524 11176 31580
rect 11112 31520 11176 31524
rect 11192 31580 11256 31584
rect 11192 31524 11196 31580
rect 11196 31524 11252 31580
rect 11252 31524 11256 31580
rect 11192 31520 11256 31524
rect 17618 31580 17682 31584
rect 17618 31524 17622 31580
rect 17622 31524 17678 31580
rect 17678 31524 17682 31580
rect 17618 31520 17682 31524
rect 17698 31580 17762 31584
rect 17698 31524 17702 31580
rect 17702 31524 17758 31580
rect 17758 31524 17762 31580
rect 17698 31520 17762 31524
rect 17778 31580 17842 31584
rect 17778 31524 17782 31580
rect 17782 31524 17838 31580
rect 17838 31524 17842 31580
rect 17778 31520 17842 31524
rect 17858 31580 17922 31584
rect 17858 31524 17862 31580
rect 17862 31524 17918 31580
rect 17918 31524 17922 31580
rect 17858 31520 17922 31524
rect 10732 31376 10796 31380
rect 10732 31320 10782 31376
rect 10782 31320 10796 31376
rect 10732 31316 10796 31320
rect 7618 31036 7682 31040
rect 7618 30980 7622 31036
rect 7622 30980 7678 31036
rect 7678 30980 7682 31036
rect 7618 30976 7682 30980
rect 7698 31036 7762 31040
rect 7698 30980 7702 31036
rect 7702 30980 7758 31036
rect 7758 30980 7762 31036
rect 7698 30976 7762 30980
rect 7778 31036 7842 31040
rect 7778 30980 7782 31036
rect 7782 30980 7838 31036
rect 7838 30980 7842 31036
rect 7778 30976 7842 30980
rect 7858 31036 7922 31040
rect 7858 30980 7862 31036
rect 7862 30980 7918 31036
rect 7918 30980 7922 31036
rect 7858 30976 7922 30980
rect 14285 31036 14349 31040
rect 14285 30980 14289 31036
rect 14289 30980 14345 31036
rect 14345 30980 14349 31036
rect 14285 30976 14349 30980
rect 14365 31036 14429 31040
rect 14365 30980 14369 31036
rect 14369 30980 14425 31036
rect 14425 30980 14429 31036
rect 14365 30976 14429 30980
rect 14445 31036 14509 31040
rect 14445 30980 14449 31036
rect 14449 30980 14505 31036
rect 14505 30980 14509 31036
rect 14445 30976 14509 30980
rect 14525 31036 14589 31040
rect 14525 30980 14529 31036
rect 14529 30980 14585 31036
rect 14585 30980 14589 31036
rect 14525 30976 14589 30980
rect 14044 30636 14108 30700
rect 4285 30492 4349 30496
rect 4285 30436 4289 30492
rect 4289 30436 4345 30492
rect 4345 30436 4349 30492
rect 4285 30432 4349 30436
rect 4365 30492 4429 30496
rect 4365 30436 4369 30492
rect 4369 30436 4425 30492
rect 4425 30436 4429 30492
rect 4365 30432 4429 30436
rect 4445 30492 4509 30496
rect 4445 30436 4449 30492
rect 4449 30436 4505 30492
rect 4505 30436 4509 30492
rect 4445 30432 4509 30436
rect 4525 30492 4589 30496
rect 4525 30436 4529 30492
rect 4529 30436 4585 30492
rect 4585 30436 4589 30492
rect 4525 30432 4589 30436
rect 10952 30492 11016 30496
rect 10952 30436 10956 30492
rect 10956 30436 11012 30492
rect 11012 30436 11016 30492
rect 10952 30432 11016 30436
rect 11032 30492 11096 30496
rect 11032 30436 11036 30492
rect 11036 30436 11092 30492
rect 11092 30436 11096 30492
rect 11032 30432 11096 30436
rect 11112 30492 11176 30496
rect 11112 30436 11116 30492
rect 11116 30436 11172 30492
rect 11172 30436 11176 30492
rect 11112 30432 11176 30436
rect 11192 30492 11256 30496
rect 11192 30436 11196 30492
rect 11196 30436 11252 30492
rect 11252 30436 11256 30492
rect 11192 30432 11256 30436
rect 17618 30492 17682 30496
rect 17618 30436 17622 30492
rect 17622 30436 17678 30492
rect 17678 30436 17682 30492
rect 17618 30432 17682 30436
rect 17698 30492 17762 30496
rect 17698 30436 17702 30492
rect 17702 30436 17758 30492
rect 17758 30436 17762 30492
rect 17698 30432 17762 30436
rect 17778 30492 17842 30496
rect 17778 30436 17782 30492
rect 17782 30436 17838 30492
rect 17838 30436 17842 30492
rect 17778 30432 17842 30436
rect 17858 30492 17922 30496
rect 17858 30436 17862 30492
rect 17862 30436 17918 30492
rect 17918 30436 17922 30492
rect 17858 30432 17922 30436
rect 7618 29948 7682 29952
rect 7618 29892 7622 29948
rect 7622 29892 7678 29948
rect 7678 29892 7682 29948
rect 7618 29888 7682 29892
rect 7698 29948 7762 29952
rect 7698 29892 7702 29948
rect 7702 29892 7758 29948
rect 7758 29892 7762 29948
rect 7698 29888 7762 29892
rect 7778 29948 7842 29952
rect 7778 29892 7782 29948
rect 7782 29892 7838 29948
rect 7838 29892 7842 29948
rect 7778 29888 7842 29892
rect 7858 29948 7922 29952
rect 7858 29892 7862 29948
rect 7862 29892 7918 29948
rect 7918 29892 7922 29948
rect 7858 29888 7922 29892
rect 14285 29948 14349 29952
rect 14285 29892 14289 29948
rect 14289 29892 14345 29948
rect 14345 29892 14349 29948
rect 14285 29888 14349 29892
rect 14365 29948 14429 29952
rect 14365 29892 14369 29948
rect 14369 29892 14425 29948
rect 14425 29892 14429 29948
rect 14365 29888 14429 29892
rect 14445 29948 14509 29952
rect 14445 29892 14449 29948
rect 14449 29892 14505 29948
rect 14505 29892 14509 29948
rect 14445 29888 14509 29892
rect 14525 29948 14589 29952
rect 14525 29892 14529 29948
rect 14529 29892 14585 29948
rect 14585 29892 14589 29948
rect 14525 29888 14589 29892
rect 12020 29684 12084 29748
rect 4285 29404 4349 29408
rect 4285 29348 4289 29404
rect 4289 29348 4345 29404
rect 4345 29348 4349 29404
rect 4285 29344 4349 29348
rect 4365 29404 4429 29408
rect 4365 29348 4369 29404
rect 4369 29348 4425 29404
rect 4425 29348 4429 29404
rect 4365 29344 4429 29348
rect 4445 29404 4509 29408
rect 4445 29348 4449 29404
rect 4449 29348 4505 29404
rect 4505 29348 4509 29404
rect 4445 29344 4509 29348
rect 4525 29404 4589 29408
rect 4525 29348 4529 29404
rect 4529 29348 4585 29404
rect 4585 29348 4589 29404
rect 4525 29344 4589 29348
rect 10952 29404 11016 29408
rect 10952 29348 10956 29404
rect 10956 29348 11012 29404
rect 11012 29348 11016 29404
rect 10952 29344 11016 29348
rect 11032 29404 11096 29408
rect 11032 29348 11036 29404
rect 11036 29348 11092 29404
rect 11092 29348 11096 29404
rect 11032 29344 11096 29348
rect 11112 29404 11176 29408
rect 11112 29348 11116 29404
rect 11116 29348 11172 29404
rect 11172 29348 11176 29404
rect 11112 29344 11176 29348
rect 11192 29404 11256 29408
rect 11192 29348 11196 29404
rect 11196 29348 11252 29404
rect 11252 29348 11256 29404
rect 11192 29344 11256 29348
rect 17618 29404 17682 29408
rect 17618 29348 17622 29404
rect 17622 29348 17678 29404
rect 17678 29348 17682 29404
rect 17618 29344 17682 29348
rect 17698 29404 17762 29408
rect 17698 29348 17702 29404
rect 17702 29348 17758 29404
rect 17758 29348 17762 29404
rect 17698 29344 17762 29348
rect 17778 29404 17842 29408
rect 17778 29348 17782 29404
rect 17782 29348 17838 29404
rect 17838 29348 17842 29404
rect 17778 29344 17842 29348
rect 17858 29404 17922 29408
rect 17858 29348 17862 29404
rect 17862 29348 17918 29404
rect 17918 29348 17922 29404
rect 17858 29344 17922 29348
rect 8340 29140 8404 29204
rect 7618 28860 7682 28864
rect 7618 28804 7622 28860
rect 7622 28804 7678 28860
rect 7678 28804 7682 28860
rect 7618 28800 7682 28804
rect 7698 28860 7762 28864
rect 7698 28804 7702 28860
rect 7702 28804 7758 28860
rect 7758 28804 7762 28860
rect 7698 28800 7762 28804
rect 7778 28860 7842 28864
rect 7778 28804 7782 28860
rect 7782 28804 7838 28860
rect 7838 28804 7842 28860
rect 7778 28800 7842 28804
rect 7858 28860 7922 28864
rect 7858 28804 7862 28860
rect 7862 28804 7918 28860
rect 7918 28804 7922 28860
rect 7858 28800 7922 28804
rect 11468 28928 11532 28932
rect 11468 28872 11518 28928
rect 11518 28872 11532 28928
rect 11468 28868 11532 28872
rect 14285 28860 14349 28864
rect 14285 28804 14289 28860
rect 14289 28804 14345 28860
rect 14345 28804 14349 28860
rect 14285 28800 14349 28804
rect 14365 28860 14429 28864
rect 14365 28804 14369 28860
rect 14369 28804 14425 28860
rect 14425 28804 14429 28860
rect 14365 28800 14429 28804
rect 14445 28860 14509 28864
rect 14445 28804 14449 28860
rect 14449 28804 14505 28860
rect 14505 28804 14509 28860
rect 14445 28800 14509 28804
rect 14525 28860 14589 28864
rect 14525 28804 14529 28860
rect 14529 28804 14585 28860
rect 14585 28804 14589 28860
rect 14525 28800 14589 28804
rect 4285 28316 4349 28320
rect 4285 28260 4289 28316
rect 4289 28260 4345 28316
rect 4345 28260 4349 28316
rect 4285 28256 4349 28260
rect 4365 28316 4429 28320
rect 4365 28260 4369 28316
rect 4369 28260 4425 28316
rect 4425 28260 4429 28316
rect 4365 28256 4429 28260
rect 4445 28316 4509 28320
rect 4445 28260 4449 28316
rect 4449 28260 4505 28316
rect 4505 28260 4509 28316
rect 4445 28256 4509 28260
rect 4525 28316 4589 28320
rect 4525 28260 4529 28316
rect 4529 28260 4585 28316
rect 4585 28260 4589 28316
rect 4525 28256 4589 28260
rect 10952 28316 11016 28320
rect 10952 28260 10956 28316
rect 10956 28260 11012 28316
rect 11012 28260 11016 28316
rect 10952 28256 11016 28260
rect 11032 28316 11096 28320
rect 11032 28260 11036 28316
rect 11036 28260 11092 28316
rect 11092 28260 11096 28316
rect 11032 28256 11096 28260
rect 11112 28316 11176 28320
rect 11112 28260 11116 28316
rect 11116 28260 11172 28316
rect 11172 28260 11176 28316
rect 11112 28256 11176 28260
rect 11192 28316 11256 28320
rect 11192 28260 11196 28316
rect 11196 28260 11252 28316
rect 11252 28260 11256 28316
rect 11192 28256 11256 28260
rect 17618 28316 17682 28320
rect 17618 28260 17622 28316
rect 17622 28260 17678 28316
rect 17678 28260 17682 28316
rect 17618 28256 17682 28260
rect 17698 28316 17762 28320
rect 17698 28260 17702 28316
rect 17702 28260 17758 28316
rect 17758 28260 17762 28316
rect 17698 28256 17762 28260
rect 17778 28316 17842 28320
rect 17778 28260 17782 28316
rect 17782 28260 17838 28316
rect 17838 28260 17842 28316
rect 17778 28256 17842 28260
rect 17858 28316 17922 28320
rect 17858 28260 17862 28316
rect 17862 28260 17918 28316
rect 17918 28260 17922 28316
rect 17858 28256 17922 28260
rect 7618 27772 7682 27776
rect 7618 27716 7622 27772
rect 7622 27716 7678 27772
rect 7678 27716 7682 27772
rect 7618 27712 7682 27716
rect 7698 27772 7762 27776
rect 7698 27716 7702 27772
rect 7702 27716 7758 27772
rect 7758 27716 7762 27772
rect 7698 27712 7762 27716
rect 7778 27772 7842 27776
rect 7778 27716 7782 27772
rect 7782 27716 7838 27772
rect 7838 27716 7842 27772
rect 7778 27712 7842 27716
rect 7858 27772 7922 27776
rect 7858 27716 7862 27772
rect 7862 27716 7918 27772
rect 7918 27716 7922 27772
rect 7858 27712 7922 27716
rect 14285 27772 14349 27776
rect 14285 27716 14289 27772
rect 14289 27716 14345 27772
rect 14345 27716 14349 27772
rect 14285 27712 14349 27716
rect 14365 27772 14429 27776
rect 14365 27716 14369 27772
rect 14369 27716 14425 27772
rect 14425 27716 14429 27772
rect 14365 27712 14429 27716
rect 14445 27772 14509 27776
rect 14445 27716 14449 27772
rect 14449 27716 14505 27772
rect 14505 27716 14509 27772
rect 14445 27712 14509 27716
rect 14525 27772 14589 27776
rect 14525 27716 14529 27772
rect 14529 27716 14585 27772
rect 14585 27716 14589 27772
rect 14525 27712 14589 27716
rect 4285 27228 4349 27232
rect 4285 27172 4289 27228
rect 4289 27172 4345 27228
rect 4345 27172 4349 27228
rect 4285 27168 4349 27172
rect 4365 27228 4429 27232
rect 4365 27172 4369 27228
rect 4369 27172 4425 27228
rect 4425 27172 4429 27228
rect 4365 27168 4429 27172
rect 4445 27228 4509 27232
rect 4445 27172 4449 27228
rect 4449 27172 4505 27228
rect 4505 27172 4509 27228
rect 4445 27168 4509 27172
rect 4525 27228 4589 27232
rect 4525 27172 4529 27228
rect 4529 27172 4585 27228
rect 4585 27172 4589 27228
rect 4525 27168 4589 27172
rect 10952 27228 11016 27232
rect 10952 27172 10956 27228
rect 10956 27172 11012 27228
rect 11012 27172 11016 27228
rect 10952 27168 11016 27172
rect 11032 27228 11096 27232
rect 11032 27172 11036 27228
rect 11036 27172 11092 27228
rect 11092 27172 11096 27228
rect 11032 27168 11096 27172
rect 11112 27228 11176 27232
rect 11112 27172 11116 27228
rect 11116 27172 11172 27228
rect 11172 27172 11176 27228
rect 11112 27168 11176 27172
rect 11192 27228 11256 27232
rect 11192 27172 11196 27228
rect 11196 27172 11252 27228
rect 11252 27172 11256 27228
rect 11192 27168 11256 27172
rect 17618 27228 17682 27232
rect 17618 27172 17622 27228
rect 17622 27172 17678 27228
rect 17678 27172 17682 27228
rect 17618 27168 17682 27172
rect 17698 27228 17762 27232
rect 17698 27172 17702 27228
rect 17702 27172 17758 27228
rect 17758 27172 17762 27228
rect 17698 27168 17762 27172
rect 17778 27228 17842 27232
rect 17778 27172 17782 27228
rect 17782 27172 17838 27228
rect 17838 27172 17842 27228
rect 17778 27168 17842 27172
rect 17858 27228 17922 27232
rect 17858 27172 17862 27228
rect 17862 27172 17918 27228
rect 17918 27172 17922 27228
rect 17858 27168 17922 27172
rect 7618 26684 7682 26688
rect 7618 26628 7622 26684
rect 7622 26628 7678 26684
rect 7678 26628 7682 26684
rect 7618 26624 7682 26628
rect 7698 26684 7762 26688
rect 7698 26628 7702 26684
rect 7702 26628 7758 26684
rect 7758 26628 7762 26684
rect 7698 26624 7762 26628
rect 7778 26684 7842 26688
rect 7778 26628 7782 26684
rect 7782 26628 7838 26684
rect 7838 26628 7842 26684
rect 7778 26624 7842 26628
rect 7858 26684 7922 26688
rect 7858 26628 7862 26684
rect 7862 26628 7918 26684
rect 7918 26628 7922 26684
rect 7858 26624 7922 26628
rect 14285 26684 14349 26688
rect 14285 26628 14289 26684
rect 14289 26628 14345 26684
rect 14345 26628 14349 26684
rect 14285 26624 14349 26628
rect 14365 26684 14429 26688
rect 14365 26628 14369 26684
rect 14369 26628 14425 26684
rect 14425 26628 14429 26684
rect 14365 26624 14429 26628
rect 14445 26684 14509 26688
rect 14445 26628 14449 26684
rect 14449 26628 14505 26684
rect 14505 26628 14509 26684
rect 14445 26624 14509 26628
rect 14525 26684 14589 26688
rect 14525 26628 14529 26684
rect 14529 26628 14585 26684
rect 14585 26628 14589 26684
rect 14525 26624 14589 26628
rect 5396 26556 5460 26620
rect 9628 26420 9692 26484
rect 4285 26140 4349 26144
rect 4285 26084 4289 26140
rect 4289 26084 4345 26140
rect 4345 26084 4349 26140
rect 4285 26080 4349 26084
rect 4365 26140 4429 26144
rect 4365 26084 4369 26140
rect 4369 26084 4425 26140
rect 4425 26084 4429 26140
rect 4365 26080 4429 26084
rect 4445 26140 4509 26144
rect 4445 26084 4449 26140
rect 4449 26084 4505 26140
rect 4505 26084 4509 26140
rect 4445 26080 4509 26084
rect 4525 26140 4589 26144
rect 4525 26084 4529 26140
rect 4529 26084 4585 26140
rect 4585 26084 4589 26140
rect 4525 26080 4589 26084
rect 10952 26140 11016 26144
rect 10952 26084 10956 26140
rect 10956 26084 11012 26140
rect 11012 26084 11016 26140
rect 10952 26080 11016 26084
rect 11032 26140 11096 26144
rect 11032 26084 11036 26140
rect 11036 26084 11092 26140
rect 11092 26084 11096 26140
rect 11032 26080 11096 26084
rect 11112 26140 11176 26144
rect 11112 26084 11116 26140
rect 11116 26084 11172 26140
rect 11172 26084 11176 26140
rect 11112 26080 11176 26084
rect 11192 26140 11256 26144
rect 11192 26084 11196 26140
rect 11196 26084 11252 26140
rect 11252 26084 11256 26140
rect 11192 26080 11256 26084
rect 17618 26140 17682 26144
rect 17618 26084 17622 26140
rect 17622 26084 17678 26140
rect 17678 26084 17682 26140
rect 17618 26080 17682 26084
rect 17698 26140 17762 26144
rect 17698 26084 17702 26140
rect 17702 26084 17758 26140
rect 17758 26084 17762 26140
rect 17698 26080 17762 26084
rect 17778 26140 17842 26144
rect 17778 26084 17782 26140
rect 17782 26084 17838 26140
rect 17838 26084 17842 26140
rect 17778 26080 17842 26084
rect 17858 26140 17922 26144
rect 17858 26084 17862 26140
rect 17862 26084 17918 26140
rect 17918 26084 17922 26140
rect 17858 26080 17922 26084
rect 7618 25596 7682 25600
rect 7618 25540 7622 25596
rect 7622 25540 7678 25596
rect 7678 25540 7682 25596
rect 7618 25536 7682 25540
rect 7698 25596 7762 25600
rect 7698 25540 7702 25596
rect 7702 25540 7758 25596
rect 7758 25540 7762 25596
rect 7698 25536 7762 25540
rect 7778 25596 7842 25600
rect 7778 25540 7782 25596
rect 7782 25540 7838 25596
rect 7838 25540 7842 25596
rect 7778 25536 7842 25540
rect 7858 25596 7922 25600
rect 7858 25540 7862 25596
rect 7862 25540 7918 25596
rect 7918 25540 7922 25596
rect 7858 25536 7922 25540
rect 14285 25596 14349 25600
rect 14285 25540 14289 25596
rect 14289 25540 14345 25596
rect 14345 25540 14349 25596
rect 14285 25536 14349 25540
rect 14365 25596 14429 25600
rect 14365 25540 14369 25596
rect 14369 25540 14425 25596
rect 14425 25540 14429 25596
rect 14365 25536 14429 25540
rect 14445 25596 14509 25600
rect 14445 25540 14449 25596
rect 14449 25540 14505 25596
rect 14505 25540 14509 25596
rect 14445 25536 14509 25540
rect 14525 25596 14589 25600
rect 14525 25540 14529 25596
rect 14529 25540 14585 25596
rect 14585 25540 14589 25596
rect 14525 25536 14589 25540
rect 4285 25052 4349 25056
rect 4285 24996 4289 25052
rect 4289 24996 4345 25052
rect 4345 24996 4349 25052
rect 4285 24992 4349 24996
rect 4365 25052 4429 25056
rect 4365 24996 4369 25052
rect 4369 24996 4425 25052
rect 4425 24996 4429 25052
rect 4365 24992 4429 24996
rect 4445 25052 4509 25056
rect 4445 24996 4449 25052
rect 4449 24996 4505 25052
rect 4505 24996 4509 25052
rect 4445 24992 4509 24996
rect 4525 25052 4589 25056
rect 4525 24996 4529 25052
rect 4529 24996 4585 25052
rect 4585 24996 4589 25052
rect 4525 24992 4589 24996
rect 10952 25052 11016 25056
rect 10952 24996 10956 25052
rect 10956 24996 11012 25052
rect 11012 24996 11016 25052
rect 10952 24992 11016 24996
rect 11032 25052 11096 25056
rect 11032 24996 11036 25052
rect 11036 24996 11092 25052
rect 11092 24996 11096 25052
rect 11032 24992 11096 24996
rect 11112 25052 11176 25056
rect 11112 24996 11116 25052
rect 11116 24996 11172 25052
rect 11172 24996 11176 25052
rect 11112 24992 11176 24996
rect 11192 25052 11256 25056
rect 11192 24996 11196 25052
rect 11196 24996 11252 25052
rect 11252 24996 11256 25052
rect 11192 24992 11256 24996
rect 17618 25052 17682 25056
rect 17618 24996 17622 25052
rect 17622 24996 17678 25052
rect 17678 24996 17682 25052
rect 17618 24992 17682 24996
rect 17698 25052 17762 25056
rect 17698 24996 17702 25052
rect 17702 24996 17758 25052
rect 17758 24996 17762 25052
rect 17698 24992 17762 24996
rect 17778 25052 17842 25056
rect 17778 24996 17782 25052
rect 17782 24996 17838 25052
rect 17838 24996 17842 25052
rect 17778 24992 17842 24996
rect 17858 25052 17922 25056
rect 17858 24996 17862 25052
rect 17862 24996 17918 25052
rect 17918 24996 17922 25052
rect 17858 24992 17922 24996
rect 7618 24508 7682 24512
rect 7618 24452 7622 24508
rect 7622 24452 7678 24508
rect 7678 24452 7682 24508
rect 7618 24448 7682 24452
rect 7698 24508 7762 24512
rect 7698 24452 7702 24508
rect 7702 24452 7758 24508
rect 7758 24452 7762 24508
rect 7698 24448 7762 24452
rect 7778 24508 7842 24512
rect 7778 24452 7782 24508
rect 7782 24452 7838 24508
rect 7838 24452 7842 24508
rect 7778 24448 7842 24452
rect 7858 24508 7922 24512
rect 7858 24452 7862 24508
rect 7862 24452 7918 24508
rect 7918 24452 7922 24508
rect 7858 24448 7922 24452
rect 14285 24508 14349 24512
rect 14285 24452 14289 24508
rect 14289 24452 14345 24508
rect 14345 24452 14349 24508
rect 14285 24448 14349 24452
rect 14365 24508 14429 24512
rect 14365 24452 14369 24508
rect 14369 24452 14425 24508
rect 14425 24452 14429 24508
rect 14365 24448 14429 24452
rect 14445 24508 14509 24512
rect 14445 24452 14449 24508
rect 14449 24452 14505 24508
rect 14505 24452 14509 24508
rect 14445 24448 14509 24452
rect 14525 24508 14589 24512
rect 14525 24452 14529 24508
rect 14529 24452 14585 24508
rect 14585 24452 14589 24508
rect 14525 24448 14589 24452
rect 10548 24244 10612 24308
rect 4285 23964 4349 23968
rect 4285 23908 4289 23964
rect 4289 23908 4345 23964
rect 4345 23908 4349 23964
rect 4285 23904 4349 23908
rect 4365 23964 4429 23968
rect 4365 23908 4369 23964
rect 4369 23908 4425 23964
rect 4425 23908 4429 23964
rect 4365 23904 4429 23908
rect 4445 23964 4509 23968
rect 4445 23908 4449 23964
rect 4449 23908 4505 23964
rect 4505 23908 4509 23964
rect 4445 23904 4509 23908
rect 4525 23964 4589 23968
rect 4525 23908 4529 23964
rect 4529 23908 4585 23964
rect 4585 23908 4589 23964
rect 4525 23904 4589 23908
rect 10952 23964 11016 23968
rect 10952 23908 10956 23964
rect 10956 23908 11012 23964
rect 11012 23908 11016 23964
rect 10952 23904 11016 23908
rect 11032 23964 11096 23968
rect 11032 23908 11036 23964
rect 11036 23908 11092 23964
rect 11092 23908 11096 23964
rect 11032 23904 11096 23908
rect 11112 23964 11176 23968
rect 11112 23908 11116 23964
rect 11116 23908 11172 23964
rect 11172 23908 11176 23964
rect 11112 23904 11176 23908
rect 11192 23964 11256 23968
rect 11192 23908 11196 23964
rect 11196 23908 11252 23964
rect 11252 23908 11256 23964
rect 11192 23904 11256 23908
rect 17618 23964 17682 23968
rect 17618 23908 17622 23964
rect 17622 23908 17678 23964
rect 17678 23908 17682 23964
rect 17618 23904 17682 23908
rect 17698 23964 17762 23968
rect 17698 23908 17702 23964
rect 17702 23908 17758 23964
rect 17758 23908 17762 23964
rect 17698 23904 17762 23908
rect 17778 23964 17842 23968
rect 17778 23908 17782 23964
rect 17782 23908 17838 23964
rect 17838 23908 17842 23964
rect 17778 23904 17842 23908
rect 17858 23964 17922 23968
rect 17858 23908 17862 23964
rect 17862 23908 17918 23964
rect 17918 23908 17922 23964
rect 17858 23904 17922 23908
rect 7618 23420 7682 23424
rect 7618 23364 7622 23420
rect 7622 23364 7678 23420
rect 7678 23364 7682 23420
rect 7618 23360 7682 23364
rect 7698 23420 7762 23424
rect 7698 23364 7702 23420
rect 7702 23364 7758 23420
rect 7758 23364 7762 23420
rect 7698 23360 7762 23364
rect 7778 23420 7842 23424
rect 7778 23364 7782 23420
rect 7782 23364 7838 23420
rect 7838 23364 7842 23420
rect 7778 23360 7842 23364
rect 7858 23420 7922 23424
rect 7858 23364 7862 23420
rect 7862 23364 7918 23420
rect 7918 23364 7922 23420
rect 7858 23360 7922 23364
rect 14285 23420 14349 23424
rect 14285 23364 14289 23420
rect 14289 23364 14345 23420
rect 14345 23364 14349 23420
rect 14285 23360 14349 23364
rect 14365 23420 14429 23424
rect 14365 23364 14369 23420
rect 14369 23364 14425 23420
rect 14425 23364 14429 23420
rect 14365 23360 14429 23364
rect 14445 23420 14509 23424
rect 14445 23364 14449 23420
rect 14449 23364 14505 23420
rect 14505 23364 14509 23420
rect 14445 23360 14509 23364
rect 14525 23420 14589 23424
rect 14525 23364 14529 23420
rect 14529 23364 14585 23420
rect 14585 23364 14589 23420
rect 14525 23360 14589 23364
rect 4285 22876 4349 22880
rect 4285 22820 4289 22876
rect 4289 22820 4345 22876
rect 4345 22820 4349 22876
rect 4285 22816 4349 22820
rect 4365 22876 4429 22880
rect 4365 22820 4369 22876
rect 4369 22820 4425 22876
rect 4425 22820 4429 22876
rect 4365 22816 4429 22820
rect 4445 22876 4509 22880
rect 4445 22820 4449 22876
rect 4449 22820 4505 22876
rect 4505 22820 4509 22876
rect 4445 22816 4509 22820
rect 4525 22876 4589 22880
rect 4525 22820 4529 22876
rect 4529 22820 4585 22876
rect 4585 22820 4589 22876
rect 4525 22816 4589 22820
rect 10952 22876 11016 22880
rect 10952 22820 10956 22876
rect 10956 22820 11012 22876
rect 11012 22820 11016 22876
rect 10952 22816 11016 22820
rect 11032 22876 11096 22880
rect 11032 22820 11036 22876
rect 11036 22820 11092 22876
rect 11092 22820 11096 22876
rect 11032 22816 11096 22820
rect 11112 22876 11176 22880
rect 11112 22820 11116 22876
rect 11116 22820 11172 22876
rect 11172 22820 11176 22876
rect 11112 22816 11176 22820
rect 11192 22876 11256 22880
rect 11192 22820 11196 22876
rect 11196 22820 11252 22876
rect 11252 22820 11256 22876
rect 11192 22816 11256 22820
rect 17618 22876 17682 22880
rect 17618 22820 17622 22876
rect 17622 22820 17678 22876
rect 17678 22820 17682 22876
rect 17618 22816 17682 22820
rect 17698 22876 17762 22880
rect 17698 22820 17702 22876
rect 17702 22820 17758 22876
rect 17758 22820 17762 22876
rect 17698 22816 17762 22820
rect 17778 22876 17842 22880
rect 17778 22820 17782 22876
rect 17782 22820 17838 22876
rect 17838 22820 17842 22876
rect 17778 22816 17842 22820
rect 17858 22876 17922 22880
rect 17858 22820 17862 22876
rect 17862 22820 17918 22876
rect 17918 22820 17922 22876
rect 17858 22816 17922 22820
rect 11468 22672 11532 22676
rect 11468 22616 11482 22672
rect 11482 22616 11532 22672
rect 11468 22612 11532 22616
rect 7618 22332 7682 22336
rect 7618 22276 7622 22332
rect 7622 22276 7678 22332
rect 7678 22276 7682 22332
rect 7618 22272 7682 22276
rect 7698 22332 7762 22336
rect 7698 22276 7702 22332
rect 7702 22276 7758 22332
rect 7758 22276 7762 22332
rect 7698 22272 7762 22276
rect 7778 22332 7842 22336
rect 7778 22276 7782 22332
rect 7782 22276 7838 22332
rect 7838 22276 7842 22332
rect 7778 22272 7842 22276
rect 7858 22332 7922 22336
rect 7858 22276 7862 22332
rect 7862 22276 7918 22332
rect 7918 22276 7922 22332
rect 7858 22272 7922 22276
rect 14285 22332 14349 22336
rect 14285 22276 14289 22332
rect 14289 22276 14345 22332
rect 14345 22276 14349 22332
rect 14285 22272 14349 22276
rect 14365 22332 14429 22336
rect 14365 22276 14369 22332
rect 14369 22276 14425 22332
rect 14425 22276 14429 22332
rect 14365 22272 14429 22276
rect 14445 22332 14509 22336
rect 14445 22276 14449 22332
rect 14449 22276 14505 22332
rect 14505 22276 14509 22332
rect 14445 22272 14509 22276
rect 14525 22332 14589 22336
rect 14525 22276 14529 22332
rect 14529 22276 14585 22332
rect 14585 22276 14589 22332
rect 14525 22272 14589 22276
rect 4285 21788 4349 21792
rect 4285 21732 4289 21788
rect 4289 21732 4345 21788
rect 4345 21732 4349 21788
rect 4285 21728 4349 21732
rect 4365 21788 4429 21792
rect 4365 21732 4369 21788
rect 4369 21732 4425 21788
rect 4425 21732 4429 21788
rect 4365 21728 4429 21732
rect 4445 21788 4509 21792
rect 4445 21732 4449 21788
rect 4449 21732 4505 21788
rect 4505 21732 4509 21788
rect 4445 21728 4509 21732
rect 4525 21788 4589 21792
rect 4525 21732 4529 21788
rect 4529 21732 4585 21788
rect 4585 21732 4589 21788
rect 4525 21728 4589 21732
rect 10952 21788 11016 21792
rect 10952 21732 10956 21788
rect 10956 21732 11012 21788
rect 11012 21732 11016 21788
rect 10952 21728 11016 21732
rect 11032 21788 11096 21792
rect 11032 21732 11036 21788
rect 11036 21732 11092 21788
rect 11092 21732 11096 21788
rect 11032 21728 11096 21732
rect 11112 21788 11176 21792
rect 11112 21732 11116 21788
rect 11116 21732 11172 21788
rect 11172 21732 11176 21788
rect 11112 21728 11176 21732
rect 11192 21788 11256 21792
rect 11192 21732 11196 21788
rect 11196 21732 11252 21788
rect 11252 21732 11256 21788
rect 11192 21728 11256 21732
rect 17618 21788 17682 21792
rect 17618 21732 17622 21788
rect 17622 21732 17678 21788
rect 17678 21732 17682 21788
rect 17618 21728 17682 21732
rect 17698 21788 17762 21792
rect 17698 21732 17702 21788
rect 17702 21732 17758 21788
rect 17758 21732 17762 21788
rect 17698 21728 17762 21732
rect 17778 21788 17842 21792
rect 17778 21732 17782 21788
rect 17782 21732 17838 21788
rect 17838 21732 17842 21788
rect 17778 21728 17842 21732
rect 17858 21788 17922 21792
rect 17858 21732 17862 21788
rect 17862 21732 17918 21788
rect 17918 21732 17922 21788
rect 17858 21728 17922 21732
rect 7618 21244 7682 21248
rect 7618 21188 7622 21244
rect 7622 21188 7678 21244
rect 7678 21188 7682 21244
rect 7618 21184 7682 21188
rect 7698 21244 7762 21248
rect 7698 21188 7702 21244
rect 7702 21188 7758 21244
rect 7758 21188 7762 21244
rect 7698 21184 7762 21188
rect 7778 21244 7842 21248
rect 7778 21188 7782 21244
rect 7782 21188 7838 21244
rect 7838 21188 7842 21244
rect 7778 21184 7842 21188
rect 7858 21244 7922 21248
rect 7858 21188 7862 21244
rect 7862 21188 7918 21244
rect 7918 21188 7922 21244
rect 7858 21184 7922 21188
rect 14285 21244 14349 21248
rect 14285 21188 14289 21244
rect 14289 21188 14345 21244
rect 14345 21188 14349 21244
rect 14285 21184 14349 21188
rect 14365 21244 14429 21248
rect 14365 21188 14369 21244
rect 14369 21188 14425 21244
rect 14425 21188 14429 21244
rect 14365 21184 14429 21188
rect 14445 21244 14509 21248
rect 14445 21188 14449 21244
rect 14449 21188 14505 21244
rect 14505 21188 14509 21244
rect 14445 21184 14509 21188
rect 14525 21244 14589 21248
rect 14525 21188 14529 21244
rect 14529 21188 14585 21244
rect 14585 21188 14589 21244
rect 14525 21184 14589 21188
rect 4285 20700 4349 20704
rect 4285 20644 4289 20700
rect 4289 20644 4345 20700
rect 4345 20644 4349 20700
rect 4285 20640 4349 20644
rect 4365 20700 4429 20704
rect 4365 20644 4369 20700
rect 4369 20644 4425 20700
rect 4425 20644 4429 20700
rect 4365 20640 4429 20644
rect 4445 20700 4509 20704
rect 4445 20644 4449 20700
rect 4449 20644 4505 20700
rect 4505 20644 4509 20700
rect 4445 20640 4509 20644
rect 4525 20700 4589 20704
rect 4525 20644 4529 20700
rect 4529 20644 4585 20700
rect 4585 20644 4589 20700
rect 4525 20640 4589 20644
rect 10952 20700 11016 20704
rect 10952 20644 10956 20700
rect 10956 20644 11012 20700
rect 11012 20644 11016 20700
rect 10952 20640 11016 20644
rect 11032 20700 11096 20704
rect 11032 20644 11036 20700
rect 11036 20644 11092 20700
rect 11092 20644 11096 20700
rect 11032 20640 11096 20644
rect 11112 20700 11176 20704
rect 11112 20644 11116 20700
rect 11116 20644 11172 20700
rect 11172 20644 11176 20700
rect 11112 20640 11176 20644
rect 11192 20700 11256 20704
rect 11192 20644 11196 20700
rect 11196 20644 11252 20700
rect 11252 20644 11256 20700
rect 11192 20640 11256 20644
rect 17618 20700 17682 20704
rect 17618 20644 17622 20700
rect 17622 20644 17678 20700
rect 17678 20644 17682 20700
rect 17618 20640 17682 20644
rect 17698 20700 17762 20704
rect 17698 20644 17702 20700
rect 17702 20644 17758 20700
rect 17758 20644 17762 20700
rect 17698 20640 17762 20644
rect 17778 20700 17842 20704
rect 17778 20644 17782 20700
rect 17782 20644 17838 20700
rect 17838 20644 17842 20700
rect 17778 20640 17842 20644
rect 17858 20700 17922 20704
rect 17858 20644 17862 20700
rect 17862 20644 17918 20700
rect 17918 20644 17922 20700
rect 17858 20640 17922 20644
rect 7618 20156 7682 20160
rect 7618 20100 7622 20156
rect 7622 20100 7678 20156
rect 7678 20100 7682 20156
rect 7618 20096 7682 20100
rect 7698 20156 7762 20160
rect 7698 20100 7702 20156
rect 7702 20100 7758 20156
rect 7758 20100 7762 20156
rect 7698 20096 7762 20100
rect 7778 20156 7842 20160
rect 7778 20100 7782 20156
rect 7782 20100 7838 20156
rect 7838 20100 7842 20156
rect 7778 20096 7842 20100
rect 7858 20156 7922 20160
rect 7858 20100 7862 20156
rect 7862 20100 7918 20156
rect 7918 20100 7922 20156
rect 7858 20096 7922 20100
rect 14285 20156 14349 20160
rect 14285 20100 14289 20156
rect 14289 20100 14345 20156
rect 14345 20100 14349 20156
rect 14285 20096 14349 20100
rect 14365 20156 14429 20160
rect 14365 20100 14369 20156
rect 14369 20100 14425 20156
rect 14425 20100 14429 20156
rect 14365 20096 14429 20100
rect 14445 20156 14509 20160
rect 14445 20100 14449 20156
rect 14449 20100 14505 20156
rect 14505 20100 14509 20156
rect 14445 20096 14509 20100
rect 14525 20156 14589 20160
rect 14525 20100 14529 20156
rect 14529 20100 14585 20156
rect 14585 20100 14589 20156
rect 14525 20096 14589 20100
rect 4285 19612 4349 19616
rect 4285 19556 4289 19612
rect 4289 19556 4345 19612
rect 4345 19556 4349 19612
rect 4285 19552 4349 19556
rect 4365 19612 4429 19616
rect 4365 19556 4369 19612
rect 4369 19556 4425 19612
rect 4425 19556 4429 19612
rect 4365 19552 4429 19556
rect 4445 19612 4509 19616
rect 4445 19556 4449 19612
rect 4449 19556 4505 19612
rect 4505 19556 4509 19612
rect 4445 19552 4509 19556
rect 4525 19612 4589 19616
rect 4525 19556 4529 19612
rect 4529 19556 4585 19612
rect 4585 19556 4589 19612
rect 4525 19552 4589 19556
rect 10952 19612 11016 19616
rect 10952 19556 10956 19612
rect 10956 19556 11012 19612
rect 11012 19556 11016 19612
rect 10952 19552 11016 19556
rect 11032 19612 11096 19616
rect 11032 19556 11036 19612
rect 11036 19556 11092 19612
rect 11092 19556 11096 19612
rect 11032 19552 11096 19556
rect 11112 19612 11176 19616
rect 11112 19556 11116 19612
rect 11116 19556 11172 19612
rect 11172 19556 11176 19612
rect 11112 19552 11176 19556
rect 11192 19612 11256 19616
rect 11192 19556 11196 19612
rect 11196 19556 11252 19612
rect 11252 19556 11256 19612
rect 11192 19552 11256 19556
rect 17618 19612 17682 19616
rect 17618 19556 17622 19612
rect 17622 19556 17678 19612
rect 17678 19556 17682 19612
rect 17618 19552 17682 19556
rect 17698 19612 17762 19616
rect 17698 19556 17702 19612
rect 17702 19556 17758 19612
rect 17758 19556 17762 19612
rect 17698 19552 17762 19556
rect 17778 19612 17842 19616
rect 17778 19556 17782 19612
rect 17782 19556 17838 19612
rect 17838 19556 17842 19612
rect 17778 19552 17842 19556
rect 17858 19612 17922 19616
rect 17858 19556 17862 19612
rect 17862 19556 17918 19612
rect 17918 19556 17922 19612
rect 17858 19552 17922 19556
rect 7618 19068 7682 19072
rect 7618 19012 7622 19068
rect 7622 19012 7678 19068
rect 7678 19012 7682 19068
rect 7618 19008 7682 19012
rect 7698 19068 7762 19072
rect 7698 19012 7702 19068
rect 7702 19012 7758 19068
rect 7758 19012 7762 19068
rect 7698 19008 7762 19012
rect 7778 19068 7842 19072
rect 7778 19012 7782 19068
rect 7782 19012 7838 19068
rect 7838 19012 7842 19068
rect 7778 19008 7842 19012
rect 7858 19068 7922 19072
rect 7858 19012 7862 19068
rect 7862 19012 7918 19068
rect 7918 19012 7922 19068
rect 7858 19008 7922 19012
rect 14285 19068 14349 19072
rect 14285 19012 14289 19068
rect 14289 19012 14345 19068
rect 14345 19012 14349 19068
rect 14285 19008 14349 19012
rect 14365 19068 14429 19072
rect 14365 19012 14369 19068
rect 14369 19012 14425 19068
rect 14425 19012 14429 19068
rect 14365 19008 14429 19012
rect 14445 19068 14509 19072
rect 14445 19012 14449 19068
rect 14449 19012 14505 19068
rect 14505 19012 14509 19068
rect 14445 19008 14509 19012
rect 14525 19068 14589 19072
rect 14525 19012 14529 19068
rect 14529 19012 14585 19068
rect 14585 19012 14589 19068
rect 14525 19008 14589 19012
rect 4285 18524 4349 18528
rect 4285 18468 4289 18524
rect 4289 18468 4345 18524
rect 4345 18468 4349 18524
rect 4285 18464 4349 18468
rect 4365 18524 4429 18528
rect 4365 18468 4369 18524
rect 4369 18468 4425 18524
rect 4425 18468 4429 18524
rect 4365 18464 4429 18468
rect 4445 18524 4509 18528
rect 4445 18468 4449 18524
rect 4449 18468 4505 18524
rect 4505 18468 4509 18524
rect 4445 18464 4509 18468
rect 4525 18524 4589 18528
rect 4525 18468 4529 18524
rect 4529 18468 4585 18524
rect 4585 18468 4589 18524
rect 4525 18464 4589 18468
rect 10952 18524 11016 18528
rect 10952 18468 10956 18524
rect 10956 18468 11012 18524
rect 11012 18468 11016 18524
rect 10952 18464 11016 18468
rect 11032 18524 11096 18528
rect 11032 18468 11036 18524
rect 11036 18468 11092 18524
rect 11092 18468 11096 18524
rect 11032 18464 11096 18468
rect 11112 18524 11176 18528
rect 11112 18468 11116 18524
rect 11116 18468 11172 18524
rect 11172 18468 11176 18524
rect 11112 18464 11176 18468
rect 11192 18524 11256 18528
rect 11192 18468 11196 18524
rect 11196 18468 11252 18524
rect 11252 18468 11256 18524
rect 11192 18464 11256 18468
rect 17618 18524 17682 18528
rect 17618 18468 17622 18524
rect 17622 18468 17678 18524
rect 17678 18468 17682 18524
rect 17618 18464 17682 18468
rect 17698 18524 17762 18528
rect 17698 18468 17702 18524
rect 17702 18468 17758 18524
rect 17758 18468 17762 18524
rect 17698 18464 17762 18468
rect 17778 18524 17842 18528
rect 17778 18468 17782 18524
rect 17782 18468 17838 18524
rect 17838 18468 17842 18524
rect 17778 18464 17842 18468
rect 17858 18524 17922 18528
rect 17858 18468 17862 18524
rect 17862 18468 17918 18524
rect 17918 18468 17922 18524
rect 17858 18464 17922 18468
rect 7618 17980 7682 17984
rect 7618 17924 7622 17980
rect 7622 17924 7678 17980
rect 7678 17924 7682 17980
rect 7618 17920 7682 17924
rect 7698 17980 7762 17984
rect 7698 17924 7702 17980
rect 7702 17924 7758 17980
rect 7758 17924 7762 17980
rect 7698 17920 7762 17924
rect 7778 17980 7842 17984
rect 7778 17924 7782 17980
rect 7782 17924 7838 17980
rect 7838 17924 7842 17980
rect 7778 17920 7842 17924
rect 7858 17980 7922 17984
rect 7858 17924 7862 17980
rect 7862 17924 7918 17980
rect 7918 17924 7922 17980
rect 7858 17920 7922 17924
rect 14285 17980 14349 17984
rect 14285 17924 14289 17980
rect 14289 17924 14345 17980
rect 14345 17924 14349 17980
rect 14285 17920 14349 17924
rect 14365 17980 14429 17984
rect 14365 17924 14369 17980
rect 14369 17924 14425 17980
rect 14425 17924 14429 17980
rect 14365 17920 14429 17924
rect 14445 17980 14509 17984
rect 14445 17924 14449 17980
rect 14449 17924 14505 17980
rect 14505 17924 14509 17980
rect 14445 17920 14509 17924
rect 14525 17980 14589 17984
rect 14525 17924 14529 17980
rect 14529 17924 14585 17980
rect 14585 17924 14589 17980
rect 14525 17920 14589 17924
rect 4285 17436 4349 17440
rect 4285 17380 4289 17436
rect 4289 17380 4345 17436
rect 4345 17380 4349 17436
rect 4285 17376 4349 17380
rect 4365 17436 4429 17440
rect 4365 17380 4369 17436
rect 4369 17380 4425 17436
rect 4425 17380 4429 17436
rect 4365 17376 4429 17380
rect 4445 17436 4509 17440
rect 4445 17380 4449 17436
rect 4449 17380 4505 17436
rect 4505 17380 4509 17436
rect 4445 17376 4509 17380
rect 4525 17436 4589 17440
rect 4525 17380 4529 17436
rect 4529 17380 4585 17436
rect 4585 17380 4589 17436
rect 4525 17376 4589 17380
rect 10952 17436 11016 17440
rect 10952 17380 10956 17436
rect 10956 17380 11012 17436
rect 11012 17380 11016 17436
rect 10952 17376 11016 17380
rect 11032 17436 11096 17440
rect 11032 17380 11036 17436
rect 11036 17380 11092 17436
rect 11092 17380 11096 17436
rect 11032 17376 11096 17380
rect 11112 17436 11176 17440
rect 11112 17380 11116 17436
rect 11116 17380 11172 17436
rect 11172 17380 11176 17436
rect 11112 17376 11176 17380
rect 11192 17436 11256 17440
rect 11192 17380 11196 17436
rect 11196 17380 11252 17436
rect 11252 17380 11256 17436
rect 11192 17376 11256 17380
rect 17618 17436 17682 17440
rect 17618 17380 17622 17436
rect 17622 17380 17678 17436
rect 17678 17380 17682 17436
rect 17618 17376 17682 17380
rect 17698 17436 17762 17440
rect 17698 17380 17702 17436
rect 17702 17380 17758 17436
rect 17758 17380 17762 17436
rect 17698 17376 17762 17380
rect 17778 17436 17842 17440
rect 17778 17380 17782 17436
rect 17782 17380 17838 17436
rect 17838 17380 17842 17436
rect 17778 17376 17842 17380
rect 17858 17436 17922 17440
rect 17858 17380 17862 17436
rect 17862 17380 17918 17436
rect 17918 17380 17922 17436
rect 17858 17376 17922 17380
rect 1716 17232 1780 17236
rect 1716 17176 1730 17232
rect 1730 17176 1780 17232
rect 1716 17172 1780 17176
rect 7618 16892 7682 16896
rect 7618 16836 7622 16892
rect 7622 16836 7678 16892
rect 7678 16836 7682 16892
rect 7618 16832 7682 16836
rect 7698 16892 7762 16896
rect 7698 16836 7702 16892
rect 7702 16836 7758 16892
rect 7758 16836 7762 16892
rect 7698 16832 7762 16836
rect 7778 16892 7842 16896
rect 7778 16836 7782 16892
rect 7782 16836 7838 16892
rect 7838 16836 7842 16892
rect 7778 16832 7842 16836
rect 7858 16892 7922 16896
rect 7858 16836 7862 16892
rect 7862 16836 7918 16892
rect 7918 16836 7922 16892
rect 7858 16832 7922 16836
rect 14285 16892 14349 16896
rect 14285 16836 14289 16892
rect 14289 16836 14345 16892
rect 14345 16836 14349 16892
rect 14285 16832 14349 16836
rect 14365 16892 14429 16896
rect 14365 16836 14369 16892
rect 14369 16836 14425 16892
rect 14425 16836 14429 16892
rect 14365 16832 14429 16836
rect 14445 16892 14509 16896
rect 14445 16836 14449 16892
rect 14449 16836 14505 16892
rect 14505 16836 14509 16892
rect 14445 16832 14509 16836
rect 14525 16892 14589 16896
rect 14525 16836 14529 16892
rect 14529 16836 14585 16892
rect 14585 16836 14589 16892
rect 14525 16832 14589 16836
rect 4285 16348 4349 16352
rect 4285 16292 4289 16348
rect 4289 16292 4345 16348
rect 4345 16292 4349 16348
rect 4285 16288 4349 16292
rect 4365 16348 4429 16352
rect 4365 16292 4369 16348
rect 4369 16292 4425 16348
rect 4425 16292 4429 16348
rect 4365 16288 4429 16292
rect 4445 16348 4509 16352
rect 4445 16292 4449 16348
rect 4449 16292 4505 16348
rect 4505 16292 4509 16348
rect 4445 16288 4509 16292
rect 4525 16348 4589 16352
rect 4525 16292 4529 16348
rect 4529 16292 4585 16348
rect 4585 16292 4589 16348
rect 4525 16288 4589 16292
rect 10952 16348 11016 16352
rect 10952 16292 10956 16348
rect 10956 16292 11012 16348
rect 11012 16292 11016 16348
rect 10952 16288 11016 16292
rect 11032 16348 11096 16352
rect 11032 16292 11036 16348
rect 11036 16292 11092 16348
rect 11092 16292 11096 16348
rect 11032 16288 11096 16292
rect 11112 16348 11176 16352
rect 11112 16292 11116 16348
rect 11116 16292 11172 16348
rect 11172 16292 11176 16348
rect 11112 16288 11176 16292
rect 11192 16348 11256 16352
rect 11192 16292 11196 16348
rect 11196 16292 11252 16348
rect 11252 16292 11256 16348
rect 11192 16288 11256 16292
rect 17618 16348 17682 16352
rect 17618 16292 17622 16348
rect 17622 16292 17678 16348
rect 17678 16292 17682 16348
rect 17618 16288 17682 16292
rect 17698 16348 17762 16352
rect 17698 16292 17702 16348
rect 17702 16292 17758 16348
rect 17758 16292 17762 16348
rect 17698 16288 17762 16292
rect 17778 16348 17842 16352
rect 17778 16292 17782 16348
rect 17782 16292 17838 16348
rect 17838 16292 17842 16348
rect 17778 16288 17842 16292
rect 17858 16348 17922 16352
rect 17858 16292 17862 16348
rect 17862 16292 17918 16348
rect 17918 16292 17922 16348
rect 17858 16288 17922 16292
rect 7618 15804 7682 15808
rect 7618 15748 7622 15804
rect 7622 15748 7678 15804
rect 7678 15748 7682 15804
rect 7618 15744 7682 15748
rect 7698 15804 7762 15808
rect 7698 15748 7702 15804
rect 7702 15748 7758 15804
rect 7758 15748 7762 15804
rect 7698 15744 7762 15748
rect 7778 15804 7842 15808
rect 7778 15748 7782 15804
rect 7782 15748 7838 15804
rect 7838 15748 7842 15804
rect 7778 15744 7842 15748
rect 7858 15804 7922 15808
rect 7858 15748 7862 15804
rect 7862 15748 7918 15804
rect 7918 15748 7922 15804
rect 7858 15744 7922 15748
rect 14285 15804 14349 15808
rect 14285 15748 14289 15804
rect 14289 15748 14345 15804
rect 14345 15748 14349 15804
rect 14285 15744 14349 15748
rect 14365 15804 14429 15808
rect 14365 15748 14369 15804
rect 14369 15748 14425 15804
rect 14425 15748 14429 15804
rect 14365 15744 14429 15748
rect 14445 15804 14509 15808
rect 14445 15748 14449 15804
rect 14449 15748 14505 15804
rect 14505 15748 14509 15804
rect 14445 15744 14509 15748
rect 14525 15804 14589 15808
rect 14525 15748 14529 15804
rect 14529 15748 14585 15804
rect 14585 15748 14589 15804
rect 14525 15744 14589 15748
rect 4285 15260 4349 15264
rect 4285 15204 4289 15260
rect 4289 15204 4345 15260
rect 4345 15204 4349 15260
rect 4285 15200 4349 15204
rect 4365 15260 4429 15264
rect 4365 15204 4369 15260
rect 4369 15204 4425 15260
rect 4425 15204 4429 15260
rect 4365 15200 4429 15204
rect 4445 15260 4509 15264
rect 4445 15204 4449 15260
rect 4449 15204 4505 15260
rect 4505 15204 4509 15260
rect 4445 15200 4509 15204
rect 4525 15260 4589 15264
rect 4525 15204 4529 15260
rect 4529 15204 4585 15260
rect 4585 15204 4589 15260
rect 4525 15200 4589 15204
rect 10952 15260 11016 15264
rect 10952 15204 10956 15260
rect 10956 15204 11012 15260
rect 11012 15204 11016 15260
rect 10952 15200 11016 15204
rect 11032 15260 11096 15264
rect 11032 15204 11036 15260
rect 11036 15204 11092 15260
rect 11092 15204 11096 15260
rect 11032 15200 11096 15204
rect 11112 15260 11176 15264
rect 11112 15204 11116 15260
rect 11116 15204 11172 15260
rect 11172 15204 11176 15260
rect 11112 15200 11176 15204
rect 11192 15260 11256 15264
rect 11192 15204 11196 15260
rect 11196 15204 11252 15260
rect 11252 15204 11256 15260
rect 11192 15200 11256 15204
rect 17618 15260 17682 15264
rect 17618 15204 17622 15260
rect 17622 15204 17678 15260
rect 17678 15204 17682 15260
rect 17618 15200 17682 15204
rect 17698 15260 17762 15264
rect 17698 15204 17702 15260
rect 17702 15204 17758 15260
rect 17758 15204 17762 15260
rect 17698 15200 17762 15204
rect 17778 15260 17842 15264
rect 17778 15204 17782 15260
rect 17782 15204 17838 15260
rect 17838 15204 17842 15260
rect 17778 15200 17842 15204
rect 17858 15260 17922 15264
rect 17858 15204 17862 15260
rect 17862 15204 17918 15260
rect 17918 15204 17922 15260
rect 17858 15200 17922 15204
rect 7618 14716 7682 14720
rect 7618 14660 7622 14716
rect 7622 14660 7678 14716
rect 7678 14660 7682 14716
rect 7618 14656 7682 14660
rect 7698 14716 7762 14720
rect 7698 14660 7702 14716
rect 7702 14660 7758 14716
rect 7758 14660 7762 14716
rect 7698 14656 7762 14660
rect 7778 14716 7842 14720
rect 7778 14660 7782 14716
rect 7782 14660 7838 14716
rect 7838 14660 7842 14716
rect 7778 14656 7842 14660
rect 7858 14716 7922 14720
rect 7858 14660 7862 14716
rect 7862 14660 7918 14716
rect 7918 14660 7922 14716
rect 7858 14656 7922 14660
rect 14285 14716 14349 14720
rect 14285 14660 14289 14716
rect 14289 14660 14345 14716
rect 14345 14660 14349 14716
rect 14285 14656 14349 14660
rect 14365 14716 14429 14720
rect 14365 14660 14369 14716
rect 14369 14660 14425 14716
rect 14425 14660 14429 14716
rect 14365 14656 14429 14660
rect 14445 14716 14509 14720
rect 14445 14660 14449 14716
rect 14449 14660 14505 14716
rect 14505 14660 14509 14716
rect 14445 14656 14509 14660
rect 14525 14716 14589 14720
rect 14525 14660 14529 14716
rect 14529 14660 14585 14716
rect 14585 14660 14589 14716
rect 14525 14656 14589 14660
rect 4285 14172 4349 14176
rect 4285 14116 4289 14172
rect 4289 14116 4345 14172
rect 4345 14116 4349 14172
rect 4285 14112 4349 14116
rect 4365 14172 4429 14176
rect 4365 14116 4369 14172
rect 4369 14116 4425 14172
rect 4425 14116 4429 14172
rect 4365 14112 4429 14116
rect 4445 14172 4509 14176
rect 4445 14116 4449 14172
rect 4449 14116 4505 14172
rect 4505 14116 4509 14172
rect 4445 14112 4509 14116
rect 4525 14172 4589 14176
rect 4525 14116 4529 14172
rect 4529 14116 4585 14172
rect 4585 14116 4589 14172
rect 4525 14112 4589 14116
rect 10952 14172 11016 14176
rect 10952 14116 10956 14172
rect 10956 14116 11012 14172
rect 11012 14116 11016 14172
rect 10952 14112 11016 14116
rect 11032 14172 11096 14176
rect 11032 14116 11036 14172
rect 11036 14116 11092 14172
rect 11092 14116 11096 14172
rect 11032 14112 11096 14116
rect 11112 14172 11176 14176
rect 11112 14116 11116 14172
rect 11116 14116 11172 14172
rect 11172 14116 11176 14172
rect 11112 14112 11176 14116
rect 11192 14172 11256 14176
rect 11192 14116 11196 14172
rect 11196 14116 11252 14172
rect 11252 14116 11256 14172
rect 11192 14112 11256 14116
rect 17618 14172 17682 14176
rect 17618 14116 17622 14172
rect 17622 14116 17678 14172
rect 17678 14116 17682 14172
rect 17618 14112 17682 14116
rect 17698 14172 17762 14176
rect 17698 14116 17702 14172
rect 17702 14116 17758 14172
rect 17758 14116 17762 14172
rect 17698 14112 17762 14116
rect 17778 14172 17842 14176
rect 17778 14116 17782 14172
rect 17782 14116 17838 14172
rect 17838 14116 17842 14172
rect 17778 14112 17842 14116
rect 17858 14172 17922 14176
rect 17858 14116 17862 14172
rect 17862 14116 17918 14172
rect 17918 14116 17922 14172
rect 17858 14112 17922 14116
rect 7618 13628 7682 13632
rect 7618 13572 7622 13628
rect 7622 13572 7678 13628
rect 7678 13572 7682 13628
rect 7618 13568 7682 13572
rect 7698 13628 7762 13632
rect 7698 13572 7702 13628
rect 7702 13572 7758 13628
rect 7758 13572 7762 13628
rect 7698 13568 7762 13572
rect 7778 13628 7842 13632
rect 7778 13572 7782 13628
rect 7782 13572 7838 13628
rect 7838 13572 7842 13628
rect 7778 13568 7842 13572
rect 7858 13628 7922 13632
rect 7858 13572 7862 13628
rect 7862 13572 7918 13628
rect 7918 13572 7922 13628
rect 7858 13568 7922 13572
rect 14285 13628 14349 13632
rect 14285 13572 14289 13628
rect 14289 13572 14345 13628
rect 14345 13572 14349 13628
rect 14285 13568 14349 13572
rect 14365 13628 14429 13632
rect 14365 13572 14369 13628
rect 14369 13572 14425 13628
rect 14425 13572 14429 13628
rect 14365 13568 14429 13572
rect 14445 13628 14509 13632
rect 14445 13572 14449 13628
rect 14449 13572 14505 13628
rect 14505 13572 14509 13628
rect 14445 13568 14509 13572
rect 14525 13628 14589 13632
rect 14525 13572 14529 13628
rect 14529 13572 14585 13628
rect 14585 13572 14589 13628
rect 14525 13568 14589 13572
rect 4285 13084 4349 13088
rect 4285 13028 4289 13084
rect 4289 13028 4345 13084
rect 4345 13028 4349 13084
rect 4285 13024 4349 13028
rect 4365 13084 4429 13088
rect 4365 13028 4369 13084
rect 4369 13028 4425 13084
rect 4425 13028 4429 13084
rect 4365 13024 4429 13028
rect 4445 13084 4509 13088
rect 4445 13028 4449 13084
rect 4449 13028 4505 13084
rect 4505 13028 4509 13084
rect 4445 13024 4509 13028
rect 4525 13084 4589 13088
rect 4525 13028 4529 13084
rect 4529 13028 4585 13084
rect 4585 13028 4589 13084
rect 4525 13024 4589 13028
rect 10952 13084 11016 13088
rect 10952 13028 10956 13084
rect 10956 13028 11012 13084
rect 11012 13028 11016 13084
rect 10952 13024 11016 13028
rect 11032 13084 11096 13088
rect 11032 13028 11036 13084
rect 11036 13028 11092 13084
rect 11092 13028 11096 13084
rect 11032 13024 11096 13028
rect 11112 13084 11176 13088
rect 11112 13028 11116 13084
rect 11116 13028 11172 13084
rect 11172 13028 11176 13084
rect 11112 13024 11176 13028
rect 11192 13084 11256 13088
rect 11192 13028 11196 13084
rect 11196 13028 11252 13084
rect 11252 13028 11256 13084
rect 11192 13024 11256 13028
rect 17618 13084 17682 13088
rect 17618 13028 17622 13084
rect 17622 13028 17678 13084
rect 17678 13028 17682 13084
rect 17618 13024 17682 13028
rect 17698 13084 17762 13088
rect 17698 13028 17702 13084
rect 17702 13028 17758 13084
rect 17758 13028 17762 13084
rect 17698 13024 17762 13028
rect 17778 13084 17842 13088
rect 17778 13028 17782 13084
rect 17782 13028 17838 13084
rect 17838 13028 17842 13084
rect 17778 13024 17842 13028
rect 17858 13084 17922 13088
rect 17858 13028 17862 13084
rect 17862 13028 17918 13084
rect 17918 13028 17922 13084
rect 17858 13024 17922 13028
rect 7618 12540 7682 12544
rect 7618 12484 7622 12540
rect 7622 12484 7678 12540
rect 7678 12484 7682 12540
rect 7618 12480 7682 12484
rect 7698 12540 7762 12544
rect 7698 12484 7702 12540
rect 7702 12484 7758 12540
rect 7758 12484 7762 12540
rect 7698 12480 7762 12484
rect 7778 12540 7842 12544
rect 7778 12484 7782 12540
rect 7782 12484 7838 12540
rect 7838 12484 7842 12540
rect 7778 12480 7842 12484
rect 7858 12540 7922 12544
rect 7858 12484 7862 12540
rect 7862 12484 7918 12540
rect 7918 12484 7922 12540
rect 7858 12480 7922 12484
rect 14285 12540 14349 12544
rect 14285 12484 14289 12540
rect 14289 12484 14345 12540
rect 14345 12484 14349 12540
rect 14285 12480 14349 12484
rect 14365 12540 14429 12544
rect 14365 12484 14369 12540
rect 14369 12484 14425 12540
rect 14425 12484 14429 12540
rect 14365 12480 14429 12484
rect 14445 12540 14509 12544
rect 14445 12484 14449 12540
rect 14449 12484 14505 12540
rect 14505 12484 14509 12540
rect 14445 12480 14509 12484
rect 14525 12540 14589 12544
rect 14525 12484 14529 12540
rect 14529 12484 14585 12540
rect 14585 12484 14589 12540
rect 14525 12480 14589 12484
rect 4285 11996 4349 12000
rect 4285 11940 4289 11996
rect 4289 11940 4345 11996
rect 4345 11940 4349 11996
rect 4285 11936 4349 11940
rect 4365 11996 4429 12000
rect 4365 11940 4369 11996
rect 4369 11940 4425 11996
rect 4425 11940 4429 11996
rect 4365 11936 4429 11940
rect 4445 11996 4509 12000
rect 4445 11940 4449 11996
rect 4449 11940 4505 11996
rect 4505 11940 4509 11996
rect 4445 11936 4509 11940
rect 4525 11996 4589 12000
rect 4525 11940 4529 11996
rect 4529 11940 4585 11996
rect 4585 11940 4589 11996
rect 4525 11936 4589 11940
rect 10952 11996 11016 12000
rect 10952 11940 10956 11996
rect 10956 11940 11012 11996
rect 11012 11940 11016 11996
rect 10952 11936 11016 11940
rect 11032 11996 11096 12000
rect 11032 11940 11036 11996
rect 11036 11940 11092 11996
rect 11092 11940 11096 11996
rect 11032 11936 11096 11940
rect 11112 11996 11176 12000
rect 11112 11940 11116 11996
rect 11116 11940 11172 11996
rect 11172 11940 11176 11996
rect 11112 11936 11176 11940
rect 11192 11996 11256 12000
rect 11192 11940 11196 11996
rect 11196 11940 11252 11996
rect 11252 11940 11256 11996
rect 11192 11936 11256 11940
rect 17618 11996 17682 12000
rect 17618 11940 17622 11996
rect 17622 11940 17678 11996
rect 17678 11940 17682 11996
rect 17618 11936 17682 11940
rect 17698 11996 17762 12000
rect 17698 11940 17702 11996
rect 17702 11940 17758 11996
rect 17758 11940 17762 11996
rect 17698 11936 17762 11940
rect 17778 11996 17842 12000
rect 17778 11940 17782 11996
rect 17782 11940 17838 11996
rect 17838 11940 17842 11996
rect 17778 11936 17842 11940
rect 17858 11996 17922 12000
rect 17858 11940 17862 11996
rect 17862 11940 17918 11996
rect 17918 11940 17922 11996
rect 17858 11936 17922 11940
rect 7618 11452 7682 11456
rect 7618 11396 7622 11452
rect 7622 11396 7678 11452
rect 7678 11396 7682 11452
rect 7618 11392 7682 11396
rect 7698 11452 7762 11456
rect 7698 11396 7702 11452
rect 7702 11396 7758 11452
rect 7758 11396 7762 11452
rect 7698 11392 7762 11396
rect 7778 11452 7842 11456
rect 7778 11396 7782 11452
rect 7782 11396 7838 11452
rect 7838 11396 7842 11452
rect 7778 11392 7842 11396
rect 7858 11452 7922 11456
rect 7858 11396 7862 11452
rect 7862 11396 7918 11452
rect 7918 11396 7922 11452
rect 7858 11392 7922 11396
rect 14285 11452 14349 11456
rect 14285 11396 14289 11452
rect 14289 11396 14345 11452
rect 14345 11396 14349 11452
rect 14285 11392 14349 11396
rect 14365 11452 14429 11456
rect 14365 11396 14369 11452
rect 14369 11396 14425 11452
rect 14425 11396 14429 11452
rect 14365 11392 14429 11396
rect 14445 11452 14509 11456
rect 14445 11396 14449 11452
rect 14449 11396 14505 11452
rect 14505 11396 14509 11452
rect 14445 11392 14509 11396
rect 14525 11452 14589 11456
rect 14525 11396 14529 11452
rect 14529 11396 14585 11452
rect 14585 11396 14589 11452
rect 14525 11392 14589 11396
rect 4285 10908 4349 10912
rect 4285 10852 4289 10908
rect 4289 10852 4345 10908
rect 4345 10852 4349 10908
rect 4285 10848 4349 10852
rect 4365 10908 4429 10912
rect 4365 10852 4369 10908
rect 4369 10852 4425 10908
rect 4425 10852 4429 10908
rect 4365 10848 4429 10852
rect 4445 10908 4509 10912
rect 4445 10852 4449 10908
rect 4449 10852 4505 10908
rect 4505 10852 4509 10908
rect 4445 10848 4509 10852
rect 4525 10908 4589 10912
rect 4525 10852 4529 10908
rect 4529 10852 4585 10908
rect 4585 10852 4589 10908
rect 4525 10848 4589 10852
rect 10952 10908 11016 10912
rect 10952 10852 10956 10908
rect 10956 10852 11012 10908
rect 11012 10852 11016 10908
rect 10952 10848 11016 10852
rect 11032 10908 11096 10912
rect 11032 10852 11036 10908
rect 11036 10852 11092 10908
rect 11092 10852 11096 10908
rect 11032 10848 11096 10852
rect 11112 10908 11176 10912
rect 11112 10852 11116 10908
rect 11116 10852 11172 10908
rect 11172 10852 11176 10908
rect 11112 10848 11176 10852
rect 11192 10908 11256 10912
rect 11192 10852 11196 10908
rect 11196 10852 11252 10908
rect 11252 10852 11256 10908
rect 11192 10848 11256 10852
rect 17618 10908 17682 10912
rect 17618 10852 17622 10908
rect 17622 10852 17678 10908
rect 17678 10852 17682 10908
rect 17618 10848 17682 10852
rect 17698 10908 17762 10912
rect 17698 10852 17702 10908
rect 17702 10852 17758 10908
rect 17758 10852 17762 10908
rect 17698 10848 17762 10852
rect 17778 10908 17842 10912
rect 17778 10852 17782 10908
rect 17782 10852 17838 10908
rect 17838 10852 17842 10908
rect 17778 10848 17842 10852
rect 17858 10908 17922 10912
rect 17858 10852 17862 10908
rect 17862 10852 17918 10908
rect 17918 10852 17922 10908
rect 17858 10848 17922 10852
rect 7618 10364 7682 10368
rect 7618 10308 7622 10364
rect 7622 10308 7678 10364
rect 7678 10308 7682 10364
rect 7618 10304 7682 10308
rect 7698 10364 7762 10368
rect 7698 10308 7702 10364
rect 7702 10308 7758 10364
rect 7758 10308 7762 10364
rect 7698 10304 7762 10308
rect 7778 10364 7842 10368
rect 7778 10308 7782 10364
rect 7782 10308 7838 10364
rect 7838 10308 7842 10364
rect 7778 10304 7842 10308
rect 7858 10364 7922 10368
rect 7858 10308 7862 10364
rect 7862 10308 7918 10364
rect 7918 10308 7922 10364
rect 7858 10304 7922 10308
rect 14285 10364 14349 10368
rect 14285 10308 14289 10364
rect 14289 10308 14345 10364
rect 14345 10308 14349 10364
rect 14285 10304 14349 10308
rect 14365 10364 14429 10368
rect 14365 10308 14369 10364
rect 14369 10308 14425 10364
rect 14425 10308 14429 10364
rect 14365 10304 14429 10308
rect 14445 10364 14509 10368
rect 14445 10308 14449 10364
rect 14449 10308 14505 10364
rect 14505 10308 14509 10364
rect 14445 10304 14509 10308
rect 14525 10364 14589 10368
rect 14525 10308 14529 10364
rect 14529 10308 14585 10364
rect 14585 10308 14589 10364
rect 14525 10304 14589 10308
rect 4285 9820 4349 9824
rect 4285 9764 4289 9820
rect 4289 9764 4345 9820
rect 4345 9764 4349 9820
rect 4285 9760 4349 9764
rect 4365 9820 4429 9824
rect 4365 9764 4369 9820
rect 4369 9764 4425 9820
rect 4425 9764 4429 9820
rect 4365 9760 4429 9764
rect 4445 9820 4509 9824
rect 4445 9764 4449 9820
rect 4449 9764 4505 9820
rect 4505 9764 4509 9820
rect 4445 9760 4509 9764
rect 4525 9820 4589 9824
rect 4525 9764 4529 9820
rect 4529 9764 4585 9820
rect 4585 9764 4589 9820
rect 4525 9760 4589 9764
rect 10952 9820 11016 9824
rect 10952 9764 10956 9820
rect 10956 9764 11012 9820
rect 11012 9764 11016 9820
rect 10952 9760 11016 9764
rect 11032 9820 11096 9824
rect 11032 9764 11036 9820
rect 11036 9764 11092 9820
rect 11092 9764 11096 9820
rect 11032 9760 11096 9764
rect 11112 9820 11176 9824
rect 11112 9764 11116 9820
rect 11116 9764 11172 9820
rect 11172 9764 11176 9820
rect 11112 9760 11176 9764
rect 11192 9820 11256 9824
rect 11192 9764 11196 9820
rect 11196 9764 11252 9820
rect 11252 9764 11256 9820
rect 11192 9760 11256 9764
rect 17618 9820 17682 9824
rect 17618 9764 17622 9820
rect 17622 9764 17678 9820
rect 17678 9764 17682 9820
rect 17618 9760 17682 9764
rect 17698 9820 17762 9824
rect 17698 9764 17702 9820
rect 17702 9764 17758 9820
rect 17758 9764 17762 9820
rect 17698 9760 17762 9764
rect 17778 9820 17842 9824
rect 17778 9764 17782 9820
rect 17782 9764 17838 9820
rect 17838 9764 17842 9820
rect 17778 9760 17842 9764
rect 17858 9820 17922 9824
rect 17858 9764 17862 9820
rect 17862 9764 17918 9820
rect 17918 9764 17922 9820
rect 17858 9760 17922 9764
rect 7618 9276 7682 9280
rect 7618 9220 7622 9276
rect 7622 9220 7678 9276
rect 7678 9220 7682 9276
rect 7618 9216 7682 9220
rect 7698 9276 7762 9280
rect 7698 9220 7702 9276
rect 7702 9220 7758 9276
rect 7758 9220 7762 9276
rect 7698 9216 7762 9220
rect 7778 9276 7842 9280
rect 7778 9220 7782 9276
rect 7782 9220 7838 9276
rect 7838 9220 7842 9276
rect 7778 9216 7842 9220
rect 7858 9276 7922 9280
rect 7858 9220 7862 9276
rect 7862 9220 7918 9276
rect 7918 9220 7922 9276
rect 7858 9216 7922 9220
rect 14285 9276 14349 9280
rect 14285 9220 14289 9276
rect 14289 9220 14345 9276
rect 14345 9220 14349 9276
rect 14285 9216 14349 9220
rect 14365 9276 14429 9280
rect 14365 9220 14369 9276
rect 14369 9220 14425 9276
rect 14425 9220 14429 9276
rect 14365 9216 14429 9220
rect 14445 9276 14509 9280
rect 14445 9220 14449 9276
rect 14449 9220 14505 9276
rect 14505 9220 14509 9276
rect 14445 9216 14509 9220
rect 14525 9276 14589 9280
rect 14525 9220 14529 9276
rect 14529 9220 14585 9276
rect 14585 9220 14589 9276
rect 14525 9216 14589 9220
rect 4285 8732 4349 8736
rect 4285 8676 4289 8732
rect 4289 8676 4345 8732
rect 4345 8676 4349 8732
rect 4285 8672 4349 8676
rect 4365 8732 4429 8736
rect 4365 8676 4369 8732
rect 4369 8676 4425 8732
rect 4425 8676 4429 8732
rect 4365 8672 4429 8676
rect 4445 8732 4509 8736
rect 4445 8676 4449 8732
rect 4449 8676 4505 8732
rect 4505 8676 4509 8732
rect 4445 8672 4509 8676
rect 4525 8732 4589 8736
rect 4525 8676 4529 8732
rect 4529 8676 4585 8732
rect 4585 8676 4589 8732
rect 4525 8672 4589 8676
rect 10952 8732 11016 8736
rect 10952 8676 10956 8732
rect 10956 8676 11012 8732
rect 11012 8676 11016 8732
rect 10952 8672 11016 8676
rect 11032 8732 11096 8736
rect 11032 8676 11036 8732
rect 11036 8676 11092 8732
rect 11092 8676 11096 8732
rect 11032 8672 11096 8676
rect 11112 8732 11176 8736
rect 11112 8676 11116 8732
rect 11116 8676 11172 8732
rect 11172 8676 11176 8732
rect 11112 8672 11176 8676
rect 11192 8732 11256 8736
rect 11192 8676 11196 8732
rect 11196 8676 11252 8732
rect 11252 8676 11256 8732
rect 11192 8672 11256 8676
rect 17618 8732 17682 8736
rect 17618 8676 17622 8732
rect 17622 8676 17678 8732
rect 17678 8676 17682 8732
rect 17618 8672 17682 8676
rect 17698 8732 17762 8736
rect 17698 8676 17702 8732
rect 17702 8676 17758 8732
rect 17758 8676 17762 8732
rect 17698 8672 17762 8676
rect 17778 8732 17842 8736
rect 17778 8676 17782 8732
rect 17782 8676 17838 8732
rect 17838 8676 17842 8732
rect 17778 8672 17842 8676
rect 17858 8732 17922 8736
rect 17858 8676 17862 8732
rect 17862 8676 17918 8732
rect 17918 8676 17922 8732
rect 17858 8672 17922 8676
rect 7618 8188 7682 8192
rect 7618 8132 7622 8188
rect 7622 8132 7678 8188
rect 7678 8132 7682 8188
rect 7618 8128 7682 8132
rect 7698 8188 7762 8192
rect 7698 8132 7702 8188
rect 7702 8132 7758 8188
rect 7758 8132 7762 8188
rect 7698 8128 7762 8132
rect 7778 8188 7842 8192
rect 7778 8132 7782 8188
rect 7782 8132 7838 8188
rect 7838 8132 7842 8188
rect 7778 8128 7842 8132
rect 7858 8188 7922 8192
rect 7858 8132 7862 8188
rect 7862 8132 7918 8188
rect 7918 8132 7922 8188
rect 7858 8128 7922 8132
rect 14285 8188 14349 8192
rect 14285 8132 14289 8188
rect 14289 8132 14345 8188
rect 14345 8132 14349 8188
rect 14285 8128 14349 8132
rect 14365 8188 14429 8192
rect 14365 8132 14369 8188
rect 14369 8132 14425 8188
rect 14425 8132 14429 8188
rect 14365 8128 14429 8132
rect 14445 8188 14509 8192
rect 14445 8132 14449 8188
rect 14449 8132 14505 8188
rect 14505 8132 14509 8188
rect 14445 8128 14509 8132
rect 14525 8188 14589 8192
rect 14525 8132 14529 8188
rect 14529 8132 14585 8188
rect 14585 8132 14589 8188
rect 14525 8128 14589 8132
rect 4285 7644 4349 7648
rect 4285 7588 4289 7644
rect 4289 7588 4345 7644
rect 4345 7588 4349 7644
rect 4285 7584 4349 7588
rect 4365 7644 4429 7648
rect 4365 7588 4369 7644
rect 4369 7588 4425 7644
rect 4425 7588 4429 7644
rect 4365 7584 4429 7588
rect 4445 7644 4509 7648
rect 4445 7588 4449 7644
rect 4449 7588 4505 7644
rect 4505 7588 4509 7644
rect 4445 7584 4509 7588
rect 4525 7644 4589 7648
rect 4525 7588 4529 7644
rect 4529 7588 4585 7644
rect 4585 7588 4589 7644
rect 4525 7584 4589 7588
rect 10952 7644 11016 7648
rect 10952 7588 10956 7644
rect 10956 7588 11012 7644
rect 11012 7588 11016 7644
rect 10952 7584 11016 7588
rect 11032 7644 11096 7648
rect 11032 7588 11036 7644
rect 11036 7588 11092 7644
rect 11092 7588 11096 7644
rect 11032 7584 11096 7588
rect 11112 7644 11176 7648
rect 11112 7588 11116 7644
rect 11116 7588 11172 7644
rect 11172 7588 11176 7644
rect 11112 7584 11176 7588
rect 11192 7644 11256 7648
rect 11192 7588 11196 7644
rect 11196 7588 11252 7644
rect 11252 7588 11256 7644
rect 11192 7584 11256 7588
rect 17618 7644 17682 7648
rect 17618 7588 17622 7644
rect 17622 7588 17678 7644
rect 17678 7588 17682 7644
rect 17618 7584 17682 7588
rect 17698 7644 17762 7648
rect 17698 7588 17702 7644
rect 17702 7588 17758 7644
rect 17758 7588 17762 7644
rect 17698 7584 17762 7588
rect 17778 7644 17842 7648
rect 17778 7588 17782 7644
rect 17782 7588 17838 7644
rect 17838 7588 17842 7644
rect 17778 7584 17842 7588
rect 17858 7644 17922 7648
rect 17858 7588 17862 7644
rect 17862 7588 17918 7644
rect 17918 7588 17922 7644
rect 17858 7584 17922 7588
rect 7618 7100 7682 7104
rect 7618 7044 7622 7100
rect 7622 7044 7678 7100
rect 7678 7044 7682 7100
rect 7618 7040 7682 7044
rect 7698 7100 7762 7104
rect 7698 7044 7702 7100
rect 7702 7044 7758 7100
rect 7758 7044 7762 7100
rect 7698 7040 7762 7044
rect 7778 7100 7842 7104
rect 7778 7044 7782 7100
rect 7782 7044 7838 7100
rect 7838 7044 7842 7100
rect 7778 7040 7842 7044
rect 7858 7100 7922 7104
rect 7858 7044 7862 7100
rect 7862 7044 7918 7100
rect 7918 7044 7922 7100
rect 7858 7040 7922 7044
rect 14285 7100 14349 7104
rect 14285 7044 14289 7100
rect 14289 7044 14345 7100
rect 14345 7044 14349 7100
rect 14285 7040 14349 7044
rect 14365 7100 14429 7104
rect 14365 7044 14369 7100
rect 14369 7044 14425 7100
rect 14425 7044 14429 7100
rect 14365 7040 14429 7044
rect 14445 7100 14509 7104
rect 14445 7044 14449 7100
rect 14449 7044 14505 7100
rect 14505 7044 14509 7100
rect 14445 7040 14509 7044
rect 14525 7100 14589 7104
rect 14525 7044 14529 7100
rect 14529 7044 14585 7100
rect 14585 7044 14589 7100
rect 14525 7040 14589 7044
rect 4285 6556 4349 6560
rect 4285 6500 4289 6556
rect 4289 6500 4345 6556
rect 4345 6500 4349 6556
rect 4285 6496 4349 6500
rect 4365 6556 4429 6560
rect 4365 6500 4369 6556
rect 4369 6500 4425 6556
rect 4425 6500 4429 6556
rect 4365 6496 4429 6500
rect 4445 6556 4509 6560
rect 4445 6500 4449 6556
rect 4449 6500 4505 6556
rect 4505 6500 4509 6556
rect 4445 6496 4509 6500
rect 4525 6556 4589 6560
rect 4525 6500 4529 6556
rect 4529 6500 4585 6556
rect 4585 6500 4589 6556
rect 4525 6496 4589 6500
rect 10952 6556 11016 6560
rect 10952 6500 10956 6556
rect 10956 6500 11012 6556
rect 11012 6500 11016 6556
rect 10952 6496 11016 6500
rect 11032 6556 11096 6560
rect 11032 6500 11036 6556
rect 11036 6500 11092 6556
rect 11092 6500 11096 6556
rect 11032 6496 11096 6500
rect 11112 6556 11176 6560
rect 11112 6500 11116 6556
rect 11116 6500 11172 6556
rect 11172 6500 11176 6556
rect 11112 6496 11176 6500
rect 11192 6556 11256 6560
rect 11192 6500 11196 6556
rect 11196 6500 11252 6556
rect 11252 6500 11256 6556
rect 11192 6496 11256 6500
rect 17618 6556 17682 6560
rect 17618 6500 17622 6556
rect 17622 6500 17678 6556
rect 17678 6500 17682 6556
rect 17618 6496 17682 6500
rect 17698 6556 17762 6560
rect 17698 6500 17702 6556
rect 17702 6500 17758 6556
rect 17758 6500 17762 6556
rect 17698 6496 17762 6500
rect 17778 6556 17842 6560
rect 17778 6500 17782 6556
rect 17782 6500 17838 6556
rect 17838 6500 17842 6556
rect 17778 6496 17842 6500
rect 17858 6556 17922 6560
rect 17858 6500 17862 6556
rect 17862 6500 17918 6556
rect 17918 6500 17922 6556
rect 17858 6496 17922 6500
rect 7618 6012 7682 6016
rect 7618 5956 7622 6012
rect 7622 5956 7678 6012
rect 7678 5956 7682 6012
rect 7618 5952 7682 5956
rect 7698 6012 7762 6016
rect 7698 5956 7702 6012
rect 7702 5956 7758 6012
rect 7758 5956 7762 6012
rect 7698 5952 7762 5956
rect 7778 6012 7842 6016
rect 7778 5956 7782 6012
rect 7782 5956 7838 6012
rect 7838 5956 7842 6012
rect 7778 5952 7842 5956
rect 7858 6012 7922 6016
rect 7858 5956 7862 6012
rect 7862 5956 7918 6012
rect 7918 5956 7922 6012
rect 7858 5952 7922 5956
rect 14285 6012 14349 6016
rect 14285 5956 14289 6012
rect 14289 5956 14345 6012
rect 14345 5956 14349 6012
rect 14285 5952 14349 5956
rect 14365 6012 14429 6016
rect 14365 5956 14369 6012
rect 14369 5956 14425 6012
rect 14425 5956 14429 6012
rect 14365 5952 14429 5956
rect 14445 6012 14509 6016
rect 14445 5956 14449 6012
rect 14449 5956 14505 6012
rect 14505 5956 14509 6012
rect 14445 5952 14509 5956
rect 14525 6012 14589 6016
rect 14525 5956 14529 6012
rect 14529 5956 14585 6012
rect 14585 5956 14589 6012
rect 14525 5952 14589 5956
rect 4285 5468 4349 5472
rect 4285 5412 4289 5468
rect 4289 5412 4345 5468
rect 4345 5412 4349 5468
rect 4285 5408 4349 5412
rect 4365 5468 4429 5472
rect 4365 5412 4369 5468
rect 4369 5412 4425 5468
rect 4425 5412 4429 5468
rect 4365 5408 4429 5412
rect 4445 5468 4509 5472
rect 4445 5412 4449 5468
rect 4449 5412 4505 5468
rect 4505 5412 4509 5468
rect 4445 5408 4509 5412
rect 4525 5468 4589 5472
rect 4525 5412 4529 5468
rect 4529 5412 4585 5468
rect 4585 5412 4589 5468
rect 4525 5408 4589 5412
rect 10952 5468 11016 5472
rect 10952 5412 10956 5468
rect 10956 5412 11012 5468
rect 11012 5412 11016 5468
rect 10952 5408 11016 5412
rect 11032 5468 11096 5472
rect 11032 5412 11036 5468
rect 11036 5412 11092 5468
rect 11092 5412 11096 5468
rect 11032 5408 11096 5412
rect 11112 5468 11176 5472
rect 11112 5412 11116 5468
rect 11116 5412 11172 5468
rect 11172 5412 11176 5468
rect 11112 5408 11176 5412
rect 11192 5468 11256 5472
rect 11192 5412 11196 5468
rect 11196 5412 11252 5468
rect 11252 5412 11256 5468
rect 11192 5408 11256 5412
rect 17618 5468 17682 5472
rect 17618 5412 17622 5468
rect 17622 5412 17678 5468
rect 17678 5412 17682 5468
rect 17618 5408 17682 5412
rect 17698 5468 17762 5472
rect 17698 5412 17702 5468
rect 17702 5412 17758 5468
rect 17758 5412 17762 5468
rect 17698 5408 17762 5412
rect 17778 5468 17842 5472
rect 17778 5412 17782 5468
rect 17782 5412 17838 5468
rect 17838 5412 17842 5468
rect 17778 5408 17842 5412
rect 17858 5468 17922 5472
rect 17858 5412 17862 5468
rect 17862 5412 17918 5468
rect 17918 5412 17922 5468
rect 17858 5408 17922 5412
rect 7618 4924 7682 4928
rect 7618 4868 7622 4924
rect 7622 4868 7678 4924
rect 7678 4868 7682 4924
rect 7618 4864 7682 4868
rect 7698 4924 7762 4928
rect 7698 4868 7702 4924
rect 7702 4868 7758 4924
rect 7758 4868 7762 4924
rect 7698 4864 7762 4868
rect 7778 4924 7842 4928
rect 7778 4868 7782 4924
rect 7782 4868 7838 4924
rect 7838 4868 7842 4924
rect 7778 4864 7842 4868
rect 7858 4924 7922 4928
rect 7858 4868 7862 4924
rect 7862 4868 7918 4924
rect 7918 4868 7922 4924
rect 7858 4864 7922 4868
rect 14285 4924 14349 4928
rect 14285 4868 14289 4924
rect 14289 4868 14345 4924
rect 14345 4868 14349 4924
rect 14285 4864 14349 4868
rect 14365 4924 14429 4928
rect 14365 4868 14369 4924
rect 14369 4868 14425 4924
rect 14425 4868 14429 4924
rect 14365 4864 14429 4868
rect 14445 4924 14509 4928
rect 14445 4868 14449 4924
rect 14449 4868 14505 4924
rect 14505 4868 14509 4924
rect 14445 4864 14509 4868
rect 14525 4924 14589 4928
rect 14525 4868 14529 4924
rect 14529 4868 14585 4924
rect 14585 4868 14589 4924
rect 14525 4864 14589 4868
rect 4285 4380 4349 4384
rect 4285 4324 4289 4380
rect 4289 4324 4345 4380
rect 4345 4324 4349 4380
rect 4285 4320 4349 4324
rect 4365 4380 4429 4384
rect 4365 4324 4369 4380
rect 4369 4324 4425 4380
rect 4425 4324 4429 4380
rect 4365 4320 4429 4324
rect 4445 4380 4509 4384
rect 4445 4324 4449 4380
rect 4449 4324 4505 4380
rect 4505 4324 4509 4380
rect 4445 4320 4509 4324
rect 4525 4380 4589 4384
rect 4525 4324 4529 4380
rect 4529 4324 4585 4380
rect 4585 4324 4589 4380
rect 4525 4320 4589 4324
rect 10952 4380 11016 4384
rect 10952 4324 10956 4380
rect 10956 4324 11012 4380
rect 11012 4324 11016 4380
rect 10952 4320 11016 4324
rect 11032 4380 11096 4384
rect 11032 4324 11036 4380
rect 11036 4324 11092 4380
rect 11092 4324 11096 4380
rect 11032 4320 11096 4324
rect 11112 4380 11176 4384
rect 11112 4324 11116 4380
rect 11116 4324 11172 4380
rect 11172 4324 11176 4380
rect 11112 4320 11176 4324
rect 11192 4380 11256 4384
rect 11192 4324 11196 4380
rect 11196 4324 11252 4380
rect 11252 4324 11256 4380
rect 11192 4320 11256 4324
rect 17618 4380 17682 4384
rect 17618 4324 17622 4380
rect 17622 4324 17678 4380
rect 17678 4324 17682 4380
rect 17618 4320 17682 4324
rect 17698 4380 17762 4384
rect 17698 4324 17702 4380
rect 17702 4324 17758 4380
rect 17758 4324 17762 4380
rect 17698 4320 17762 4324
rect 17778 4380 17842 4384
rect 17778 4324 17782 4380
rect 17782 4324 17838 4380
rect 17838 4324 17842 4380
rect 17778 4320 17842 4324
rect 17858 4380 17922 4384
rect 17858 4324 17862 4380
rect 17862 4324 17918 4380
rect 17918 4324 17922 4380
rect 17858 4320 17922 4324
rect 7618 3836 7682 3840
rect 7618 3780 7622 3836
rect 7622 3780 7678 3836
rect 7678 3780 7682 3836
rect 7618 3776 7682 3780
rect 7698 3836 7762 3840
rect 7698 3780 7702 3836
rect 7702 3780 7758 3836
rect 7758 3780 7762 3836
rect 7698 3776 7762 3780
rect 7778 3836 7842 3840
rect 7778 3780 7782 3836
rect 7782 3780 7838 3836
rect 7838 3780 7842 3836
rect 7778 3776 7842 3780
rect 7858 3836 7922 3840
rect 7858 3780 7862 3836
rect 7862 3780 7918 3836
rect 7918 3780 7922 3836
rect 7858 3776 7922 3780
rect 14285 3836 14349 3840
rect 14285 3780 14289 3836
rect 14289 3780 14345 3836
rect 14345 3780 14349 3836
rect 14285 3776 14349 3780
rect 14365 3836 14429 3840
rect 14365 3780 14369 3836
rect 14369 3780 14425 3836
rect 14425 3780 14429 3836
rect 14365 3776 14429 3780
rect 14445 3836 14509 3840
rect 14445 3780 14449 3836
rect 14449 3780 14505 3836
rect 14505 3780 14509 3836
rect 14445 3776 14509 3780
rect 14525 3836 14589 3840
rect 14525 3780 14529 3836
rect 14529 3780 14585 3836
rect 14585 3780 14589 3836
rect 14525 3776 14589 3780
rect 4285 3292 4349 3296
rect 4285 3236 4289 3292
rect 4289 3236 4345 3292
rect 4345 3236 4349 3292
rect 4285 3232 4349 3236
rect 4365 3292 4429 3296
rect 4365 3236 4369 3292
rect 4369 3236 4425 3292
rect 4425 3236 4429 3292
rect 4365 3232 4429 3236
rect 4445 3292 4509 3296
rect 4445 3236 4449 3292
rect 4449 3236 4505 3292
rect 4505 3236 4509 3292
rect 4445 3232 4509 3236
rect 4525 3292 4589 3296
rect 4525 3236 4529 3292
rect 4529 3236 4585 3292
rect 4585 3236 4589 3292
rect 4525 3232 4589 3236
rect 10952 3292 11016 3296
rect 10952 3236 10956 3292
rect 10956 3236 11012 3292
rect 11012 3236 11016 3292
rect 10952 3232 11016 3236
rect 11032 3292 11096 3296
rect 11032 3236 11036 3292
rect 11036 3236 11092 3292
rect 11092 3236 11096 3292
rect 11032 3232 11096 3236
rect 11112 3292 11176 3296
rect 11112 3236 11116 3292
rect 11116 3236 11172 3292
rect 11172 3236 11176 3292
rect 11112 3232 11176 3236
rect 11192 3292 11256 3296
rect 11192 3236 11196 3292
rect 11196 3236 11252 3292
rect 11252 3236 11256 3292
rect 11192 3232 11256 3236
rect 17618 3292 17682 3296
rect 17618 3236 17622 3292
rect 17622 3236 17678 3292
rect 17678 3236 17682 3292
rect 17618 3232 17682 3236
rect 17698 3292 17762 3296
rect 17698 3236 17702 3292
rect 17702 3236 17758 3292
rect 17758 3236 17762 3292
rect 17698 3232 17762 3236
rect 17778 3292 17842 3296
rect 17778 3236 17782 3292
rect 17782 3236 17838 3292
rect 17838 3236 17842 3292
rect 17778 3232 17842 3236
rect 17858 3292 17922 3296
rect 17858 3236 17862 3292
rect 17862 3236 17918 3292
rect 17918 3236 17922 3292
rect 17858 3232 17922 3236
rect 7618 2748 7682 2752
rect 7618 2692 7622 2748
rect 7622 2692 7678 2748
rect 7678 2692 7682 2748
rect 7618 2688 7682 2692
rect 7698 2748 7762 2752
rect 7698 2692 7702 2748
rect 7702 2692 7758 2748
rect 7758 2692 7762 2748
rect 7698 2688 7762 2692
rect 7778 2748 7842 2752
rect 7778 2692 7782 2748
rect 7782 2692 7838 2748
rect 7838 2692 7842 2748
rect 7778 2688 7842 2692
rect 7858 2748 7922 2752
rect 7858 2692 7862 2748
rect 7862 2692 7918 2748
rect 7918 2692 7922 2748
rect 7858 2688 7922 2692
rect 14285 2748 14349 2752
rect 14285 2692 14289 2748
rect 14289 2692 14345 2748
rect 14345 2692 14349 2748
rect 14285 2688 14349 2692
rect 14365 2748 14429 2752
rect 14365 2692 14369 2748
rect 14369 2692 14425 2748
rect 14425 2692 14429 2748
rect 14365 2688 14429 2692
rect 14445 2748 14509 2752
rect 14445 2692 14449 2748
rect 14449 2692 14505 2748
rect 14505 2692 14509 2748
rect 14445 2688 14509 2692
rect 14525 2748 14589 2752
rect 14525 2692 14529 2748
rect 14529 2692 14585 2748
rect 14585 2692 14589 2748
rect 14525 2688 14589 2692
rect 4285 2204 4349 2208
rect 4285 2148 4289 2204
rect 4289 2148 4345 2204
rect 4345 2148 4349 2204
rect 4285 2144 4349 2148
rect 4365 2204 4429 2208
rect 4365 2148 4369 2204
rect 4369 2148 4425 2204
rect 4425 2148 4429 2204
rect 4365 2144 4429 2148
rect 4445 2204 4509 2208
rect 4445 2148 4449 2204
rect 4449 2148 4505 2204
rect 4505 2148 4509 2204
rect 4445 2144 4509 2148
rect 4525 2204 4589 2208
rect 4525 2148 4529 2204
rect 4529 2148 4585 2204
rect 4585 2148 4589 2204
rect 4525 2144 4589 2148
rect 10952 2204 11016 2208
rect 10952 2148 10956 2204
rect 10956 2148 11012 2204
rect 11012 2148 11016 2204
rect 10952 2144 11016 2148
rect 11032 2204 11096 2208
rect 11032 2148 11036 2204
rect 11036 2148 11092 2204
rect 11092 2148 11096 2204
rect 11032 2144 11096 2148
rect 11112 2204 11176 2208
rect 11112 2148 11116 2204
rect 11116 2148 11172 2204
rect 11172 2148 11176 2204
rect 11112 2144 11176 2148
rect 11192 2204 11256 2208
rect 11192 2148 11196 2204
rect 11196 2148 11252 2204
rect 11252 2148 11256 2204
rect 11192 2144 11256 2148
rect 17618 2204 17682 2208
rect 17618 2148 17622 2204
rect 17622 2148 17678 2204
rect 17678 2148 17682 2204
rect 17618 2144 17682 2148
rect 17698 2204 17762 2208
rect 17698 2148 17702 2204
rect 17702 2148 17758 2204
rect 17758 2148 17762 2204
rect 17698 2144 17762 2148
rect 17778 2204 17842 2208
rect 17778 2148 17782 2204
rect 17782 2148 17838 2204
rect 17838 2148 17842 2204
rect 17778 2144 17842 2148
rect 17858 2204 17922 2208
rect 17858 2148 17862 2204
rect 17862 2148 17918 2204
rect 17918 2148 17922 2204
rect 17858 2144 17922 2148
<< metal4 >>
rect 5395 79660 5461 79661
rect 5395 79596 5396 79660
rect 5460 79596 5461 79660
rect 5395 79595 5461 79596
rect 4277 77280 4597 77840
rect 4277 77216 4285 77280
rect 4349 77216 4365 77280
rect 4429 77216 4445 77280
rect 4509 77216 4525 77280
rect 4589 77216 4597 77280
rect 4277 76192 4597 77216
rect 5211 76396 5277 76397
rect 5211 76332 5212 76396
rect 5276 76332 5277 76396
rect 5211 76331 5277 76332
rect 4277 76128 4285 76192
rect 4349 76128 4365 76192
rect 4429 76128 4445 76192
rect 4509 76128 4525 76192
rect 4589 76128 4597 76192
rect 4277 75104 4597 76128
rect 4843 75988 4909 75989
rect 4843 75924 4844 75988
rect 4908 75924 4909 75988
rect 4843 75923 4909 75924
rect 4277 75040 4285 75104
rect 4349 75040 4365 75104
rect 4429 75040 4445 75104
rect 4509 75040 4525 75104
rect 4589 75040 4597 75104
rect 2451 74764 2517 74765
rect 2451 74700 2452 74764
rect 2516 74700 2517 74764
rect 2451 74699 2517 74700
rect 1715 50692 1781 50693
rect 1715 50628 1716 50692
rect 1780 50628 1781 50692
rect 1715 50627 1781 50628
rect 1718 17237 1778 50627
rect 2267 50012 2333 50013
rect 2267 49948 2268 50012
rect 2332 49948 2333 50012
rect 2267 49947 2333 49948
rect 2270 45933 2330 49947
rect 2267 45932 2333 45933
rect 2267 45868 2268 45932
rect 2332 45868 2333 45932
rect 2267 45867 2333 45868
rect 2454 42805 2514 74699
rect 4277 74016 4597 75040
rect 4277 73952 4285 74016
rect 4349 73952 4365 74016
rect 4429 73952 4445 74016
rect 4509 73952 4525 74016
rect 4589 73952 4597 74016
rect 4277 72928 4597 73952
rect 4277 72864 4285 72928
rect 4349 72864 4365 72928
rect 4429 72864 4445 72928
rect 4509 72864 4525 72928
rect 4589 72864 4597 72928
rect 4277 71840 4597 72864
rect 4277 71776 4285 71840
rect 4349 71776 4365 71840
rect 4429 71776 4445 71840
rect 4509 71776 4525 71840
rect 4589 71776 4597 71840
rect 4107 71500 4173 71501
rect 4107 71436 4108 71500
rect 4172 71436 4173 71500
rect 4107 71435 4173 71436
rect 2635 68780 2701 68781
rect 2635 68716 2636 68780
rect 2700 68716 2701 68780
rect 2635 68715 2701 68716
rect 2451 42804 2517 42805
rect 2451 42740 2452 42804
rect 2516 42740 2517 42804
rect 2451 42739 2517 42740
rect 2638 33149 2698 68715
rect 3371 62932 3437 62933
rect 3371 62868 3372 62932
rect 3436 62868 3437 62932
rect 3371 62867 3437 62868
rect 3374 60621 3434 62867
rect 3371 60620 3437 60621
rect 3371 60556 3372 60620
rect 3436 60556 3437 60620
rect 3371 60555 3437 60556
rect 3371 59396 3437 59397
rect 3371 59332 3372 59396
rect 3436 59332 3437 59396
rect 3371 59331 3437 59332
rect 3187 55996 3253 55997
rect 3187 55932 3188 55996
rect 3252 55932 3253 55996
rect 3187 55931 3253 55932
rect 3003 55044 3069 55045
rect 3003 54980 3004 55044
rect 3068 54980 3069 55044
rect 3003 54979 3069 54980
rect 3006 51373 3066 54979
rect 3003 51372 3069 51373
rect 3003 51308 3004 51372
rect 3068 51308 3069 51372
rect 3003 51307 3069 51308
rect 3190 46749 3250 55931
rect 3374 51509 3434 59331
rect 3555 58716 3621 58717
rect 3555 58652 3556 58716
rect 3620 58652 3621 58716
rect 3555 58651 3621 58652
rect 3558 51645 3618 58651
rect 3739 55724 3805 55725
rect 3739 55660 3740 55724
rect 3804 55660 3805 55724
rect 3739 55659 3805 55660
rect 3555 51644 3621 51645
rect 3555 51580 3556 51644
rect 3620 51580 3621 51644
rect 3555 51579 3621 51580
rect 3371 51508 3437 51509
rect 3371 51444 3372 51508
rect 3436 51444 3437 51508
rect 3371 51443 3437 51444
rect 3742 48245 3802 55659
rect 3923 55452 3989 55453
rect 3923 55388 3924 55452
rect 3988 55388 3989 55452
rect 3923 55387 3989 55388
rect 3926 51373 3986 55387
rect 3923 51372 3989 51373
rect 3923 51308 3924 51372
rect 3988 51308 3989 51372
rect 3923 51307 3989 51308
rect 3739 48244 3805 48245
rect 3739 48180 3740 48244
rect 3804 48180 3805 48244
rect 3739 48179 3805 48180
rect 3923 47564 3989 47565
rect 3923 47500 3924 47564
rect 3988 47500 3989 47564
rect 3923 47499 3989 47500
rect 3187 46748 3253 46749
rect 3187 46684 3188 46748
rect 3252 46684 3253 46748
rect 3187 46683 3253 46684
rect 3926 44437 3986 47499
rect 3923 44436 3989 44437
rect 3923 44372 3924 44436
rect 3988 44372 3989 44436
rect 3923 44371 3989 44372
rect 3926 40221 3986 44371
rect 3923 40220 3989 40221
rect 3923 40156 3924 40220
rect 3988 40156 3989 40220
rect 3923 40155 3989 40156
rect 4110 39949 4170 71435
rect 4277 70752 4597 71776
rect 4277 70688 4285 70752
rect 4349 70688 4365 70752
rect 4429 70688 4445 70752
rect 4509 70688 4525 70752
rect 4589 70688 4597 70752
rect 4277 69664 4597 70688
rect 4659 70548 4725 70549
rect 4659 70484 4660 70548
rect 4724 70484 4725 70548
rect 4659 70483 4725 70484
rect 4277 69600 4285 69664
rect 4349 69600 4365 69664
rect 4429 69600 4445 69664
rect 4509 69600 4525 69664
rect 4589 69600 4597 69664
rect 4277 68912 4597 69600
rect 4277 68676 4319 68912
rect 4555 68676 4597 68912
rect 4277 68576 4597 68676
rect 4277 68512 4285 68576
rect 4349 68512 4365 68576
rect 4429 68512 4445 68576
rect 4509 68512 4525 68576
rect 4589 68512 4597 68576
rect 4277 67488 4597 68512
rect 4277 67424 4285 67488
rect 4349 67424 4365 67488
rect 4429 67424 4445 67488
rect 4509 67424 4525 67488
rect 4589 67424 4597 67488
rect 4277 66400 4597 67424
rect 4277 66336 4285 66400
rect 4349 66336 4365 66400
rect 4429 66336 4445 66400
rect 4509 66336 4525 66400
rect 4589 66336 4597 66400
rect 4277 65312 4597 66336
rect 4277 65248 4285 65312
rect 4349 65248 4365 65312
rect 4429 65248 4445 65312
rect 4509 65248 4525 65312
rect 4589 65248 4597 65312
rect 4277 64224 4597 65248
rect 4277 64160 4285 64224
rect 4349 64160 4365 64224
rect 4429 64160 4445 64224
rect 4509 64160 4525 64224
rect 4589 64160 4597 64224
rect 4277 63136 4597 64160
rect 4277 63072 4285 63136
rect 4349 63072 4365 63136
rect 4429 63072 4445 63136
rect 4509 63072 4525 63136
rect 4589 63072 4597 63136
rect 4277 62048 4597 63072
rect 4277 61984 4285 62048
rect 4349 61984 4365 62048
rect 4429 61984 4445 62048
rect 4509 61984 4525 62048
rect 4589 61984 4597 62048
rect 4277 60960 4597 61984
rect 4277 60896 4285 60960
rect 4349 60896 4365 60960
rect 4429 60896 4445 60960
rect 4509 60896 4525 60960
rect 4589 60896 4597 60960
rect 4277 59872 4597 60896
rect 4277 59808 4285 59872
rect 4349 59808 4365 59872
rect 4429 59808 4445 59872
rect 4509 59808 4525 59872
rect 4589 59808 4597 59872
rect 4277 58784 4597 59808
rect 4277 58720 4285 58784
rect 4349 58720 4365 58784
rect 4429 58720 4445 58784
rect 4509 58720 4525 58784
rect 4589 58720 4597 58784
rect 4277 57696 4597 58720
rect 4277 57632 4285 57696
rect 4349 57632 4365 57696
rect 4429 57632 4445 57696
rect 4509 57632 4525 57696
rect 4589 57632 4597 57696
rect 4277 56608 4597 57632
rect 4277 56544 4285 56608
rect 4349 56544 4365 56608
rect 4429 56544 4445 56608
rect 4509 56544 4525 56608
rect 4589 56544 4597 56608
rect 4277 55520 4597 56544
rect 4277 55456 4285 55520
rect 4349 55456 4365 55520
rect 4429 55456 4445 55520
rect 4509 55456 4525 55520
rect 4589 55456 4597 55520
rect 4277 54432 4597 55456
rect 4277 54368 4285 54432
rect 4349 54368 4365 54432
rect 4429 54368 4445 54432
rect 4509 54368 4525 54432
rect 4589 54368 4597 54432
rect 4277 53344 4597 54368
rect 4277 53280 4285 53344
rect 4349 53280 4365 53344
rect 4429 53280 4445 53344
rect 4509 53280 4525 53344
rect 4589 53280 4597 53344
rect 4277 52256 4597 53280
rect 4277 52192 4285 52256
rect 4349 52192 4365 52256
rect 4429 52192 4445 52256
rect 4509 52192 4525 52256
rect 4589 52192 4597 52256
rect 4277 51168 4597 52192
rect 4277 51104 4285 51168
rect 4349 51104 4365 51168
rect 4429 51104 4445 51168
rect 4509 51104 4525 51168
rect 4589 51104 4597 51168
rect 4277 50080 4597 51104
rect 4277 50016 4285 50080
rect 4349 50016 4365 50080
rect 4429 50016 4445 50080
rect 4509 50016 4525 50080
rect 4589 50016 4597 50080
rect 4277 48992 4597 50016
rect 4277 48928 4285 48992
rect 4349 48928 4365 48992
rect 4429 48928 4445 48992
rect 4509 48928 4525 48992
rect 4589 48928 4597 48992
rect 4277 47904 4597 48928
rect 4277 47840 4285 47904
rect 4349 47840 4365 47904
rect 4429 47840 4445 47904
rect 4509 47840 4525 47904
rect 4589 47840 4597 47904
rect 4277 46816 4597 47840
rect 4277 46752 4285 46816
rect 4349 46752 4365 46816
rect 4429 46752 4445 46816
rect 4509 46752 4525 46816
rect 4589 46752 4597 46816
rect 4277 45728 4597 46752
rect 4277 45664 4285 45728
rect 4349 45664 4365 45728
rect 4429 45664 4445 45728
rect 4509 45664 4525 45728
rect 4589 45664 4597 45728
rect 4277 44640 4597 45664
rect 4662 45117 4722 70483
rect 4846 45933 4906 75923
rect 5027 75444 5093 75445
rect 5027 75380 5028 75444
rect 5092 75380 5093 75444
rect 5027 75379 5093 75380
rect 5030 46069 5090 75379
rect 5214 55725 5274 76331
rect 5211 55724 5277 55725
rect 5211 55660 5212 55724
rect 5276 55660 5277 55724
rect 5211 55659 5277 55660
rect 5398 52050 5458 79595
rect 7610 77824 7930 77840
rect 7610 77760 7618 77824
rect 7682 77760 7698 77824
rect 7762 77760 7778 77824
rect 7842 77760 7858 77824
rect 7922 77760 7930 77824
rect 7610 76736 7930 77760
rect 7610 76672 7618 76736
rect 7682 76672 7698 76736
rect 7762 76672 7778 76736
rect 7842 76672 7858 76736
rect 7922 76672 7930 76736
rect 7610 75648 7930 76672
rect 7610 75584 7618 75648
rect 7682 75584 7698 75648
rect 7762 75584 7778 75648
rect 7842 75584 7858 75648
rect 7922 75584 7930 75648
rect 7610 74560 7930 75584
rect 7610 74496 7618 74560
rect 7682 74496 7698 74560
rect 7762 74496 7778 74560
rect 7842 74496 7858 74560
rect 7922 74496 7930 74560
rect 7235 73812 7301 73813
rect 7235 73748 7236 73812
rect 7300 73748 7301 73812
rect 7235 73747 7301 73748
rect 6867 69732 6933 69733
rect 6867 69668 6868 69732
rect 6932 69668 6933 69732
rect 6867 69667 6933 69668
rect 5579 56132 5645 56133
rect 5579 56068 5580 56132
rect 5644 56068 5645 56132
rect 5579 56067 5645 56068
rect 5582 52189 5642 56067
rect 5947 55724 6013 55725
rect 5947 55660 5948 55724
rect 6012 55660 6013 55724
rect 5947 55659 6013 55660
rect 5763 54092 5829 54093
rect 5763 54028 5764 54092
rect 5828 54028 5829 54092
rect 5763 54027 5829 54028
rect 5579 52188 5645 52189
rect 5579 52124 5580 52188
rect 5644 52124 5645 52188
rect 5579 52123 5645 52124
rect 5398 51990 5642 52050
rect 5211 51236 5277 51237
rect 5211 51172 5212 51236
rect 5276 51172 5277 51236
rect 5211 51171 5277 51172
rect 5027 46068 5093 46069
rect 5027 46004 5028 46068
rect 5092 46004 5093 46068
rect 5027 46003 5093 46004
rect 4843 45932 4909 45933
rect 4843 45868 4844 45932
rect 4908 45868 4909 45932
rect 4843 45867 4909 45868
rect 4659 45116 4725 45117
rect 4659 45052 4660 45116
rect 4724 45052 4725 45116
rect 4659 45051 4725 45052
rect 4277 44576 4285 44640
rect 4349 44576 4365 44640
rect 4429 44576 4445 44640
rect 4509 44576 4525 44640
rect 4589 44576 4597 44640
rect 4277 43552 4597 44576
rect 4277 43488 4285 43552
rect 4349 43488 4365 43552
rect 4429 43488 4445 43552
rect 4509 43488 4525 43552
rect 4589 43488 4597 43552
rect 4277 42464 4597 43488
rect 5214 43210 5274 51171
rect 5582 50690 5642 51990
rect 5766 50965 5826 54027
rect 5950 53141 6010 55659
rect 6131 55044 6197 55045
rect 6131 54980 6132 55044
rect 6196 54980 6197 55044
rect 6131 54979 6197 54980
rect 5947 53140 6013 53141
rect 5947 53076 5948 53140
rect 6012 53076 6013 53140
rect 5947 53075 6013 53076
rect 5950 51509 6010 53075
rect 5947 51508 6013 51509
rect 5947 51444 5948 51508
rect 6012 51444 6013 51508
rect 5947 51443 6013 51444
rect 5947 51236 6013 51237
rect 5947 51172 5948 51236
rect 6012 51172 6013 51236
rect 5947 51171 6013 51172
rect 5763 50964 5829 50965
rect 5763 50900 5764 50964
rect 5828 50900 5829 50964
rect 5763 50899 5829 50900
rect 5950 50829 6010 51171
rect 5947 50828 6013 50829
rect 5947 50764 5948 50828
rect 6012 50764 6013 50828
rect 5947 50763 6013 50764
rect 5398 50630 5642 50690
rect 5398 49197 5458 50630
rect 6134 50421 6194 54979
rect 6683 54364 6749 54365
rect 6683 54300 6684 54364
rect 6748 54300 6749 54364
rect 6683 54299 6749 54300
rect 6499 53956 6565 53957
rect 6499 53892 6500 53956
rect 6564 53892 6565 53956
rect 6499 53891 6565 53892
rect 6315 53004 6381 53005
rect 6315 52940 6316 53004
rect 6380 52940 6381 53004
rect 6315 52939 6381 52940
rect 6131 50420 6197 50421
rect 6131 50356 6132 50420
rect 6196 50356 6197 50420
rect 6131 50355 6197 50356
rect 6131 50148 6197 50149
rect 6131 50084 6132 50148
rect 6196 50084 6197 50148
rect 6131 50083 6197 50084
rect 5395 49196 5461 49197
rect 5395 49132 5396 49196
rect 5460 49132 5461 49196
rect 5395 49131 5461 49132
rect 5395 48924 5461 48925
rect 5395 48860 5396 48924
rect 5460 48860 5461 48924
rect 5395 48859 5461 48860
rect 5398 43893 5458 48859
rect 5763 48380 5829 48381
rect 5763 48316 5764 48380
rect 5828 48316 5829 48380
rect 5763 48315 5829 48316
rect 5395 43892 5461 43893
rect 5395 43828 5396 43892
rect 5460 43828 5461 43892
rect 5395 43827 5461 43828
rect 5214 43150 5458 43210
rect 4277 42400 4285 42464
rect 4349 42400 4365 42464
rect 4429 42400 4445 42464
rect 4509 42400 4525 42464
rect 4589 42400 4597 42464
rect 4277 42246 4597 42400
rect 4277 42010 4319 42246
rect 4555 42010 4597 42246
rect 4277 41376 4597 42010
rect 4277 41312 4285 41376
rect 4349 41312 4365 41376
rect 4429 41312 4445 41376
rect 4509 41312 4525 41376
rect 4589 41312 4597 41376
rect 4277 40288 4597 41312
rect 4277 40224 4285 40288
rect 4349 40224 4365 40288
rect 4429 40224 4445 40288
rect 4509 40224 4525 40288
rect 4589 40224 4597 40288
rect 4107 39948 4173 39949
rect 4107 39884 4108 39948
rect 4172 39884 4173 39948
rect 4107 39883 4173 39884
rect 4277 39200 4597 40224
rect 4277 39136 4285 39200
rect 4349 39136 4365 39200
rect 4429 39136 4445 39200
rect 4509 39136 4525 39200
rect 4589 39136 4597 39200
rect 4277 38112 4597 39136
rect 4277 38048 4285 38112
rect 4349 38048 4365 38112
rect 4429 38048 4445 38112
rect 4509 38048 4525 38112
rect 4589 38048 4597 38112
rect 4277 37024 4597 38048
rect 4277 36960 4285 37024
rect 4349 36960 4365 37024
rect 4429 36960 4445 37024
rect 4509 36960 4525 37024
rect 4589 36960 4597 37024
rect 4277 35936 4597 36960
rect 4277 35872 4285 35936
rect 4349 35872 4365 35936
rect 4429 35872 4445 35936
rect 4509 35872 4525 35936
rect 4589 35872 4597 35936
rect 4277 34848 4597 35872
rect 4277 34784 4285 34848
rect 4349 34784 4365 34848
rect 4429 34784 4445 34848
rect 4509 34784 4525 34848
rect 4589 34784 4597 34848
rect 4277 33760 4597 34784
rect 4277 33696 4285 33760
rect 4349 33696 4365 33760
rect 4429 33696 4445 33760
rect 4509 33696 4525 33760
rect 4589 33696 4597 33760
rect 2635 33148 2701 33149
rect 2635 33084 2636 33148
rect 2700 33084 2701 33148
rect 2635 33083 2701 33084
rect 4277 32672 4597 33696
rect 4277 32608 4285 32672
rect 4349 32608 4365 32672
rect 4429 32608 4445 32672
rect 4509 32608 4525 32672
rect 4589 32608 4597 32672
rect 4277 31584 4597 32608
rect 4277 31520 4285 31584
rect 4349 31520 4365 31584
rect 4429 31520 4445 31584
rect 4509 31520 4525 31584
rect 4589 31520 4597 31584
rect 4277 30496 4597 31520
rect 4277 30432 4285 30496
rect 4349 30432 4365 30496
rect 4429 30432 4445 30496
rect 4509 30432 4525 30496
rect 4589 30432 4597 30496
rect 4277 29408 4597 30432
rect 4277 29344 4285 29408
rect 4349 29344 4365 29408
rect 4429 29344 4445 29408
rect 4509 29344 4525 29408
rect 4589 29344 4597 29408
rect 4277 28320 4597 29344
rect 4277 28256 4285 28320
rect 4349 28256 4365 28320
rect 4429 28256 4445 28320
rect 4509 28256 4525 28320
rect 4589 28256 4597 28320
rect 4277 27232 4597 28256
rect 4277 27168 4285 27232
rect 4349 27168 4365 27232
rect 4429 27168 4445 27232
rect 4509 27168 4525 27232
rect 4589 27168 4597 27232
rect 4277 26144 4597 27168
rect 5398 26621 5458 43150
rect 5579 41988 5645 41989
rect 5579 41924 5580 41988
rect 5644 41924 5645 41988
rect 5579 41923 5645 41924
rect 5582 40901 5642 41923
rect 5766 41445 5826 48315
rect 6134 45525 6194 50083
rect 6318 47701 6378 52939
rect 6315 47700 6381 47701
rect 6315 47636 6316 47700
rect 6380 47636 6381 47700
rect 6315 47635 6381 47636
rect 6502 47021 6562 53891
rect 6686 51645 6746 54299
rect 6683 51644 6749 51645
rect 6683 51580 6684 51644
rect 6748 51580 6749 51644
rect 6683 51579 6749 51580
rect 6683 51372 6749 51373
rect 6683 51308 6684 51372
rect 6748 51308 6749 51372
rect 6683 51307 6749 51308
rect 6686 50690 6746 51307
rect 6870 50829 6930 69667
rect 7051 63612 7117 63613
rect 7051 63548 7052 63612
rect 7116 63548 7117 63612
rect 7051 63547 7117 63548
rect 7054 51373 7114 63547
rect 7238 63069 7298 73747
rect 7610 73472 7930 74496
rect 7610 73408 7618 73472
rect 7682 73408 7698 73472
rect 7762 73408 7778 73472
rect 7842 73408 7858 73472
rect 7922 73408 7930 73472
rect 7610 72384 7930 73408
rect 10944 77280 11264 77840
rect 10944 77216 10952 77280
rect 11016 77216 11032 77280
rect 11096 77216 11112 77280
rect 11176 77216 11192 77280
rect 11256 77216 11264 77280
rect 10944 76192 11264 77216
rect 10944 76128 10952 76192
rect 11016 76128 11032 76192
rect 11096 76128 11112 76192
rect 11176 76128 11192 76192
rect 11256 76128 11264 76192
rect 10944 75104 11264 76128
rect 10944 75040 10952 75104
rect 11016 75040 11032 75104
rect 11096 75040 11112 75104
rect 11176 75040 11192 75104
rect 11256 75040 11264 75104
rect 10944 74016 11264 75040
rect 10944 73952 10952 74016
rect 11016 73952 11032 74016
rect 11096 73952 11112 74016
rect 11176 73952 11192 74016
rect 11256 73952 11264 74016
rect 10731 73268 10797 73269
rect 10731 73204 10732 73268
rect 10796 73204 10797 73268
rect 10731 73203 10797 73204
rect 7610 72320 7618 72384
rect 7682 72320 7698 72384
rect 7762 72320 7778 72384
rect 7842 72320 7858 72384
rect 7922 72320 7930 72384
rect 7610 71296 7930 72320
rect 7610 71232 7618 71296
rect 7682 71232 7698 71296
rect 7762 71232 7778 71296
rect 7842 71232 7858 71296
rect 7922 71232 7930 71296
rect 7610 70208 7930 71232
rect 9627 70684 9693 70685
rect 9627 70620 9628 70684
rect 9692 70620 9693 70684
rect 9627 70619 9693 70620
rect 8155 70412 8221 70413
rect 8155 70348 8156 70412
rect 8220 70348 8221 70412
rect 8155 70347 8221 70348
rect 7610 70144 7618 70208
rect 7682 70144 7698 70208
rect 7762 70144 7778 70208
rect 7842 70144 7858 70208
rect 7922 70144 7930 70208
rect 7610 69120 7930 70144
rect 7610 69056 7618 69120
rect 7682 69056 7698 69120
rect 7762 69056 7778 69120
rect 7842 69056 7858 69120
rect 7922 69056 7930 69120
rect 7610 68032 7930 69056
rect 7610 67968 7618 68032
rect 7682 67968 7698 68032
rect 7762 67968 7778 68032
rect 7842 67968 7858 68032
rect 7922 67968 7930 68032
rect 7610 66944 7930 67968
rect 7610 66880 7618 66944
rect 7682 66880 7698 66944
rect 7762 66880 7778 66944
rect 7842 66880 7858 66944
rect 7922 66880 7930 66944
rect 7610 65856 7930 66880
rect 7610 65792 7618 65856
rect 7682 65792 7698 65856
rect 7762 65792 7778 65856
rect 7842 65792 7858 65856
rect 7922 65792 7930 65856
rect 7610 64768 7930 65792
rect 7610 64704 7618 64768
rect 7682 64704 7698 64768
rect 7762 64704 7778 64768
rect 7842 64704 7858 64768
rect 7922 64704 7930 64768
rect 7419 64564 7485 64565
rect 7419 64500 7420 64564
rect 7484 64500 7485 64564
rect 7419 64499 7485 64500
rect 7235 63068 7301 63069
rect 7235 63004 7236 63068
rect 7300 63004 7301 63068
rect 7235 63003 7301 63004
rect 7235 58988 7301 58989
rect 7235 58924 7236 58988
rect 7300 58924 7301 58988
rect 7235 58923 7301 58924
rect 7238 54093 7298 58923
rect 7235 54092 7301 54093
rect 7235 54028 7236 54092
rect 7300 54028 7301 54092
rect 7235 54027 7301 54028
rect 7235 53956 7301 53957
rect 7235 53892 7236 53956
rect 7300 53892 7301 53956
rect 7235 53891 7301 53892
rect 7051 51372 7117 51373
rect 7051 51308 7052 51372
rect 7116 51308 7117 51372
rect 7051 51307 7117 51308
rect 7051 51236 7117 51237
rect 7051 51172 7052 51236
rect 7116 51172 7117 51236
rect 7051 51171 7117 51172
rect 6867 50828 6933 50829
rect 6867 50764 6868 50828
rect 6932 50764 6933 50828
rect 6867 50763 6933 50764
rect 6686 50630 6930 50690
rect 6683 50556 6749 50557
rect 6683 50492 6684 50556
rect 6748 50492 6749 50556
rect 6683 50491 6749 50492
rect 6686 49330 6746 50491
rect 6870 49877 6930 50630
rect 6867 49876 6933 49877
rect 6867 49812 6868 49876
rect 6932 49812 6933 49876
rect 6867 49811 6933 49812
rect 6870 49605 6930 49811
rect 6867 49604 6933 49605
rect 6867 49540 6868 49604
rect 6932 49540 6933 49604
rect 6867 49539 6933 49540
rect 6686 49270 6930 49330
rect 6870 48378 6930 49270
rect 6870 48318 6976 48378
rect 6916 47970 6976 48318
rect 6870 47910 6976 47970
rect 6683 47836 6749 47837
rect 6683 47772 6684 47836
rect 6748 47772 6749 47836
rect 6683 47771 6749 47772
rect 6499 47020 6565 47021
rect 6499 46956 6500 47020
rect 6564 46956 6565 47020
rect 6499 46955 6565 46956
rect 6131 45524 6197 45525
rect 6131 45460 6132 45524
rect 6196 45460 6197 45524
rect 6131 45459 6197 45460
rect 6134 42805 6194 45459
rect 6315 43076 6381 43077
rect 6315 43012 6316 43076
rect 6380 43012 6381 43076
rect 6315 43011 6381 43012
rect 6131 42804 6197 42805
rect 6131 42740 6132 42804
rect 6196 42740 6197 42804
rect 6131 42739 6197 42740
rect 5763 41444 5829 41445
rect 5763 41380 5764 41444
rect 5828 41380 5829 41444
rect 5763 41379 5829 41380
rect 5763 41172 5829 41173
rect 5763 41108 5764 41172
rect 5828 41108 5829 41172
rect 5763 41107 5829 41108
rect 5579 40900 5645 40901
rect 5579 40836 5580 40900
rect 5644 40836 5645 40900
rect 5579 40835 5645 40836
rect 5766 36413 5826 41107
rect 6318 39813 6378 43011
rect 6686 42125 6746 47771
rect 6870 42941 6930 47910
rect 7054 46477 7114 51171
rect 7051 46476 7117 46477
rect 7051 46412 7052 46476
rect 7116 46412 7117 46476
rect 7051 46411 7117 46412
rect 7051 45660 7117 45661
rect 7051 45596 7052 45660
rect 7116 45596 7117 45660
rect 7051 45595 7117 45596
rect 6867 42940 6933 42941
rect 6867 42876 6868 42940
rect 6932 42876 6933 42940
rect 6867 42875 6933 42876
rect 6683 42124 6749 42125
rect 6683 42060 6684 42124
rect 6748 42060 6749 42124
rect 6683 42059 6749 42060
rect 6683 41444 6749 41445
rect 6683 41380 6684 41444
rect 6748 41380 6749 41444
rect 6683 41379 6749 41380
rect 6686 41309 6746 41379
rect 6683 41308 6749 41309
rect 6683 41244 6684 41308
rect 6748 41244 6749 41308
rect 6683 41243 6749 41244
rect 6315 39812 6381 39813
rect 6315 39748 6316 39812
rect 6380 39748 6381 39812
rect 6315 39747 6381 39748
rect 6867 38180 6933 38181
rect 6867 38116 6868 38180
rect 6932 38116 6933 38180
rect 6867 38115 6933 38116
rect 5763 36412 5829 36413
rect 5763 36348 5764 36412
rect 5828 36348 5829 36412
rect 5763 36347 5829 36348
rect 6870 33693 6930 38115
rect 6867 33692 6933 33693
rect 6867 33628 6868 33692
rect 6932 33628 6933 33692
rect 6867 33627 6933 33628
rect 7054 31789 7114 45595
rect 7238 37093 7298 53891
rect 7422 51237 7482 64499
rect 7610 63680 7930 64704
rect 7610 63616 7618 63680
rect 7682 63616 7698 63680
rect 7762 63616 7778 63680
rect 7842 63616 7858 63680
rect 7922 63616 7930 63680
rect 7610 62592 7930 63616
rect 7610 62528 7618 62592
rect 7682 62528 7698 62592
rect 7762 62528 7778 62592
rect 7842 62528 7858 62592
rect 7922 62528 7930 62592
rect 7610 61504 7930 62528
rect 7610 61440 7618 61504
rect 7682 61440 7698 61504
rect 7762 61440 7778 61504
rect 7842 61440 7858 61504
rect 7922 61440 7930 61504
rect 7610 60416 7930 61440
rect 7610 60352 7618 60416
rect 7682 60352 7698 60416
rect 7762 60352 7778 60416
rect 7842 60352 7858 60416
rect 7922 60352 7930 60416
rect 7610 59328 7930 60352
rect 7610 59264 7618 59328
rect 7682 59264 7698 59328
rect 7762 59264 7778 59328
rect 7842 59264 7858 59328
rect 7922 59264 7930 59328
rect 7610 58240 7930 59264
rect 7610 58176 7618 58240
rect 7682 58176 7698 58240
rect 7762 58176 7778 58240
rect 7842 58176 7858 58240
rect 7922 58176 7930 58240
rect 7610 57152 7930 58176
rect 7610 57088 7618 57152
rect 7682 57088 7698 57152
rect 7762 57088 7778 57152
rect 7842 57088 7858 57152
rect 7922 57088 7930 57152
rect 7610 56064 7930 57088
rect 7610 56000 7618 56064
rect 7682 56000 7698 56064
rect 7762 56000 7778 56064
rect 7842 56000 7858 56064
rect 7922 56000 7930 56064
rect 7610 55579 7930 56000
rect 7610 55343 7652 55579
rect 7888 55343 7930 55579
rect 7610 54976 7930 55343
rect 7610 54912 7618 54976
rect 7682 54912 7698 54976
rect 7762 54912 7778 54976
rect 7842 54912 7858 54976
rect 7922 54912 7930 54976
rect 7610 53888 7930 54912
rect 7610 53824 7618 53888
rect 7682 53824 7698 53888
rect 7762 53824 7778 53888
rect 7842 53824 7858 53888
rect 7922 53824 7930 53888
rect 7610 52800 7930 53824
rect 7610 52736 7618 52800
rect 7682 52736 7698 52800
rect 7762 52736 7778 52800
rect 7842 52736 7858 52800
rect 7922 52736 7930 52800
rect 7610 51712 7930 52736
rect 7610 51648 7618 51712
rect 7682 51648 7698 51712
rect 7762 51648 7778 51712
rect 7842 51648 7858 51712
rect 7922 51648 7930 51712
rect 7419 51236 7485 51237
rect 7419 51172 7420 51236
rect 7484 51172 7485 51236
rect 7419 51171 7485 51172
rect 7419 51100 7485 51101
rect 7419 51036 7420 51100
rect 7484 51036 7485 51100
rect 7419 51035 7485 51036
rect 7235 37092 7301 37093
rect 7235 37028 7236 37092
rect 7300 37028 7301 37092
rect 7235 37027 7301 37028
rect 7422 32605 7482 51035
rect 7610 50624 7930 51648
rect 7610 50560 7618 50624
rect 7682 50560 7698 50624
rect 7762 50560 7778 50624
rect 7842 50560 7858 50624
rect 7922 50560 7930 50624
rect 7610 49536 7930 50560
rect 7610 49472 7618 49536
rect 7682 49472 7698 49536
rect 7762 49472 7778 49536
rect 7842 49472 7858 49536
rect 7922 49472 7930 49536
rect 7610 48448 7930 49472
rect 7610 48384 7618 48448
rect 7682 48384 7698 48448
rect 7762 48384 7778 48448
rect 7842 48384 7858 48448
rect 7922 48384 7930 48448
rect 7610 47360 7930 48384
rect 7610 47296 7618 47360
rect 7682 47296 7698 47360
rect 7762 47296 7778 47360
rect 7842 47296 7858 47360
rect 7922 47296 7930 47360
rect 7610 46272 7930 47296
rect 7610 46208 7618 46272
rect 7682 46208 7698 46272
rect 7762 46208 7778 46272
rect 7842 46208 7858 46272
rect 7922 46208 7930 46272
rect 7610 45184 7930 46208
rect 7610 45120 7618 45184
rect 7682 45120 7698 45184
rect 7762 45120 7778 45184
rect 7842 45120 7858 45184
rect 7922 45120 7930 45184
rect 7610 44096 7930 45120
rect 7610 44032 7618 44096
rect 7682 44032 7698 44096
rect 7762 44032 7778 44096
rect 7842 44032 7858 44096
rect 7922 44032 7930 44096
rect 7610 43008 7930 44032
rect 7610 42944 7618 43008
rect 7682 42944 7698 43008
rect 7762 42944 7778 43008
rect 7842 42944 7858 43008
rect 7922 42944 7930 43008
rect 7610 41920 7930 42944
rect 7610 41856 7618 41920
rect 7682 41856 7698 41920
rect 7762 41856 7778 41920
rect 7842 41856 7858 41920
rect 7922 41856 7930 41920
rect 7610 40832 7930 41856
rect 7610 40768 7618 40832
rect 7682 40768 7698 40832
rect 7762 40768 7778 40832
rect 7842 40768 7858 40832
rect 7922 40768 7930 40832
rect 7610 39744 7930 40768
rect 7610 39680 7618 39744
rect 7682 39680 7698 39744
rect 7762 39680 7778 39744
rect 7842 39680 7858 39744
rect 7922 39680 7930 39744
rect 7610 38656 7930 39680
rect 7610 38592 7618 38656
rect 7682 38592 7698 38656
rect 7762 38592 7778 38656
rect 7842 38592 7858 38656
rect 7922 38592 7930 38656
rect 7610 37568 7930 38592
rect 7610 37504 7618 37568
rect 7682 37504 7698 37568
rect 7762 37504 7778 37568
rect 7842 37504 7858 37568
rect 7922 37504 7930 37568
rect 7610 36480 7930 37504
rect 7610 36416 7618 36480
rect 7682 36416 7698 36480
rect 7762 36416 7778 36480
rect 7842 36416 7858 36480
rect 7922 36416 7930 36480
rect 7610 35392 7930 36416
rect 7610 35328 7618 35392
rect 7682 35328 7698 35392
rect 7762 35328 7778 35392
rect 7842 35328 7858 35392
rect 7922 35328 7930 35392
rect 7610 34304 7930 35328
rect 7610 34240 7618 34304
rect 7682 34240 7698 34304
rect 7762 34240 7778 34304
rect 7842 34240 7858 34304
rect 7922 34240 7930 34304
rect 7610 33216 7930 34240
rect 7610 33152 7618 33216
rect 7682 33152 7698 33216
rect 7762 33152 7778 33216
rect 7842 33152 7858 33216
rect 7922 33152 7930 33216
rect 7419 32604 7485 32605
rect 7419 32540 7420 32604
rect 7484 32540 7485 32604
rect 7419 32539 7485 32540
rect 7610 32128 7930 33152
rect 8158 32877 8218 70347
rect 8339 63068 8405 63069
rect 8339 63004 8340 63068
rect 8404 63004 8405 63068
rect 8339 63003 8405 63004
rect 8342 52050 8402 63003
rect 9259 60076 9325 60077
rect 9259 60012 9260 60076
rect 9324 60012 9325 60076
rect 9259 60011 9325 60012
rect 9075 56404 9141 56405
rect 9075 56340 9076 56404
rect 9140 56340 9141 56404
rect 9075 56339 9141 56340
rect 8891 56268 8957 56269
rect 8891 56204 8892 56268
rect 8956 56204 8957 56268
rect 8891 56203 8957 56204
rect 8523 55860 8589 55861
rect 8523 55796 8524 55860
rect 8588 55796 8589 55860
rect 8523 55795 8589 55796
rect 8526 52733 8586 55795
rect 8707 55452 8773 55453
rect 8707 55388 8708 55452
rect 8772 55388 8773 55452
rect 8707 55387 8773 55388
rect 8523 52732 8589 52733
rect 8523 52668 8524 52732
rect 8588 52668 8589 52732
rect 8523 52667 8589 52668
rect 8342 51990 8586 52050
rect 8339 51372 8405 51373
rect 8339 51308 8340 51372
rect 8404 51308 8405 51372
rect 8339 51307 8405 51308
rect 8342 50149 8402 51307
rect 8339 50148 8405 50149
rect 8339 50084 8340 50148
rect 8404 50084 8405 50148
rect 8339 50083 8405 50084
rect 8342 46885 8402 50083
rect 8339 46884 8405 46885
rect 8339 46820 8340 46884
rect 8404 46820 8405 46884
rect 8339 46819 8405 46820
rect 8526 43349 8586 51990
rect 8710 51237 8770 55387
rect 8894 55181 8954 56203
rect 8891 55180 8957 55181
rect 8891 55116 8892 55180
rect 8956 55116 8957 55180
rect 8891 55115 8957 55116
rect 8707 51236 8773 51237
rect 8707 51172 8708 51236
rect 8772 51172 8773 51236
rect 8707 51171 8773 51172
rect 8894 51098 8954 55115
rect 9078 51101 9138 56339
rect 9262 55045 9322 60011
rect 9443 57356 9509 57357
rect 9443 57292 9444 57356
rect 9508 57292 9509 57356
rect 9443 57291 9509 57292
rect 9259 55044 9325 55045
rect 9259 54980 9260 55044
rect 9324 54980 9325 55044
rect 9259 54979 9325 54980
rect 9446 53685 9506 57291
rect 9443 53684 9509 53685
rect 9443 53620 9444 53684
rect 9508 53620 9509 53684
rect 9443 53619 9509 53620
rect 9259 51236 9325 51237
rect 9259 51172 9260 51236
rect 9324 51172 9325 51236
rect 9259 51171 9325 51172
rect 8710 51038 8954 51098
rect 9075 51100 9141 51101
rect 8710 48381 8770 51038
rect 9075 51036 9076 51100
rect 9140 51036 9141 51100
rect 9075 51035 9141 51036
rect 9075 50692 9141 50693
rect 9075 50628 9076 50692
rect 9140 50628 9141 50692
rect 9075 50627 9141 50628
rect 8891 49196 8957 49197
rect 8891 49132 8892 49196
rect 8956 49132 8957 49196
rect 8891 49131 8957 49132
rect 8707 48380 8773 48381
rect 8707 48316 8708 48380
rect 8772 48316 8773 48380
rect 8707 48315 8773 48316
rect 8707 45796 8773 45797
rect 8707 45732 8708 45796
rect 8772 45732 8773 45796
rect 8707 45731 8773 45732
rect 8523 43348 8589 43349
rect 8523 43284 8524 43348
rect 8588 43284 8589 43348
rect 8523 43283 8589 43284
rect 8339 42804 8405 42805
rect 8339 42740 8340 42804
rect 8404 42740 8405 42804
rect 8339 42739 8405 42740
rect 8342 41309 8402 42739
rect 8710 42261 8770 45731
rect 8894 45661 8954 49131
rect 8891 45660 8957 45661
rect 8891 45596 8892 45660
rect 8956 45596 8957 45660
rect 8891 45595 8957 45596
rect 9078 44301 9138 50627
rect 9262 49877 9322 51171
rect 9446 50965 9506 53619
rect 9443 50964 9509 50965
rect 9443 50900 9444 50964
rect 9508 50900 9509 50964
rect 9443 50899 9509 50900
rect 9443 50692 9509 50693
rect 9443 50628 9444 50692
rect 9508 50628 9509 50692
rect 9443 50627 9509 50628
rect 9259 49876 9325 49877
rect 9259 49812 9260 49876
rect 9324 49812 9325 49876
rect 9259 49811 9325 49812
rect 9259 49468 9325 49469
rect 9259 49404 9260 49468
rect 9324 49404 9325 49468
rect 9259 49403 9325 49404
rect 9262 44437 9322 49403
rect 9259 44436 9325 44437
rect 9259 44372 9260 44436
rect 9324 44372 9325 44436
rect 9259 44371 9325 44372
rect 9075 44300 9141 44301
rect 9075 44236 9076 44300
rect 9140 44236 9141 44300
rect 9075 44235 9141 44236
rect 9078 42941 9138 44235
rect 9075 42940 9141 42941
rect 9075 42876 9076 42940
rect 9140 42876 9141 42940
rect 9075 42875 9141 42876
rect 8707 42260 8773 42261
rect 8707 42196 8708 42260
rect 8772 42196 8773 42260
rect 8707 42195 8773 42196
rect 8339 41308 8405 41309
rect 8339 41244 8340 41308
rect 8404 41244 8405 41308
rect 8339 41243 8405 41244
rect 8339 40628 8405 40629
rect 8339 40564 8340 40628
rect 8404 40564 8405 40628
rect 8339 40563 8405 40564
rect 8155 32876 8221 32877
rect 8155 32812 8156 32876
rect 8220 32812 8221 32876
rect 8155 32811 8221 32812
rect 7610 32064 7618 32128
rect 7682 32064 7698 32128
rect 7762 32064 7778 32128
rect 7842 32064 7858 32128
rect 7922 32064 7930 32128
rect 7051 31788 7117 31789
rect 7051 31724 7052 31788
rect 7116 31724 7117 31788
rect 7051 31723 7117 31724
rect 7610 31040 7930 32064
rect 7610 30976 7618 31040
rect 7682 30976 7698 31040
rect 7762 30976 7778 31040
rect 7842 30976 7858 31040
rect 7922 30976 7930 31040
rect 7610 29952 7930 30976
rect 7610 29888 7618 29952
rect 7682 29888 7698 29952
rect 7762 29888 7778 29952
rect 7842 29888 7858 29952
rect 7922 29888 7930 29952
rect 7610 28912 7930 29888
rect 8342 29205 8402 40563
rect 8710 38453 8770 42195
rect 9262 41445 9322 44371
rect 9446 44165 9506 50627
rect 9630 50013 9690 70619
rect 10363 65924 10429 65925
rect 10363 65860 10364 65924
rect 10428 65860 10429 65924
rect 10363 65859 10429 65860
rect 9811 64020 9877 64021
rect 9811 63956 9812 64020
rect 9876 63956 9877 64020
rect 9811 63955 9877 63956
rect 9814 60757 9874 63955
rect 9995 62252 10061 62253
rect 9995 62188 9996 62252
rect 10060 62188 10061 62252
rect 9995 62187 10061 62188
rect 9811 60756 9877 60757
rect 9811 60692 9812 60756
rect 9876 60692 9877 60756
rect 9811 60691 9877 60692
rect 9811 54908 9877 54909
rect 9811 54844 9812 54908
rect 9876 54844 9877 54908
rect 9811 54843 9877 54844
rect 9627 50012 9693 50013
rect 9627 49948 9628 50012
rect 9692 49948 9693 50012
rect 9627 49947 9693 49948
rect 9627 49876 9693 49877
rect 9627 49812 9628 49876
rect 9692 49812 9693 49876
rect 9627 49811 9693 49812
rect 9443 44164 9509 44165
rect 9443 44100 9444 44164
rect 9508 44100 9509 44164
rect 9443 44099 9509 44100
rect 9259 41444 9325 41445
rect 9259 41380 9260 41444
rect 9324 41380 9325 41444
rect 9259 41379 9325 41380
rect 8707 38452 8773 38453
rect 8707 38388 8708 38452
rect 8772 38388 8773 38452
rect 8707 38387 8773 38388
rect 8339 29204 8405 29205
rect 8339 29140 8340 29204
rect 8404 29140 8405 29204
rect 8339 29139 8405 29140
rect 7610 28864 7652 28912
rect 7888 28864 7930 28912
rect 7610 28800 7618 28864
rect 7922 28800 7930 28864
rect 7610 28676 7652 28800
rect 7888 28676 7930 28800
rect 7610 27776 7930 28676
rect 7610 27712 7618 27776
rect 7682 27712 7698 27776
rect 7762 27712 7778 27776
rect 7842 27712 7858 27776
rect 7922 27712 7930 27776
rect 7610 26688 7930 27712
rect 7610 26624 7618 26688
rect 7682 26624 7698 26688
rect 7762 26624 7778 26688
rect 7842 26624 7858 26688
rect 7922 26624 7930 26688
rect 5395 26620 5461 26621
rect 5395 26556 5396 26620
rect 5460 26556 5461 26620
rect 5395 26555 5461 26556
rect 4277 26080 4285 26144
rect 4349 26080 4365 26144
rect 4429 26080 4445 26144
rect 4509 26080 4525 26144
rect 4589 26080 4597 26144
rect 4277 25056 4597 26080
rect 4277 24992 4285 25056
rect 4349 24992 4365 25056
rect 4429 24992 4445 25056
rect 4509 24992 4525 25056
rect 4589 24992 4597 25056
rect 4277 23968 4597 24992
rect 4277 23904 4285 23968
rect 4349 23904 4365 23968
rect 4429 23904 4445 23968
rect 4509 23904 4525 23968
rect 4589 23904 4597 23968
rect 4277 22880 4597 23904
rect 4277 22816 4285 22880
rect 4349 22816 4365 22880
rect 4429 22816 4445 22880
rect 4509 22816 4525 22880
rect 4589 22816 4597 22880
rect 4277 21792 4597 22816
rect 4277 21728 4285 21792
rect 4349 21728 4365 21792
rect 4429 21728 4445 21792
rect 4509 21728 4525 21792
rect 4589 21728 4597 21792
rect 4277 20704 4597 21728
rect 4277 20640 4285 20704
rect 4349 20640 4365 20704
rect 4429 20640 4445 20704
rect 4509 20640 4525 20704
rect 4589 20640 4597 20704
rect 4277 19616 4597 20640
rect 4277 19552 4285 19616
rect 4349 19552 4365 19616
rect 4429 19552 4445 19616
rect 4509 19552 4525 19616
rect 4589 19552 4597 19616
rect 4277 18528 4597 19552
rect 4277 18464 4285 18528
rect 4349 18464 4365 18528
rect 4429 18464 4445 18528
rect 4509 18464 4525 18528
rect 4589 18464 4597 18528
rect 4277 17440 4597 18464
rect 4277 17376 4285 17440
rect 4349 17376 4365 17440
rect 4429 17376 4445 17440
rect 4509 17376 4525 17440
rect 4589 17376 4597 17440
rect 1715 17236 1781 17237
rect 1715 17172 1716 17236
rect 1780 17172 1781 17236
rect 1715 17171 1781 17172
rect 4277 16352 4597 17376
rect 4277 16288 4285 16352
rect 4349 16288 4365 16352
rect 4429 16288 4445 16352
rect 4509 16288 4525 16352
rect 4589 16288 4597 16352
rect 4277 15579 4597 16288
rect 4277 15343 4319 15579
rect 4555 15343 4597 15579
rect 4277 15264 4597 15343
rect 4277 15200 4285 15264
rect 4349 15200 4365 15264
rect 4429 15200 4445 15264
rect 4509 15200 4525 15264
rect 4589 15200 4597 15264
rect 4277 14176 4597 15200
rect 4277 14112 4285 14176
rect 4349 14112 4365 14176
rect 4429 14112 4445 14176
rect 4509 14112 4525 14176
rect 4589 14112 4597 14176
rect 4277 13088 4597 14112
rect 4277 13024 4285 13088
rect 4349 13024 4365 13088
rect 4429 13024 4445 13088
rect 4509 13024 4525 13088
rect 4589 13024 4597 13088
rect 4277 12000 4597 13024
rect 4277 11936 4285 12000
rect 4349 11936 4365 12000
rect 4429 11936 4445 12000
rect 4509 11936 4525 12000
rect 4589 11936 4597 12000
rect 4277 10912 4597 11936
rect 4277 10848 4285 10912
rect 4349 10848 4365 10912
rect 4429 10848 4445 10912
rect 4509 10848 4525 10912
rect 4589 10848 4597 10912
rect 4277 9824 4597 10848
rect 4277 9760 4285 9824
rect 4349 9760 4365 9824
rect 4429 9760 4445 9824
rect 4509 9760 4525 9824
rect 4589 9760 4597 9824
rect 4277 8736 4597 9760
rect 4277 8672 4285 8736
rect 4349 8672 4365 8736
rect 4429 8672 4445 8736
rect 4509 8672 4525 8736
rect 4589 8672 4597 8736
rect 4277 7648 4597 8672
rect 4277 7584 4285 7648
rect 4349 7584 4365 7648
rect 4429 7584 4445 7648
rect 4509 7584 4525 7648
rect 4589 7584 4597 7648
rect 4277 6560 4597 7584
rect 4277 6496 4285 6560
rect 4349 6496 4365 6560
rect 4429 6496 4445 6560
rect 4509 6496 4525 6560
rect 4589 6496 4597 6560
rect 4277 5472 4597 6496
rect 4277 5408 4285 5472
rect 4349 5408 4365 5472
rect 4429 5408 4445 5472
rect 4509 5408 4525 5472
rect 4589 5408 4597 5472
rect 4277 4384 4597 5408
rect 4277 4320 4285 4384
rect 4349 4320 4365 4384
rect 4429 4320 4445 4384
rect 4509 4320 4525 4384
rect 4589 4320 4597 4384
rect 4277 3296 4597 4320
rect 4277 3232 4285 3296
rect 4349 3232 4365 3296
rect 4429 3232 4445 3296
rect 4509 3232 4525 3296
rect 4589 3232 4597 3296
rect 4277 2208 4597 3232
rect 4277 2144 4285 2208
rect 4349 2144 4365 2208
rect 4429 2144 4445 2208
rect 4509 2144 4525 2208
rect 4589 2144 4597 2208
rect 4277 2128 4597 2144
rect 7610 25600 7930 26624
rect 9630 26485 9690 49811
rect 9814 45797 9874 54843
rect 9811 45796 9877 45797
rect 9811 45732 9812 45796
rect 9876 45732 9877 45796
rect 9811 45731 9877 45732
rect 9811 45524 9877 45525
rect 9811 45460 9812 45524
rect 9876 45460 9877 45524
rect 9811 45459 9877 45460
rect 9814 36821 9874 45459
rect 9998 43893 10058 62187
rect 10179 62116 10245 62117
rect 10179 62052 10180 62116
rect 10244 62052 10245 62116
rect 10179 62051 10245 62052
rect 9995 43892 10061 43893
rect 9995 43828 9996 43892
rect 10060 43828 10061 43892
rect 9995 43827 10061 43828
rect 10182 43349 10242 62051
rect 10366 57493 10426 65859
rect 10547 65244 10613 65245
rect 10547 65180 10548 65244
rect 10612 65180 10613 65244
rect 10547 65179 10613 65180
rect 10550 61301 10610 65179
rect 10547 61300 10613 61301
rect 10547 61236 10548 61300
rect 10612 61236 10613 61300
rect 10547 61235 10613 61236
rect 10547 61164 10613 61165
rect 10547 61100 10548 61164
rect 10612 61100 10613 61164
rect 10547 61099 10613 61100
rect 10363 57492 10429 57493
rect 10363 57428 10364 57492
rect 10428 57428 10429 57492
rect 10363 57427 10429 57428
rect 10363 56404 10429 56405
rect 10363 56340 10364 56404
rect 10428 56340 10429 56404
rect 10363 56339 10429 56340
rect 10366 52869 10426 56339
rect 10363 52868 10429 52869
rect 10363 52804 10364 52868
rect 10428 52804 10429 52868
rect 10363 52803 10429 52804
rect 10363 52596 10429 52597
rect 10363 52532 10364 52596
rect 10428 52532 10429 52596
rect 10363 52531 10429 52532
rect 10366 45933 10426 52531
rect 10550 51781 10610 61099
rect 10547 51780 10613 51781
rect 10547 51716 10548 51780
rect 10612 51716 10613 51780
rect 10547 51715 10613 51716
rect 10547 50964 10613 50965
rect 10547 50900 10548 50964
rect 10612 50900 10613 50964
rect 10547 50899 10613 50900
rect 10550 49877 10610 50899
rect 10547 49876 10613 49877
rect 10547 49812 10548 49876
rect 10612 49812 10613 49876
rect 10547 49811 10613 49812
rect 10547 49740 10613 49741
rect 10547 49676 10548 49740
rect 10612 49676 10613 49740
rect 10547 49675 10613 49676
rect 10363 45932 10429 45933
rect 10363 45868 10364 45932
rect 10428 45868 10429 45932
rect 10363 45867 10429 45868
rect 10179 43348 10245 43349
rect 10179 43284 10180 43348
rect 10244 43284 10245 43348
rect 10179 43283 10245 43284
rect 9995 42940 10061 42941
rect 9995 42876 9996 42940
rect 10060 42876 10061 42940
rect 9995 42875 10061 42876
rect 10363 42940 10429 42941
rect 10363 42876 10364 42940
rect 10428 42876 10429 42940
rect 10363 42875 10429 42876
rect 9998 39133 10058 42875
rect 9995 39132 10061 39133
rect 9995 39068 9996 39132
rect 10060 39068 10061 39132
rect 9995 39067 10061 39068
rect 9811 36820 9877 36821
rect 9811 36756 9812 36820
rect 9876 36756 9877 36820
rect 9811 36755 9877 36756
rect 10366 34101 10426 42875
rect 10363 34100 10429 34101
rect 10363 34036 10364 34100
rect 10428 34036 10429 34100
rect 10363 34035 10429 34036
rect 9627 26484 9693 26485
rect 9627 26420 9628 26484
rect 9692 26420 9693 26484
rect 9627 26419 9693 26420
rect 7610 25536 7618 25600
rect 7682 25536 7698 25600
rect 7762 25536 7778 25600
rect 7842 25536 7858 25600
rect 7922 25536 7930 25600
rect 7610 24512 7930 25536
rect 7610 24448 7618 24512
rect 7682 24448 7698 24512
rect 7762 24448 7778 24512
rect 7842 24448 7858 24512
rect 7922 24448 7930 24512
rect 7610 23424 7930 24448
rect 10550 24309 10610 49675
rect 10734 31381 10794 73203
rect 10944 72928 11264 73952
rect 10944 72864 10952 72928
rect 11016 72864 11032 72928
rect 11096 72864 11112 72928
rect 11176 72864 11192 72928
rect 11256 72864 11264 72928
rect 10944 71840 11264 72864
rect 10944 71776 10952 71840
rect 11016 71776 11032 71840
rect 11096 71776 11112 71840
rect 11176 71776 11192 71840
rect 11256 71776 11264 71840
rect 10944 70752 11264 71776
rect 10944 70688 10952 70752
rect 11016 70688 11032 70752
rect 11096 70688 11112 70752
rect 11176 70688 11192 70752
rect 11256 70688 11264 70752
rect 10944 69664 11264 70688
rect 10944 69600 10952 69664
rect 11016 69600 11032 69664
rect 11096 69600 11112 69664
rect 11176 69600 11192 69664
rect 11256 69600 11264 69664
rect 10944 68912 11264 69600
rect 14277 77824 14597 77840
rect 14277 77760 14285 77824
rect 14349 77760 14365 77824
rect 14429 77760 14445 77824
rect 14509 77760 14525 77824
rect 14589 77760 14597 77824
rect 14277 76736 14597 77760
rect 14963 77484 15029 77485
rect 14963 77420 14964 77484
rect 15028 77420 15029 77484
rect 14963 77419 15029 77420
rect 14277 76672 14285 76736
rect 14349 76672 14365 76736
rect 14429 76672 14445 76736
rect 14509 76672 14525 76736
rect 14589 76672 14597 76736
rect 14277 75648 14597 76672
rect 14277 75584 14285 75648
rect 14349 75584 14365 75648
rect 14429 75584 14445 75648
rect 14509 75584 14525 75648
rect 14589 75584 14597 75648
rect 14277 74560 14597 75584
rect 14277 74496 14285 74560
rect 14349 74496 14365 74560
rect 14429 74496 14445 74560
rect 14509 74496 14525 74560
rect 14589 74496 14597 74560
rect 14277 73472 14597 74496
rect 14277 73408 14285 73472
rect 14349 73408 14365 73472
rect 14429 73408 14445 73472
rect 14509 73408 14525 73472
rect 14589 73408 14597 73472
rect 14277 72384 14597 73408
rect 14277 72320 14285 72384
rect 14349 72320 14365 72384
rect 14429 72320 14445 72384
rect 14509 72320 14525 72384
rect 14589 72320 14597 72384
rect 14277 71296 14597 72320
rect 14277 71232 14285 71296
rect 14349 71232 14365 71296
rect 14429 71232 14445 71296
rect 14509 71232 14525 71296
rect 14589 71232 14597 71296
rect 14277 70208 14597 71232
rect 14277 70144 14285 70208
rect 14349 70144 14365 70208
rect 14429 70144 14445 70208
rect 14509 70144 14525 70208
rect 14589 70144 14597 70208
rect 14277 69120 14597 70144
rect 14277 69056 14285 69120
rect 14349 69056 14365 69120
rect 14429 69056 14445 69120
rect 14509 69056 14525 69120
rect 14589 69056 14597 69120
rect 12019 69052 12085 69053
rect 12019 68988 12020 69052
rect 12084 68988 12085 69052
rect 12019 68987 12085 68988
rect 10944 68676 10986 68912
rect 11222 68676 11264 68912
rect 10944 68576 11264 68676
rect 10944 68512 10952 68576
rect 11016 68512 11032 68576
rect 11096 68512 11112 68576
rect 11176 68512 11192 68576
rect 11256 68512 11264 68576
rect 10944 67488 11264 68512
rect 10944 67424 10952 67488
rect 11016 67424 11032 67488
rect 11096 67424 11112 67488
rect 11176 67424 11192 67488
rect 11256 67424 11264 67488
rect 10944 66400 11264 67424
rect 10944 66336 10952 66400
rect 11016 66336 11032 66400
rect 11096 66336 11112 66400
rect 11176 66336 11192 66400
rect 11256 66336 11264 66400
rect 10944 65312 11264 66336
rect 11467 65788 11533 65789
rect 11467 65724 11468 65788
rect 11532 65724 11533 65788
rect 11467 65723 11533 65724
rect 10944 65248 10952 65312
rect 11016 65248 11032 65312
rect 11096 65248 11112 65312
rect 11176 65248 11192 65312
rect 11256 65248 11264 65312
rect 10944 64224 11264 65248
rect 10944 64160 10952 64224
rect 11016 64160 11032 64224
rect 11096 64160 11112 64224
rect 11176 64160 11192 64224
rect 11256 64160 11264 64224
rect 10944 63136 11264 64160
rect 10944 63072 10952 63136
rect 11016 63072 11032 63136
rect 11096 63072 11112 63136
rect 11176 63072 11192 63136
rect 11256 63072 11264 63136
rect 10944 62048 11264 63072
rect 10944 61984 10952 62048
rect 11016 61984 11032 62048
rect 11096 61984 11112 62048
rect 11176 61984 11192 62048
rect 11256 61984 11264 62048
rect 10944 60960 11264 61984
rect 10944 60896 10952 60960
rect 11016 60896 11032 60960
rect 11096 60896 11112 60960
rect 11176 60896 11192 60960
rect 11256 60896 11264 60960
rect 10944 59872 11264 60896
rect 10944 59808 10952 59872
rect 11016 59808 11032 59872
rect 11096 59808 11112 59872
rect 11176 59808 11192 59872
rect 11256 59808 11264 59872
rect 10944 58784 11264 59808
rect 10944 58720 10952 58784
rect 11016 58720 11032 58784
rect 11096 58720 11112 58784
rect 11176 58720 11192 58784
rect 11256 58720 11264 58784
rect 10944 57696 11264 58720
rect 10944 57632 10952 57696
rect 11016 57632 11032 57696
rect 11096 57632 11112 57696
rect 11176 57632 11192 57696
rect 11256 57632 11264 57696
rect 10944 56608 11264 57632
rect 10944 56544 10952 56608
rect 11016 56544 11032 56608
rect 11096 56544 11112 56608
rect 11176 56544 11192 56608
rect 11256 56544 11264 56608
rect 10944 55520 11264 56544
rect 10944 55456 10952 55520
rect 11016 55456 11032 55520
rect 11096 55456 11112 55520
rect 11176 55456 11192 55520
rect 11256 55456 11264 55520
rect 10944 54432 11264 55456
rect 10944 54368 10952 54432
rect 11016 54368 11032 54432
rect 11096 54368 11112 54432
rect 11176 54368 11192 54432
rect 11256 54368 11264 54432
rect 10944 53344 11264 54368
rect 10944 53280 10952 53344
rect 11016 53280 11032 53344
rect 11096 53280 11112 53344
rect 11176 53280 11192 53344
rect 11256 53280 11264 53344
rect 10944 52256 11264 53280
rect 10944 52192 10952 52256
rect 11016 52192 11032 52256
rect 11096 52192 11112 52256
rect 11176 52192 11192 52256
rect 11256 52192 11264 52256
rect 10944 51168 11264 52192
rect 10944 51104 10952 51168
rect 11016 51104 11032 51168
rect 11096 51104 11112 51168
rect 11176 51104 11192 51168
rect 11256 51104 11264 51168
rect 10944 50080 11264 51104
rect 11470 50690 11530 65723
rect 12022 62389 12082 68987
rect 14043 68372 14109 68373
rect 14043 68308 14044 68372
rect 14108 68308 14109 68372
rect 14043 68307 14109 68308
rect 13859 68100 13925 68101
rect 13859 68036 13860 68100
rect 13924 68036 13925 68100
rect 13859 68035 13925 68036
rect 12019 62388 12085 62389
rect 12019 62324 12020 62388
rect 12084 62324 12085 62388
rect 12019 62323 12085 62324
rect 12203 62252 12269 62253
rect 12203 62188 12204 62252
rect 12268 62188 12269 62252
rect 12203 62187 12269 62188
rect 11835 57764 11901 57765
rect 11835 57700 11836 57764
rect 11900 57700 11901 57764
rect 11835 57699 11901 57700
rect 11651 55316 11717 55317
rect 11651 55252 11652 55316
rect 11716 55252 11717 55316
rect 11651 55251 11717 55252
rect 11654 50829 11714 55251
rect 11838 54229 11898 57699
rect 12019 55180 12085 55181
rect 12019 55116 12020 55180
rect 12084 55116 12085 55180
rect 12019 55115 12085 55116
rect 11835 54228 11901 54229
rect 11835 54164 11836 54228
rect 11900 54164 11901 54228
rect 11835 54163 11901 54164
rect 11835 53956 11901 53957
rect 11835 53892 11836 53956
rect 11900 53892 11901 53956
rect 11835 53891 11901 53892
rect 11651 50828 11717 50829
rect 11651 50764 11652 50828
rect 11716 50764 11717 50828
rect 11651 50763 11717 50764
rect 11470 50630 11714 50690
rect 11467 50556 11533 50557
rect 11467 50492 11468 50556
rect 11532 50492 11533 50556
rect 11467 50491 11533 50492
rect 10944 50016 10952 50080
rect 11016 50016 11032 50080
rect 11096 50016 11112 50080
rect 11176 50016 11192 50080
rect 11256 50016 11264 50080
rect 10944 48992 11264 50016
rect 10944 48928 10952 48992
rect 11016 48928 11032 48992
rect 11096 48928 11112 48992
rect 11176 48928 11192 48992
rect 11256 48928 11264 48992
rect 10944 47904 11264 48928
rect 10944 47840 10952 47904
rect 11016 47840 11032 47904
rect 11096 47840 11112 47904
rect 11176 47840 11192 47904
rect 11256 47840 11264 47904
rect 10944 46816 11264 47840
rect 10944 46752 10952 46816
rect 11016 46752 11032 46816
rect 11096 46752 11112 46816
rect 11176 46752 11192 46816
rect 11256 46752 11264 46816
rect 10944 45728 11264 46752
rect 10944 45664 10952 45728
rect 11016 45664 11032 45728
rect 11096 45664 11112 45728
rect 11176 45664 11192 45728
rect 11256 45664 11264 45728
rect 10944 44640 11264 45664
rect 10944 44576 10952 44640
rect 11016 44576 11032 44640
rect 11096 44576 11112 44640
rect 11176 44576 11192 44640
rect 11256 44576 11264 44640
rect 10944 43552 11264 44576
rect 10944 43488 10952 43552
rect 11016 43488 11032 43552
rect 11096 43488 11112 43552
rect 11176 43488 11192 43552
rect 11256 43488 11264 43552
rect 10944 42464 11264 43488
rect 10944 42400 10952 42464
rect 11016 42400 11032 42464
rect 11096 42400 11112 42464
rect 11176 42400 11192 42464
rect 11256 42400 11264 42464
rect 10944 42246 11264 42400
rect 10944 42010 10986 42246
rect 11222 42010 11264 42246
rect 10944 41376 11264 42010
rect 10944 41312 10952 41376
rect 11016 41312 11032 41376
rect 11096 41312 11112 41376
rect 11176 41312 11192 41376
rect 11256 41312 11264 41376
rect 10944 40288 11264 41312
rect 10944 40224 10952 40288
rect 11016 40224 11032 40288
rect 11096 40224 11112 40288
rect 11176 40224 11192 40288
rect 11256 40224 11264 40288
rect 10944 39200 11264 40224
rect 11470 39949 11530 50491
rect 11654 45797 11714 50630
rect 11651 45796 11717 45797
rect 11651 45732 11652 45796
rect 11716 45732 11717 45796
rect 11651 45731 11717 45732
rect 11651 42260 11717 42261
rect 11651 42196 11652 42260
rect 11716 42196 11717 42260
rect 11651 42195 11717 42196
rect 11654 39949 11714 42195
rect 11467 39948 11533 39949
rect 11467 39884 11468 39948
rect 11532 39884 11533 39948
rect 11467 39883 11533 39884
rect 11651 39948 11717 39949
rect 11651 39884 11652 39948
rect 11716 39884 11717 39948
rect 11651 39883 11717 39884
rect 11838 39810 11898 53891
rect 10944 39136 10952 39200
rect 11016 39136 11032 39200
rect 11096 39136 11112 39200
rect 11176 39136 11192 39200
rect 11256 39136 11264 39200
rect 10944 38112 11264 39136
rect 10944 38048 10952 38112
rect 11016 38048 11032 38112
rect 11096 38048 11112 38112
rect 11176 38048 11192 38112
rect 11256 38048 11264 38112
rect 10944 37024 11264 38048
rect 10944 36960 10952 37024
rect 11016 36960 11032 37024
rect 11096 36960 11112 37024
rect 11176 36960 11192 37024
rect 11256 36960 11264 37024
rect 10944 35936 11264 36960
rect 10944 35872 10952 35936
rect 11016 35872 11032 35936
rect 11096 35872 11112 35936
rect 11176 35872 11192 35936
rect 11256 35872 11264 35936
rect 10944 34848 11264 35872
rect 10944 34784 10952 34848
rect 11016 34784 11032 34848
rect 11096 34784 11112 34848
rect 11176 34784 11192 34848
rect 11256 34784 11264 34848
rect 10944 33760 11264 34784
rect 10944 33696 10952 33760
rect 11016 33696 11032 33760
rect 11096 33696 11112 33760
rect 11176 33696 11192 33760
rect 11256 33696 11264 33760
rect 10944 32672 11264 33696
rect 11654 39750 11898 39810
rect 11654 33149 11714 39750
rect 11651 33148 11717 33149
rect 11651 33084 11652 33148
rect 11716 33084 11717 33148
rect 11651 33083 11717 33084
rect 10944 32608 10952 32672
rect 11016 32608 11032 32672
rect 11096 32608 11112 32672
rect 11176 32608 11192 32672
rect 11256 32608 11264 32672
rect 10944 31584 11264 32608
rect 10944 31520 10952 31584
rect 11016 31520 11032 31584
rect 11096 31520 11112 31584
rect 11176 31520 11192 31584
rect 11256 31520 11264 31584
rect 10731 31380 10797 31381
rect 10731 31316 10732 31380
rect 10796 31316 10797 31380
rect 10731 31315 10797 31316
rect 10944 30496 11264 31520
rect 10944 30432 10952 30496
rect 11016 30432 11032 30496
rect 11096 30432 11112 30496
rect 11176 30432 11192 30496
rect 11256 30432 11264 30496
rect 10944 29408 11264 30432
rect 12022 29749 12082 55115
rect 12206 46205 12266 62187
rect 12571 56676 12637 56677
rect 12571 56612 12572 56676
rect 12636 56612 12637 56676
rect 12571 56611 12637 56612
rect 12387 56540 12453 56541
rect 12387 56476 12388 56540
rect 12452 56476 12453 56540
rect 12387 56475 12453 56476
rect 12390 54909 12450 56475
rect 12574 55181 12634 56611
rect 12571 55180 12637 55181
rect 12571 55116 12572 55180
rect 12636 55116 12637 55180
rect 12571 55115 12637 55116
rect 12387 54908 12453 54909
rect 12387 54844 12388 54908
rect 12452 54844 12453 54908
rect 12387 54843 12453 54844
rect 12387 54228 12453 54229
rect 12387 54164 12388 54228
rect 12452 54164 12453 54228
rect 12387 54163 12453 54164
rect 12390 47970 12450 54163
rect 13123 53820 13189 53821
rect 13123 53756 13124 53820
rect 13188 53756 13189 53820
rect 13123 53755 13189 53756
rect 12571 52732 12637 52733
rect 12571 52668 12572 52732
rect 12636 52668 12637 52732
rect 12571 52667 12637 52668
rect 12574 49333 12634 52667
rect 12755 51508 12821 51509
rect 12755 51444 12756 51508
rect 12820 51444 12821 51508
rect 12755 51443 12821 51444
rect 12571 49332 12637 49333
rect 12571 49268 12572 49332
rect 12636 49268 12637 49332
rect 12571 49267 12637 49268
rect 12758 48789 12818 51443
rect 12939 51100 13005 51101
rect 12939 51036 12940 51100
rect 13004 51036 13005 51100
rect 12939 51035 13005 51036
rect 12755 48788 12821 48789
rect 12755 48724 12756 48788
rect 12820 48724 12821 48788
rect 12755 48723 12821 48724
rect 12942 48381 13002 51035
rect 13126 49197 13186 53755
rect 13491 52732 13557 52733
rect 13491 52668 13492 52732
rect 13556 52668 13557 52732
rect 13491 52667 13557 52668
rect 13307 52460 13373 52461
rect 13307 52396 13308 52460
rect 13372 52396 13373 52460
rect 13307 52395 13373 52396
rect 13310 50285 13370 52395
rect 13494 50965 13554 52667
rect 13491 50964 13557 50965
rect 13491 50900 13492 50964
rect 13556 50900 13557 50964
rect 13491 50899 13557 50900
rect 13675 50964 13741 50965
rect 13675 50900 13676 50964
rect 13740 50900 13741 50964
rect 13675 50899 13741 50900
rect 13491 50692 13557 50693
rect 13491 50628 13492 50692
rect 13556 50628 13557 50692
rect 13491 50627 13557 50628
rect 13307 50284 13373 50285
rect 13307 50220 13308 50284
rect 13372 50220 13373 50284
rect 13307 50219 13373 50220
rect 13307 50148 13373 50149
rect 13307 50084 13308 50148
rect 13372 50084 13373 50148
rect 13307 50083 13373 50084
rect 13123 49196 13189 49197
rect 13123 49132 13124 49196
rect 13188 49132 13189 49196
rect 13123 49131 13189 49132
rect 12939 48380 13005 48381
rect 12939 48316 12940 48380
rect 13004 48316 13005 48380
rect 12939 48315 13005 48316
rect 12390 47910 12634 47970
rect 12387 47700 12453 47701
rect 12387 47636 12388 47700
rect 12452 47636 12453 47700
rect 12387 47635 12453 47636
rect 12203 46204 12269 46205
rect 12203 46140 12204 46204
rect 12268 46140 12269 46204
rect 12203 46139 12269 46140
rect 12390 45930 12450 47635
rect 12574 47293 12634 47910
rect 12755 47428 12821 47429
rect 12755 47364 12756 47428
rect 12820 47364 12821 47428
rect 12755 47363 12821 47364
rect 12571 47292 12637 47293
rect 12571 47228 12572 47292
rect 12636 47228 12637 47292
rect 12571 47227 12637 47228
rect 12571 46204 12637 46205
rect 12571 46140 12572 46204
rect 12636 46140 12637 46204
rect 12571 46139 12637 46140
rect 12206 45870 12450 45930
rect 12206 45253 12266 45870
rect 12387 45796 12453 45797
rect 12387 45732 12388 45796
rect 12452 45732 12453 45796
rect 12387 45731 12453 45732
rect 12203 45252 12269 45253
rect 12203 45188 12204 45252
rect 12268 45188 12269 45252
rect 12203 45187 12269 45188
rect 12390 45114 12450 45731
rect 12206 45054 12450 45114
rect 12206 38997 12266 45054
rect 12574 39405 12634 46139
rect 12571 39404 12637 39405
rect 12571 39340 12572 39404
rect 12636 39340 12637 39404
rect 12571 39339 12637 39340
rect 12203 38996 12269 38997
rect 12203 38932 12204 38996
rect 12268 38932 12269 38996
rect 12203 38931 12269 38932
rect 12758 38725 12818 47363
rect 13310 46341 13370 50083
rect 13494 49197 13554 50627
rect 13491 49196 13557 49197
rect 13491 49132 13492 49196
rect 13556 49132 13557 49196
rect 13491 49131 13557 49132
rect 13307 46340 13373 46341
rect 13307 46276 13308 46340
rect 13372 46276 13373 46340
rect 13307 46275 13373 46276
rect 13678 43757 13738 50899
rect 13675 43756 13741 43757
rect 13675 43692 13676 43756
rect 13740 43692 13741 43756
rect 13675 43691 13741 43692
rect 13675 41172 13741 41173
rect 13675 41108 13676 41172
rect 13740 41108 13741 41172
rect 13675 41107 13741 41108
rect 13491 41036 13557 41037
rect 13491 40972 13492 41036
rect 13556 40972 13557 41036
rect 13491 40971 13557 40972
rect 13494 39541 13554 40971
rect 13491 39540 13557 39541
rect 13491 39476 13492 39540
rect 13556 39476 13557 39540
rect 13491 39475 13557 39476
rect 12755 38724 12821 38725
rect 12755 38660 12756 38724
rect 12820 38660 12821 38724
rect 12755 38659 12821 38660
rect 13678 35053 13738 41107
rect 13675 35052 13741 35053
rect 13675 34988 13676 35052
rect 13740 34988 13741 35052
rect 13675 34987 13741 34988
rect 13862 31925 13922 68035
rect 14046 61029 14106 68307
rect 14277 68032 14597 69056
rect 14277 67968 14285 68032
rect 14349 67968 14365 68032
rect 14429 67968 14445 68032
rect 14509 67968 14525 68032
rect 14589 67968 14597 68032
rect 14277 66944 14597 67968
rect 14277 66880 14285 66944
rect 14349 66880 14365 66944
rect 14429 66880 14445 66944
rect 14509 66880 14525 66944
rect 14589 66880 14597 66944
rect 14277 65856 14597 66880
rect 14779 65924 14845 65925
rect 14779 65860 14780 65924
rect 14844 65860 14845 65924
rect 14779 65859 14845 65860
rect 14277 65792 14285 65856
rect 14349 65792 14365 65856
rect 14429 65792 14445 65856
rect 14509 65792 14525 65856
rect 14589 65792 14597 65856
rect 14277 64768 14597 65792
rect 14277 64704 14285 64768
rect 14349 64704 14365 64768
rect 14429 64704 14445 64768
rect 14509 64704 14525 64768
rect 14589 64704 14597 64768
rect 14277 63680 14597 64704
rect 14277 63616 14285 63680
rect 14349 63616 14365 63680
rect 14429 63616 14445 63680
rect 14509 63616 14525 63680
rect 14589 63616 14597 63680
rect 14277 62592 14597 63616
rect 14277 62528 14285 62592
rect 14349 62528 14365 62592
rect 14429 62528 14445 62592
rect 14509 62528 14525 62592
rect 14589 62528 14597 62592
rect 14277 61504 14597 62528
rect 14277 61440 14285 61504
rect 14349 61440 14365 61504
rect 14429 61440 14445 61504
rect 14509 61440 14525 61504
rect 14589 61440 14597 61504
rect 14043 61028 14109 61029
rect 14043 60964 14044 61028
rect 14108 60964 14109 61028
rect 14043 60963 14109 60964
rect 14043 60756 14109 60757
rect 14043 60692 14044 60756
rect 14108 60692 14109 60756
rect 14043 60691 14109 60692
rect 13859 31924 13925 31925
rect 13859 31860 13860 31924
rect 13924 31860 13925 31924
rect 13859 31859 13925 31860
rect 14046 30701 14106 60691
rect 14277 60416 14597 61440
rect 14782 61301 14842 65859
rect 14779 61300 14845 61301
rect 14779 61236 14780 61300
rect 14844 61236 14845 61300
rect 14779 61235 14845 61236
rect 14779 60756 14845 60757
rect 14779 60692 14780 60756
rect 14844 60692 14845 60756
rect 14779 60691 14845 60692
rect 14277 60352 14285 60416
rect 14349 60352 14365 60416
rect 14429 60352 14445 60416
rect 14509 60352 14525 60416
rect 14589 60352 14597 60416
rect 14277 59328 14597 60352
rect 14277 59264 14285 59328
rect 14349 59264 14365 59328
rect 14429 59264 14445 59328
rect 14509 59264 14525 59328
rect 14589 59264 14597 59328
rect 14277 58240 14597 59264
rect 14277 58176 14285 58240
rect 14349 58176 14365 58240
rect 14429 58176 14445 58240
rect 14509 58176 14525 58240
rect 14589 58176 14597 58240
rect 14277 57152 14597 58176
rect 14277 57088 14285 57152
rect 14349 57088 14365 57152
rect 14429 57088 14445 57152
rect 14509 57088 14525 57152
rect 14589 57088 14597 57152
rect 14277 56064 14597 57088
rect 14277 56000 14285 56064
rect 14349 56000 14365 56064
rect 14429 56000 14445 56064
rect 14509 56000 14525 56064
rect 14589 56000 14597 56064
rect 14277 55579 14597 56000
rect 14277 55343 14319 55579
rect 14555 55343 14597 55579
rect 14277 54976 14597 55343
rect 14277 54912 14285 54976
rect 14349 54912 14365 54976
rect 14429 54912 14445 54976
rect 14509 54912 14525 54976
rect 14589 54912 14597 54976
rect 14277 53888 14597 54912
rect 14277 53824 14285 53888
rect 14349 53824 14365 53888
rect 14429 53824 14445 53888
rect 14509 53824 14525 53888
rect 14589 53824 14597 53888
rect 14277 52800 14597 53824
rect 14277 52736 14285 52800
rect 14349 52736 14365 52800
rect 14429 52736 14445 52800
rect 14509 52736 14525 52800
rect 14589 52736 14597 52800
rect 14277 51712 14597 52736
rect 14277 51648 14285 51712
rect 14349 51648 14365 51712
rect 14429 51648 14445 51712
rect 14509 51648 14525 51712
rect 14589 51648 14597 51712
rect 14277 50624 14597 51648
rect 14782 51101 14842 60691
rect 14966 53410 15026 77419
rect 17610 77280 17930 77840
rect 17610 77216 17618 77280
rect 17682 77216 17698 77280
rect 17762 77216 17778 77280
rect 17842 77216 17858 77280
rect 17922 77216 17930 77280
rect 17610 76192 17930 77216
rect 17610 76128 17618 76192
rect 17682 76128 17698 76192
rect 17762 76128 17778 76192
rect 17842 76128 17858 76192
rect 17922 76128 17930 76192
rect 17610 75104 17930 76128
rect 17610 75040 17618 75104
rect 17682 75040 17698 75104
rect 17762 75040 17778 75104
rect 17842 75040 17858 75104
rect 17922 75040 17930 75104
rect 17610 74016 17930 75040
rect 17610 73952 17618 74016
rect 17682 73952 17698 74016
rect 17762 73952 17778 74016
rect 17842 73952 17858 74016
rect 17922 73952 17930 74016
rect 17610 72928 17930 73952
rect 17610 72864 17618 72928
rect 17682 72864 17698 72928
rect 17762 72864 17778 72928
rect 17842 72864 17858 72928
rect 17922 72864 17930 72928
rect 17610 71840 17930 72864
rect 17610 71776 17618 71840
rect 17682 71776 17698 71840
rect 17762 71776 17778 71840
rect 17842 71776 17858 71840
rect 17922 71776 17930 71840
rect 16619 71364 16685 71365
rect 16619 71300 16620 71364
rect 16684 71300 16685 71364
rect 16619 71299 16685 71300
rect 15331 61300 15397 61301
rect 15331 61236 15332 61300
rect 15396 61236 15397 61300
rect 15331 61235 15397 61236
rect 14966 53350 15210 53410
rect 14963 52868 15029 52869
rect 14963 52804 14964 52868
rect 15028 52804 15029 52868
rect 14963 52803 15029 52804
rect 14779 51100 14845 51101
rect 14779 51036 14780 51100
rect 14844 51036 14845 51100
rect 14779 51035 14845 51036
rect 14779 50964 14845 50965
rect 14779 50900 14780 50964
rect 14844 50900 14845 50964
rect 14779 50899 14845 50900
rect 14277 50560 14285 50624
rect 14349 50560 14365 50624
rect 14429 50560 14445 50624
rect 14509 50560 14525 50624
rect 14589 50560 14597 50624
rect 14277 49536 14597 50560
rect 14277 49472 14285 49536
rect 14349 49472 14365 49536
rect 14429 49472 14445 49536
rect 14509 49472 14525 49536
rect 14589 49472 14597 49536
rect 14277 48448 14597 49472
rect 14277 48384 14285 48448
rect 14349 48384 14365 48448
rect 14429 48384 14445 48448
rect 14509 48384 14525 48448
rect 14589 48384 14597 48448
rect 14277 47360 14597 48384
rect 14277 47296 14285 47360
rect 14349 47296 14365 47360
rect 14429 47296 14445 47360
rect 14509 47296 14525 47360
rect 14589 47296 14597 47360
rect 14277 46272 14597 47296
rect 14277 46208 14285 46272
rect 14349 46208 14365 46272
rect 14429 46208 14445 46272
rect 14509 46208 14525 46272
rect 14589 46208 14597 46272
rect 14277 45184 14597 46208
rect 14277 45120 14285 45184
rect 14349 45120 14365 45184
rect 14429 45120 14445 45184
rect 14509 45120 14525 45184
rect 14589 45120 14597 45184
rect 14277 44096 14597 45120
rect 14277 44032 14285 44096
rect 14349 44032 14365 44096
rect 14429 44032 14445 44096
rect 14509 44032 14525 44096
rect 14589 44032 14597 44096
rect 14277 43008 14597 44032
rect 14277 42944 14285 43008
rect 14349 42944 14365 43008
rect 14429 42944 14445 43008
rect 14509 42944 14525 43008
rect 14589 42944 14597 43008
rect 14277 41920 14597 42944
rect 14277 41856 14285 41920
rect 14349 41856 14365 41920
rect 14429 41856 14445 41920
rect 14509 41856 14525 41920
rect 14589 41856 14597 41920
rect 14277 40832 14597 41856
rect 14782 41173 14842 50899
rect 14779 41172 14845 41173
rect 14779 41108 14780 41172
rect 14844 41108 14845 41172
rect 14779 41107 14845 41108
rect 14779 41036 14845 41037
rect 14779 40972 14780 41036
rect 14844 40972 14845 41036
rect 14779 40971 14845 40972
rect 14277 40768 14285 40832
rect 14349 40768 14365 40832
rect 14429 40768 14445 40832
rect 14509 40768 14525 40832
rect 14589 40768 14597 40832
rect 14277 39744 14597 40768
rect 14277 39680 14285 39744
rect 14349 39680 14365 39744
rect 14429 39680 14445 39744
rect 14509 39680 14525 39744
rect 14589 39680 14597 39744
rect 14277 38656 14597 39680
rect 14277 38592 14285 38656
rect 14349 38592 14365 38656
rect 14429 38592 14445 38656
rect 14509 38592 14525 38656
rect 14589 38592 14597 38656
rect 14277 37568 14597 38592
rect 14277 37504 14285 37568
rect 14349 37504 14365 37568
rect 14429 37504 14445 37568
rect 14509 37504 14525 37568
rect 14589 37504 14597 37568
rect 14277 36480 14597 37504
rect 14782 37229 14842 40971
rect 14779 37228 14845 37229
rect 14779 37164 14780 37228
rect 14844 37164 14845 37228
rect 14779 37163 14845 37164
rect 14277 36416 14285 36480
rect 14349 36416 14365 36480
rect 14429 36416 14445 36480
rect 14509 36416 14525 36480
rect 14589 36416 14597 36480
rect 14277 35392 14597 36416
rect 14277 35328 14285 35392
rect 14349 35328 14365 35392
rect 14429 35328 14445 35392
rect 14509 35328 14525 35392
rect 14589 35328 14597 35392
rect 14277 34304 14597 35328
rect 14277 34240 14285 34304
rect 14349 34240 14365 34304
rect 14429 34240 14445 34304
rect 14509 34240 14525 34304
rect 14589 34240 14597 34304
rect 14277 33216 14597 34240
rect 14277 33152 14285 33216
rect 14349 33152 14365 33216
rect 14429 33152 14445 33216
rect 14509 33152 14525 33216
rect 14589 33152 14597 33216
rect 14277 32128 14597 33152
rect 14966 32333 15026 52803
rect 15150 52594 15210 53350
rect 15334 52869 15394 61235
rect 15331 52868 15397 52869
rect 15331 52804 15332 52868
rect 15396 52804 15397 52868
rect 15331 52803 15397 52804
rect 15150 52534 15394 52594
rect 15147 51100 15213 51101
rect 15147 51036 15148 51100
rect 15212 51036 15213 51100
rect 15147 51035 15213 51036
rect 15150 41037 15210 51035
rect 15334 46749 15394 52534
rect 15331 46748 15397 46749
rect 15331 46684 15332 46748
rect 15396 46684 15397 46748
rect 15331 46683 15397 46684
rect 15331 45660 15397 45661
rect 15331 45596 15332 45660
rect 15396 45596 15397 45660
rect 15331 45595 15397 45596
rect 15334 43213 15394 45595
rect 15699 45116 15765 45117
rect 15699 45052 15700 45116
rect 15764 45052 15765 45116
rect 15699 45051 15765 45052
rect 15515 43892 15581 43893
rect 15515 43828 15516 43892
rect 15580 43828 15581 43892
rect 15515 43827 15581 43828
rect 15331 43212 15397 43213
rect 15331 43148 15332 43212
rect 15396 43148 15397 43212
rect 15331 43147 15397 43148
rect 15331 41580 15397 41581
rect 15331 41516 15332 41580
rect 15396 41516 15397 41580
rect 15331 41515 15397 41516
rect 15334 41309 15394 41515
rect 15331 41308 15397 41309
rect 15331 41244 15332 41308
rect 15396 41244 15397 41308
rect 15331 41243 15397 41244
rect 15147 41036 15213 41037
rect 15147 40972 15148 41036
rect 15212 40972 15213 41036
rect 15518 41034 15578 43827
rect 15147 40971 15213 40972
rect 15334 40974 15578 41034
rect 15147 38316 15213 38317
rect 15147 38252 15148 38316
rect 15212 38252 15213 38316
rect 15147 38251 15213 38252
rect 15150 34101 15210 38251
rect 15334 37501 15394 40974
rect 15515 40764 15581 40765
rect 15515 40700 15516 40764
rect 15580 40700 15581 40764
rect 15515 40699 15581 40700
rect 15518 39269 15578 40699
rect 15515 39268 15581 39269
rect 15515 39204 15516 39268
rect 15580 39204 15581 39268
rect 15515 39203 15581 39204
rect 15331 37500 15397 37501
rect 15331 37436 15332 37500
rect 15396 37436 15397 37500
rect 15331 37435 15397 37436
rect 15702 35733 15762 45051
rect 16435 43484 16501 43485
rect 16435 43420 16436 43484
rect 16500 43420 16501 43484
rect 16435 43419 16501 43420
rect 16067 42804 16133 42805
rect 16067 42740 16068 42804
rect 16132 42740 16133 42804
rect 16067 42739 16133 42740
rect 15883 41172 15949 41173
rect 15883 41108 15884 41172
rect 15948 41108 15949 41172
rect 15883 41107 15949 41108
rect 15886 38589 15946 41107
rect 16070 39541 16130 42739
rect 16438 41581 16498 43419
rect 16435 41580 16501 41581
rect 16435 41516 16436 41580
rect 16500 41516 16501 41580
rect 16435 41515 16501 41516
rect 16435 40356 16501 40357
rect 16435 40292 16436 40356
rect 16500 40292 16501 40356
rect 16435 40291 16501 40292
rect 16067 39540 16133 39541
rect 16067 39476 16068 39540
rect 16132 39476 16133 39540
rect 16067 39475 16133 39476
rect 15883 38588 15949 38589
rect 15883 38524 15884 38588
rect 15948 38524 15949 38588
rect 15883 38523 15949 38524
rect 15699 35732 15765 35733
rect 15699 35668 15700 35732
rect 15764 35668 15765 35732
rect 15699 35667 15765 35668
rect 16438 34509 16498 40291
rect 16435 34508 16501 34509
rect 16435 34444 16436 34508
rect 16500 34444 16501 34508
rect 16435 34443 16501 34444
rect 15147 34100 15213 34101
rect 15147 34036 15148 34100
rect 15212 34036 15213 34100
rect 15147 34035 15213 34036
rect 16622 33421 16682 71299
rect 17610 70752 17930 71776
rect 17610 70688 17618 70752
rect 17682 70688 17698 70752
rect 17762 70688 17778 70752
rect 17842 70688 17858 70752
rect 17922 70688 17930 70752
rect 17610 69664 17930 70688
rect 17610 69600 17618 69664
rect 17682 69600 17698 69664
rect 17762 69600 17778 69664
rect 17842 69600 17858 69664
rect 17922 69600 17930 69664
rect 17610 68912 17930 69600
rect 17610 68676 17652 68912
rect 17888 68676 17930 68912
rect 17610 68576 17930 68676
rect 17610 68512 17618 68576
rect 17682 68512 17698 68576
rect 17762 68512 17778 68576
rect 17842 68512 17858 68576
rect 17922 68512 17930 68576
rect 17610 67488 17930 68512
rect 17610 67424 17618 67488
rect 17682 67424 17698 67488
rect 17762 67424 17778 67488
rect 17842 67424 17858 67488
rect 17922 67424 17930 67488
rect 17610 66400 17930 67424
rect 17610 66336 17618 66400
rect 17682 66336 17698 66400
rect 17762 66336 17778 66400
rect 17842 66336 17858 66400
rect 17922 66336 17930 66400
rect 17610 65312 17930 66336
rect 17610 65248 17618 65312
rect 17682 65248 17698 65312
rect 17762 65248 17778 65312
rect 17842 65248 17858 65312
rect 17922 65248 17930 65312
rect 17610 64224 17930 65248
rect 17610 64160 17618 64224
rect 17682 64160 17698 64224
rect 17762 64160 17778 64224
rect 17842 64160 17858 64224
rect 17922 64160 17930 64224
rect 17610 63136 17930 64160
rect 17610 63072 17618 63136
rect 17682 63072 17698 63136
rect 17762 63072 17778 63136
rect 17842 63072 17858 63136
rect 17922 63072 17930 63136
rect 17610 62048 17930 63072
rect 17610 61984 17618 62048
rect 17682 61984 17698 62048
rect 17762 61984 17778 62048
rect 17842 61984 17858 62048
rect 17922 61984 17930 62048
rect 17610 60960 17930 61984
rect 17610 60896 17618 60960
rect 17682 60896 17698 60960
rect 17762 60896 17778 60960
rect 17842 60896 17858 60960
rect 17922 60896 17930 60960
rect 17610 59872 17930 60896
rect 17610 59808 17618 59872
rect 17682 59808 17698 59872
rect 17762 59808 17778 59872
rect 17842 59808 17858 59872
rect 17922 59808 17930 59872
rect 17610 58784 17930 59808
rect 17610 58720 17618 58784
rect 17682 58720 17698 58784
rect 17762 58720 17778 58784
rect 17842 58720 17858 58784
rect 17922 58720 17930 58784
rect 17610 57696 17930 58720
rect 17610 57632 17618 57696
rect 17682 57632 17698 57696
rect 17762 57632 17778 57696
rect 17842 57632 17858 57696
rect 17922 57632 17930 57696
rect 17610 56608 17930 57632
rect 17610 56544 17618 56608
rect 17682 56544 17698 56608
rect 17762 56544 17778 56608
rect 17842 56544 17858 56608
rect 17922 56544 17930 56608
rect 17610 55520 17930 56544
rect 17610 55456 17618 55520
rect 17682 55456 17698 55520
rect 17762 55456 17778 55520
rect 17842 55456 17858 55520
rect 17922 55456 17930 55520
rect 17610 54432 17930 55456
rect 17610 54368 17618 54432
rect 17682 54368 17698 54432
rect 17762 54368 17778 54432
rect 17842 54368 17858 54432
rect 17922 54368 17930 54432
rect 17171 53412 17237 53413
rect 17171 53348 17172 53412
rect 17236 53348 17237 53412
rect 17171 53347 17237 53348
rect 16987 46476 17053 46477
rect 16987 46412 16988 46476
rect 17052 46412 17053 46476
rect 16987 46411 17053 46412
rect 16803 41852 16869 41853
rect 16803 41788 16804 41852
rect 16868 41788 16869 41852
rect 16803 41787 16869 41788
rect 16806 41445 16866 41787
rect 16990 41717 17050 46411
rect 16987 41716 17053 41717
rect 16987 41652 16988 41716
rect 17052 41652 17053 41716
rect 16987 41651 17053 41652
rect 16803 41444 16869 41445
rect 16803 41380 16804 41444
rect 16868 41380 16869 41444
rect 16803 41379 16869 41380
rect 16987 41444 17053 41445
rect 16987 41380 16988 41444
rect 17052 41380 17053 41444
rect 16987 41379 17053 41380
rect 16806 41309 16866 41379
rect 16803 41308 16869 41309
rect 16803 41244 16804 41308
rect 16868 41244 16869 41308
rect 16803 41243 16869 41244
rect 16990 41170 17050 41379
rect 16806 41110 17050 41170
rect 16806 37229 16866 41110
rect 17174 40490 17234 53347
rect 17610 53344 17930 54368
rect 17610 53280 17618 53344
rect 17682 53280 17698 53344
rect 17762 53280 17778 53344
rect 17842 53280 17858 53344
rect 17922 53280 17930 53344
rect 17355 52324 17421 52325
rect 17355 52260 17356 52324
rect 17420 52260 17421 52324
rect 17355 52259 17421 52260
rect 16990 40430 17234 40490
rect 16803 37228 16869 37229
rect 16803 37164 16804 37228
rect 16868 37164 16869 37228
rect 16803 37163 16869 37164
rect 16990 33557 17050 40430
rect 17171 40084 17237 40085
rect 17171 40020 17172 40084
rect 17236 40020 17237 40084
rect 17171 40019 17237 40020
rect 16987 33556 17053 33557
rect 16987 33492 16988 33556
rect 17052 33492 17053 33556
rect 16987 33491 17053 33492
rect 16619 33420 16685 33421
rect 16619 33356 16620 33420
rect 16684 33356 16685 33420
rect 16619 33355 16685 33356
rect 17174 32877 17234 40019
rect 17358 33013 17418 52259
rect 17610 52256 17930 53280
rect 17610 52192 17618 52256
rect 17682 52192 17698 52256
rect 17762 52192 17778 52256
rect 17842 52192 17858 52256
rect 17922 52192 17930 52256
rect 17610 51168 17930 52192
rect 17610 51104 17618 51168
rect 17682 51104 17698 51168
rect 17762 51104 17778 51168
rect 17842 51104 17858 51168
rect 17922 51104 17930 51168
rect 17610 50080 17930 51104
rect 17610 50016 17618 50080
rect 17682 50016 17698 50080
rect 17762 50016 17778 50080
rect 17842 50016 17858 50080
rect 17922 50016 17930 50080
rect 17610 48992 17930 50016
rect 17610 48928 17618 48992
rect 17682 48928 17698 48992
rect 17762 48928 17778 48992
rect 17842 48928 17858 48992
rect 17922 48928 17930 48992
rect 17610 47904 17930 48928
rect 17610 47840 17618 47904
rect 17682 47840 17698 47904
rect 17762 47840 17778 47904
rect 17842 47840 17858 47904
rect 17922 47840 17930 47904
rect 17610 46816 17930 47840
rect 17610 46752 17618 46816
rect 17682 46752 17698 46816
rect 17762 46752 17778 46816
rect 17842 46752 17858 46816
rect 17922 46752 17930 46816
rect 17610 45728 17930 46752
rect 17610 45664 17618 45728
rect 17682 45664 17698 45728
rect 17762 45664 17778 45728
rect 17842 45664 17858 45728
rect 17922 45664 17930 45728
rect 17610 44640 17930 45664
rect 17610 44576 17618 44640
rect 17682 44576 17698 44640
rect 17762 44576 17778 44640
rect 17842 44576 17858 44640
rect 17922 44576 17930 44640
rect 17610 43552 17930 44576
rect 17610 43488 17618 43552
rect 17682 43488 17698 43552
rect 17762 43488 17778 43552
rect 17842 43488 17858 43552
rect 17922 43488 17930 43552
rect 17610 42464 17930 43488
rect 17610 42400 17618 42464
rect 17682 42400 17698 42464
rect 17762 42400 17778 42464
rect 17842 42400 17858 42464
rect 17922 42400 17930 42464
rect 17610 42246 17930 42400
rect 17610 42010 17652 42246
rect 17888 42010 17930 42246
rect 17610 41376 17930 42010
rect 17610 41312 17618 41376
rect 17682 41312 17698 41376
rect 17762 41312 17778 41376
rect 17842 41312 17858 41376
rect 17922 41312 17930 41376
rect 17610 40288 17930 41312
rect 17610 40224 17618 40288
rect 17682 40224 17698 40288
rect 17762 40224 17778 40288
rect 17842 40224 17858 40288
rect 17922 40224 17930 40288
rect 17610 39200 17930 40224
rect 17610 39136 17618 39200
rect 17682 39136 17698 39200
rect 17762 39136 17778 39200
rect 17842 39136 17858 39200
rect 17922 39136 17930 39200
rect 17610 38112 17930 39136
rect 17610 38048 17618 38112
rect 17682 38048 17698 38112
rect 17762 38048 17778 38112
rect 17842 38048 17858 38112
rect 17922 38048 17930 38112
rect 17610 37024 17930 38048
rect 17610 36960 17618 37024
rect 17682 36960 17698 37024
rect 17762 36960 17778 37024
rect 17842 36960 17858 37024
rect 17922 36960 17930 37024
rect 17610 35936 17930 36960
rect 17610 35872 17618 35936
rect 17682 35872 17698 35936
rect 17762 35872 17778 35936
rect 17842 35872 17858 35936
rect 17922 35872 17930 35936
rect 17610 34848 17930 35872
rect 17610 34784 17618 34848
rect 17682 34784 17698 34848
rect 17762 34784 17778 34848
rect 17842 34784 17858 34848
rect 17922 34784 17930 34848
rect 17610 33760 17930 34784
rect 17610 33696 17618 33760
rect 17682 33696 17698 33760
rect 17762 33696 17778 33760
rect 17842 33696 17858 33760
rect 17922 33696 17930 33760
rect 17355 33012 17421 33013
rect 17355 32948 17356 33012
rect 17420 32948 17421 33012
rect 17355 32947 17421 32948
rect 17171 32876 17237 32877
rect 17171 32812 17172 32876
rect 17236 32812 17237 32876
rect 17171 32811 17237 32812
rect 17610 32672 17930 33696
rect 17610 32608 17618 32672
rect 17682 32608 17698 32672
rect 17762 32608 17778 32672
rect 17842 32608 17858 32672
rect 17922 32608 17930 32672
rect 14963 32332 15029 32333
rect 14963 32268 14964 32332
rect 15028 32268 15029 32332
rect 14963 32267 15029 32268
rect 14277 32064 14285 32128
rect 14349 32064 14365 32128
rect 14429 32064 14445 32128
rect 14509 32064 14525 32128
rect 14589 32064 14597 32128
rect 14277 31040 14597 32064
rect 14277 30976 14285 31040
rect 14349 30976 14365 31040
rect 14429 30976 14445 31040
rect 14509 30976 14525 31040
rect 14589 30976 14597 31040
rect 14043 30700 14109 30701
rect 14043 30636 14044 30700
rect 14108 30636 14109 30700
rect 14043 30635 14109 30636
rect 14277 29952 14597 30976
rect 14277 29888 14285 29952
rect 14349 29888 14365 29952
rect 14429 29888 14445 29952
rect 14509 29888 14525 29952
rect 14589 29888 14597 29952
rect 12019 29748 12085 29749
rect 12019 29684 12020 29748
rect 12084 29684 12085 29748
rect 12019 29683 12085 29684
rect 10944 29344 10952 29408
rect 11016 29344 11032 29408
rect 11096 29344 11112 29408
rect 11176 29344 11192 29408
rect 11256 29344 11264 29408
rect 10944 28320 11264 29344
rect 11467 28932 11533 28933
rect 11467 28868 11468 28932
rect 11532 28868 11533 28932
rect 11467 28867 11533 28868
rect 14277 28912 14597 29888
rect 10944 28256 10952 28320
rect 11016 28256 11032 28320
rect 11096 28256 11112 28320
rect 11176 28256 11192 28320
rect 11256 28256 11264 28320
rect 10944 27232 11264 28256
rect 10944 27168 10952 27232
rect 11016 27168 11032 27232
rect 11096 27168 11112 27232
rect 11176 27168 11192 27232
rect 11256 27168 11264 27232
rect 10944 26144 11264 27168
rect 10944 26080 10952 26144
rect 11016 26080 11032 26144
rect 11096 26080 11112 26144
rect 11176 26080 11192 26144
rect 11256 26080 11264 26144
rect 10944 25056 11264 26080
rect 10944 24992 10952 25056
rect 11016 24992 11032 25056
rect 11096 24992 11112 25056
rect 11176 24992 11192 25056
rect 11256 24992 11264 25056
rect 10547 24308 10613 24309
rect 10547 24244 10548 24308
rect 10612 24244 10613 24308
rect 10547 24243 10613 24244
rect 7610 23360 7618 23424
rect 7682 23360 7698 23424
rect 7762 23360 7778 23424
rect 7842 23360 7858 23424
rect 7922 23360 7930 23424
rect 7610 22336 7930 23360
rect 7610 22272 7618 22336
rect 7682 22272 7698 22336
rect 7762 22272 7778 22336
rect 7842 22272 7858 22336
rect 7922 22272 7930 22336
rect 7610 21248 7930 22272
rect 7610 21184 7618 21248
rect 7682 21184 7698 21248
rect 7762 21184 7778 21248
rect 7842 21184 7858 21248
rect 7922 21184 7930 21248
rect 7610 20160 7930 21184
rect 7610 20096 7618 20160
rect 7682 20096 7698 20160
rect 7762 20096 7778 20160
rect 7842 20096 7858 20160
rect 7922 20096 7930 20160
rect 7610 19072 7930 20096
rect 7610 19008 7618 19072
rect 7682 19008 7698 19072
rect 7762 19008 7778 19072
rect 7842 19008 7858 19072
rect 7922 19008 7930 19072
rect 7610 17984 7930 19008
rect 7610 17920 7618 17984
rect 7682 17920 7698 17984
rect 7762 17920 7778 17984
rect 7842 17920 7858 17984
rect 7922 17920 7930 17984
rect 7610 16896 7930 17920
rect 7610 16832 7618 16896
rect 7682 16832 7698 16896
rect 7762 16832 7778 16896
rect 7842 16832 7858 16896
rect 7922 16832 7930 16896
rect 7610 15808 7930 16832
rect 7610 15744 7618 15808
rect 7682 15744 7698 15808
rect 7762 15744 7778 15808
rect 7842 15744 7858 15808
rect 7922 15744 7930 15808
rect 7610 14720 7930 15744
rect 7610 14656 7618 14720
rect 7682 14656 7698 14720
rect 7762 14656 7778 14720
rect 7842 14656 7858 14720
rect 7922 14656 7930 14720
rect 7610 13632 7930 14656
rect 7610 13568 7618 13632
rect 7682 13568 7698 13632
rect 7762 13568 7778 13632
rect 7842 13568 7858 13632
rect 7922 13568 7930 13632
rect 7610 12544 7930 13568
rect 7610 12480 7618 12544
rect 7682 12480 7698 12544
rect 7762 12480 7778 12544
rect 7842 12480 7858 12544
rect 7922 12480 7930 12544
rect 7610 11456 7930 12480
rect 7610 11392 7618 11456
rect 7682 11392 7698 11456
rect 7762 11392 7778 11456
rect 7842 11392 7858 11456
rect 7922 11392 7930 11456
rect 7610 10368 7930 11392
rect 7610 10304 7618 10368
rect 7682 10304 7698 10368
rect 7762 10304 7778 10368
rect 7842 10304 7858 10368
rect 7922 10304 7930 10368
rect 7610 9280 7930 10304
rect 7610 9216 7618 9280
rect 7682 9216 7698 9280
rect 7762 9216 7778 9280
rect 7842 9216 7858 9280
rect 7922 9216 7930 9280
rect 7610 8192 7930 9216
rect 7610 8128 7618 8192
rect 7682 8128 7698 8192
rect 7762 8128 7778 8192
rect 7842 8128 7858 8192
rect 7922 8128 7930 8192
rect 7610 7104 7930 8128
rect 7610 7040 7618 7104
rect 7682 7040 7698 7104
rect 7762 7040 7778 7104
rect 7842 7040 7858 7104
rect 7922 7040 7930 7104
rect 7610 6016 7930 7040
rect 7610 5952 7618 6016
rect 7682 5952 7698 6016
rect 7762 5952 7778 6016
rect 7842 5952 7858 6016
rect 7922 5952 7930 6016
rect 7610 4928 7930 5952
rect 7610 4864 7618 4928
rect 7682 4864 7698 4928
rect 7762 4864 7778 4928
rect 7842 4864 7858 4928
rect 7922 4864 7930 4928
rect 7610 3840 7930 4864
rect 7610 3776 7618 3840
rect 7682 3776 7698 3840
rect 7762 3776 7778 3840
rect 7842 3776 7858 3840
rect 7922 3776 7930 3840
rect 7610 2752 7930 3776
rect 7610 2688 7618 2752
rect 7682 2688 7698 2752
rect 7762 2688 7778 2752
rect 7842 2688 7858 2752
rect 7922 2688 7930 2752
rect 7610 2128 7930 2688
rect 10944 23968 11264 24992
rect 10944 23904 10952 23968
rect 11016 23904 11032 23968
rect 11096 23904 11112 23968
rect 11176 23904 11192 23968
rect 11256 23904 11264 23968
rect 10944 22880 11264 23904
rect 10944 22816 10952 22880
rect 11016 22816 11032 22880
rect 11096 22816 11112 22880
rect 11176 22816 11192 22880
rect 11256 22816 11264 22880
rect 10944 21792 11264 22816
rect 11470 22677 11530 28867
rect 14277 28864 14319 28912
rect 14555 28864 14597 28912
rect 14277 28800 14285 28864
rect 14589 28800 14597 28864
rect 14277 28676 14319 28800
rect 14555 28676 14597 28800
rect 14277 27776 14597 28676
rect 14277 27712 14285 27776
rect 14349 27712 14365 27776
rect 14429 27712 14445 27776
rect 14509 27712 14525 27776
rect 14589 27712 14597 27776
rect 14277 26688 14597 27712
rect 14277 26624 14285 26688
rect 14349 26624 14365 26688
rect 14429 26624 14445 26688
rect 14509 26624 14525 26688
rect 14589 26624 14597 26688
rect 14277 25600 14597 26624
rect 14277 25536 14285 25600
rect 14349 25536 14365 25600
rect 14429 25536 14445 25600
rect 14509 25536 14525 25600
rect 14589 25536 14597 25600
rect 14277 24512 14597 25536
rect 14277 24448 14285 24512
rect 14349 24448 14365 24512
rect 14429 24448 14445 24512
rect 14509 24448 14525 24512
rect 14589 24448 14597 24512
rect 14277 23424 14597 24448
rect 14277 23360 14285 23424
rect 14349 23360 14365 23424
rect 14429 23360 14445 23424
rect 14509 23360 14525 23424
rect 14589 23360 14597 23424
rect 11467 22676 11533 22677
rect 11467 22612 11468 22676
rect 11532 22612 11533 22676
rect 11467 22611 11533 22612
rect 10944 21728 10952 21792
rect 11016 21728 11032 21792
rect 11096 21728 11112 21792
rect 11176 21728 11192 21792
rect 11256 21728 11264 21792
rect 10944 20704 11264 21728
rect 10944 20640 10952 20704
rect 11016 20640 11032 20704
rect 11096 20640 11112 20704
rect 11176 20640 11192 20704
rect 11256 20640 11264 20704
rect 10944 19616 11264 20640
rect 10944 19552 10952 19616
rect 11016 19552 11032 19616
rect 11096 19552 11112 19616
rect 11176 19552 11192 19616
rect 11256 19552 11264 19616
rect 10944 18528 11264 19552
rect 10944 18464 10952 18528
rect 11016 18464 11032 18528
rect 11096 18464 11112 18528
rect 11176 18464 11192 18528
rect 11256 18464 11264 18528
rect 10944 17440 11264 18464
rect 10944 17376 10952 17440
rect 11016 17376 11032 17440
rect 11096 17376 11112 17440
rect 11176 17376 11192 17440
rect 11256 17376 11264 17440
rect 10944 16352 11264 17376
rect 10944 16288 10952 16352
rect 11016 16288 11032 16352
rect 11096 16288 11112 16352
rect 11176 16288 11192 16352
rect 11256 16288 11264 16352
rect 10944 15579 11264 16288
rect 10944 15343 10986 15579
rect 11222 15343 11264 15579
rect 10944 15264 11264 15343
rect 10944 15200 10952 15264
rect 11016 15200 11032 15264
rect 11096 15200 11112 15264
rect 11176 15200 11192 15264
rect 11256 15200 11264 15264
rect 10944 14176 11264 15200
rect 10944 14112 10952 14176
rect 11016 14112 11032 14176
rect 11096 14112 11112 14176
rect 11176 14112 11192 14176
rect 11256 14112 11264 14176
rect 10944 13088 11264 14112
rect 10944 13024 10952 13088
rect 11016 13024 11032 13088
rect 11096 13024 11112 13088
rect 11176 13024 11192 13088
rect 11256 13024 11264 13088
rect 10944 12000 11264 13024
rect 10944 11936 10952 12000
rect 11016 11936 11032 12000
rect 11096 11936 11112 12000
rect 11176 11936 11192 12000
rect 11256 11936 11264 12000
rect 10944 10912 11264 11936
rect 10944 10848 10952 10912
rect 11016 10848 11032 10912
rect 11096 10848 11112 10912
rect 11176 10848 11192 10912
rect 11256 10848 11264 10912
rect 10944 9824 11264 10848
rect 10944 9760 10952 9824
rect 11016 9760 11032 9824
rect 11096 9760 11112 9824
rect 11176 9760 11192 9824
rect 11256 9760 11264 9824
rect 10944 8736 11264 9760
rect 10944 8672 10952 8736
rect 11016 8672 11032 8736
rect 11096 8672 11112 8736
rect 11176 8672 11192 8736
rect 11256 8672 11264 8736
rect 10944 7648 11264 8672
rect 10944 7584 10952 7648
rect 11016 7584 11032 7648
rect 11096 7584 11112 7648
rect 11176 7584 11192 7648
rect 11256 7584 11264 7648
rect 10944 6560 11264 7584
rect 10944 6496 10952 6560
rect 11016 6496 11032 6560
rect 11096 6496 11112 6560
rect 11176 6496 11192 6560
rect 11256 6496 11264 6560
rect 10944 5472 11264 6496
rect 10944 5408 10952 5472
rect 11016 5408 11032 5472
rect 11096 5408 11112 5472
rect 11176 5408 11192 5472
rect 11256 5408 11264 5472
rect 10944 4384 11264 5408
rect 10944 4320 10952 4384
rect 11016 4320 11032 4384
rect 11096 4320 11112 4384
rect 11176 4320 11192 4384
rect 11256 4320 11264 4384
rect 10944 3296 11264 4320
rect 10944 3232 10952 3296
rect 11016 3232 11032 3296
rect 11096 3232 11112 3296
rect 11176 3232 11192 3296
rect 11256 3232 11264 3296
rect 10944 2208 11264 3232
rect 10944 2144 10952 2208
rect 11016 2144 11032 2208
rect 11096 2144 11112 2208
rect 11176 2144 11192 2208
rect 11256 2144 11264 2208
rect 10944 2128 11264 2144
rect 14277 22336 14597 23360
rect 14277 22272 14285 22336
rect 14349 22272 14365 22336
rect 14429 22272 14445 22336
rect 14509 22272 14525 22336
rect 14589 22272 14597 22336
rect 14277 21248 14597 22272
rect 14277 21184 14285 21248
rect 14349 21184 14365 21248
rect 14429 21184 14445 21248
rect 14509 21184 14525 21248
rect 14589 21184 14597 21248
rect 14277 20160 14597 21184
rect 14277 20096 14285 20160
rect 14349 20096 14365 20160
rect 14429 20096 14445 20160
rect 14509 20096 14525 20160
rect 14589 20096 14597 20160
rect 14277 19072 14597 20096
rect 14277 19008 14285 19072
rect 14349 19008 14365 19072
rect 14429 19008 14445 19072
rect 14509 19008 14525 19072
rect 14589 19008 14597 19072
rect 14277 17984 14597 19008
rect 14277 17920 14285 17984
rect 14349 17920 14365 17984
rect 14429 17920 14445 17984
rect 14509 17920 14525 17984
rect 14589 17920 14597 17984
rect 14277 16896 14597 17920
rect 14277 16832 14285 16896
rect 14349 16832 14365 16896
rect 14429 16832 14445 16896
rect 14509 16832 14525 16896
rect 14589 16832 14597 16896
rect 14277 15808 14597 16832
rect 14277 15744 14285 15808
rect 14349 15744 14365 15808
rect 14429 15744 14445 15808
rect 14509 15744 14525 15808
rect 14589 15744 14597 15808
rect 14277 14720 14597 15744
rect 14277 14656 14285 14720
rect 14349 14656 14365 14720
rect 14429 14656 14445 14720
rect 14509 14656 14525 14720
rect 14589 14656 14597 14720
rect 14277 13632 14597 14656
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 12544 14597 13568
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 11456 14597 12480
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 10368 14597 11392
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 9280 14597 10304
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 8192 14597 9216
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 7104 14597 8128
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 6016 14597 7040
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 4928 14597 5952
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 3840 14597 4864
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 2752 14597 3776
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2128 14597 2688
rect 17610 31584 17930 32608
rect 17610 31520 17618 31584
rect 17682 31520 17698 31584
rect 17762 31520 17778 31584
rect 17842 31520 17858 31584
rect 17922 31520 17930 31584
rect 17610 30496 17930 31520
rect 17610 30432 17618 30496
rect 17682 30432 17698 30496
rect 17762 30432 17778 30496
rect 17842 30432 17858 30496
rect 17922 30432 17930 30496
rect 17610 29408 17930 30432
rect 17610 29344 17618 29408
rect 17682 29344 17698 29408
rect 17762 29344 17778 29408
rect 17842 29344 17858 29408
rect 17922 29344 17930 29408
rect 17610 28320 17930 29344
rect 17610 28256 17618 28320
rect 17682 28256 17698 28320
rect 17762 28256 17778 28320
rect 17842 28256 17858 28320
rect 17922 28256 17930 28320
rect 17610 27232 17930 28256
rect 17610 27168 17618 27232
rect 17682 27168 17698 27232
rect 17762 27168 17778 27232
rect 17842 27168 17858 27232
rect 17922 27168 17930 27232
rect 17610 26144 17930 27168
rect 17610 26080 17618 26144
rect 17682 26080 17698 26144
rect 17762 26080 17778 26144
rect 17842 26080 17858 26144
rect 17922 26080 17930 26144
rect 17610 25056 17930 26080
rect 17610 24992 17618 25056
rect 17682 24992 17698 25056
rect 17762 24992 17778 25056
rect 17842 24992 17858 25056
rect 17922 24992 17930 25056
rect 17610 23968 17930 24992
rect 17610 23904 17618 23968
rect 17682 23904 17698 23968
rect 17762 23904 17778 23968
rect 17842 23904 17858 23968
rect 17922 23904 17930 23968
rect 17610 22880 17930 23904
rect 17610 22816 17618 22880
rect 17682 22816 17698 22880
rect 17762 22816 17778 22880
rect 17842 22816 17858 22880
rect 17922 22816 17930 22880
rect 17610 21792 17930 22816
rect 17610 21728 17618 21792
rect 17682 21728 17698 21792
rect 17762 21728 17778 21792
rect 17842 21728 17858 21792
rect 17922 21728 17930 21792
rect 17610 20704 17930 21728
rect 17610 20640 17618 20704
rect 17682 20640 17698 20704
rect 17762 20640 17778 20704
rect 17842 20640 17858 20704
rect 17922 20640 17930 20704
rect 17610 19616 17930 20640
rect 17610 19552 17618 19616
rect 17682 19552 17698 19616
rect 17762 19552 17778 19616
rect 17842 19552 17858 19616
rect 17922 19552 17930 19616
rect 17610 18528 17930 19552
rect 17610 18464 17618 18528
rect 17682 18464 17698 18528
rect 17762 18464 17778 18528
rect 17842 18464 17858 18528
rect 17922 18464 17930 18528
rect 17610 17440 17930 18464
rect 17610 17376 17618 17440
rect 17682 17376 17698 17440
rect 17762 17376 17778 17440
rect 17842 17376 17858 17440
rect 17922 17376 17930 17440
rect 17610 16352 17930 17376
rect 17610 16288 17618 16352
rect 17682 16288 17698 16352
rect 17762 16288 17778 16352
rect 17842 16288 17858 16352
rect 17922 16288 17930 16352
rect 17610 15579 17930 16288
rect 17610 15343 17652 15579
rect 17888 15343 17930 15579
rect 17610 15264 17930 15343
rect 17610 15200 17618 15264
rect 17682 15200 17698 15264
rect 17762 15200 17778 15264
rect 17842 15200 17858 15264
rect 17922 15200 17930 15264
rect 17610 14176 17930 15200
rect 17610 14112 17618 14176
rect 17682 14112 17698 14176
rect 17762 14112 17778 14176
rect 17842 14112 17858 14176
rect 17922 14112 17930 14176
rect 17610 13088 17930 14112
rect 17610 13024 17618 13088
rect 17682 13024 17698 13088
rect 17762 13024 17778 13088
rect 17842 13024 17858 13088
rect 17922 13024 17930 13088
rect 17610 12000 17930 13024
rect 17610 11936 17618 12000
rect 17682 11936 17698 12000
rect 17762 11936 17778 12000
rect 17842 11936 17858 12000
rect 17922 11936 17930 12000
rect 17610 10912 17930 11936
rect 17610 10848 17618 10912
rect 17682 10848 17698 10912
rect 17762 10848 17778 10912
rect 17842 10848 17858 10912
rect 17922 10848 17930 10912
rect 17610 9824 17930 10848
rect 17610 9760 17618 9824
rect 17682 9760 17698 9824
rect 17762 9760 17778 9824
rect 17842 9760 17858 9824
rect 17922 9760 17930 9824
rect 17610 8736 17930 9760
rect 17610 8672 17618 8736
rect 17682 8672 17698 8736
rect 17762 8672 17778 8736
rect 17842 8672 17858 8736
rect 17922 8672 17930 8736
rect 17610 7648 17930 8672
rect 17610 7584 17618 7648
rect 17682 7584 17698 7648
rect 17762 7584 17778 7648
rect 17842 7584 17858 7648
rect 17922 7584 17930 7648
rect 17610 6560 17930 7584
rect 17610 6496 17618 6560
rect 17682 6496 17698 6560
rect 17762 6496 17778 6560
rect 17842 6496 17858 6560
rect 17922 6496 17930 6560
rect 17610 5472 17930 6496
rect 17610 5408 17618 5472
rect 17682 5408 17698 5472
rect 17762 5408 17778 5472
rect 17842 5408 17858 5472
rect 17922 5408 17930 5472
rect 17610 4384 17930 5408
rect 17610 4320 17618 4384
rect 17682 4320 17698 4384
rect 17762 4320 17778 4384
rect 17842 4320 17858 4384
rect 17922 4320 17930 4384
rect 17610 3296 17930 4320
rect 17610 3232 17618 3296
rect 17682 3232 17698 3296
rect 17762 3232 17778 3296
rect 17842 3232 17858 3296
rect 17922 3232 17930 3296
rect 17610 2208 17930 3232
rect 17610 2144 17618 2208
rect 17682 2144 17698 2208
rect 17762 2144 17778 2208
rect 17842 2144 17858 2208
rect 17922 2144 17930 2208
rect 17610 2128 17930 2144
<< via4 >>
rect 4319 68676 4555 68912
rect 4319 42010 4555 42246
rect 7652 55343 7888 55579
rect 7652 28864 7888 28912
rect 7652 28800 7682 28864
rect 7682 28800 7698 28864
rect 7698 28800 7762 28864
rect 7762 28800 7778 28864
rect 7778 28800 7842 28864
rect 7842 28800 7858 28864
rect 7858 28800 7888 28864
rect 7652 28676 7888 28800
rect 4319 15343 4555 15579
rect 10986 68676 11222 68912
rect 10986 42010 11222 42246
rect 14319 55343 14555 55579
rect 17652 68676 17888 68912
rect 17652 42010 17888 42246
rect 14319 28864 14555 28912
rect 14319 28800 14349 28864
rect 14349 28800 14365 28864
rect 14365 28800 14429 28864
rect 14429 28800 14445 28864
rect 14445 28800 14509 28864
rect 14509 28800 14525 28864
rect 14525 28800 14555 28864
rect 14319 28676 14555 28800
rect 10986 15343 11222 15579
rect 17652 15343 17888 15579
<< metal5 >>
rect 1104 68912 18860 68954
rect 1104 68676 4319 68912
rect 4555 68676 10986 68912
rect 11222 68676 17652 68912
rect 17888 68676 18860 68912
rect 1104 68634 18860 68676
rect 1104 55579 18860 55621
rect 1104 55343 7652 55579
rect 7888 55343 14319 55579
rect 14555 55343 18860 55579
rect 1104 55301 18860 55343
rect 1104 42246 18860 42288
rect 1104 42010 4319 42246
rect 4555 42010 10986 42246
rect 11222 42010 17652 42246
rect 17888 42010 18860 42246
rect 1104 41968 18860 42010
rect 1104 28912 18860 28955
rect 1104 28676 7652 28912
rect 7888 28676 14319 28912
rect 14555 28676 18860 28912
rect 1104 28634 18860 28676
rect 1104 15579 18860 15621
rect 1104 15343 4319 15579
rect 4555 15343 10986 15579
rect 11222 15343 17652 15579
rect 17888 15343 18860 15579
rect 1104 15301 18860 15343
use sky130_fd_sc_hd__decap_3  PHY_0 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 1104 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606120353
transform 1 0 1104 0 1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 1380 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606120353
transform 1 0 2484 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606120353
transform 1 0 1380 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1606120353
transform 1 0 2484 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 3956 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1606120353
transform 1 0 3956 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 3588 0 -1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1606120353
transform 1 0 4048 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1606120353
transform 1 0 5152 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1606120353
transform 1 0 3588 0 1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_1_32
timestamp 1606120353
transform 1 0 4048 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1606120353
transform 1 0 5152 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1606120353
transform 1 0 6808 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 6256 0 -1 2720
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1606120353
transform 1 0 6900 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_56
timestamp 1606120353
transform 1 0 6256 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__CLK /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 9108 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1606120353
transform 1 0 8004 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_68
timestamp 1606120353
transform 1 0 7360 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_80
timestamp 1606120353
transform 1 0 8464 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1228_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 9752 0 -1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1606120353
transform 1 0 9660 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1606120353
transform 1 0 9568 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__D
timestamp 1606120353
transform 1 0 9476 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 9292 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1606120353
transform 1 0 9660 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_105
timestamp 1606120353
transform 1 0 10764 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1606120353
transform 1 0 12512 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 11500 0 -1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_0_121
timestamp 1606120353
transform 1 0 12236 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1606120353
transform 1 0 12604 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_117
timestamp 1606120353
transform 1 0 11868 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_129
timestamp 1606120353
transform 1 0 12972 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1606120353
transform 1 0 15180 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1606120353
transform 1 0 13708 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1606120353
transform 1 0 14812 0 -1 2720
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_1_141
timestamp 1606120353
transform 1 0 14076 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_154
timestamp 1606120353
transform 1 0 15272 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1606120353
transform 1 0 15364 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1606120353
transform 1 0 15456 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1606120353
transform 1 0 16560 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_166
timestamp 1606120353
transform 1 0 16376 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606120353
transform -1 0 18860 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606120353
transform -1 0 18860 0 1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1606120353
transform 1 0 18216 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1606120353
transform 1 0 17664 0 -1 2720
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1606120353
transform 1 0 18308 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_1_178
timestamp 1606120353
transform 1 0 17480 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606120353
transform 1 0 1104 0 -1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__D
timestamp 1606120353
transform 1 0 1564 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1606120353
transform 1 0 1380 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_2_7
timestamp 1606120353
transform 1 0 1748 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_19
timestamp 1606120353
transform 1 0 2852 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_31
timestamp 1606120353
transform 1 0 3956 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_43
timestamp 1606120353
transform 1 0 5060 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1606120353
transform 1 0 6716 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_2_55
timestamp 1606120353
transform 1 0 6164 0 -1 3808
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_2_62
timestamp 1606120353
transform 1 0 6808 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_74
timestamp 1606120353
transform 1 0 7912 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_86
timestamp 1606120353
transform 1 0 9016 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__CLK
timestamp 1606120353
transform 1 0 10212 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_2_98 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 10120 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_2_101
timestamp 1606120353
transform 1 0 10396 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1606120353
transform 1 0 12328 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_2_113
timestamp 1606120353
transform 1 0 11500 0 -1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_2_121
timestamp 1606120353
transform 1 0 12236 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1606120353
transform 1 0 12420 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_135
timestamp 1606120353
transform 1 0 13524 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_147
timestamp 1606120353
transform 1 0 14628 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_159
timestamp 1606120353
transform 1 0 15732 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_171
timestamp 1606120353
transform 1 0 16836 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606120353
transform -1 0 18860 0 -1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1606120353
transform 1 0 17940 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_2_184
timestamp 1606120353
transform 1 0 18032 0 -1 3808
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1232_
timestamp 1606120353
transform 1 0 1380 0 1 3808
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606120353
transform 1 0 1104 0 1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_3_22
timestamp 1606120353
transform 1 0 3128 0 1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1606120353
transform 1 0 3956 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_3_30
timestamp 1606120353
transform 1 0 3864 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1606120353
transform 1 0 4048 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1606120353
transform 1 0 5152 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_56
timestamp 1606120353
transform 1 0 6256 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_68
timestamp 1606120353
transform 1 0 7360 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_80
timestamp 1606120353
transform 1 0 8464 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1229_
timestamp 1606120353
transform 1 0 10212 0 1 3808
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1606120353
transform 1 0 9568 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__D
timestamp 1606120353
transform 1 0 10028 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_3_93
timestamp 1606120353
transform 1 0 9660 0 1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_3_118
timestamp 1606120353
transform 1 0 11960 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_130
timestamp 1606120353
transform 1 0 13064 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1606120353
transform 1 0 15180 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A
timestamp 1606120353
transform 1 0 14168 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__B
timestamp 1606120353
transform 1 0 14536 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_144
timestamp 1606120353
transform 1 0 14352 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_3_148
timestamp 1606120353
transform 1 0 14720 0 1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_3_152
timestamp 1606120353
transform 1 0 15088 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_3_154
timestamp 1606120353
transform 1 0 15272 0 1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__A
timestamp 1606120353
transform 1 0 15732 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_3_158
timestamp 1606120353
transform 1 0 15640 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_3_161
timestamp 1606120353
transform 1 0 15916 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_173
timestamp 1606120353
transform 1 0 17020 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606120353
transform -1 0 18860 0 1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_3_185
timestamp 1606120353
transform 1 0 18124 0 1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1606120353
transform 1 0 18492 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606120353
transform 1 0 1104 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__CLK
timestamp 1606120353
transform 1 0 1564 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1606120353
transform 1 0 1380 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_4_7
timestamp 1606120353
transform 1 0 1748 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_19
timestamp 1606120353
transform 1 0 2852 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_31
timestamp 1606120353
transform 1 0 3956 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_43
timestamp 1606120353
transform 1 0 5060 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1606120353
transform 1 0 6716 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_4_55
timestamp 1606120353
transform 1 0 6164 0 -1 4896
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_4_62
timestamp 1606120353
transform 1 0 6808 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_74
timestamp 1606120353
transform 1 0 7912 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_86
timestamp 1606120353
transform 1 0 9016 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_98
timestamp 1606120353
transform 1 0 10120 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_110
timestamp 1606120353
transform 1 0 11224 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1606120353
transform 1 0 12328 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1606120353
transform 1 0 12420 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__nand2_4  _0982_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 14168 0 -1 4896
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__B1
timestamp 1606120353
transform 1 0 15272 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__B
timestamp 1606120353
transform 1 0 13616 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A
timestamp 1606120353
transform 1 0 13984 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_4_135
timestamp 1606120353
transform 1 0 13524 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1606120353
transform 1 0 13800 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_4_151
timestamp 1606120353
transform 1 0 14996 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _0953_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 15732 0 -1 4896
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A1
timestamp 1606120353
transform 1 0 16744 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_4_156
timestamp 1606120353
transform 1 0 15456 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_4_168
timestamp 1606120353
transform 1 0 16560 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_4_172
timestamp 1606120353
transform 1 0 16928 0 -1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606120353
transform -1 0 18860 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1606120353
transform 1 0 17940 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_4_180
timestamp 1606120353
transform 1 0 17664 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_4_184
timestamp 1606120353
transform 1 0 18032 0 -1 4896
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606120353
transform 1 0 1104 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__D
timestamp 1606120353
transform 1 0 2116 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__CLK
timestamp 1606120353
transform 1 0 2484 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3
timestamp 1606120353
transform 1 0 1380 0 1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_5_13
timestamp 1606120353
transform 1 0 2300 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_5_17
timestamp 1606120353
transform 1 0 2668 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1606120353
transform 1 0 3956 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_5_29
timestamp 1606120353
transform 1 0 3772 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_5_32
timestamp 1606120353
transform 1 0 4048 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_44
timestamp 1606120353
transform 1 0 5152 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_5_56
timestamp 1606120353
transform 1 0 6256 0 1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_5_64
timestamp 1606120353
transform 1 0 6992 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__D
timestamp 1606120353
transform 1 0 7268 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__CLK
timestamp 1606120353
transform 1 0 7636 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_69
timestamp 1606120353
transform 1 0 7452 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_5_73
timestamp 1606120353
transform 1 0 7820 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_5_85
timestamp 1606120353
transform 1 0 8924 0 1 4896
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1606120353
transform 1 0 9568 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__D
timestamp 1606120353
transform 1 0 9844 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__CLK
timestamp 1606120353
transform 1 0 10212 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_5_91
timestamp 1606120353
transform 1 0 9476 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_5_93
timestamp 1606120353
transform 1 0 9660 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_97
timestamp 1606120353
transform 1 0 10028 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_5_101
timestamp 1606120353
transform 1 0 10396 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A
timestamp 1606120353
transform 1 0 12420 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A1
timestamp 1606120353
transform 1 0 13064 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp 1606120353
transform 1 0 11500 0 1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_5_121
timestamp 1606120353
transform 1 0 12236 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_5_125
timestamp 1606120353
transform 1 0 12604 0 1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_5_129
timestamp 1606120353
transform 1 0 12972 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_5_132
timestamp 1606120353
transform 1 0 13248 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0948_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 15272 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__nand2_4  _0969_
timestamp 1606120353
transform 1 0 13616 0 1 4896
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1606120353
transform 1 0 15180 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A2
timestamp 1606120353
transform 1 0 14996 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__A
timestamp 1606120353
transform 1 0 13432 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A1
timestamp 1606120353
transform 1 0 14628 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_145
timestamp 1606120353
transform 1 0 14444 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_149
timestamp 1606120353
transform 1 0 14812 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A2
timestamp 1606120353
transform 1 0 16560 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__B1
timestamp 1606120353
transform 1 0 16928 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1606120353
transform 1 0 16376 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_170
timestamp 1606120353
transform 1 0 16744 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_5_174
timestamp 1606120353
transform 1 0 17112 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606120353
transform -1 0 18860 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_5_186
timestamp 1606120353
transform 1 0 18216 0 1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1233_
timestamp 1606120353
transform 1 0 2116 0 -1 5984
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606120353
transform 1 0 1104 0 -1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606120353
transform 1 0 1104 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1606120353
transform 1 0 1380 0 -1 5984
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606120353
transform 1 0 1380 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1606120353
transform 1 0 2484 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1606120353
transform 1 0 3956 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1606120353
transform 1 0 3864 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_42
timestamp 1606120353
transform 1 0 4968 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1606120353
transform 1 0 3588 0 1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_7_32
timestamp 1606120353
transform 1 0 4048 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_44
timestamp 1606120353
transform 1 0 5152 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1606120353
transform 1 0 6716 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_6_54
timestamp 1606120353
transform 1 0 6072 0 -1 5984
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_6_60
timestamp 1606120353
transform 1 0 6624 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_6_62
timestamp 1606120353
transform 1 0 6808 0 -1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_6_66
timestamp 1606120353
transform 1 0 7176 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_7_56
timestamp 1606120353
transform 1 0 6256 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1230_
timestamp 1606120353
transform 1 0 7268 0 -1 5984
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_8  FILLER_6_86
timestamp 1606120353
transform 1 0 9016 0 -1 5984
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_7_68
timestamp 1606120353
transform 1 0 7360 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_80
timestamp 1606120353
transform 1 0 8464 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_7_97
timestamp 1606120353
transform 1 0 10028 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_7_93
timestamp 1606120353
transform 1 0 9660 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__CLK
timestamp 1606120353
transform 1 0 10212 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__D
timestamp 1606120353
transform 1 0 9844 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1606120353
transform 1 0 9568 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_7_108
timestamp 1606120353
transform 1 0 11040 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_7_105
timestamp 1606120353
transform 1 0 10764 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_7_101
timestamp 1606120353
transform 1 0 10396 0 1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__B1_N
timestamp 1606120353
transform 1 0 10856 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A2
timestamp 1606120353
transform 1 0 11224 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1231_
timestamp 1606120353
transform 1 0 9752 0 -1 5984
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  FILLER_6_117
timestamp 1606120353
transform 1 0 11868 0 -1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_6_113
timestamp 1606120353
transform 1 0 11500 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__B1
timestamp 1606120353
transform 1 0 12144 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A1
timestamp 1606120353
transform 1 0 11684 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_7_129
timestamp 1606120353
transform 1 0 12972 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_7_125
timestamp 1606120353
transform 1 0 12604 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_6_132
timestamp 1606120353
transform 1 0 13248 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A2
timestamp 1606120353
transform 1 0 12788 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A1_N
timestamp 1606120353
transform 1 0 13156 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1606120353
transform 1 0 12328 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _0899_
timestamp 1606120353
transform 1 0 12420 0 -1 5984
box 0 -48 828 592
use sky130_fd_sc_hd__a21bo_4  _0980_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 11408 0 1 5984
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_6_140
timestamp 1606120353
transform 1 0 13984 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_6_136
timestamp 1606120353
transform 1 0 13616 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__B1
timestamp 1606120353
transform 1 0 14168 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__B2
timestamp 1606120353
transform 1 0 13800 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A2_N
timestamp 1606120353
transform 1 0 13432 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_7_154
timestamp 1606120353
transform 1 0 15272 0 1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_7_149
timestamp 1606120353
transform 1 0 14812 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_7_145
timestamp 1606120353
transform 1 0 14444 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_6_144
timestamp 1606120353
transform 1 0 14352 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__B1
timestamp 1606120353
transform 1 0 14996 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__B2
timestamp 1606120353
transform 1 0 14628 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1606120353
transform 1 0 15180 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _0949_
timestamp 1606120353
transform 1 0 14536 0 -1 5984
box 0 -48 828 592
use sky130_fd_sc_hd__a21o_4  _0970_
timestamp 1606120353
transform 1 0 13340 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp 1606120353
transform 1 0 16284 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_7_161
timestamp 1606120353
transform 1 0 15916 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_7_158
timestamp 1606120353
transform 1 0 15640 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_6_155
timestamp 1606120353
transform 1 0 15364 0 -1 5984
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A1
timestamp 1606120353
transform 1 0 15916 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__B1
timestamp 1606120353
transform 1 0 15732 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A2
timestamp 1606120353
transform 1 0 16100 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_6_175
timestamp 1606120353
transform 1 0 17204 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A2
timestamp 1606120353
transform 1 0 16560 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0955_
timestamp 1606120353
transform 1 0 16744 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__a21o_4  _0952_
timestamp 1606120353
transform 1 0 16100 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606120353
transform -1 0 18860 0 -1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606120353
transform -1 0 18860 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1606120353
transform 1 0 17940 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__B1
timestamp 1606120353
transform 1 0 17388 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_6_179
timestamp 1606120353
transform 1 0 17572 0 -1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_6_184
timestamp 1606120353
transform 1 0 18032 0 -1 5984
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_7_182
timestamp 1606120353
transform 1 0 17848 0 1 5984
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606120353
transform 1 0 1104 0 -1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1606120353
transform 1 0 1380 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1606120353
transform 1 0 2484 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_27
timestamp 1606120353
transform 1 0 3588 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_8_39
timestamp 1606120353
transform 1 0 4692 0 -1 7072
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1606120353
transform 1 0 6716 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__CLK
timestamp 1606120353
transform 1 0 5612 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_47
timestamp 1606120353
transform 1 0 5428 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_8_51
timestamp 1606120353
transform 1 0 5796 0 -1 7072
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_8_59
timestamp 1606120353
transform 1 0 6532 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_8_62
timestamp 1606120353
transform 1 0 6808 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_74
timestamp 1606120353
transform 1 0 7912 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_8_86
timestamp 1606120353
transform 1 0 9016 0 -1 7072
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1237_
timestamp 1606120353
transform 1 0 9844 0 -1 7072
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_1  FILLER_8_94
timestamp 1606120353
transform 1 0 9752 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__a2bb2oi_4  _0968_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 13156 0 -1 7072
box 0 -48 1932 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1606120353
transform 1 0 12328 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A2
timestamp 1606120353
transform 1 0 12972 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__B1
timestamp 1606120353
transform 1 0 12604 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A2
timestamp 1606120353
transform 1 0 12144 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_8_114
timestamp 1606120353
transform 1 0 11592 0 -1 7072
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_8_123
timestamp 1606120353
transform 1 0 12420 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_127
timestamp 1606120353
transform 1 0 12788 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_8_152
timestamp 1606120353
transform 1 0 15088 0 -1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__a21o_4  _0940_
timestamp 1606120353
transform 1 0 16100 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A1
timestamp 1606120353
transform 1 0 15364 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__B1
timestamp 1606120353
transform 1 0 15732 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_157
timestamp 1606120353
transform 1 0 15548 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_161
timestamp 1606120353
transform 1 0 15916 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_175
timestamp 1606120353
transform 1 0 17204 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606120353
transform -1 0 18860 0 -1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1606120353
transform 1 0 17940 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A1
timestamp 1606120353
transform 1 0 17388 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_8_179
timestamp 1606120353
transform 1 0 17572 0 -1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_8_184
timestamp 1606120353
transform 1 0 18032 0 -1 7072
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606120353
transform 1 0 1104 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606120353
transform 1 0 1380 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1606120353
transform 1 0 2484 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1606120353
transform 1 0 3956 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1606120353
transform 1 0 3588 0 1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_9_32
timestamp 1606120353
transform 1 0 4048 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_9_44
timestamp 1606120353
transform 1 0 5152 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1234_
timestamp 1606120353
transform 1 0 5612 0 1 7072
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__D
timestamp 1606120353
transform 1 0 5428 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__D
timestamp 1606120353
transform 1 0 8740 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__CLK
timestamp 1606120353
transform 1 0 9108 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_9_68
timestamp 1606120353
transform 1 0 7360 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_9_80
timestamp 1606120353
transform 1 0 8464 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_9_85
timestamp 1606120353
transform 1 0 8924 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0965_
timestamp 1606120353
transform 1 0 11040 0 1 7072
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1606120353
transform 1 0 9568 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A2
timestamp 1606120353
transform 1 0 10856 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A1
timestamp 1606120353
transform 1 0 10488 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_9_89
timestamp 1606120353
transform 1 0 9292 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_9_93
timestamp 1606120353
transform 1 0 9660 0 1 7072
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_9_101
timestamp 1606120353
transform 1 0 10396 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_9_104
timestamp 1606120353
transform 1 0 10672 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0913_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 12972 0 1 7072
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A1
timestamp 1606120353
transform 1 0 12420 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A1
timestamp 1606120353
transform 1 0 12788 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_121
timestamp 1606120353
transform 1 0 12236 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_125
timestamp 1606120353
transform 1 0 12604 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1606120353
transform 1 0 15180 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A2
timestamp 1606120353
transform 1 0 14996 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A1_N
timestamp 1606120353
transform 1 0 14352 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_142
timestamp 1606120353
transform 1 0 14168 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_9_146
timestamp 1606120353
transform 1 0 14536 0 1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_9_150
timestamp 1606120353
transform 1 0 14904 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_9_154
timestamp 1606120353
transform 1 0 15272 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__o21ai_4  _0951_
timestamp 1606120353
transform 1 0 15364 0 1 7072
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILLER_9_168
timestamp 1606120353
transform 1 0 16560 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606120353
transform -1 0 18860 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_9_180
timestamp 1606120353
transform 1 0 17664 0 1 7072
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1606120353
transform 1 0 18400 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606120353
transform 1 0 1104 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1606120353
transform 1 0 1380 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1606120353
transform 1 0 2484 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_27
timestamp 1606120353
transform 1 0 3588 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_39
timestamp 1606120353
transform 1 0 4692 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1606120353
transform 1 0 6716 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_10_51
timestamp 1606120353
transform 1 0 5796 0 -1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp 1606120353
transform 1 0 6532 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_10_62
timestamp 1606120353
transform 1 0 6808 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1236_
timestamp 1606120353
transform 1 0 8740 0 -1 8160
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_8  FILLER_10_74
timestamp 1606120353
transform 1 0 7912 0 -1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_10_82
timestamp 1606120353
transform 1 0 8648 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__B1_N
timestamp 1606120353
transform 1 0 11040 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_10_102
timestamp 1606120353
transform 1 0 10488 0 -1 8160
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_10_110
timestamp 1606120353
transform 1 0 11224 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0950_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 12420 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1606120353
transform 1 0 12328 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__C
timestamp 1606120353
transform 1 0 11408 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_10_114
timestamp 1606120353
transform 1 0 11592 0 -1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__a2bb2oi_4  _0981_
timestamp 1606120353
transform 1 0 14260 0 -1 8160
box 0 -48 1932 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__B1
timestamp 1606120353
transform 1 0 13708 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A2_N
timestamp 1606120353
transform 1 0 14076 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_10_135
timestamp 1606120353
transform 1 0 13524 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_10_139
timestamp 1606120353
transform 1 0 13892 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A
timestamp 1606120353
transform 1 0 16376 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_10_164
timestamp 1606120353
transform 1 0 16192 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_10_168
timestamp 1606120353
transform 1 0 16560 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606120353
transform -1 0 18860 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1606120353
transform 1 0 17940 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_10_180
timestamp 1606120353
transform 1 0 17664 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_10_184
timestamp 1606120353
transform 1 0 18032 0 -1 8160
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606120353
transform 1 0 1104 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1606120353
transform 1 0 1380 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1606120353
transform 1 0 2484 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1606120353
transform 1 0 3956 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1606120353
transform 1 0 3588 0 1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_11_32
timestamp 1606120353
transform 1 0 4048 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_44
timestamp 1606120353
transform 1 0 5152 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_56
timestamp 1606120353
transform 1 0 6256 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A
timestamp 1606120353
transform 1 0 9016 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__CLK
timestamp 1606120353
transform 1 0 8648 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_11_68
timestamp 1606120353
transform 1 0 7360 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_11_80
timestamp 1606120353
transform 1 0 8464 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_84
timestamp 1606120353
transform 1 0 8832 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_88
timestamp 1606120353
transform 1 0 9200 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0945_
timestamp 1606120353
transform 1 0 9844 0 1 8160
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1606120353
transform 1 0 9568 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__D
timestamp 1606120353
transform 1 0 9384 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A
timestamp 1606120353
transform 1 0 11224 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__D
timestamp 1606120353
transform 1 0 10856 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_93
timestamp 1606120353
transform 1 0 9660 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_104
timestamp 1606120353
transform 1 0 10672 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_108
timestamp 1606120353
transform 1 0 11040 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _0978_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 11408 0 1 8160
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__B1
timestamp 1606120353
transform 1 0 13156 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_129
timestamp 1606120353
transform 1 0 12972 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_11_141
timestamp 1606120353
transform 1 0 14076 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_11_137
timestamp 1606120353
transform 1 0 13708 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_133
timestamp 1606120353
transform 1 0 13340 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A2
timestamp 1606120353
transform 1 0 13892 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A1
timestamp 1606120353
transform 1 0 13524 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_11_150
timestamp 1606120353
transform 1 0 14904 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_11_146
timestamp 1606120353
transform 1 0 14536 0 1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__A2
timestamp 1606120353
transform 1 0 14352 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A2
timestamp 1606120353
transform 1 0 14996 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1606120353
transform 1 0 15180 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__a21o_4  _0983_
timestamp 1606120353
transform 1 0 15272 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__A1
timestamp 1606120353
transform 1 0 16560 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A1
timestamp 1606120353
transform 1 0 16928 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1606120353
transform 1 0 16376 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_170
timestamp 1606120353
transform 1 0 16744 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_11_174
timestamp 1606120353
transform 1 0 17112 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606120353
transform -1 0 18860 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_11_186
timestamp 1606120353
transform 1 0 18216 0 1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606120353
transform 1 0 1104 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__CLK
timestamp 1606120353
transform 1 0 1564 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__CLK
timestamp 1606120353
transform 1 0 1932 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1606120353
transform 1 0 1380 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_7
timestamp 1606120353
transform 1 0 1748 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_12_11
timestamp 1606120353
transform 1 0 2116 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_23
timestamp 1606120353
transform 1 0 3220 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_35
timestamp 1606120353
transform 1 0 4324 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1606120353
transform 1 0 6716 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_12_47
timestamp 1606120353
transform 1 0 5428 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_12_59
timestamp 1606120353
transform 1 0 6532 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_12_62
timestamp 1606120353
transform 1 0 6808 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_74
timestamp 1606120353
transform 1 0 7912 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_12_86
timestamp 1606120353
transform 1 0 9016 0 -1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1238_
timestamp 1606120353
transform 1 0 9476 0 -1 9248
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_1  FILLER_12_90
timestamp 1606120353
transform 1 0 9384 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_12_110
timestamp 1606120353
transform 1 0 11224 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0946_
timestamp 1606120353
transform 1 0 12420 0 -1 9248
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1606120353
transform 1 0 12328 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__B
timestamp 1606120353
transform 1 0 11408 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__D
timestamp 1606120353
transform 1 0 11776 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_114
timestamp 1606120353
transform 1 0 11592 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_12_118
timestamp 1606120353
transform 1 0 11960 0 -1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__a21o_4  _0973_
timestamp 1606120353
transform 1 0 14352 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__B
timestamp 1606120353
transform 1 0 13800 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__C
timestamp 1606120353
transform 1 0 14168 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_136
timestamp 1606120353
transform 1 0 13616 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_140
timestamp 1606120353
transform 1 0 13984 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0917_
timestamp 1606120353
transform 1 0 16192 0 -1 9248
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__B1
timestamp 1606120353
transform 1 0 15640 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__B1
timestamp 1606120353
transform 1 0 16008 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_156
timestamp 1606120353
transform 1 0 15456 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_160
timestamp 1606120353
transform 1 0 15824 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_12_173
timestamp 1606120353
transform 1 0 17020 0 -1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606120353
transform -1 0 18860 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1606120353
transform 1 0 17940 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_12_181
timestamp 1606120353
transform 1 0 17756 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_12_184
timestamp 1606120353
transform 1 0 18032 0 -1 9248
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1606120353
transform 1 0 1380 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_13_11
timestamp 1606120353
transform 1 0 2116 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1606120353
transform 1 0 1748 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1606120353
transform 1 0 1380 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__D
timestamp 1606120353
transform 1 0 1932 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__D
timestamp 1606120353
transform 1 0 1564 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606120353
transform 1 0 1104 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606120353
transform 1 0 1104 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__D
timestamp 1606120353
transform 1 0 2300 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1606120353
transform 1 0 2484 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1246_
timestamp 1606120353
transform 1 0 1472 0 -1 10336
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_2  FILLER_14_33
timestamp 1606120353
transform 1 0 4140 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_14_23
timestamp 1606120353
transform 1 0 3220 0 -1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1606120353
transform 1 0 3588 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__CLK
timestamp 1606120353
transform 1 0 3956 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1606120353
transform 1 0 3956 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_14_37
timestamp 1606120353
transform 1 0 4508 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__CLK
timestamp 1606120353
transform 1 0 4692 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__D
timestamp 1606120353
transform 1 0 4324 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1606120353
transform 1 0 4876 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_13_44
timestamp 1606120353
transform 1 0 5152 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_13_32
timestamp 1606120353
transform 1 0 4048 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1606120353
transform 1 0 6716 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_13_56
timestamp 1606120353
transform 1 0 6256 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_14_53
timestamp 1606120353
transform 1 0 5980 0 -1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_14_62
timestamp 1606120353
transform 1 0 6808 0 -1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_14_70
timestamp 1606120353
transform 1 0 7544 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_74
timestamp 1606120353
transform 1 0 7912 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_13_68
timestamp 1606120353
transform 1 0 7360 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A
timestamp 1606120353
transform 1 0 7728 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _0979_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 7728 0 -1 10336
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILLER_14_81
timestamp 1606120353
transform 1 0 8556 0 -1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_13_82
timestamp 1606120353
transform 1 0 8648 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_13_78
timestamp 1606120353
transform 1 0 8280 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__C
timestamp 1606120353
transform 1 0 8464 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__B
timestamp 1606120353
transform 1 0 8096 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_87
timestamp 1606120353
transform 1 0 9108 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1241__CLK
timestamp 1606120353
transform 1 0 8924 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_13_99
timestamp 1606120353
transform 1 0 10212 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_13_93
timestamp 1606120353
transform 1 0 9660 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_13_91
timestamp 1606120353
transform 1 0 9476 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__D
timestamp 1606120353
transform 1 0 10028 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1241__D
timestamp 1606120353
transform 1 0 9292 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1606120353
transform 1 0 9568 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_14_108
timestamp 1606120353
transform 1 0 11040 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_105
timestamp 1606120353
transform 1 0 10764 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__C
timestamp 1606120353
transform 1 0 11224 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__B
timestamp 1606120353
transform 1 0 10580 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A
timestamp 1606120353
transform 1 0 10948 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1241_
timestamp 1606120353
transform 1 0 9292 0 -1 10336
box 0 -48 1748 592
use sky130_fd_sc_hd__nand4_4  _0963_
timestamp 1606120353
transform 1 0 11132 0 1 9248
box 0 -48 1564 592
use sky130_fd_sc_hd__decap_4  FILLER_14_112
timestamp 1606120353
transform 1 0 11408 0 -1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_14_118
timestamp 1606120353
transform 1 0 11960 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__D
timestamp 1606120353
transform 1 0 11776 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__B
timestamp 1606120353
transform 1 0 12144 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1606120353
transform 1 0 12328 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_14_123
timestamp 1606120353
transform 1 0 12420 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_126
timestamp 1606120353
transform 1 0 12696 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__B
timestamp 1606120353
transform 1 0 12604 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_14_127
timestamp 1606120353
transform 1 0 12788 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_13_130
timestamp 1606120353
transform 1 0 13064 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__A
timestamp 1606120353
transform 1 0 12880 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0912_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 12880 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_14_131
timestamp 1606120353
transform 1 0 13156 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A
timestamp 1606120353
transform 1 0 13248 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_135
timestamp 1606120353
transform 1 0 13524 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_143
timestamp 1606120353
transform 1 0 14260 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__C
timestamp 1606120353
transform 1 0 13708 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A
timestamp 1606120353
transform 1 0 13340 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _0931_
timestamp 1606120353
transform 1 0 13432 0 1 9248
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_13_154
timestamp 1606120353
transform 1 0 15272 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 1606120353
transform 1 0 14996 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_147
timestamp 1606120353
transform 1 0 14628 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__A2_N
timestamp 1606120353
transform 1 0 14812 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__A1_N
timestamp 1606120353
transform 1 0 14444 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1606120353
transform 1 0 15180 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__a2bb2oi_4  _0971_
timestamp 1606120353
transform 1 0 13892 0 -1 10336
box 0 -48 1932 592
use sky130_fd_sc_hd__fill_2  FILLER_14_164
timestamp 1606120353
transform 1 0 16192 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_160
timestamp 1606120353
transform 1 0 15824 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_162
timestamp 1606120353
transform 1 0 16008 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_158
timestamp 1606120353
transform 1 0 15640 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A1
timestamp 1606120353
transform 1 0 16192 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__B1
timestamp 1606120353
transform 1 0 15824 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__B2
timestamp 1606120353
transform 1 0 15456 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__B1
timestamp 1606120353
transform 1 0 16008 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_14_172
timestamp 1606120353
transform 1 0 16928 0 -1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_14_168
timestamp 1606120353
transform 1 0 16560 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1606120353
transform 1 0 16376 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A1
timestamp 1606120353
transform 1 0 16376 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__B1
timestamp 1606120353
transform 1 0 16744 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A2
timestamp 1606120353
transform 1 0 16560 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0933_
timestamp 1606120353
transform 1 0 16744 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606120353
transform -1 0 18860 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606120353
transform -1 0 18860 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1606120353
transform 1 0 17940 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_13_182
timestamp 1606120353
transform 1 0 17848 0 1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_14_180
timestamp 1606120353
transform 1 0 17664 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_14_184
timestamp 1606120353
transform 1 0 18032 0 -1 10336
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1283_
timestamp 1606120353
transform 1 0 1380 0 1 10336
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606120353
transform 1 0 1104 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_15_22
timestamp 1606120353
transform 1 0 3128 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1220_
timestamp 1606120353
transform 1 0 4324 0 1 10336
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1606120353
transform 1 0 3956 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__D
timestamp 1606120353
transform 1 0 3772 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__CLK
timestamp 1606120353
transform 1 0 3312 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_15_26
timestamp 1606120353
transform 1 0 3496 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_15_32
timestamp 1606120353
transform 1 0 4048 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_15_54
timestamp 1606120353
transform 1 0 6072 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_15_66
timestamp 1606120353
transform 1 0 7176 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__and3_4  _0964_
timestamp 1606120353
transform 1 0 8004 0 1 10336
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__A
timestamp 1606120353
transform 1 0 7820 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__B
timestamp 1606120353
transform 1 0 9016 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__C
timestamp 1606120353
transform 1 0 7452 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1606120353
transform 1 0 7636 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_84
timestamp 1606120353
transform 1 0 8832 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_88
timestamp 1606120353
transform 1 0 9200 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1240_
timestamp 1606120353
transform 1 0 9660 0 1 10336
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1606120353
transform 1 0 9568 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1240__D
timestamp 1606120353
transform 1 0 9384 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _0972_
timestamp 1606120353
transform 1 0 12880 0 1 10336
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A
timestamp 1606120353
transform 1 0 12420 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__C
timestamp 1606120353
transform 1 0 11592 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__C
timestamp 1606120353
transform 1 0 12052 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_112
timestamp 1606120353
transform 1 0 11408 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_15_116
timestamp 1606120353
transform 1 0 11776 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_15_121
timestamp 1606120353
transform 1 0 12236 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_15_125
timestamp 1606120353
transform 1 0 12604 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1606120353
transform 1 0 15180 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__A2
timestamp 1606120353
transform 1 0 14996 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__D
timestamp 1606120353
transform 1 0 14628 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_145
timestamp 1606120353
transform 1 0 14444 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_149
timestamp 1606120353
transform 1 0 14812 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_154
timestamp 1606120353
transform 1 0 15272 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0932_
timestamp 1606120353
transform 1 0 15640 0 1 10336
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__A1
timestamp 1606120353
transform 1 0 15456 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_15_171
timestamp 1606120353
transform 1 0 16836 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606120353
transform -1 0 18860 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_15_183
timestamp 1606120353
transform 1 0 17940 0 1 10336
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_15_189
timestamp 1606120353
transform 1 0 18492 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1285_
timestamp 1606120353
transform 1 0 1472 0 -1 11424
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606120353
transform 1 0 1104 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1606120353
transform 1 0 1380 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1222_
timestamp 1606120353
transform 1 0 4140 0 -1 11424
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__CLK
timestamp 1606120353
transform 1 0 3956 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_16_23
timestamp 1606120353
transform 1 0 3220 0 -1 11424
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1606120353
transform 1 0 6716 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__CLK
timestamp 1606120353
transform 1 0 7084 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_16_52
timestamp 1606120353
transform 1 0 5888 0 -1 11424
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_16_60
timestamp 1606120353
transform 1 0 6624 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_16_62
timestamp 1606120353
transform 1 0 6808 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__B
timestamp 1606120353
transform 1 0 8004 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__CLK
timestamp 1606120353
transform 1 0 7452 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_67
timestamp 1606120353
transform 1 0 7268 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_16_71
timestamp 1606120353
transform 1 0 7636 0 -1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_16_77
timestamp 1606120353
transform 1 0 8188 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__nand4_4  _0977_
timestamp 1606120353
transform 1 0 10028 0 -1 11424
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A
timestamp 1606120353
transform 1 0 9844 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1240__CLK
timestamp 1606120353
transform 1 0 9476 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_89
timestamp 1606120353
transform 1 0 9292 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1606120353
transform 1 0 9660 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _0927_
timestamp 1606120353
transform 1 0 12420 0 -1 11424
box 0 -48 1564 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1606120353
transform 1 0 12328 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A
timestamp 1606120353
transform 1 0 11776 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A2
timestamp 1606120353
transform 1 0 12144 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_114
timestamp 1606120353
transform 1 0 11592 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_118
timestamp 1606120353
transform 1 0 11960 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0947_
timestamp 1606120353
transform 1 0 14720 0 -1 11424
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A2
timestamp 1606120353
transform 1 0 14536 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__B1_N
timestamp 1606120353
transform 1 0 14168 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_140
timestamp 1606120353
transform 1 0 13984 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_144
timestamp 1606120353
transform 1 0 14352 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A2
timestamp 1606120353
transform 1 0 16100 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A1
timestamp 1606120353
transform 1 0 16468 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_161
timestamp 1606120353
transform 1 0 15916 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_165
timestamp 1606120353
transform 1 0 16284 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_16_169
timestamp 1606120353
transform 1 0 16652 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606120353
transform -1 0 18860 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1606120353
transform 1 0 17940 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_16_181
timestamp 1606120353
transform 1 0 17756 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_16_184
timestamp 1606120353
transform 1 0 18032 0 -1 11424
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1243_
timestamp 1606120353
transform 1 0 1380 0 1 11424
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606120353
transform 1 0 1104 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_17_22
timestamp 1606120353
transform 1 0 3128 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1235_
timestamp 1606120353
transform 1 0 4324 0 1 11424
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1606120353
transform 1 0 3956 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__D
timestamp 1606120353
transform 1 0 3772 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__D
timestamp 1606120353
transform 1 0 3404 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_27
timestamp 1606120353
transform 1 0 3588 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_17_32
timestamp 1606120353
transform 1 0 4048 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1212_
timestamp 1606120353
transform 1 0 7084 0 1 11424
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__D
timestamp 1606120353
transform 1 0 6900 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__D
timestamp 1606120353
transform 1 0 6532 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_17_54
timestamp 1606120353
transform 1 0 6072 0 1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_17_58
timestamp 1606120353
transform 1 0 6440 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_17_61
timestamp 1606120353
transform 1 0 6716 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_17_84
timestamp 1606120353
transform 1 0 8832 0 1 11424
box 0 -48 736 592
use sky130_fd_sc_hd__nand4_4  _0962_
timestamp 1606120353
transform 1 0 10948 0 1 11424
box 0 -48 1564 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1606120353
transform 1 0 9568 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__D
timestamp 1606120353
transform 1 0 10764 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A1
timestamp 1606120353
transform 1 0 10396 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__C
timestamp 1606120353
transform 1 0 10028 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_17_93
timestamp 1606120353
transform 1 0 9660 0 1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_17_99
timestamp 1606120353
transform 1 0 10212 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_103
timestamp 1606120353
transform 1 0 10580 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A
timestamp 1606120353
transform 1 0 13156 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__C
timestamp 1606120353
transform 1 0 12788 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_17_124
timestamp 1606120353
transform 1 0 12512 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_17_129
timestamp 1606120353
transform 1 0 12972 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0987_
timestamp 1606120353
transform 1 0 13340 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1606120353
transform 1 0 15180 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__D
timestamp 1606120353
transform 1 0 14628 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__B1
timestamp 1606120353
transform 1 0 14996 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_145
timestamp 1606120353
transform 1 0 14444 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_149
timestamp 1606120353
transform 1 0 14812 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_17_154
timestamp 1606120353
transform 1 0 15272 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _0954_
timestamp 1606120353
transform 1 0 15548 0 1 11424
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__B1
timestamp 1606120353
transform 1 0 16928 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A1
timestamp 1606120353
transform 1 0 17296 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_170
timestamp 1606120353
transform 1 0 16744 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_174
timestamp 1606120353
transform 1 0 17112 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606120353
transform -1 0 18860 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_17_178
timestamp 1606120353
transform 1 0 17480 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1248_
timestamp 1606120353
transform 1 0 1380 0 -1 12512
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606120353
transform 1 0 1104 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_18_22
timestamp 1606120353
transform 1 0 3128 0 -1 12512
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1242_
timestamp 1606120353
transform 1 0 4232 0 -1 12512
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__CLK
timestamp 1606120353
transform 1 0 4048 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_30
timestamp 1606120353
transform 1 0 3864 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1214_
timestamp 1606120353
transform 1 0 6808 0 -1 12512
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1606120353
transform 1 0 6716 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_18_53
timestamp 1606120353
transform 1 0 5980 0 -1 12512
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_18_81
timestamp 1606120353
transform 1 0 8556 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__o21a_4  _0906_
timestamp 1606120353
transform 1 0 10488 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A2
timestamp 1606120353
transform 1 0 10304 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__B1
timestamp 1606120353
transform 1 0 9936 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_18_93
timestamp 1606120353
transform 1 0 9660 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_18_98
timestamp 1606120353
transform 1 0 10120 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_118
timestamp 1606120353
transform 1 0 11960 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_114
timestamp 1606120353
transform 1 0 11592 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__B
timestamp 1606120353
transform 1 0 12144 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__B
timestamp 1606120353
transform 1 0 11776 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_127
timestamp 1606120353
transform 1 0 12788 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_123
timestamp 1606120353
transform 1 0 12420 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__C
timestamp 1606120353
transform 1 0 12972 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__B
timestamp 1606120353
transform 1 0 12604 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1606120353
transform 1 0 12328 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__nand4_4  _0986_
timestamp 1606120353
transform 1 0 13156 0 -1 12512
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A2_N
timestamp 1606120353
transform 1 0 14904 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_148
timestamp 1606120353
transform 1 0 14720 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_18_152
timestamp 1606120353
transform 1 0 15088 0 -1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__a21o_4  _0997_
timestamp 1606120353
transform 1 0 16100 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A2
timestamp 1606120353
transform 1 0 15548 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A1
timestamp 1606120353
transform 1 0 15916 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_18_156
timestamp 1606120353
transform 1 0 15456 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_18_159
timestamp 1606120353
transform 1 0 15732 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_18_175
timestamp 1606120353
transform 1 0 17204 0 -1 12512
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606120353
transform -1 0 18860 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1606120353
transform 1 0 17940 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_18_184
timestamp 1606120353
transform 1 0 18032 0 -1 12512
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1606120353
transform 1 0 1380 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 1606120353
transform 1 0 2116 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 1606120353
transform 1 0 1748 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1606120353
transform 1 0 1380 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__CLK
timestamp 1606120353
transform 1 0 1564 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__D
timestamp 1606120353
transform 1 0 1932 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__D
timestamp 1606120353
transform 1 0 1564 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606120353
transform 1 0 1104 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606120353
transform 1 0 1104 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_20_19
timestamp 1606120353
transform 1 0 2852 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_19_22
timestamp 1606120353
transform 1 0 3128 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_19_19
timestamp 1606120353
transform 1 0 2852 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_19_15
timestamp 1606120353
transform 1 0 2484 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__CLK
timestamp 1606120353
transform 1 0 2300 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__D
timestamp 1606120353
transform 1 0 2944 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_20_7
timestamp 1606120353
transform 1 0 1748 0 -1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1245_
timestamp 1606120353
transform 1 0 2944 0 -1 13600
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1244_
timestamp 1606120353
transform 1 0 4048 0 1 12512
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1606120353
transform 1 0 3956 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__D
timestamp 1606120353
transform 1 0 3772 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__CLK
timestamp 1606120353
transform 1 0 3312 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__CLK
timestamp 1606120353
transform 1 0 4876 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_19_26
timestamp 1606120353
transform 1 0 3496 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_20_39
timestamp 1606120353
transform 1 0 4692 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_20_43
timestamp 1606120353
transform 1 0 5060 0 -1 13600
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1606120353
transform 1 0 6716 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__CLK
timestamp 1606120353
transform 1 0 5704 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_19_51
timestamp 1606120353
transform 1 0 5796 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_19_63
timestamp 1606120353
transform 1 0 6900 0 1 12512
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_20_49
timestamp 1606120353
transform 1 0 5612 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_20_52
timestamp 1606120353
transform 1 0 5888 0 -1 13600
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_20_60
timestamp 1606120353
transform 1 0 6624 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_20_62
timestamp 1606120353
transform 1 0 6808 0 -1 13600
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1239_
timestamp 1606120353
transform 1 0 7544 0 -1 13600
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__D
timestamp 1606120353
transform 1 0 7544 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__CLK
timestamp 1606120353
transform 1 0 7912 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_19_69
timestamp 1606120353
transform 1 0 7452 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_19_72
timestamp 1606120353
transform 1 0 7728 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_19_76
timestamp 1606120353
transform 1 0 8096 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_19_88
timestamp 1606120353
transform 1 0 9200 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1606120353
transform 1 0 9568 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__B
timestamp 1606120353
transform 1 0 9384 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_20_89
timestamp 1606120353
transform 1 0 9292 0 -1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A
timestamp 1606120353
transform 1 0 9936 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__C
timestamp 1606120353
transform 1 0 9752 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_19_93
timestamp 1606120353
transform 1 0 9660 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_20_93
timestamp 1606120353
transform 1 0 9660 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_20_96
timestamp 1606120353
transform 1 0 9936 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__B
timestamp 1606120353
transform 1 0 10120 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_98
timestamp 1606120353
transform 1 0 10120 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_19_102
timestamp 1606120353
transform 1 0 10488 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A
timestamp 1606120353
transform 1 0 10304 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__nand3_4  _0995_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 10304 0 -1 13600
box 0 -48 1288 592
use sky130_fd_sc_hd__nand3_4  _0992_
timestamp 1606120353
transform 1 0 10580 0 1 12512
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_1  FILLER_20_121
timestamp 1606120353
transform 1 0 12236 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_20_118
timestamp 1606120353
transform 1 0 11960 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_20_114
timestamp 1606120353
transform 1 0 11592 0 -1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_19_121
timestamp 1606120353
transform 1 0 12236 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_117
timestamp 1606120353
transform 1 0 11868 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__B
timestamp 1606120353
transform 1 0 12052 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__C
timestamp 1606120353
transform 1 0 12052 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_20_123
timestamp 1606120353
transform 1 0 12420 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A
timestamp 1606120353
transform 1 0 12420 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1606120353
transform 1 0 12328 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__or3_4  _0994_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 12512 0 -1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__nand3_4  _0996_
timestamp 1606120353
transform 1 0 12604 0 1 12512
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_20_137
timestamp 1606120353
transform 1 0 13708 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_133
timestamp 1606120353
transform 1 0 13340 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_143
timestamp 1606120353
transform 1 0 14260 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_139
timestamp 1606120353
transform 1 0 13892 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A
timestamp 1606120353
transform 1 0 13892 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__B1
timestamp 1606120353
transform 1 0 13524 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__B2
timestamp 1606120353
transform 1 0 14076 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_19_147
timestamp 1606120353
transform 1 0 14628 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A1_N
timestamp 1606120353
transform 1 0 14444 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__B1
timestamp 1606120353
transform 1 0 14996 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1606120353
transform 1 0 15180 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__a21o_4  _0999_
timestamp 1606120353
transform 1 0 15272 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__a2bb2oi_4  _0985_
timestamp 1606120353
transform 1 0 14076 0 -1 13600
box 0 -48 1932 592
use sky130_fd_sc_hd__decap_4  FILLER_20_162
timestamp 1606120353
transform 1 0 16008 0 -1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_20_169
timestamp 1606120353
transform 1 0 16652 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_20_166
timestamp 1606120353
transform 1 0 16376 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_19_170
timestamp 1606120353
transform 1 0 16744 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1606120353
transform 1 0 16376 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A2
timestamp 1606120353
transform 1 0 16468 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A2
timestamp 1606120353
transform 1 0 16560 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_20_173
timestamp 1606120353
transform 1 0 17020 0 -1 13600
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_19_174
timestamp 1606120353
transform 1 0 17112 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A1
timestamp 1606120353
transform 1 0 17296 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A1
timestamp 1606120353
transform 1 0 16836 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__B1
timestamp 1606120353
transform 1 0 16928 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606120353
transform -1 0 18860 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606120353
transform -1 0 18860 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1606120353
transform 1 0 17940 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_19_178
timestamp 1606120353
transform 1 0 17480 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_20_181
timestamp 1606120353
transform 1 0 17756 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_20_184
timestamp 1606120353
transform 1 0 18032 0 -1 13600
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606120353
transform 1 0 1104 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__D
timestamp 1606120353
transform 1 0 2300 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__CLK
timestamp 1606120353
transform 1 0 2668 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1606120353
transform 1 0 1380 0 1 13600
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_21_11
timestamp 1606120353
transform 1 0 2116 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_15
timestamp 1606120353
transform 1 0 2484 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_21_19
timestamp 1606120353
transform 1 0 2852 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1606120353
transform 1 0 3956 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_21_32
timestamp 1606120353
transform 1 0 4048 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_21_44
timestamp 1606120353
transform 1 0 5152 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1221_
timestamp 1606120353
transform 1 0 5704 0 1 13600
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__D
timestamp 1606120353
transform 1 0 5520 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1606120353
transform 1 0 7452 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_21_81
timestamp 1606120353
transform 1 0 8556 0 1 13600
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _0961_
timestamp 1606120353
transform 1 0 11040 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1606120353
transform 1 0 9568 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__A
timestamp 1606120353
transform 1 0 10764 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__C
timestamp 1606120353
transform 1 0 10304 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_21_89
timestamp 1606120353
transform 1 0 9292 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_21_93
timestamp 1606120353
transform 1 0 9660 0 1 13600
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_21_99
timestamp 1606120353
transform 1 0 10212 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_21_102
timestamp 1606120353
transform 1 0 10488 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_21_107
timestamp 1606120353
transform 1 0 10948 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__nand4_4  _0930_
timestamp 1606120353
transform 1 0 12052 0 1 13600
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__D
timestamp 1606120353
transform 1 0 11868 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__A
timestamp 1606120353
transform 1 0 11500 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_111
timestamp 1606120353
transform 1 0 11316 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_115
timestamp 1606120353
transform 1 0 11684 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0984_
timestamp 1606120353
transform 1 0 15272 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1606120353
transform 1 0 15180 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A
timestamp 1606120353
transform 1 0 14996 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A2
timestamp 1606120353
transform 1 0 13984 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__B1
timestamp 1606120353
transform 1 0 14352 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_21_136
timestamp 1606120353
transform 1 0 13616 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_21_142
timestamp 1606120353
transform 1 0 14168 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_21_146
timestamp 1606120353
transform 1 0 14536 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_21_150
timestamp 1606120353
transform 1 0 14904 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__a21o_4  _0998_
timestamp 1606120353
transform 1 0 16468 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__B1
timestamp 1606120353
transform 1 0 16284 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__B1
timestamp 1606120353
transform 1 0 15916 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_21_157
timestamp 1606120353
transform 1 0 15548 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_21_163
timestamp 1606120353
transform 1 0 16100 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606120353
transform -1 0 18860 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_21_179
timestamp 1606120353
transform 1 0 17572 0 1 13600
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_21_187
timestamp 1606120353
transform 1 0 18308 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1247_
timestamp 1606120353
transform 1 0 2300 0 -1 14688
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606120353
transform 1 0 1104 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1606120353
transform 1 0 1380 0 -1 14688
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_22_11
timestamp 1606120353
transform 1 0 2116 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__CLK
timestamp 1606120353
transform 1 0 4876 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_22_32
timestamp 1606120353
transform 1 0 4048 0 -1 14688
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_22_40
timestamp 1606120353
transform 1 0 4784 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_22_43
timestamp 1606120353
transform 1 0 5060 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1606120353
transform 1 0 6716 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_22_55
timestamp 1606120353
transform 1 0 6164 0 -1 14688
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_22_62
timestamp 1606120353
transform 1 0 6808 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_22_74
timestamp 1606120353
transform 1 0 7912 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_22_86
timestamp 1606120353
transform 1 0 9016 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__inv_8  _0908_
timestamp 1606120353
transform 1 0 10764 0 -1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__decap_6  FILLER_22_98
timestamp 1606120353
transform 1 0 10120 0 -1 14688
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_22_104
timestamp 1606120353
transform 1 0 10672 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_22_114
timestamp 1606120353
transform 1 0 11592 0 -1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_22_121
timestamp 1606120353
transform 1 0 12236 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_22_118
timestamp 1606120353
transform 1 0 11960 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A
timestamp 1606120353
transform 1 0 12052 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1606120353
transform 1 0 12328 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_22_127
timestamp 1606120353
transform 1 0 12788 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_123
timestamp 1606120353
transform 1 0 12420 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__B
timestamp 1606120353
transform 1 0 12604 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_22_131
timestamp 1606120353
transform 1 0 13156 0 -1 14688
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__C
timestamp 1606120353
transform 1 0 12972 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0991_
timestamp 1606120353
transform 1 0 13984 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A1
timestamp 1606120353
transform 1 0 13800 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_22_137
timestamp 1606120353
transform 1 0 13708 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_22_152
timestamp 1606120353
transform 1 0 15088 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__a21o_4  _1001_
timestamp 1606120353
transform 1 0 15916 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A2
timestamp 1606120353
transform 1 0 15732 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A1
timestamp 1606120353
transform 1 0 15364 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_157
timestamp 1606120353
transform 1 0 15548 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_22_173
timestamp 1606120353
transform 1 0 17020 0 -1 14688
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606120353
transform -1 0 18860 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1606120353
transform 1 0 17940 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_22_181
timestamp 1606120353
transform 1 0 17756 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_22_184
timestamp 1606120353
transform 1 0 18032 0 -1 14688
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606120353
transform 1 0 1104 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1606120353
transform 1 0 1380 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_23_15
timestamp 1606120353
transform 1 0 2484 0 1 14688
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1223_
timestamp 1606120353
transform 1 0 4876 0 1 14688
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1606120353
transform 1 0 3956 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__D
timestamp 1606120353
transform 1 0 3496 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__D
timestamp 1606120353
transform 1 0 4692 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__CLK
timestamp 1606120353
transform 1 0 4232 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_23_23
timestamp 1606120353
transform 1 0 3220 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_23_28
timestamp 1606120353
transform 1 0 3680 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_23_32
timestamp 1606120353
transform 1 0 4048 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_23_36
timestamp 1606120353
transform 1 0 4416 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_23_60
timestamp 1606120353
transform 1 0 6624 0 1 14688
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_23_66
timestamp 1606120353
transform 1 0 7176 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__D
timestamp 1606120353
transform 1 0 7268 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__CLK
timestamp 1606120353
transform 1 0 7636 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_69
timestamp 1606120353
transform 1 0 7452 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_23_73
timestamp 1606120353
transform 1 0 7820 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_23_85
timestamp 1606120353
transform 1 0 8924 0 1 14688
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_23_91
timestamp 1606120353
transform 1 0 9476 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1606120353
transform 1 0 9568 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_23_93
timestamp 1606120353
transform 1 0 9660 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__D
timestamp 1606120353
transform 1 0 9844 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_97
timestamp 1606120353
transform 1 0 10028 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__CLK
timestamp 1606120353
transform 1 0 10212 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_101
timestamp 1606120353
transform 1 0 10396 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_23_107
timestamp 1606120353
transform 1 0 10948 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A2
timestamp 1606120353
transform 1 0 10764 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A1
timestamp 1606120353
transform 1 0 11132 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0993_
timestamp 1606120353
transform 1 0 11316 0 1 14688
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A
timestamp 1606120353
transform 1 0 12972 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_124
timestamp 1606120353
transform 1 0 12512 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_23_128
timestamp 1606120353
transform 1 0 12880 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_23_131
timestamp 1606120353
transform 1 0 13156 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_23_135
timestamp 1606120353
transform 1 0 13524 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_23_138
timestamp 1606120353
transform 1 0 13800 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__B1
timestamp 1606120353
transform 1 0 13616 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A2
timestamp 1606120353
transform 1 0 13984 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0957_
timestamp 1606120353
transform 1 0 14168 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_23_145
timestamp 1606120353
transform 1 0 14444 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__A
timestamp 1606120353
transform 1 0 14628 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_149
timestamp 1606120353
transform 1 0 14812 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__B
timestamp 1606120353
transform 1 0 14996 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1606120353
transform 1 0 15180 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_23_154
timestamp 1606120353
transform 1 0 15272 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _1002_
timestamp 1606120353
transform 1 0 16100 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A
timestamp 1606120353
transform 1 0 15824 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__B1
timestamp 1606120353
transform 1 0 15456 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_158
timestamp 1606120353
transform 1 0 15640 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_23_162
timestamp 1606120353
transform 1 0 16008 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1606120353
transform 1 0 17204 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606120353
transform -1 0 18860 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__A1
timestamp 1606120353
transform 1 0 17388 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_23_179
timestamp 1606120353
transform 1 0 17572 0 1 14688
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_23_187
timestamp 1606120353
transform 1 0 18308 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606120353
transform 1 0 1104 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__D
timestamp 1606120353
transform 1 0 1564 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__CLK
timestamp 1606120353
transform 1 0 1932 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__CLK
timestamp 1606120353
transform 1 0 2760 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1606120353
transform 1 0 1380 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1606120353
transform 1 0 1748 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_24_11
timestamp 1606120353
transform 1 0 2116 0 -1 15776
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_24_17
timestamp 1606120353
transform 1 0 2668 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_24_20
timestamp 1606120353
transform 1 0 2944 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1249_
timestamp 1606120353
transform 1 0 3496 0 -1 15776
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__CLK
timestamp 1606120353
transform 1 0 3312 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1606120353
transform 1 0 6716 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_24_45
timestamp 1606120353
transform 1 0 5244 0 -1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_24_57
timestamp 1606120353
transform 1 0 6348 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_24_62
timestamp 1606120353
transform 1 0 6808 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_24_66
timestamp 1606120353
transform 1 0 7176 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1215_
timestamp 1606120353
transform 1 0 7268 0 -1 15776
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_8  FILLER_24_86
timestamp 1606120353
transform 1 0 9016 0 -1 15776
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1213_
timestamp 1606120353
transform 1 0 9752 0 -1 15776
box 0 -48 1748 592
use sky130_fd_sc_hd__buf_1  _0967_
timestamp 1606120353
transform 1 0 12972 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1606120353
transform 1 0 12328 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__B1
timestamp 1606120353
transform 1 0 11684 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_113
timestamp 1606120353
transform 1 0 11500 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_24_117
timestamp 1606120353
transform 1 0 11868 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_24_121
timestamp 1606120353
transform 1 0 12236 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_24_123
timestamp 1606120353
transform 1 0 12420 0 -1 15776
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_24_132
timestamp 1606120353
transform 1 0 13248 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0959_
timestamp 1606120353
transform 1 0 13984 0 -1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__B1
timestamp 1606120353
transform 1 0 15272 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A1
timestamp 1606120353
transform 1 0 13800 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A1
timestamp 1606120353
transform 1 0 13432 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_136
timestamp 1606120353
transform 1 0 13616 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_152
timestamp 1606120353
transform 1 0 15088 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__nand2_4  _0975_
timestamp 1606120353
transform 1 0 15824 0 -1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__A2
timestamp 1606120353
transform 1 0 16836 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A1
timestamp 1606120353
transform 1 0 15640 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_156
timestamp 1606120353
transform 1 0 15456 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_169
timestamp 1606120353
transform 1 0 16652 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_24_173
timestamp 1606120353
transform 1 0 17020 0 -1 15776
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606120353
transform -1 0 18860 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1606120353
transform 1 0 17940 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_24_181
timestamp 1606120353
transform 1 0 17756 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_24_184
timestamp 1606120353
transform 1 0 18032 0 -1 15776
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1250_
timestamp 1606120353
transform 1 0 1472 0 1 15776
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606120353
transform 1 0 1104 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1606120353
transform 1 0 1380 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1284_
timestamp 1606120353
transform 1 0 4048 0 1 15776
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1606120353
transform 1 0 3956 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__D
timestamp 1606120353
transform 1 0 3772 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__D
timestamp 1606120353
transform 1 0 3404 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_23
timestamp 1606120353
transform 1 0 3220 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_27
timestamp 1606120353
transform 1 0 3588 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_25_51
timestamp 1606120353
transform 1 0 5796 0 1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_25_63
timestamp 1606120353
transform 1 0 6900 0 1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_25_75
timestamp 1606120353
transform 1 0 8004 0 1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_25_87
timestamp 1606120353
transform 1 0 9108 0 1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__a21bo_4  _1004_
timestamp 1606120353
transform 1 0 11040 0 1 15776
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1606120353
transform 1 0 9568 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A2
timestamp 1606120353
transform 1 0 10856 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A1
timestamp 1606120353
transform 1 0 10488 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_25_91
timestamp 1606120353
transform 1 0 9476 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_25_93
timestamp 1606120353
transform 1 0 9660 0 1 15776
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_25_101
timestamp 1606120353
transform 1 0 10396 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_25_104
timestamp 1606120353
transform 1 0 10672 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0989_
timestamp 1606120353
transform 1 0 12972 0 1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A
timestamp 1606120353
transform 1 0 12788 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_25_121
timestamp 1606120353
transform 1 0 12236 0 1 15776
box 0 -48 552 592
use sky130_fd_sc_hd__a21o_4  _0976_
timestamp 1606120353
transform 1 0 15272 0 1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1606120353
transform 1 0 15180 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__B1
timestamp 1606120353
transform 1 0 13984 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A2
timestamp 1606120353
transform 1 0 14352 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A2
timestamp 1606120353
transform 1 0 14996 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_138
timestamp 1606120353
transform 1 0 13800 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_142
timestamp 1606120353
transform 1 0 14168 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_25_146
timestamp 1606120353
transform 1 0 14536 0 1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_25_150
timestamp 1606120353
transform 1 0 14904 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A
timestamp 1606120353
transform 1 0 16560 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1606120353
transform 1 0 16376 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_25_170
timestamp 1606120353
transform 1 0 16744 0 1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606120353
transform -1 0 18860 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_25_182
timestamp 1606120353
transform 1 0 17848 0 1 15776
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1606120353
transform 1 0 1380 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_26_11
timestamp 1606120353
transform 1 0 2116 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_7
timestamp 1606120353
transform 1 0 1748 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1606120353
transform 1 0 1380 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__D
timestamp 1606120353
transform 1 0 1932 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__D
timestamp 1606120353
transform 1 0 1564 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606120353
transform 1 0 1104 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606120353
transform 1 0 1104 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_26_15
timestamp 1606120353
transform 1 0 2484 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__CLK
timestamp 1606120353
transform 1 0 2300 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1287_
timestamp 1606120353
transform 1 0 1472 0 1 16864
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1286_
timestamp 1606120353
transform 1 0 2760 0 -1 16864
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1224_
timestamp 1606120353
transform 1 0 4692 0 1 16864
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1606120353
transform 1 0 3956 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__D
timestamp 1606120353
transform 1 0 4508 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__CLK
timestamp 1606120353
transform 1 0 4692 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_37
timestamp 1606120353
transform 1 0 4508 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1606120353
transform 1 0 4876 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_27_23
timestamp 1606120353
transform 1 0 3220 0 1 16864
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_27_32
timestamp 1606120353
transform 1 0 4048 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_27_36
timestamp 1606120353
transform 1 0 4416 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1606120353
transform 1 0 6716 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_26_53
timestamp 1606120353
transform 1 0 5980 0 -1 16864
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_26_62
timestamp 1606120353
transform 1 0 6808 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_27_58
timestamp 1606120353
transform 1 0 6440 0 1 16864
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_27_66
timestamp 1606120353
transform 1 0 7176 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__D
timestamp 1606120353
transform 1 0 7268 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__CLK
timestamp 1606120353
transform 1 0 7636 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_26_74
timestamp 1606120353
transform 1 0 7912 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_26_86
timestamp 1606120353
transform 1 0 9016 0 -1 16864
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_27_69
timestamp 1606120353
transform 1 0 7452 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_27_73
timestamp 1606120353
transform 1 0 7820 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_27_85
timestamp 1606120353
transform 1 0 8924 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_27_89
timestamp 1606120353
transform 1 0 9292 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_26_92
timestamp 1606120353
transform 1 0 9568 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__CLK
timestamp 1606120353
transform 1 0 9660 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__D
timestamp 1606120353
transform 1 0 9384 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1606120353
transform 1 0 9568 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_26_110
timestamp 1606120353
transform 1 0 11224 0 -1 16864
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_26_107
timestamp 1606120353
transform 1 0 10948 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__B1_N
timestamp 1606120353
transform 1 0 11040 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_26_95
timestamp 1606120353
transform 1 0 9844 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1252_
timestamp 1606120353
transform 1 0 9660 0 1 16864
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_2  FILLER_27_116
timestamp 1606120353
transform 1 0 11776 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_112
timestamp 1606120353
transform 1 0 11408 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_118
timestamp 1606120353
transform 1 0 11960 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A
timestamp 1606120353
transform 1 0 12144 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__C
timestamp 1606120353
transform 1 0 11960 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A
timestamp 1606120353
transform 1 0 11592 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_131
timestamp 1606120353
transform 1 0 13156 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_127
timestamp 1606120353
transform 1 0 12788 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_123
timestamp 1606120353
transform 1 0 12420 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__D
timestamp 1606120353
transform 1 0 12604 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__C1
timestamp 1606120353
transform 1 0 12972 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1606120353
transform 1 0 12328 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__nand4_4  _0988_
timestamp 1606120353
transform 1 0 12144 0 1 16864
box 0 -48 1564 592
use sky130_fd_sc_hd__fill_2  FILLER_27_141
timestamp 1606120353
transform 1 0 14076 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_137
timestamp 1606120353
transform 1 0 13708 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_26_135
timestamp 1606120353
transform 1 0 13524 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A1
timestamp 1606120353
transform 1 0 14260 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__B1
timestamp 1606120353
transform 1 0 13892 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A2
timestamp 1606120353
transform 1 0 13340 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_149
timestamp 1606120353
transform 1 0 14812 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_145
timestamp 1606120353
transform 1 0 14444 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_26_148
timestamp 1606120353
transform 1 0 14720 0 -1 16864
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__A2
timestamp 1606120353
transform 1 0 14628 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__B1
timestamp 1606120353
transform 1 0 15272 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A
timestamp 1606120353
transform 1 0 14996 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1606120353
transform 1 0 15180 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__a21o_4  _1003_
timestamp 1606120353
transform 1 0 15272 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__a21o_4  _0958_
timestamp 1606120353
transform 1 0 13616 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__inv_8  _0934_
timestamp 1606120353
transform 1 0 15824 0 -1 16864
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__A1
timestamp 1606120353
transform 1 0 15640 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_156
timestamp 1606120353
transform 1 0 15456 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_26_169
timestamp 1606120353
transform 1 0 16652 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_27_166
timestamp 1606120353
transform 1 0 16376 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606120353
transform -1 0 18860 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606120353
transform -1 0 18860 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1606120353
transform 1 0 17940 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_26_181
timestamp 1606120353
transform 1 0 17756 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_26_184
timestamp 1606120353
transform 1 0 18032 0 -1 16864
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_27_178
timestamp 1606120353
transform 1 0 17480 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1251_
timestamp 1606120353
transform 1 0 1472 0 -1 17952
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606120353
transform 1 0 1104 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1606120353
transform 1 0 1380 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__CLK
timestamp 1606120353
transform 1 0 4140 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_28_23
timestamp 1606120353
transform 1 0 3220 0 -1 17952
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_28_31
timestamp 1606120353
transform 1 0 3956 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_28_35
timestamp 1606120353
transform 1 0 4324 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1606120353
transform 1 0 6716 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_28_47
timestamp 1606120353
transform 1 0 5428 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_28_59
timestamp 1606120353
transform 1 0 6532 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_28_62
timestamp 1606120353
transform 1 0 6808 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_28_66
timestamp 1606120353
transform 1 0 7176 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1216_
timestamp 1606120353
transform 1 0 7268 0 -1 17952
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_12  FILLER_28_86
timestamp 1606120353
transform 1 0 9016 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A
timestamp 1606120353
transform 1 0 10764 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_28_98
timestamp 1606120353
transform 1 0 10120 0 -1 17952
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_28_104
timestamp 1606120353
transform 1 0 10672 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_28_107
timestamp 1606120353
transform 1 0 10948 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _0904_
timestamp 1606120353
transform 1 0 11316 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__a211o_4  _0990_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 12972 0 -1 17952
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1606120353
transform 1 0 12328 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__B
timestamp 1606120353
transform 1 0 11776 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__B
timestamp 1606120353
transform 1 0 12144 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__A2
timestamp 1606120353
transform 1 0 12788 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_114
timestamp 1606120353
transform 1 0 11592 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_118
timestamp 1606120353
transform 1 0 11960 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_28_123
timestamp 1606120353
transform 1 0 12420 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _0938_
timestamp 1606120353
transform 1 0 14996 0 -1 17952
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__B2
timestamp 1606120353
transform 1 0 14812 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__B1
timestamp 1606120353
transform 1 0 14444 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_143
timestamp 1606120353
transform 1 0 14260 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_147
timestamp 1606120353
transform 1 0 14628 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A1
timestamp 1606120353
transform 1 0 16008 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__B1
timestamp 1606120353
transform 1 0 16376 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__B1
timestamp 1606120353
transform 1 0 16744 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_160
timestamp 1606120353
transform 1 0 15824 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_164
timestamp 1606120353
transform 1 0 16192 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_168
timestamp 1606120353
transform 1 0 16560 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_28_172
timestamp 1606120353
transform 1 0 16928 0 -1 17952
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606120353
transform -1 0 18860 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1606120353
transform 1 0 17940 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_28_180
timestamp 1606120353
transform 1 0 17664 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_28_184
timestamp 1606120353
transform 1 0 18032 0 -1 17952
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606120353
transform 1 0 1104 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__CLK
timestamp 1606120353
transform 1 0 1564 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1606120353
transform 1 0 1380 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_29_7
timestamp 1606120353
transform 1 0 1748 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_29_19
timestamp 1606120353
transform 1 0 2852 0 1 17952
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1217_
timestamp 1606120353
transform 1 0 4140 0 1 17952
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1606120353
transform 1 0 3956 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__D
timestamp 1606120353
transform 1 0 3772 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_27
timestamp 1606120353
transform 1 0 3588 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_29_32
timestamp 1606120353
transform 1 0 4048 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1209_
timestamp 1606120353
transform 1 0 6624 0 1 17952
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__D
timestamp 1606120353
transform 1 0 6440 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__CLK
timestamp 1606120353
transform 1 0 6072 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_52
timestamp 1606120353
transform 1 0 5888 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_56
timestamp 1606120353
transform 1 0 6256 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_29_79
timestamp 1606120353
transform 1 0 8372 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__nor3_4  _0910_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 11224 0 1 17952
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1606120353
transform 1 0 9568 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__B
timestamp 1606120353
transform 1 0 10764 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__A
timestamp 1606120353
transform 1 0 10396 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_29_91
timestamp 1606120353
transform 1 0 9476 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_29_93
timestamp 1606120353
transform 1 0 9660 0 1 17952
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_29_103
timestamp 1606120353
transform 1 0 10580 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_29_107
timestamp 1606120353
transform 1 0 10948 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A
timestamp 1606120353
transform 1 0 12604 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__B1
timestamp 1606120353
transform 1 0 13156 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_123
timestamp 1606120353
transform 1 0 12420 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_29_127
timestamp 1606120353
transform 1 0 12788 0 1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__a2bb2oi_4  _0974_
timestamp 1606120353
transform 1 0 15272 0 1 17952
box 0 -48 1932 592
use sky130_fd_sc_hd__a21o_4  _1005_
timestamp 1606120353
transform 1 0 13340 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1606120353
transform 1 0 15180 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A2
timestamp 1606120353
transform 1 0 14996 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A2_N
timestamp 1606120353
transform 1 0 14628 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_145
timestamp 1606120353
transform 1 0 14444 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_149
timestamp 1606120353
transform 1 0 14812 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_29_175
timestamp 1606120353
transform 1 0 17204 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606120353
transform -1 0 18860 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_29_187
timestamp 1606120353
transform 1 0 18308 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606120353
transform 1 0 1104 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__D
timestamp 1606120353
transform 1 0 1564 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1606120353
transform 1 0 1380 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_30_7
timestamp 1606120353
transform 1 0 1748 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_30_19
timestamp 1606120353
transform 1 0 2852 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_clk_A
timestamp 1606120353
transform 1 0 4876 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_30_31
timestamp 1606120353
transform 1 0 3956 0 -1 19040
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_30_39
timestamp 1606120353
transform 1 0 4692 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_43
timestamp 1606120353
transform 1 0 5060 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1606120353
transform 1 0 6716 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_clk_A
timestamp 1606120353
transform 1 0 6440 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__CLK
timestamp 1606120353
transform 1 0 5244 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_30_47
timestamp 1606120353
transform 1 0 5428 0 -1 19040
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_30_55
timestamp 1606120353
transform 1 0 6164 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_30_60
timestamp 1606120353
transform 1 0 6624 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_30_62
timestamp 1606120353
transform 1 0 6808 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_30_74
timestamp 1606120353
transform 1 0 7912 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_30_86
timestamp 1606120353
transform 1 0 9016 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__nor2_4  _0909_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 10764 0 -1 19040
box 0 -48 828 592
use sky130_fd_sc_hd__decap_6  FILLER_30_98
timestamp 1606120353
transform 1 0 10120 0 -1 19040
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_30_104
timestamp 1606120353
transform 1 0 10672 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_30_114
timestamp 1606120353
transform 1 0 11592 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__C
timestamp 1606120353
transform 1 0 11776 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_118
timestamp 1606120353
transform 1 0 11960 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A1
timestamp 1606120353
transform 1 0 12144 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1606120353
transform 1 0 12328 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0926_
timestamp 1606120353
transform 1 0 12420 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_30_126
timestamp 1606120353
transform 1 0 12696 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__B1
timestamp 1606120353
transform 1 0 12880 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_130
timestamp 1606120353
transform 1 0 13064 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__B1_N
timestamp 1606120353
transform 1 0 13248 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _1006_
timestamp 1606120353
transform 1 0 13708 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A1_N
timestamp 1606120353
transform 1 0 15272 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_30_134
timestamp 1606120353
transform 1 0 13432 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1606120353
transform 1 0 14812 0 -1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_30_153
timestamp 1606120353
transform 1 0 15180 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__o21ai_4  _0939_
timestamp 1606120353
transform 1 0 15640 0 -1 19040
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_30_156
timestamp 1606120353
transform 1 0 15456 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_30_171
timestamp 1606120353
transform 1 0 16836 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606120353
transform -1 0 18860 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1606120353
transform 1 0 17940 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_30_184
timestamp 1606120353
transform 1 0 18032 0 -1 19040
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1254_
timestamp 1606120353
transform 1 0 1380 0 1 19040
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606120353
transform 1 0 1104 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_31_22
timestamp 1606120353
transform 1 0 3128 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_31_32
timestamp 1606120353
transform 1 0 4048 0 1 19040
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_31_30
timestamp 1606120353
transform 1 0 3864 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_31_26
timestamp 1606120353
transform 1 0 3496 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__CLK
timestamp 1606120353
transform 1 0 3680 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__D
timestamp 1606120353
transform 1 0 3312 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1606120353
transform 1 0 3956 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_31_38
timestamp 1606120353
transform 1 0 4600 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__D
timestamp 1606120353
transform 1 0 4692 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_clk /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 4876 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1210_
timestamp 1606120353
transform 1 0 5152 0 1 19040
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__A
timestamp 1606120353
transform 1 0 7084 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_63
timestamp 1606120353
transform 1 0 6900 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_clk
timestamp 1606120353
transform 1 0 7636 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__B
timestamp 1606120353
transform 1 0 7452 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_clk_A
timestamp 1606120353
transform 1 0 8096 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_67
timestamp 1606120353
transform 1 0 7268 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_74
timestamp 1606120353
transform 1 0 7912 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_31_78
timestamp 1606120353
transform 1 0 8280 0 1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__inv_8  _0911_
timestamp 1606120353
transform 1 0 10672 0 1 19040
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1606120353
transform 1 0 9568 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A
timestamp 1606120353
transform 1 0 10488 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_90
timestamp 1606120353
transform 1 0 9384 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_31_93
timestamp 1606120353
transform 1 0 9660 0 1 19040
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_31_101
timestamp 1606120353
transform 1 0 10396 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__a211o_4  _0937_
timestamp 1606120353
transform 1 0 12236 0 1 19040
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__C1
timestamp 1606120353
transform 1 0 12052 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A2
timestamp 1606120353
transform 1 0 11684 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1606120353
transform 1 0 11500 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_117
timestamp 1606120353
transform 1 0 11868 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_135
timestamp 1606120353
transform 1 0 13524 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A2
timestamp 1606120353
transform 1 0 13708 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1606120353
transform 1 0 13892 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A2
timestamp 1606120353
transform 1 0 14076 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_31_143
timestamp 1606120353
transform 1 0 14260 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__B1
timestamp 1606120353
transform 1 0 14536 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_148
timestamp 1606120353
transform 1 0 14720 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A2
timestamp 1606120353
transform 1 0 14904 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_31_152
timestamp 1606120353
transform 1 0 15088 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1606120353
transform 1 0 15180 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _1000_
timestamp 1606120353
transform 1 0 15272 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__o21a_4  _1063_
timestamp 1606120353
transform 1 0 16744 0 1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__A
timestamp 1606120353
transform 1 0 15732 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__A2
timestamp 1606120353
transform 1 0 16560 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__B1
timestamp 1606120353
transform 1 0 16192 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_157
timestamp 1606120353
transform 1 0 15548 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_31_161
timestamp 1606120353
transform 1 0 15916 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1606120353
transform 1 0 16376 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606120353
transform -1 0 18860 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_31_182
timestamp 1606120353
transform 1 0 17848 0 1 19040
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1253_
timestamp 1606120353
transform 1 0 3128 0 -1 20128
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606120353
transform 1 0 1104 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__CLK
timestamp 1606120353
transform 1 0 1564 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1606120353
transform 1 0 1380 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_32_7
timestamp 1606120353
transform 1 0 1748 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_32_19
timestamp 1606120353
transform 1 0 2852 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__A
timestamp 1606120353
transform 1 0 5152 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_32_41
timestamp 1606120353
transform 1 0 4876 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__and2_4  _0694_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 6808 0 -1 20128
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1606120353
transform 1 0 6716 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_clk
timestamp 1606120353
transform 1 0 6440 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__C
timestamp 1606120353
transform 1 0 6256 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_32_46
timestamp 1606120353
transform 1 0 5336 0 -1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_32_54
timestamp 1606120353
transform 1 0 6072 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__B
timestamp 1606120353
transform 1 0 7636 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_69
timestamp 1606120353
transform 1 0 7452 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_32_73
timestamp 1606120353
transform 1 0 7820 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1606120353
transform 1 0 8924 0 -1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__CLK
timestamp 1606120353
transform 1 0 9844 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1606120353
transform 1 0 9660 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1606120353
transform 1 0 10028 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_32_109
timestamp 1606120353
transform 1 0 11132 0 -1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__a21bo_4  _1008_
timestamp 1606120353
transform 1 0 12420 0 -1 20128
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1606120353
transform 1 0 12328 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A1
timestamp 1606120353
transform 1 0 12144 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_32_117
timestamp 1606120353
transform 1 0 11868 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__a21o_4  _1007_
timestamp 1606120353
transform 1 0 14904 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__A1
timestamp 1606120353
transform 1 0 13800 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A1
timestamp 1606120353
transform 1 0 14168 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A1
timestamp 1606120353
transform 1 0 14720 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_136
timestamp 1606120353
transform 1 0 13616 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_140
timestamp 1606120353
transform 1 0 13984 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_32_144
timestamp 1606120353
transform 1 0 14352 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A2
timestamp 1606120353
transform 1 0 16192 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__A1
timestamp 1606120353
transform 1 0 16744 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__B1
timestamp 1606120353
transform 1 0 17112 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_162
timestamp 1606120353
transform 1 0 16008 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_32_166
timestamp 1606120353
transform 1 0 16376 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_32_172
timestamp 1606120353
transform 1 0 16928 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_176
timestamp 1606120353
transform 1 0 17296 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606120353
transform -1 0 18860 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1606120353
transform 1 0 17940 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A2
timestamp 1606120353
transform 1 0 17480 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_32_180
timestamp 1606120353
transform 1 0 17664 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_32_184
timestamp 1606120353
transform 1 0 18032 0 -1 20128
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_33_11
timestamp 1606120353
transform 1 0 2116 0 1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_33_7
timestamp 1606120353
transform 1 0 1748 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1606120353
transform 1 0 1380 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__CLK
timestamp 1606120353
transform 1 0 1932 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__D
timestamp 1606120353
transform 1 0 1564 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1606120353
transform 1 0 1104 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1606120353
transform 1 0 1104 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_34_22
timestamp 1606120353
transform 1 0 3128 0 -1 21216
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILLER_33_19
timestamp 1606120353
transform 1 0 2852 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_clk_A
timestamp 1606120353
transform 1 0 3128 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1255_
timestamp 1606120353
transform 1 0 1380 0 -1 21216
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_2  FILLER_34_33
timestamp 1606120353
transform 1 0 4140 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_24
timestamp 1606120353
transform 1 0 3312 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_clk_A
timestamp 1606120353
transform 1 0 3680 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__D
timestamp 1606120353
transform 1 0 3496 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_clk
timestamp 1606120353
transform 1 0 3680 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_clk
timestamp 1606120353
transform 1 0 3864 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1606120353
transform 1 0 3956 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_34_43
timestamp 1606120353
transform 1 0 5060 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_34_37
timestamp 1606120353
transform 1 0 4508 0 -1 21216
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__CLK
timestamp 1606120353
transform 1 0 4324 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0569_
timestamp 1606120353
transform 1 0 5152 0 -1 21216
box 0 -48 828 592
use sky130_fd_sc_hd__dfxtp_4  _1218_
timestamp 1606120353
transform 1 0 4048 0 1 20128
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_2  FILLER_34_53
timestamp 1606120353
transform 1 0 5980 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_55
timestamp 1606120353
transform 1 0 6164 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_51
timestamp 1606120353
transform 1 0 5796 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0563__A
timestamp 1606120353
transform 1 0 6164 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__A
timestamp 1606120353
transform 1 0 5980 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_57
timestamp 1606120353
transform 1 0 6348 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__A
timestamp 1606120353
transform 1 0 6532 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__C
timestamp 1606120353
transform 1 0 6348 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1606120353
transform 1 0 6716 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__nor3_4  _0653_
timestamp 1606120353
transform 1 0 6808 0 -1 21216
box 0 -48 1196 592
use sky130_fd_sc_hd__nand3_4  _0564_
timestamp 1606120353
transform 1 0 6532 0 1 20128
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_34_75
timestamp 1606120353
transform 1 0 8004 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_73
timestamp 1606120353
transform 1 0 7820 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__B
timestamp 1606120353
transform 1 0 8004 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_34_79
timestamp 1606120353
transform 1 0 8372 0 -1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_33_84
timestamp 1606120353
transform 1 0 8832 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_77
timestamp 1606120353
transform 1 0 8188 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__B
timestamp 1606120353
transform 1 0 8188 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0568__A
timestamp 1606120353
transform 1 0 8372 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0654_
timestamp 1606120353
transform 1 0 8740 0 -1 21216
box 0 -48 828 592
use sky130_fd_sc_hd__buf_1  _0568_
timestamp 1606120353
transform 1 0 8556 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_33_88
timestamp 1606120353
transform 1 0 9200 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0654__A
timestamp 1606120353
transform 1 0 9016 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1256_
timestamp 1606120353
transform 1 0 9844 0 1 20128
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1606120353
transform 1 0 9568 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__D
timestamp 1606120353
transform 1 0 9384 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_93
timestamp 1606120353
transform 1 0 9660 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_34_92
timestamp 1606120353
transform 1 0 9568 0 -1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_34_104
timestamp 1606120353
transform 1 0 10672 0 -1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_34_116
timestamp 1606120353
transform 1 0 11776 0 -1 21216
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_33_118
timestamp 1606120353
transform 1 0 11960 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_114
timestamp 1606120353
transform 1 0 11592 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__C
timestamp 1606120353
transform 1 0 11776 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_34_127
timestamp 1606120353
transform 1 0 12788 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_34_123
timestamp 1606120353
transform 1 0 12420 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A
timestamp 1606120353
transform 1 0 12604 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__B
timestamp 1606120353
transform 1 0 12144 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1606120353
transform 1 0 12328 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0936_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 12328 0 1 20128
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_33_131
timestamp 1606120353
transform 1 0 13156 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__C
timestamp 1606120353
transform 1 0 13064 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0956_
timestamp 1606120353
transform 1 0 13248 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_34_139
timestamp 1606120353
transform 1 0 13892 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_135
timestamp 1606120353
transform 1 0 13524 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_33_139
timestamp 1606120353
transform 1 0 13892 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_33_135
timestamp 1606120353
transform 1 0 13524 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__D
timestamp 1606120353
transform 1 0 13708 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__B
timestamp 1606120353
transform 1 0 14076 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__A
timestamp 1606120353
transform 1 0 13708 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A
timestamp 1606120353
transform 1 0 13340 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_143
timestamp 1606120353
transform 1 0 14260 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_149
timestamp 1606120353
transform 1 0 14812 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_145
timestamp 1606120353
transform 1 0 14444 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A
timestamp 1606120353
transform 1 0 14628 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _1035_
timestamp 1606120353
transform 1 0 14444 0 -1 21216
box 0 -48 828 592
use sky130_fd_sc_hd__buf_1  _0925_
timestamp 1606120353
transform 1 0 14168 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_34_154
timestamp 1606120353
transform 1 0 15272 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_154
timestamp 1606120353
transform 1 0 15272 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A
timestamp 1606120353
transform 1 0 14996 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1606120353
transform 1 0 15180 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_34_158
timestamp 1606120353
transform 1 0 15640 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_165
timestamp 1606120353
transform 1 0 16284 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_161
timestamp 1606120353
transform 1 0 15916 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__B1
timestamp 1606120353
transform 1 0 15456 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__B1
timestamp 1606120353
transform 1 0 15824 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A1
timestamp 1606120353
transform 1 0 15456 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A
timestamp 1606120353
transform 1 0 16100 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0916_
timestamp 1606120353
transform 1 0 15640 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_34_175
timestamp 1606120353
transform 1 0 17204 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A1
timestamp 1606120353
transform 1 0 16468 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1056_
timestamp 1606120353
transform 1 0 16652 0 1 20128
box 0 -48 1196 592
use sky130_fd_sc_hd__o21ai_4  _1053_
timestamp 1606120353
transform 1 0 16008 0 -1 21216
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1606120353
transform -1 0 18860 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1606120353
transform -1 0 18860 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1606120353
transform 1 0 17940 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A1
timestamp 1606120353
transform 1 0 17388 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A2
timestamp 1606120353
transform 1 0 17756 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_33_182
timestamp 1606120353
transform 1 0 17848 0 1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_34_179
timestamp 1606120353
transform 1 0 17572 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_34_184
timestamp 1606120353
transform 1 0 18032 0 -1 21216
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1606120353
transform 1 0 1104 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__D
timestamp 1606120353
transform 1 0 1840 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__CLK
timestamp 1606120353
transform 1 0 2208 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1606120353
transform 1 0 1380 0 1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_35_7
timestamp 1606120353
transform 1 0 1748 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_35_10
timestamp 1606120353
transform 1 0 2024 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_35_14
timestamp 1606120353
transform 1 0 2392 0 1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1606120353
transform 1 0 3956 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_clk_A
timestamp 1606120353
transform 1 0 5152 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_clk_A
timestamp 1606120353
transform 1 0 4784 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_35_26
timestamp 1606120353
transform 1 0 3496 0 1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_35_30
timestamp 1606120353
transform 1 0 3864 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_35_32
timestamp 1606120353
transform 1 0 4048 0 1 21216
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_35_42
timestamp 1606120353
transform 1 0 4968 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0563_
timestamp 1606120353
transform 1 0 6624 0 1 21216
box 0 -48 828 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_clk
timestamp 1606120353
transform 1 0 6348 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__A
timestamp 1606120353
transform 1 0 5704 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0570__A
timestamp 1606120353
transform 1 0 6164 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_35_46
timestamp 1606120353
transform 1 0 5336 0 1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_35_52
timestamp 1606120353
transform 1 0 5888 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0565_
timestamp 1606120353
transform 1 0 8188 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0565__A
timestamp 1606120353
transform 1 0 8648 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__C
timestamp 1606120353
transform 1 0 7636 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__A
timestamp 1606120353
transform 1 0 8004 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_69
timestamp 1606120353
transform 1 0 7452 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_73
timestamp 1606120353
transform 1 0 7820 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_80
timestamp 1606120353
transform 1 0 8464 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_35_84
timestamp 1606120353
transform 1 0 8832 0 1 21216
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1606120353
transform 1 0 9568 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__A2
timestamp 1606120353
transform 1 0 9844 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__B1
timestamp 1606120353
transform 1 0 10212 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__A1
timestamp 1606120353
transform 1 0 9384 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_93
timestamp 1606120353
transform 1 0 9660 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_97
timestamp 1606120353
transform 1 0 10028 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_35_101
timestamp 1606120353
transform 1 0 10396 0 1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_35_113
timestamp 1606120353
transform 1 0 11500 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0966_
timestamp 1606120353
transform 1 0 11592 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_35_117
timestamp 1606120353
transform 1 0 11868 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A
timestamp 1606120353
transform 1 0 12052 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_121
timestamp 1606120353
transform 1 0 12236 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A1
timestamp 1606120353
transform 1 0 12420 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0960_
timestamp 1606120353
transform 1 0 12604 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_35_128
timestamp 1606120353
transform 1 0 12880 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__A
timestamp 1606120353
transform 1 0 13064 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_132
timestamp 1606120353
transform 1 0 13248 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__or3_4  _1036_
timestamp 1606120353
transform 1 0 13616 0 1 21216
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1606120353
transform 1 0 15180 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A2
timestamp 1606120353
transform 1 0 14628 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__A
timestamp 1606120353
transform 1 0 13432 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__B1
timestamp 1606120353
transform 1 0 14996 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_145
timestamp 1606120353
transform 1 0 14444 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_149
timestamp 1606120353
transform 1 0 14812 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_35_154
timestamp 1606120353
transform 1 0 15272 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _1050_
timestamp 1606120353
transform 1 0 15732 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__o21a_4  _1052_
timestamp 1606120353
transform 1 0 16744 0 1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A
timestamp 1606120353
transform 1 0 16192 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__B1
timestamp 1606120353
transform 1 0 16560 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A1
timestamp 1606120353
transform 1 0 15548 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_162
timestamp 1606120353
transform 1 0 16008 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1606120353
transform 1 0 16376 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1606120353
transform -1 0 18860 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A2
timestamp 1606120353
transform 1 0 18032 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_182
timestamp 1606120353
transform 1 0 17848 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_35_186
timestamp 1606120353
transform 1 0 18216 0 1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1257_
timestamp 1606120353
transform 1 0 1840 0 -1 22304
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1606120353
transform 1 0 1104 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1606120353
transform 1 0 1380 0 -1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_36_7
timestamp 1606120353
transform 1 0 1748 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_clk
timestamp 1606120353
transform 1 0 5152 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_clk_A
timestamp 1606120353
transform 1 0 4784 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__CLK
timestamp 1606120353
transform 1 0 4416 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__CLK
timestamp 1606120353
transform 1 0 3956 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1606120353
transform 1 0 3588 0 -1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_36_33
timestamp 1606120353
transform 1 0 4140 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_36_38
timestamp 1606120353
transform 1 0 4600 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_42
timestamp 1606120353
transform 1 0 4968 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_36_47
timestamp 1606120353
transform 1 0 5428 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0695_
timestamp 1606120353
transform 1 0 5704 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_36_53
timestamp 1606120353
transform 1 0 5980 0 -1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_36_60
timestamp 1606120353
transform 1 0 6624 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_36_57
timestamp 1606120353
transform 1 0 6348 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__D1
timestamp 1606120353
transform 1 0 6440 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_62
timestamp 1606120353
transform 1 0 6808 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__A
timestamp 1606120353
transform 1 0 6992 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1606120353
transform 1 0 6716 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_36_66
timestamp 1606120353
transform 1 0 7176 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _0651_
timestamp 1606120353
transform 1 0 7360 0 -1 22304
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__A
timestamp 1606120353
transform 1 0 8372 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_77
timestamp 1606120353
transform 1 0 8188 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_36_81
timestamp 1606120353
transform 1 0 8556 0 -1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__o21a_4  _0655_
timestamp 1606120353
transform 1 0 9660 0 -1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A2
timestamp 1606120353
transform 1 0 9476 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_89
timestamp 1606120353
transform 1 0 9292 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_36_105
timestamp 1606120353
transform 1 0 10764 0 -1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__buf_1  _0901_
timestamp 1606120353
transform 1 0 12880 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1606120353
transform 1 0 12328 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_36_117
timestamp 1606120353
transform 1 0 11868 0 -1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_36_121
timestamp 1606120353
transform 1 0 12236 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_36_123
timestamp 1606120353
transform 1 0 12420 0 -1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_36_127
timestamp 1606120353
transform 1 0 12788 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_36_131
timestamp 1606120353
transform 1 0 13156 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _1009_
timestamp 1606120353
transform 1 0 14168 0 -1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__B1
timestamp 1606120353
transform 1 0 13892 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__B1
timestamp 1606120353
transform 1 0 13340 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_36_135
timestamp 1606120353
transform 1 0 13524 0 -1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_36_141
timestamp 1606120353
transform 1 0 14076 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_36_154
timestamp 1606120353
transform 1 0 15272 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1066_
timestamp 1606120353
transform 1 0 16008 0 -1 22304
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__C1
timestamp 1606120353
transform 1 0 15824 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A2
timestamp 1606120353
transform 1 0 15456 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_158
timestamp 1606120353
transform 1 0 15640 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_175
timestamp 1606120353
transform 1 0 17204 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1606120353
transform -1 0 18860 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1606120353
transform 1 0 17940 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__A1
timestamp 1606120353
transform 1 0 17388 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_36_179
timestamp 1606120353
transform 1 0 17572 0 -1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_36_184
timestamp 1606120353
transform 1 0 18032 0 -1 22304
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1606120353
transform 1 0 1104 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1606120353
transform 1 0 1380 0 1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1606120353
transform 1 0 2484 0 1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_37_32
timestamp 1606120353
transform 1 0 4048 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_37_30
timestamp 1606120353
transform 1 0 3864 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_37_27
timestamp 1606120353
transform 1 0 3588 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_clk_A
timestamp 1606120353
transform 1 0 3680 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1606120353
transform 1 0 3956 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_37_43
timestamp 1606120353
transform 1 0 5060 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_37_36
timestamp 1606120353
transform 1 0 4416 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__D
timestamp 1606120353
transform 1 0 4600 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__D
timestamp 1606120353
transform 1 0 4232 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_clk
timestamp 1606120353
transform 1 0 4784 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1211_
timestamp 1606120353
transform 1 0 5152 0 1 22304
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0570__B
timestamp 1606120353
transform 1 0 7084 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_63
timestamp 1606120353
transform 1 0 6900 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__nand2_4  _0680_
timestamp 1606120353
transform 1 0 8004 0 1 22304
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__B
timestamp 1606120353
transform 1 0 7820 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0570__C
timestamp 1606120353
transform 1 0 7452 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__A2
timestamp 1606120353
transform 1 0 9016 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_67
timestamp 1606120353
transform 1 0 7268 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_71
timestamp 1606120353
transform 1 0 7636 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_84
timestamp 1606120353
transform 1 0 8832 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_88
timestamp 1606120353
transform 1 0 9200 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__a21oi_4  _0681_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 9660 0 1 22304
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1606120353
transform 1 0 9568 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__A1
timestamp 1606120353
transform 1 0 9384 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__B1
timestamp 1606120353
transform 1 0 11040 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_106
timestamp 1606120353
transform 1 0 10856 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1606120353
transform 1 0 11224 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0915_
timestamp 1606120353
transform 1 0 12328 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A1
timestamp 1606120353
transform 1 0 11408 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A
timestamp 1606120353
transform 1 0 12788 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A2
timestamp 1606120353
transform 1 0 13156 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A
timestamp 1606120353
transform 1 0 12144 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_37_114
timestamp 1606120353
transform 1 0 11592 0 1 22304
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_37_125
timestamp 1606120353
transform 1 0 12604 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_129
timestamp 1606120353
transform 1 0 12972 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0924_
timestamp 1606120353
transform 1 0 15272 0 1 22304
box 0 -48 644 592
use sky130_fd_sc_hd__a21o_4  _1011_
timestamp 1606120353
transform 1 0 13340 0 1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1606120353
transform 1 0 15180 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A2
timestamp 1606120353
transform 1 0 14628 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__B
timestamp 1606120353
transform 1 0 14996 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_145
timestamp 1606120353
transform 1 0 14444 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_149
timestamp 1606120353
transform 1 0 14812 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1064_
timestamp 1606120353
transform 1 0 16652 0 1 22304
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A
timestamp 1606120353
transform 1 0 16100 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__B1
timestamp 1606120353
transform 1 0 16468 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_161
timestamp 1606120353
transform 1 0 15916 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_165
timestamp 1606120353
transform 1 0 16284 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1606120353
transform -1 0 18860 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__A2
timestamp 1606120353
transform 1 0 18032 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__B1
timestamp 1606120353
transform 1 0 18400 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_182
timestamp 1606120353
transform 1 0 17848 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_186
timestamp 1606120353
transform 1 0 18216 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1606120353
transform 1 0 1380 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__D
timestamp 1606120353
transform 1 0 1564 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1606120353
transform 1 0 1104 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_38_11
timestamp 1606120353
transform 1 0 2116 0 -1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_38_7
timestamp 1606120353
transform 1 0 1748 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__CLK
timestamp 1606120353
transform 1 0 1932 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_17
timestamp 1606120353
transform 1 0 2668 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__D
timestamp 1606120353
transform 1 0 2484 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1606120353
transform 1 0 3036 0 -1 23392
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__CLK
timestamp 1606120353
transform 1 0 2852 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1219_
timestamp 1606120353
transform 1 0 3956 0 -1 23392
box 0 -48 1748 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_clk
timestamp 1606120353
transform 1 0 3680 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1606120353
transform 1 0 3588 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__nor3_4  _0570_
timestamp 1606120353
transform 1 0 6808 0 -1 23392
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1606120353
transform 1 0 6716 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__A
timestamp 1606120353
transform 1 0 5888 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A1
timestamp 1606120353
transform 1 0 6440 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_50
timestamp 1606120353
transform 1 0 5704 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_38_54
timestamp 1606120353
transform 1 0 6072 0 -1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_38_60
timestamp 1606120353
transform 1 0 6624 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__A2
timestamp 1606120353
transform 1 0 8372 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__A1
timestamp 1606120353
transform 1 0 8740 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_38_75
timestamp 1606120353
transform 1 0 8004 0 -1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_38_81
timestamp 1606120353
transform 1 0 8556 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_38_85
timestamp 1606120353
transform 1 0 8924 0 -1 23392
box 0 -48 552 592
use sky130_fd_sc_hd__o21ai_4  _0652_
timestamp 1606120353
transform 1 0 9660 0 -1 23392
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__B
timestamp 1606120353
transform 1 0 11040 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__B1
timestamp 1606120353
transform 1 0 9476 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_106
timestamp 1606120353
transform 1 0 10856 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_38_110
timestamp 1606120353
transform 1 0 11224 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__buf_1  _0900_
timestamp 1606120353
transform 1 0 12420 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1606120353
transform 1 0 12328 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A1
timestamp 1606120353
transform 1 0 13248 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A1
timestamp 1606120353
transform 1 0 12880 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_126
timestamp 1606120353
transform 1 0 12696 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_130
timestamp 1606120353
transform 1 0 13064 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _1010_
timestamp 1606120353
transform 1 0 13892 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__B
timestamp 1606120353
transform 1 0 13616 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_134
timestamp 1606120353
transform 1 0 13432 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_38_138
timestamp 1606120353
transform 1 0 13800 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_38_151
timestamp 1606120353
transform 1 0 14996 0 -1 23392
box 0 -48 736 592
use sky130_fd_sc_hd__a211o_4  _1041_
timestamp 1606120353
transform 1 0 15916 0 -1 23392
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A1
timestamp 1606120353
transform 1 0 15732 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_175
timestamp 1606120353
transform 1 0 17204 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1606120353
transform -1 0 18860 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1606120353
transform 1 0 17940 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A1
timestamp 1606120353
transform 1 0 17388 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_38_179
timestamp 1606120353
transform 1 0 17572 0 -1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_38_184
timestamp 1606120353
transform 1 0 18032 0 -1 23392
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1258_
timestamp 1606120353
transform 1 0 1472 0 1 23392
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1259_
timestamp 1606120353
transform 1 0 2484 0 -1 24480
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1606120353
transform 1 0 1104 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1606120353
transform 1 0 1104 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__D
timestamp 1606120353
transform 1 0 1564 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_39_3
timestamp 1606120353
transform 1 0 1380 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1606120353
transform 1 0 1380 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_40_7
timestamp 1606120353
transform 1 0 1748 0 -1 24480
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_39_23
timestamp 1606120353
transform 1 0 3220 0 1 23392
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1606120353
transform 1 0 3956 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_40_38
timestamp 1606120353
transform 1 0 4600 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_34
timestamp 1606120353
transform 1 0 4232 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_37
timestamp 1606120353
transform 1 0 4508 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_39_32
timestamp 1606120353
transform 1 0 4048 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_clk_A
timestamp 1606120353
transform 1 0 4416 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__B1
timestamp 1606120353
transform 1 0 4784 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__A
timestamp 1606120353
transform 1 0 4324 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__C
timestamp 1606120353
transform 1 0 4692 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_clk
timestamp 1606120353
transform 1 0 4968 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__and4_4  _0691_
timestamp 1606120353
transform 1 0 4876 0 1 23392
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_40_53
timestamp 1606120353
transform 1 0 5980 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_40_49
timestamp 1606120353
transform 1 0 5612 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_40_45
timestamp 1606120353
transform 1 0 5244 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1606120353
transform 1 0 6072 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_50
timestamp 1606120353
transform 1 0 5704 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A2
timestamp 1606120353
transform 1 0 6164 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__B
timestamp 1606120353
transform 1 0 5428 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__D
timestamp 1606120353
transform 1 0 5888 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0687_
timestamp 1606120353
transform 1 0 5704 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1606120353
transform 1 0 6348 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A2
timestamp 1606120353
transform 1 0 6532 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__C1
timestamp 1606120353
transform 1 0 6256 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1606120353
transform 1 0 6716 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _0689_
timestamp 1606120353
transform 1 0 6808 0 -1 24480
box 0 -48 828 592
use sky130_fd_sc_hd__a2111oi_4  _0688_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 6440 0 1 23392
box 0 -48 2024 592
use sky130_fd_sc_hd__fill_2  FILLER_40_75
timestamp 1606120353
transform 1 0 8004 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_71
timestamp 1606120353
transform 1 0 7636 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__A
timestamp 1606120353
transform 1 0 8188 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__C
timestamp 1606120353
transform 1 0 7820 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_88
timestamp 1606120353
transform 1 0 9200 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_84
timestamp 1606120353
transform 1 0 8832 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_80
timestamp 1606120353
transform 1 0 8464 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__B1_N
timestamp 1606120353
transform 1 0 9016 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__B1_N
timestamp 1606120353
transform 1 0 8648 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__a21boi_4  _0725_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 8372 0 -1 24480
box 0 -48 1380 592
use sky130_fd_sc_hd__fill_2  FILLER_40_98
timestamp 1606120353
transform 1 0 10120 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_94
timestamp 1606120353
transform 1 0 9752 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__A2
timestamp 1606120353
transform 1 0 9936 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__A1
timestamp 1606120353
transform 1 0 9384 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1606120353
transform 1 0 9568 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_39_108
timestamp 1606120353
transform 1 0 11040 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A
timestamp 1606120353
transform 1 0 11224 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__A1
timestamp 1606120353
transform 1 0 10304 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__nand2_4  _0679_
timestamp 1606120353
transform 1 0 10488 0 -1 24480
box 0 -48 828 592
use sky130_fd_sc_hd__a21boi_4  _0678_
timestamp 1606120353
transform 1 0 9660 0 1 23392
box 0 -48 1380 592
use sky130_fd_sc_hd__decap_6  FILLER_40_115
timestamp 1606120353
transform 1 0 11684 0 -1 24480
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_40_111
timestamp 1606120353
transform 1 0 11316 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_112
timestamp 1606120353
transform 1 0 11408 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__CLK
timestamp 1606120353
transform 1 0 11500 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__A
timestamp 1606120353
transform 1 0 11592 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0907_
timestamp 1606120353
transform 1 0 11776 0 1 23392
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILLER_40_123
timestamp 1606120353
transform 1 0 12420 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_40_121
timestamp 1606120353
transform 1 0 12236 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_39_125
timestamp 1606120353
transform 1 0 12604 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__A
timestamp 1606120353
transform 1 0 12788 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1606120353
transform 1 0 12328 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _1042_
timestamp 1606120353
transform 1 0 12696 0 -1 24480
box 0 -48 828 592
use sky130_fd_sc_hd__decap_4  FILLER_39_129
timestamp 1606120353
transform 1 0 12972 0 1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_40_139
timestamp 1606120353
transform 1 0 13892 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_135
timestamp 1606120353
transform 1 0 13524 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_39_133
timestamp 1606120353
transform 1 0 13340 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__B
timestamp 1606120353
transform 1 0 14076 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__A
timestamp 1606120353
transform 1 0 13708 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__A
timestamp 1606120353
transform 1 0 13432 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__nand2_4  _0941_
timestamp 1606120353
transform 1 0 13616 0 1 23392
box 0 -48 828 592
use sky130_fd_sc_hd__inv_8  _0920_
timestamp 1606120353
transform 1 0 14260 0 -1 24480
box 0 -48 828 592
use sky130_fd_sc_hd__decap_4  FILLER_39_154
timestamp 1606120353
transform 1 0 15272 0 1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_39_149
timestamp 1606120353
transform 1 0 14812 0 1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_39_145
timestamp 1606120353
transform 1 0 14444 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A
timestamp 1606120353
transform 1 0 14628 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1606120353
transform 1 0 15180 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_40_152
timestamp 1606120353
transform 1 0 15088 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_40_164
timestamp 1606120353
transform 1 0 16192 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_162
timestamp 1606120353
transform 1 0 16008 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_39_158
timestamp 1606120353
transform 1 0 15640 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__A
timestamp 1606120353
transform 1 0 16192 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1034_
timestamp 1606120353
transform 1 0 15732 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_40_175
timestamp 1606120353
transform 1 0 17204 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1606120353
transform 1 0 16376 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A
timestamp 1606120353
transform 1 0 16560 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _1051_
timestamp 1606120353
transform 1 0 16376 0 -1 24480
box 0 -48 828 592
use sky130_fd_sc_hd__o21a_4  _1068_
timestamp 1606120353
transform 1 0 16744 0 1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1606120353
transform -1 0 18860 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1606120353
transform -1 0 18860 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1606120353
transform 1 0 17940 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A2
timestamp 1606120353
transform 1 0 17388 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__B1
timestamp 1606120353
transform 1 0 18032 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_182
timestamp 1606120353
transform 1 0 17848 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_39_186
timestamp 1606120353
transform 1 0 18216 0 1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_40_179
timestamp 1606120353
transform 1 0 17572 0 -1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_40_184
timestamp 1606120353
transform 1 0 18032 0 -1 24480
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1288_
timestamp 1606120353
transform 1 0 1380 0 1 24480
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1606120353
transform 1 0 1104 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_41_22
timestamp 1606120353
transform 1 0 3128 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1146_
timestamp 1606120353
transform 1 0 4048 0 1 24480
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1606120353
transform 1 0 3956 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A
timestamp 1606120353
transform 1 0 3772 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__D
timestamp 1606120353
transform 1 0 3404 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_27
timestamp 1606120353
transform 1 0 3588 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_clk
timestamp 1606120353
transform 1 0 6532 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__A
timestamp 1606120353
transform 1 0 5980 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A1
timestamp 1606120353
transform 1 0 6348 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_51
timestamp 1606120353
transform 1 0 5796 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_55
timestamp 1606120353
transform 1 0 6164 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_41_62
timestamp 1606120353
transform 1 0 6808 0 1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_41_66
timestamp 1606120353
transform 1 0 7176 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__nand3_4  _0686_
timestamp 1606120353
transform 1 0 7452 0 1 24480
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__B
timestamp 1606120353
transform 1 0 7268 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__A
timestamp 1606120353
transform 1 0 9016 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_41_83
timestamp 1606120353
transform 1 0 8740 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_41_88
timestamp 1606120353
transform 1 0 9200 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1177_
timestamp 1606120353
transform 1 0 10212 0 1 24480
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1606120353
transform 1 0 9568 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__D
timestamp 1606120353
transform 1 0 10028 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__A2
timestamp 1606120353
transform 1 0 9384 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_41_93
timestamp 1606120353
transform 1 0 9660 0 1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__A
timestamp 1606120353
transform 1 0 12420 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__B
timestamp 1606120353
transform 1 0 12788 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__C
timestamp 1606120353
transform 1 0 13156 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_41_118
timestamp 1606120353
transform 1 0 11960 0 1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_41_122
timestamp 1606120353
transform 1 0 12328 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_41_125
timestamp 1606120353
transform 1 0 12604 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_129
timestamp 1606120353
transform 1 0 12972 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _1025_
timestamp 1606120353
transform 1 0 13616 0 1 24480
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1606120353
transform 1 0 15180 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__B
timestamp 1606120353
transform 1 0 14996 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__A
timestamp 1606120353
transform 1 0 14628 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_41_133
timestamp 1606120353
transform 1 0 13340 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_41_145
timestamp 1606120353
transform 1 0 14444 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_149
timestamp 1606120353
transform 1 0 14812 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_154
timestamp 1606120353
transform 1 0 15272 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1040_
timestamp 1606120353
transform 1 0 15640 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _1069_
timestamp 1606120353
transform 1 0 16652 0 1 24480
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__C
timestamp 1606120353
transform 1 0 15456 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__A
timestamp 1606120353
transform 1 0 16100 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A1
timestamp 1606120353
transform 1 0 16468 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_161
timestamp 1606120353
transform 1 0 15916 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_165
timestamp 1606120353
transform 1 0 16284 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1606120353
transform -1 0 18860 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_41_182
timestamp 1606120353
transform 1 0 17848 0 1 24480
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1606120353
transform 1 0 1104 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__CLK
timestamp 1606120353
transform 1 0 1564 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1606120353
transform 1 0 1380 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_42_7
timestamp 1606120353
transform 1 0 1748 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_42_19
timestamp 1606120353
transform 1 0 2852 0 -1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _0753_
timestamp 1606120353
transform 1 0 4140 0 -1 25568
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A2
timestamp 1606120353
transform 1 0 3956 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__B
timestamp 1606120353
transform 1 0 3588 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__CLK
timestamp 1606120353
transform 1 0 3220 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_25
timestamp 1606120353
transform 1 0 3404 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1606120353
transform 1 0 3772 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_42_42
timestamp 1606120353
transform 1 0 4968 0 -1 25568
box 0 -48 736 592
use sky130_fd_sc_hd__o21ai_4  _0690_
timestamp 1606120353
transform 1 0 7084 0 -1 25568
box 0 -48 1196 592
use sky130_fd_sc_hd__buf_1  _0698_
timestamp 1606120353
transform 1 0 5704 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1606120353
transform 1 0 6716 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__B1
timestamp 1606120353
transform 1 0 6532 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_clk_A
timestamp 1606120353
transform 1 0 6164 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_53
timestamp 1606120353
transform 1 0 5980 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_57
timestamp 1606120353
transform 1 0 6348 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_42_62
timestamp 1606120353
transform 1 0 6808 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A2
timestamp 1606120353
transform 1 0 8556 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__B1
timestamp 1606120353
transform 1 0 8924 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_42_78
timestamp 1606120353
transform 1 0 8280 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_42_83
timestamp 1606120353
transform 1 0 8740 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_87
timestamp 1606120353
transform 1 0 9108 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__a21oi_4  _0650_
timestamp 1606120353
transform 1 0 10304 0 -1 25568
box 0 -48 1196 592
use sky130_fd_sc_hd__buf_1  _0905_
timestamp 1606120353
transform 1 0 9292 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A
timestamp 1606120353
transform 1 0 9752 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__B1
timestamp 1606120353
transform 1 0 10120 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_92
timestamp 1606120353
transform 1 0 9568 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_96
timestamp 1606120353
transform 1 0 9936 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__nor3_4  _0935_
timestamp 1606120353
transform 1 0 12420 0 -1 25568
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1606120353
transform 1 0 12328 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__D
timestamp 1606120353
transform 1 0 12144 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_42_113
timestamp 1606120353
transform 1 0 11500 0 -1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_42_119
timestamp 1606120353
transform 1 0 12052 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__nor3_4  _1027_
timestamp 1606120353
transform 1 0 15088 0 -1 25568
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__C
timestamp 1606120353
transform 1 0 13800 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_136
timestamp 1606120353
transform 1 0 13616 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_42_140
timestamp 1606120353
transform 1 0 13984 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A2
timestamp 1606120353
transform 1 0 16652 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__B1
timestamp 1606120353
transform 1 0 17020 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_42_165
timestamp 1606120353
transform 1 0 16284 0 -1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_42_171
timestamp 1606120353
transform 1 0 16836 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_175
timestamp 1606120353
transform 1 0 17204 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1606120353
transform -1 0 18860 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1606120353
transform 1 0 17940 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__B1
timestamp 1606120353
transform 1 0 17388 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_42_179
timestamp 1606120353
transform 1 0 17572 0 -1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_42_184
timestamp 1606120353
transform 1 0 18032 0 -1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1606120353
transform 1 0 1104 0 1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__D
timestamp 1606120353
transform 1 0 1564 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A
timestamp 1606120353
transform 1 0 2392 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__CLK
timestamp 1606120353
transform 1 0 1932 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1606120353
transform 1 0 1380 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_7
timestamp 1606120353
transform 1 0 1748 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_43_11
timestamp 1606120353
transform 1 0 2116 0 1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_43_16
timestamp 1606120353
transform 1 0 2576 0 1 25568
box 0 -48 736 592
use sky130_fd_sc_hd__nand2_4  _0754_
timestamp 1606120353
transform 1 0 4048 0 1 25568
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1606120353
transform 1 0 3956 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__B1
timestamp 1606120353
transform 1 0 5060 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A1
timestamp 1606120353
transform 1 0 3772 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A
timestamp 1606120353
transform 1 0 3404 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_43_24
timestamp 1606120353
transform 1 0 3312 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_43_27
timestamp 1606120353
transform 1 0 3588 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_41
timestamp 1606120353
transform 1 0 4876 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__a21oi_4  _0700_
timestamp 1606120353
transform 1 0 5612 0 1 25568
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0566__A
timestamp 1606120353
transform 1 0 6992 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A1
timestamp 1606120353
transform 1 0 5428 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_45
timestamp 1606120353
transform 1 0 5244 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_62
timestamp 1606120353
transform 1 0 6808 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_43_66
timestamp 1606120353
transform 1 0 7176 0 1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__a21o_4  _0726_
timestamp 1606120353
transform 1 0 7728 0 1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__B1
timestamp 1606120353
transform 1 0 7544 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A1
timestamp 1606120353
transform 1 0 9016 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_84
timestamp 1606120353
transform 1 0 8832 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_88
timestamp 1606120353
transform 1 0 9200 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__nand3_4  _0649_
timestamp 1606120353
transform 1 0 9752 0 1 25568
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1606120353
transform 1 0 9568 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__C
timestamp 1606120353
transform 1 0 9384 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_43_93
timestamp 1606120353
transform 1 0 9660 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_43_108
timestamp 1606120353
transform 1 0 11040 0 1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__nand4_4  _1104_
timestamp 1606120353
transform 1 0 12696 0 1 25568
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__B
timestamp 1606120353
transform 1 0 12512 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__C
timestamp 1606120353
transform 1 0 12144 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__B
timestamp 1606120353
transform 1 0 11776 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A
timestamp 1606120353
transform 1 0 11316 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_43_113
timestamp 1606120353
transform 1 0 11500 0 1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_43_118
timestamp 1606120353
transform 1 0 11960 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_122
timestamp 1606120353
transform 1 0 12328 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1606120353
transform 1 0 15180 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A
timestamp 1606120353
transform 1 0 14444 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_143
timestamp 1606120353
transform 1 0 14260 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_43_147
timestamp 1606120353
transform 1 0 14628 0 1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_43_154
timestamp 1606120353
transform 1 0 15272 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1043_
timestamp 1606120353
transform 1 0 15640 0 1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _1072_
timestamp 1606120353
transform 1 0 16652 0 1 25568
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__A
timestamp 1606120353
transform 1 0 16100 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A1
timestamp 1606120353
transform 1 0 16468 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A2
timestamp 1606120353
transform 1 0 15456 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_161
timestamp 1606120353
transform 1 0 15916 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_165
timestamp 1606120353
transform 1 0 16284 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1606120353
transform -1 0 18860 0 1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A1
timestamp 1606120353
transform 1 0 18032 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A2
timestamp 1606120353
transform 1 0 18400 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_182
timestamp 1606120353
transform 1 0 17848 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_186
timestamp 1606120353
transform 1 0 18216 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1273_
timestamp 1606120353
transform 1 0 1564 0 -1 26656
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1606120353
transform 1 0 1104 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1606120353
transform 1 0 1380 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0755_
timestamp 1606120353
transform 1 0 4048 0 -1 26656
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__B1
timestamp 1606120353
transform 1 0 3864 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__CLK
timestamp 1606120353
transform 1 0 3496 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_24
timestamp 1606120353
transform 1 0 3312 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_28
timestamp 1606120353
transform 1 0 3680 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0566_
timestamp 1606120353
transform 1 0 6992 0 -1 26656
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1606120353
transform 1 0 6716 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A2
timestamp 1606120353
transform 1 0 5612 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__A2
timestamp 1606120353
transform 1 0 6532 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_44_45
timestamp 1606120353
transform 1 0 5244 0 -1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_44_51
timestamp 1606120353
transform 1 0 5796 0 -1 26656
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_44_62
timestamp 1606120353
transform 1 0 6808 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__a21oi_4  _0727_
timestamp 1606120353
transform 1 0 8556 0 -1 26656
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A1
timestamp 1606120353
transform 1 0 8004 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A2
timestamp 1606120353
transform 1 0 8372 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_73
timestamp 1606120353
transform 1 0 7820 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_77
timestamp 1606120353
transform 1 0 8188 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__B
timestamp 1606120353
transform 1 0 9936 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A
timestamp 1606120353
transform 1 0 11132 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_94
timestamp 1606120353
transform 1 0 9752 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_44_98
timestamp 1606120353
transform 1 0 10120 0 -1 26656
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_44_106
timestamp 1606120353
transform 1 0 10856 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_44_118
timestamp 1606120353
transform 1 0 11960 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_114
timestamp 1606120353
transform 1 0 11592 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__C
timestamp 1606120353
transform 1 0 12144 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__B
timestamp 1606120353
transform 1 0 11776 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1070_
timestamp 1606120353
transform 1 0 11316 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_44_128
timestamp 1606120353
transform 1 0 12880 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_44_123
timestamp 1606120353
transform 1 0 12420 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__A
timestamp 1606120353
transform 1 0 12696 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1606120353
transform 1 0 12328 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__nand3_4  _1026_
timestamp 1606120353
transform 1 0 13156 0 -1 26656
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILLER_44_145
timestamp 1606120353
transform 1 0 14444 0 -1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__o21a_4  _1086_
timestamp 1606120353
transform 1 0 16100 0 -1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__B1
timestamp 1606120353
transform 1 0 15916 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_44_157
timestamp 1606120353
transform 1 0 15548 0 -1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_44_175
timestamp 1606120353
transform 1 0 17204 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1606120353
transform -1 0 18860 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1606120353
transform 1 0 17940 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A1
timestamp 1606120353
transform 1 0 17388 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_44_179
timestamp 1606120353
transform 1 0 17572 0 -1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_44_184
timestamp 1606120353
transform 1 0 18032 0 -1 26656
box 0 -48 552 592
use sky130_fd_sc_hd__nand2_4  _0706_
timestamp 1606120353
transform 1 0 2392 0 1 26656
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1606120353
transform 1 0 1104 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__D
timestamp 1606120353
transform 1 0 1656 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__B
timestamp 1606120353
transform 1 0 2208 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_45_3
timestamp 1606120353
transform 1 0 1380 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_45_8
timestamp 1606120353
transform 1 0 1840 0 1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1145_
timestamp 1606120353
transform 1 0 4048 0 1 26656
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1606120353
transform 1 0 3956 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__A2
timestamp 1606120353
transform 1 0 3772 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__A1
timestamp 1606120353
transform 1 0 3404 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_23
timestamp 1606120353
transform 1 0 3220 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_27
timestamp 1606120353
transform 1 0 3588 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0743_
timestamp 1606120353
transform 1 0 6992 0 1 26656
box 0 -48 1196 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_clk
timestamp 1606120353
transform 1 0 6532 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0572__A
timestamp 1606120353
transform 1 0 6348 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_clk_A
timestamp 1606120353
transform 1 0 5980 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_51
timestamp 1606120353
transform 1 0 5796 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_55
timestamp 1606120353
transform 1 0 6164 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_62
timestamp 1606120353
transform 1 0 6808 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0572__B
timestamp 1606120353
transform 1 0 8372 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__A1
timestamp 1606120353
transform 1 0 8740 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_77
timestamp 1606120353
transform 1 0 8188 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_81
timestamp 1606120353
transform 1 0 8556 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_45_85
timestamp 1606120353
transform 1 0 8924 0 1 26656
box 0 -48 552 592
use sky130_fd_sc_hd__buf_1  _0929_
timestamp 1606120353
transform 1 0 10672 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1606120353
transform 1 0 9568 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A
timestamp 1606120353
transform 1 0 11132 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__A
timestamp 1606120353
transform 1 0 10304 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_45_91
timestamp 1606120353
transform 1 0 9476 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_45_93
timestamp 1606120353
transform 1 0 9660 0 1 26656
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_45_99
timestamp 1606120353
transform 1 0 10212 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_45_102
timestamp 1606120353
transform 1 0 10488 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_107
timestamp 1606120353
transform 1 0 10948 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _0942_
timestamp 1606120353
transform 1 0 11684 0 1 26656
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A
timestamp 1606120353
transform 1 0 12696 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A
timestamp 1606120353
transform 1 0 11500 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__B
timestamp 1606120353
transform 1 0 13064 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_111
timestamp 1606120353
transform 1 0 11316 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_124
timestamp 1606120353
transform 1 0 12512 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_128
timestamp 1606120353
transform 1 0 12880 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_132
timestamp 1606120353
transform 1 0 13248 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _1037_
timestamp 1606120353
transform 1 0 13616 0 1 26656
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1606120353
transform 1 0 15180 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__A
timestamp 1606120353
transform 1 0 14628 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__B
timestamp 1606120353
transform 1 0 13432 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_145
timestamp 1606120353
transform 1 0 14444 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_45_149
timestamp 1606120353
transform 1 0 14812 0 1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_45_154
timestamp 1606120353
transform 1 0 15272 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1044_
timestamp 1606120353
transform 1 0 15640 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _1081_
timestamp 1606120353
transform 1 0 16652 0 1 26656
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__A
timestamp 1606120353
transform 1 0 16100 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__A1
timestamp 1606120353
transform 1 0 16468 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__A2
timestamp 1606120353
transform 1 0 15456 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_161
timestamp 1606120353
transform 1 0 15916 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_165
timestamp 1606120353
transform 1 0 16284 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1606120353
transform -1 0 18860 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A2
timestamp 1606120353
transform 1 0 18032 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__B1
timestamp 1606120353
transform 1 0 18400 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_182
timestamp 1606120353
transform 1 0 17848 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_186
timestamp 1606120353
transform 1 0 18216 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_11
timestamp 1606120353
transform 1 0 2116 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_7
timestamp 1606120353
transform 1 0 1748 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1606120353
transform 1 0 1380 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_46_3
timestamp 1606120353
transform 1 0 1380 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0517__A
timestamp 1606120353
transform 1 0 1932 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0517__B
timestamp 1606120353
transform 1 0 1564 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1606120353
transform 1 0 1104 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1606120353
transform 1 0 1104 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_47_15
timestamp 1606120353
transform 1 0 2484 0 1 27744
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__CLK
timestamp 1606120353
transform 1 0 2300 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1289_
timestamp 1606120353
transform 1 0 1656 0 -1 27744
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__D
timestamp 1606120353
transform 1 0 3588 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_clk_A
timestamp 1606120353
transform 1 0 3404 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_25
timestamp 1606120353
transform 1 0 3404 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_23
timestamp 1606120353
transform 1 0 3220 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_27
timestamp 1606120353
transform 1 0 3588 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1606120353
transform 1 0 3956 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__A
timestamp 1606120353
transform 1 0 3772 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__B1
timestamp 1606120353
transform 1 0 3956 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1606120353
transform 1 0 3772 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0701_
timestamp 1606120353
transform 1 0 4048 0 1 27744
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILLER_47_41
timestamp 1606120353
transform 1 0 4876 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0571__A
timestamp 1606120353
transform 1 0 5152 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0707_
timestamp 1606120353
transform 1 0 4140 0 -1 27744
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_3  FILLER_47_46
timestamp 1606120353
transform 1 0 5336 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_46_55
timestamp 1606120353
transform 1 0 6164 0 -1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_46_51
timestamp 1606120353
transform 1 0 5796 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_46_46
timestamp 1606120353
transform 1 0 5336 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A1
timestamp 1606120353
transform 1 0 5980 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__B1
timestamp 1606120353
transform 1 0 5612 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_47_62
timestamp 1606120353
transform 1 0 6808 0 1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_46_66
timestamp 1606120353
transform 1 0 7176 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_46_62
timestamp 1606120353
transform 1 0 6808 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__B1
timestamp 1606120353
transform 1 0 6532 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__A
timestamp 1606120353
transform 1 0 6992 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__A2
timestamp 1606120353
transform 1 0 7176 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1606120353
transform 1 0 6716 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__a21oi_4  _0752_
timestamp 1606120353
transform 1 0 5612 0 1 27744
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_47_68
timestamp 1606120353
transform 1 0 7360 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_76
timestamp 1606120353
transform 1 0 8096 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__A1
timestamp 1606120353
transform 1 0 7544 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__nand2_4  _0572_
timestamp 1606120353
transform 1 0 7268 0 -1 27744
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_47_88
timestamp 1606120353
transform 1 0 9200 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_84
timestamp 1606120353
transform 1 0 8832 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_80
timestamp 1606120353
transform 1 0 8464 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A2
timestamp 1606120353
transform 1 0 8648 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__B1
timestamp 1606120353
transform 1 0 9016 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__B1
timestamp 1606120353
transform 1 0 8280 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_46_84
timestamp 1606120353
transform 1 0 8832 0 -1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__o21a_4  _0741_
timestamp 1606120353
transform 1 0 7728 0 1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_47_93
timestamp 1606120353
transform 1 0 9660 0 1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_46_96
timestamp 1606120353
transform 1 0 9936 0 -1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A1
timestamp 1606120353
transform 1 0 9384 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1606120353
transform 1 0 9568 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_47_104
timestamp 1606120353
transform 1 0 10672 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_47_100
timestamp 1606120353
transform 1 0 10304 0 1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_47_97
timestamp 1606120353
transform 1 0 10028 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_46_103
timestamp 1606120353
transform 1 0 10580 0 -1 27744
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0523__A
timestamp 1606120353
transform 1 0 10120 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0943_
timestamp 1606120353
transform 1 0 10304 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_47_107
timestamp 1606120353
transform 1 0 10948 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__A
timestamp 1606120353
transform 1 0 10764 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A
timestamp 1606120353
transform 1 0 11132 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_120
timestamp 1606120353
transform 1 0 12144 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_118
timestamp 1606120353
transform 1 0 11960 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_114
timestamp 1606120353
transform 1 0 11592 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__A
timestamp 1606120353
transform 1 0 11776 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__D1
timestamp 1606120353
transform 1 0 12144 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0918_
timestamp 1606120353
transform 1 0 11316 0 1 27744
box 0 -48 828 592
use sky130_fd_sc_hd__buf_1  _0902_
timestamp 1606120353
transform 1 0 11316 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_47_124
timestamp 1606120353
transform 1 0 12512 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_46_123
timestamp 1606120353
transform 1 0 12420 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__B
timestamp 1606120353
transform 1 0 12328 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__A1
timestamp 1606120353
transform 1 0 12696 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1606120353
transform 1 0 12328 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _0928_
timestamp 1606120353
transform 1 0 12512 0 -1 27744
box 0 -48 828 592
use sky130_fd_sc_hd__a2111o_4  _1032_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 12880 0 1 27744
box 0 -48 1564 592
use sky130_fd_sc_hd__fill_2  FILLER_46_137
timestamp 1606120353
transform 1 0 13708 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_133
timestamp 1606120353
transform 1 0 13340 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A
timestamp 1606120353
transform 1 0 13892 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__C1
timestamp 1606120353
transform 1 0 13524 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0944_
timestamp 1606120353
transform 1 0 14076 0 -1 27744
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_47_149
timestamp 1606120353
transform 1 0 14812 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_145
timestamp 1606120353
transform 1 0 14444 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_46_150
timestamp 1606120353
transform 1 0 14904 0 -1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__B1
timestamp 1606120353
transform 1 0 14628 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B
timestamp 1606120353
transform 1 0 15272 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A
timestamp 1606120353
transform 1 0 14996 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1606120353
transform 1 0 15180 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _1033_
timestamp 1606120353
transform 1 0 15272 0 1 27744
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_47_165
timestamp 1606120353
transform 1 0 16284 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_161
timestamp 1606120353
transform 1 0 15916 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_46_160
timestamp 1606120353
transform 1 0 15824 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_46_156
timestamp 1606120353
transform 1 0 15456 0 -1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__B1
timestamp 1606120353
transform 1 0 15916 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A
timestamp 1606120353
transform 1 0 16100 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_175
timestamp 1606120353
transform 1 0 17204 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__A1
timestamp 1606120353
transform 1 0 16468 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1084_
timestamp 1606120353
transform 1 0 16652 0 1 27744
box 0 -48 1196 592
use sky130_fd_sc_hd__o21a_4  _1080_
timestamp 1606120353
transform 1 0 16100 0 -1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_47_182
timestamp 1606120353
transform 1 0 17848 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_179
timestamp 1606120353
transform 1 0 17572 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__B1
timestamp 1606120353
transform 1 0 17756 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__A1
timestamp 1606120353
transform 1 0 17388 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_47_186
timestamp 1606120353
transform 1 0 18216 0 1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_46_184
timestamp 1606120353
transform 1 0 18032 0 -1 27744
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__A2
timestamp 1606120353
transform 1 0 18032 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1606120353
transform 1 0 17940 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1606120353
transform -1 0 18860 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1606120353
transform -1 0 18860 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__or2_4  _0517_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 1380 0 -1 28832
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1606120353
transform 1 0 1104 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__D
timestamp 1606120353
transform 1 0 2208 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__CLK
timestamp 1606120353
transform 1 0 2576 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_10
timestamp 1606120353
transform 1 0 2024 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_14
timestamp 1606120353
transform 1 0 2392 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_48_18
timestamp 1606120353
transform 1 0 2760 0 -1 28832
box 0 -48 552 592
use sky130_fd_sc_hd__inv_8  _0571_
timestamp 1606120353
transform 1 0 5152 0 -1 28832
box 0 -48 828 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_clk
timestamp 1606120353
transform 1 0 3404 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_clk_A
timestamp 1606120353
transform 1 0 4508 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_48_24
timestamp 1606120353
transform 1 0 3312 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_48_28
timestamp 1606120353
transform 1 0 3680 0 -1 28832
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_48_36
timestamp 1606120353
transform 1 0 4416 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_48_39
timestamp 1606120353
transform 1 0 4692 0 -1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_48_43
timestamp 1606120353
transform 1 0 5060 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0742_
timestamp 1606120353
transform 1 0 6900 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1606120353
transform 1 0 6716 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A2
timestamp 1606120353
transform 1 0 6164 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_53
timestamp 1606120353
transform 1 0 5980 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_48_57
timestamp 1606120353
transform 1 0 6348 0 -1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_48_62
timestamp 1606120353
transform 1 0 6808 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_48_66
timestamp 1606120353
transform 1 0 7176 0 -1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__o21ai_4  _0567_
timestamp 1606120353
transform 1 0 7912 0 -1 28832
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__C
timestamp 1606120353
transform 1 0 7636 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_48_70
timestamp 1606120353
transform 1 0 7544 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_48_73
timestamp 1606120353
transform 1 0 7820 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_48_87
timestamp 1606120353
transform 1 0 9108 0 -1 28832
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _0523_
timestamp 1606120353
transform 1 0 10120 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__A
timestamp 1606120353
transform 1 0 10580 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_48_95
timestamp 1606120353
transform 1 0 9844 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_48_101
timestamp 1606120353
transform 1 0 10396 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_48_105
timestamp 1606120353
transform 1 0 10764 0 -1 28832
box 0 -48 552 592
use sky130_fd_sc_hd__buf_1  _0903_
timestamp 1606120353
transform 1 0 11316 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__nor3_4  _0914_
timestamp 1606120353
transform 1 0 12420 0 -1 28832
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1606120353
transform 1 0 12328 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__C
timestamp 1606120353
transform 1 0 12144 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__C
timestamp 1606120353
transform 1 0 11776 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_114
timestamp 1606120353
transform 1 0 11592 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_118
timestamp 1606120353
transform 1 0 11960 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _1023_
timestamp 1606120353
transform 1 0 14352 0 -1 28832
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__A2
timestamp 1606120353
transform 1 0 13800 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_136
timestamp 1606120353
transform 1 0 13616 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_48_140
timestamp 1606120353
transform 1 0 13984 0 -1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_48_153
timestamp 1606120353
transform 1 0 15180 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1089_
timestamp 1606120353
transform 1 0 16008 0 -1 28832
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__B
timestamp 1606120353
transform 1 0 15732 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__C
timestamp 1606120353
transform 1 0 15364 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_157
timestamp 1606120353
transform 1 0 15548 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_48_161
timestamp 1606120353
transform 1 0 15916 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_48_175
timestamp 1606120353
transform 1 0 17204 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1606120353
transform -1 0 18860 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1606120353
transform 1 0 17940 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__B1
timestamp 1606120353
transform 1 0 17388 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__A2
timestamp 1606120353
transform 1 0 17756 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_179
timestamp 1606120353
transform 1 0 17572 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_48_184
timestamp 1606120353
transform 1 0 18032 0 -1 28832
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1290_
timestamp 1606120353
transform 1 0 1472 0 1 28832
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1606120353
transform 1 0 1104 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_49_3
timestamp 1606120353
transform 1 0 1380 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_49_23
timestamp 1606120353
transform 1 0 3220 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__CLK
timestamp 1606120353
transform 1 0 3404 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_49_27
timestamp 1606120353
transform 1 0 3588 0 1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_49_32
timestamp 1606120353
transform 1 0 4048 0 1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1606120353
transform 1 0 3956 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_49_36
timestamp 1606120353
transform 1 0 4416 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__C
timestamp 1606120353
transform 1 0 4508 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_39
timestamp 1606120353
transform 1 0 4692 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__B
timestamp 1606120353
transform 1 0 4876 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_43
timestamp 1606120353
transform 1 0 5060 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0699_
timestamp 1606120353
transform 1 0 5428 0 1 28832
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__D
timestamp 1606120353
transform 1 0 5244 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__A
timestamp 1606120353
transform 1 0 6808 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_49_56
timestamp 1606120353
transform 1 0 6256 0 1 28832
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILLER_49_64
timestamp 1606120353
transform 1 0 6992 0 1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__nor3_4  _0527_
timestamp 1606120353
transform 1 0 7636 0 1 28832
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__A
timestamp 1606120353
transform 1 0 9016 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__A
timestamp 1606120353
transform 1 0 7452 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_49_68
timestamp 1606120353
transform 1 0 7360 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_49_84
timestamp 1606120353
transform 1 0 8832 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_88
timestamp 1606120353
transform 1 0 9200 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0546_
timestamp 1606120353
transform 1 0 10212 0 1 28832
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1606120353
transform 1 0 9568 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__B
timestamp 1606120353
transform 1 0 9384 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__A
timestamp 1606120353
transform 1 0 10028 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_49_93
timestamp 1606120353
transform 1 0 9660 0 1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_49_108
timestamp 1606120353
transform 1 0 11040 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__nand3_4  _0922_
timestamp 1606120353
transform 1 0 12604 0 1 28832
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__C
timestamp 1606120353
transform 1 0 12420 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A
timestamp 1606120353
transform 1 0 12052 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__B
timestamp 1606120353
transform 1 0 11684 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__B
timestamp 1606120353
transform 1 0 11316 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1606120353
transform 1 0 11500 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_117
timestamp 1606120353
transform 1 0 11868 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_121
timestamp 1606120353
transform 1 0 12236 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _1062_
timestamp 1606120353
transform 1 0 15272 0 1 28832
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1606120353
transform 1 0 15180 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A
timestamp 1606120353
transform 1 0 14352 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A
timestamp 1606120353
transform 1 0 14996 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_49_139
timestamp 1606120353
transform 1 0 13892 0 1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_49_143
timestamp 1606120353
transform 1 0 14260 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_49_146
timestamp 1606120353
transform 1 0 14536 0 1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_49_150
timestamp 1606120353
transform 1 0 14904 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__o21ai_4  _1087_
timestamp 1606120353
transform 1 0 16652 0 1 28832
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A
timestamp 1606120353
transform 1 0 16100 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__A1
timestamp 1606120353
transform 1 0 16468 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_161
timestamp 1606120353
transform 1 0 15916 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_165
timestamp 1606120353
transform 1 0 16284 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1606120353
transform -1 0 18860 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_49_182
timestamp 1606120353
transform 1 0 17848 0 1 28832
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1260_
timestamp 1606120353
transform 1 0 2024 0 -1 29920
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1606120353
transform 1 0 1104 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__D
timestamp 1606120353
transform 1 0 1564 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1606120353
transform 1 0 1380 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_50_7
timestamp 1606120353
transform 1 0 1748 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_clk
timestamp 1606120353
transform 1 0 4508 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__B
timestamp 1606120353
transform 1 0 5060 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__B1
timestamp 1606120353
transform 1 0 4324 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_50_29
timestamp 1606120353
transform 1 0 3772 0 -1 29920
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILLER_50_40
timestamp 1606120353
transform 1 0 4784 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0696_
timestamp 1606120353
transform 1 0 6808 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1606120353
transform 1 0 6716 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__A
timestamp 1606120353
transform 1 0 5428 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A
timestamp 1606120353
transform 1 0 5796 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_45
timestamp 1606120353
transform 1 0 5244 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_49
timestamp 1606120353
transform 1 0 5612 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_50_53
timestamp 1606120353
transform 1 0 5980 0 -1 29920
box 0 -48 736 592
use sky130_fd_sc_hd__decap_6  FILLER_50_65
timestamp 1606120353
transform 1 0 7084 0 -1 29920
box 0 -48 552 592
use sky130_fd_sc_hd__nor3_4  _0728_
timestamp 1606120353
transform 1 0 8280 0 -1 29920
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__B
timestamp 1606120353
transform 1 0 7636 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__C
timestamp 1606120353
transform 1 0 8096 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_50_73
timestamp 1606120353
transform 1 0 7820 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _0648_
timestamp 1606120353
transform 1 0 10212 0 -1 29920
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILLER_50_91
timestamp 1606120353
transform 1 0 9476 0 -1 29920
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_50_108
timestamp 1606120353
transform 1 0 11040 0 -1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__nor3_4  _0919_
timestamp 1606120353
transform 1 0 12420 0 -1 29920
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1606120353
transform 1 0 12328 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A
timestamp 1606120353
transform 1 0 12144 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0921_
timestamp 1606120353
transform 1 0 14352 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__B
timestamp 1606120353
transform 1 0 15272 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_50_136
timestamp 1606120353
transform 1 0 13616 0 -1 29920
box 0 -48 736 592
use sky130_fd_sc_hd__decap_6  FILLER_50_147
timestamp 1606120353
transform 1 0 14628 0 -1 29920
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_50_153
timestamp 1606120353
transform 1 0 15180 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__and3_4  _1079_
timestamp 1606120353
transform 1 0 15732 0 -1 29920
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__A1
timestamp 1606120353
transform 1 0 16744 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__A2
timestamp 1606120353
transform 1 0 17112 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_50_156
timestamp 1606120353
transform 1 0 15456 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_50_168
timestamp 1606120353
transform 1 0 16560 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_172
timestamp 1606120353
transform 1 0 16928 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_176
timestamp 1606120353
transform 1 0 17296 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1606120353
transform -1 0 18860 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1606120353
transform 1 0 17940 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__B1
timestamp 1606120353
transform 1 0 17480 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_50_180
timestamp 1606120353
transform 1 0 17664 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_50_184
timestamp 1606120353
transform 1 0 18032 0 -1 29920
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1606120353
transform 1 0 1104 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__D
timestamp 1606120353
transform 1 0 1656 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__CLK
timestamp 1606120353
transform 1 0 2024 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_51_3
timestamp 1606120353
transform 1 0 1380 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_51_8
timestamp 1606120353
transform 1 0 1840 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_51_12
timestamp 1606120353
transform 1 0 2208 0 1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__nand4_4  _0828_
timestamp 1606120353
transform 1 0 5060 0 1 29920
box 0 -48 1564 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1606120353
transform 1 0 3956 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__C
timestamp 1606120353
transform 1 0 4876 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__A1
timestamp 1606120353
transform 1 0 4508 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_51_24
timestamp 1606120353
transform 1 0 3312 0 1 29920
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_51_30
timestamp 1606120353
transform 1 0 3864 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_51_32
timestamp 1606120353
transform 1 0 4048 0 1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_51_36
timestamp 1606120353
transform 1 0 4416 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_51_39
timestamp 1606120353
transform 1 0 4692 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__D
timestamp 1606120353
transform 1 0 6808 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_60
timestamp 1606120353
transform 1 0 6624 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_51_64
timestamp 1606120353
transform 1 0 6992 0 1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _0522_
timestamp 1606120353
transform 1 0 8372 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0697_
timestamp 1606120353
transform 1 0 7360 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0522__A
timestamp 1606120353
transform 1 0 8832 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__A
timestamp 1606120353
transform 1 0 7820 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_71
timestamp 1606120353
transform 1 0 7636 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_51_75
timestamp 1606120353
transform 1 0 8004 0 1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_51_82
timestamp 1606120353
transform 1 0 8648 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_51_86
timestamp 1606120353
transform 1 0 9016 0 1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _0724_
timestamp 1606120353
transform 1 0 9660 0 1 29920
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1606120353
transform 1 0 9568 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__A
timestamp 1606120353
transform 1 0 9384 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_51_102
timestamp 1606120353
transform 1 0 10488 0 1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__a21o_4  _1029_
timestamp 1606120353
transform 1 0 12604 0 1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__A1
timestamp 1606120353
transform 1 0 12420 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__A2
timestamp 1606120353
transform 1 0 12052 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_51_114
timestamp 1606120353
transform 1 0 11592 0 1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_51_118
timestamp 1606120353
transform 1 0 11960 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_51_121
timestamp 1606120353
transform 1 0 12236 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1606120353
transform 1 0 15180 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__D
timestamp 1606120353
transform 1 0 14996 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__C
timestamp 1606120353
transform 1 0 14628 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_51_137
timestamp 1606120353
transform 1 0 13708 0 1 29920
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_51_145
timestamp 1606120353
transform 1 0 14444 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_149
timestamp 1606120353
transform 1 0 14812 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_154
timestamp 1606120353
transform 1 0 15272 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1024_
timestamp 1606120353
transform 1 0 15640 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _1094_
timestamp 1606120353
transform 1 0 16652 0 1 29920
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A
timestamp 1606120353
transform 1 0 16100 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A
timestamp 1606120353
transform 1 0 16468 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__B
timestamp 1606120353
transform 1 0 15456 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_161
timestamp 1606120353
transform 1 0 15916 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_165
timestamp 1606120353
transform 1 0 16284 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1606120353
transform -1 0 18860 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__B1
timestamp 1606120353
transform 1 0 18032 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_182
timestamp 1606120353
transform 1 0 17848 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_51_186
timestamp 1606120353
transform 1 0 18216 0 1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_53_11
timestamp 1606120353
transform 1 0 2116 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_7
timestamp 1606120353
transform 1 0 1748 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1606120353
transform 1 0 1380 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_52_3
timestamp 1606120353
transform 1 0 1380 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__D
timestamp 1606120353
transform 1 0 1932 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__D
timestamp 1606120353
transform 1 0 1564 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1606120353
transform 1 0 1104 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1606120353
transform 1 0 1104 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__CLK
timestamp 1606120353
transform 1 0 2300 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1606120353
transform 1 0 2484 0 1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1261_
timestamp 1606120353
transform 1 0 1656 0 -1 31008
box 0 -48 1748 592
use sky130_fd_sc_hd__o21ai_4  _0829_
timestamp 1606120353
transform 1 0 4784 0 -1 31008
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1606120353
transform 1 0 3956 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__A2
timestamp 1606120353
transform 1 0 4600 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_52_25
timestamp 1606120353
transform 1 0 3404 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_52_37
timestamp 1606120353
transform 1 0 4508 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_53_27
timestamp 1606120353
transform 1 0 3588 0 1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_53_32
timestamp 1606120353
transform 1 0 4048 0 1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_53_44
timestamp 1606120353
transform 1 0 5152 0 1 31008
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_53_52
timestamp 1606120353
transform 1 0 5888 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_clk_A
timestamp 1606120353
transform 1 0 5704 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_53_59
timestamp 1606120353
transform 1 0 6532 0 1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_52_53
timestamp 1606120353
transform 1 0 5980 0 -1 31008
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A
timestamp 1606120353
transform 1 0 6072 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0760_
timestamp 1606120353
transform 1 0 6256 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_53_66
timestamp 1606120353
transform 1 0 7176 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_53_63
timestamp 1606120353
transform 1 0 6900 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_52_62
timestamp 1606120353
transform 1 0 6808 0 -1 31008
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A
timestamp 1606120353
transform 1 0 6992 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1606120353
transform 1 0 6716 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_52_72
timestamp 1606120353
transform 1 0 7728 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__B1
timestamp 1606120353
transform 1 0 7912 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__B
timestamp 1606120353
transform 1 0 7544 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__A1
timestamp 1606120353
transform 1 0 7360 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0683_
timestamp 1606120353
transform 1 0 7544 0 1 31008
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_53_88
timestamp 1606120353
transform 1 0 9200 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_53_83
timestamp 1606120353
transform 1 0 8740 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_53_79
timestamp 1606120353
transform 1 0 8372 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_52_88
timestamp 1606120353
transform 1 0 9200 0 -1 31008
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__A2
timestamp 1606120353
transform 1 0 8556 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__C
timestamp 1606120353
transform 1 0 9016 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_52_76
timestamp 1606120353
transform 1 0 8096 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_53_93
timestamp 1606120353
transform 1 0 9660 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_97
timestamp 1606120353
transform 1 0 10028 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_52_94
timestamp 1606120353
transform 1 0 9752 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__A
timestamp 1606120353
transform 1 0 9844 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__A2
timestamp 1606120353
transform 1 0 9384 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__A1
timestamp 1606120353
transform 1 0 10212 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1606120353
transform 1 0 9568 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_53_108
timestamp 1606120353
transform 1 0 11040 0 1 31008
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_52_105
timestamp 1606120353
transform 1 0 10764 0 -1 31008
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_52_101
timestamp 1606120353
transform 1 0 10396 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__B1_N
timestamp 1606120353
transform 1 0 10580 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__nor3_4  _0620_
timestamp 1606120353
transform 1 0 9844 0 1 31008
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_4  FILLER_52_118
timestamp 1606120353
transform 1 0 11960 0 -1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_52_113
timestamp 1606120353
transform 1 0 11500 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__A
timestamp 1606120353
transform 1 0 11776 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__B
timestamp 1606120353
transform 1 0 11592 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0610_
timestamp 1606120353
transform 1 0 11776 0 1 31008
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_53_125
timestamp 1606120353
transform 1 0 12604 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_123
timestamp 1606120353
transform 1 0 12420 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__B1
timestamp 1606120353
transform 1 0 12604 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__A
timestamp 1606120353
transform 1 0 12788 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1606120353
transform 1 0 12328 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_53_129
timestamp 1606120353
transform 1 0 12972 0 1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_52_127
timestamp 1606120353
transform 1 0 12788 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_53_141
timestamp 1606120353
transform 1 0 14076 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A
timestamp 1606120353
transform 1 0 14168 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_53_152
timestamp 1606120353
transform 1 0 15088 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_53_148
timestamp 1606120353
transform 1 0 14720 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_144
timestamp 1606120353
transform 1 0 14352 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_52_151
timestamp 1606120353
transform 1 0 14996 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__A
timestamp 1606120353
transform 1 0 15272 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__B
timestamp 1606120353
transform 1 0 14904 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__C
timestamp 1606120353
transform 1 0 14536 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1606120353
transform 1 0 15180 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _1091_
timestamp 1606120353
transform 1 0 15272 0 1 31008
box 0 -48 644 592
use sky130_fd_sc_hd__decap_12  FILLER_52_139
timestamp 1606120353
transform 1 0 13892 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_53_165
timestamp 1606120353
transform 1 0 16284 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_161
timestamp 1606120353
transform 1 0 15916 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_52_160
timestamp 1606120353
transform 1 0 15824 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_52_156
timestamp 1606120353
transform 1 0 15456 0 -1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__B
timestamp 1606120353
transform 1 0 15916 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__B
timestamp 1606120353
transform 1 0 16100 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _1099_
timestamp 1606120353
transform 1 0 16100 0 -1 31008
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_52_176
timestamp 1606120353
transform 1 0 17296 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_172
timestamp 1606120353
transform 1 0 16928 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__A1
timestamp 1606120353
transform 1 0 17112 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__A
timestamp 1606120353
transform 1 0 16468 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1096_
timestamp 1606120353
transform 1 0 16652 0 1 31008
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1606120353
transform -1 0 18860 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1606120353
transform -1 0 18860 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1606120353
transform 1 0 17940 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__A2
timestamp 1606120353
transform 1 0 17480 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_52_180
timestamp 1606120353
transform 1 0 17664 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_52_184
timestamp 1606120353
transform 1 0 18032 0 -1 31008
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_53_182
timestamp 1606120353
transform 1 0 17848 0 1 31008
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1262_
timestamp 1606120353
transform 1 0 1472 0 -1 32096
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1606120353
transform 1 0 1104 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_54_3
timestamp 1606120353
transform 1 0 1380 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A
timestamp 1606120353
transform 1 0 4416 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__A
timestamp 1606120353
transform 1 0 4968 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_54_23
timestamp 1606120353
transform 1 0 3220 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_54_35
timestamp 1606120353
transform 1 0 4324 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_54_38
timestamp 1606120353
transform 1 0 4600 0 -1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_54_44
timestamp 1606120353
transform 1 0 5152 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1606120353
transform 1 0 6716 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk
timestamp 1606120353
transform 1 0 5888 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__C
timestamp 1606120353
transform 1 0 5336 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__D
timestamp 1606120353
transform 1 0 5704 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_48
timestamp 1606120353
transform 1 0 5520 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_54_55
timestamp 1606120353
transform 1 0 6164 0 -1 32096
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_54_62
timestamp 1606120353
transform 1 0 6808 0 -1 32096
box 0 -48 736 592
use sky130_fd_sc_hd__a21oi_4  _0684_
timestamp 1606120353
transform 1 0 7544 0 -1 32096
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_6  FILLER_54_83
timestamp 1606120353
transform 1 0 8740 0 -1 32096
box 0 -48 552 592
use sky130_fd_sc_hd__a21boi_4  _0585_
timestamp 1606120353
transform 1 0 10212 0 -1 32096
box 0 -48 1380 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__D
timestamp 1606120353
transform 1 0 9292 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__B
timestamp 1606120353
transform 1 0 9844 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_54_91
timestamp 1606120353
transform 1 0 9476 0 -1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_54_97
timestamp 1606120353
transform 1 0 10028 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0547_
timestamp 1606120353
transform 1 0 12420 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1606120353
transform 1 0 12328 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_54_114
timestamp 1606120353
transform 1 0 11592 0 -1 32096
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_54_126
timestamp 1606120353
transform 1 0 12696 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__or3_4  _1078_
timestamp 1606120353
transform 1 0 14536 0 -1 32096
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILLER_54_138
timestamp 1606120353
transform 1 0 13800 0 -1 32096
box 0 -48 736 592
use sky130_fd_sc_hd__and4_4  _1093_
timestamp 1606120353
transform 1 0 16100 0 -1 32096
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__C
timestamp 1606120353
transform 1 0 15916 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__D
timestamp 1606120353
transform 1 0 15548 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__B1
timestamp 1606120353
transform 1 0 17112 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_155
timestamp 1606120353
transform 1 0 15364 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_159
timestamp 1606120353
transform 1 0 15732 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_172
timestamp 1606120353
transform 1 0 16928 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_176
timestamp 1606120353
transform 1 0 17296 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1606120353
transform -1 0 18860 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1606120353
transform 1 0 17940 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__A2
timestamp 1606120353
transform 1 0 17480 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_54_180
timestamp 1606120353
transform 1 0 17664 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_54_184
timestamp 1606120353
transform 1 0 18032 0 -1 32096
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1263_
timestamp 1606120353
transform 1 0 1472 0 1 32096
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1606120353
transform 1 0 1104 0 1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_55_3
timestamp 1606120353
transform 1 0 1380 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_55_32
timestamp 1606120353
transform 1 0 4048 0 1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_55_27
timestamp 1606120353
transform 1 0 3588 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_23
timestamp 1606120353
transform 1 0 3220 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__CLK
timestamp 1606120353
transform 1 0 3404 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__C
timestamp 1606120353
transform 1 0 3772 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1606120353
transform 1 0 3956 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_55_38
timestamp 1606120353
transform 1 0 4600 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__B
timestamp 1606120353
transform 1 0 4784 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__B
timestamp 1606120353
transform 1 0 4416 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _0833_
timestamp 1606120353
transform 1 0 4968 0 1 32096
box 0 -48 1564 592
use sky130_fd_sc_hd__decap_12  FILLER_55_59
timestamp 1606120353
transform 1 0 6532 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__buf_1  _0685_
timestamp 1606120353
transform 1 0 8188 0 1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__C
timestamp 1606120353
transform 1 0 8924 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A
timestamp 1606120353
transform 1 0 8004 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_55_71
timestamp 1606120353
transform 1 0 7636 0 1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_55_80
timestamp 1606120353
transform 1 0 8464 0 1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_55_84
timestamp 1606120353
transform 1 0 8832 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_55_87
timestamp 1606120353
transform 1 0 9108 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__a22oi_4  _0578_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 10580 0 1 32096
box 0 -48 1564 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1606120353
transform 1 0 9568 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__A1
timestamp 1606120353
transform 1 0 10396 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__B1
timestamp 1606120353
transform 1 0 10028 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__B
timestamp 1606120353
transform 1 0 9292 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_55_91
timestamp 1606120353
transform 1 0 9476 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_55_93
timestamp 1606120353
transform 1 0 9660 0 1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_55_99
timestamp 1606120353
transform 1 0 10212 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_55_120
timestamp 1606120353
transform 1 0 12144 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_55_132
timestamp 1606120353
transform 1 0 13248 0 1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_55_138
timestamp 1606120353
transform 1 0 13800 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__B1
timestamp 1606120353
transform 1 0 13616 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_55_146
timestamp 1606120353
transform 1 0 14536 0 1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_55_142
timestamp 1606120353
transform 1 0 14168 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A1
timestamp 1606120353
transform 1 0 14352 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A2
timestamp 1606120353
transform 1 0 13984 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_55_150
timestamp 1606120353
transform 1 0 14904 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__B
timestamp 1606120353
transform 1 0 14996 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1606120353
transform 1 0 15180 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _1098_
timestamp 1606120353
transform 1 0 15272 0 1 32096
box 0 -48 644 592
use sky130_fd_sc_hd__o21ai_4  _1100_
timestamp 1606120353
transform 1 0 16652 0 1 32096
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__A1
timestamp 1606120353
transform 1 0 16100 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__A1
timestamp 1606120353
transform 1 0 16468 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_161
timestamp 1606120353
transform 1 0 15916 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_165
timestamp 1606120353
transform 1 0 16284 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1606120353
transform -1 0 18860 0 1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__B1
timestamp 1606120353
transform 1 0 18032 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__B1
timestamp 1606120353
transform 1 0 18400 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_182
timestamp 1606120353
transform 1 0 17848 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_186
timestamp 1606120353
transform 1 0 18216 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1264_
timestamp 1606120353
transform 1 0 1380 0 -1 33184
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1606120353
transform 1 0 1104 0 -1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_56_22
timestamp 1606120353
transform 1 0 3128 0 -1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__nand4_4  _0854_
timestamp 1606120353
transform 1 0 4416 0 -1 33184
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__D
timestamp 1606120353
transform 1 0 4232 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__CLK
timestamp 1606120353
transform 1 0 3864 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_32
timestamp 1606120353
transform 1 0 4048 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1606120353
transform 1 0 6716 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__A
timestamp 1606120353
transform 1 0 6532 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A1
timestamp 1606120353
transform 1 0 6992 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__D
timestamp 1606120353
transform 1 0 6164 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_53
timestamp 1606120353
transform 1 0 5980 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_57
timestamp 1606120353
transform 1 0 6348 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_62
timestamp 1606120353
transform 1 0 6808 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_66
timestamp 1606120353
transform 1 0 7176 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A2
timestamp 1606120353
transform 1 0 7360 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__A
timestamp 1606120353
transform 1 0 9108 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_56_70
timestamp 1606120353
transform 1 0 7544 0 -1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_56_82
timestamp 1606120353
transform 1 0 8648 0 -1 33184
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_56_86
timestamp 1606120353
transform 1 0 9016 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__nand4_4  _0602_
timestamp 1606120353
transform 1 0 9292 0 -1 33184
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__B2
timestamp 1606120353
transform 1 0 11040 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_106
timestamp 1606120353
transform 1 0 10856 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_110
timestamp 1606120353
transform 1 0 11224 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1606120353
transform 1 0 12328 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__A2
timestamp 1606120353
transform 1 0 11408 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_56_114
timestamp 1606120353
transform 1 0 11592 0 -1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_56_123
timestamp 1606120353
transform 1 0 12420 0 -1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__a21oi_4  _1030_
timestamp 1606120353
transform 1 0 13984 0 -1 33184
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_4  FILLER_56_135
timestamp 1606120353
transform 1 0 13524 0 -1 33184
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1606120353
transform 1 0 13892 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_56_153
timestamp 1606120353
transform 1 0 15180 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1112_
timestamp 1606120353
transform 1 0 16008 0 -1 33184
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__A
timestamp 1606120353
transform 1 0 15364 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A2
timestamp 1606120353
transform 1 0 15824 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_56_157
timestamp 1606120353
transform 1 0 15548 0 -1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_56_175
timestamp 1606120353
transform 1 0 17204 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1606120353
transform -1 0 18860 0 -1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1606120353
transform 1 0 17940 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__A2
timestamp 1606120353
transform 1 0 17388 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__A2
timestamp 1606120353
transform 1 0 17756 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_179
timestamp 1606120353
transform 1 0 17572 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_56_184
timestamp 1606120353
transform 1 0 18032 0 -1 33184
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1606120353
transform 1 0 1104 0 1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__D
timestamp 1606120353
transform 1 0 1564 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__CLK
timestamp 1606120353
transform 1 0 1932 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__CLK
timestamp 1606120353
transform 1 0 2852 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1606120353
transform 1 0 1380 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_7
timestamp 1606120353
transform 1 0 1748 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_57_11
timestamp 1606120353
transform 1 0 2116 0 1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_57_21
timestamp 1606120353
transform 1 0 3036 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1265_
timestamp 1606120353
transform 1 0 4048 0 1 33184
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1606120353
transform 1 0 3956 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__D
timestamp 1606120353
transform 1 0 3220 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__D
timestamp 1606120353
transform 1 0 3772 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_57_25
timestamp 1606120353
transform 1 0 3404 0 1 33184
box 0 -48 368 592
use sky130_fd_sc_hd__nand4_4  _0846_
timestamp 1606120353
transform 1 0 6532 0 1 33184
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__B
timestamp 1606120353
transform 1 0 6348 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__C
timestamp 1606120353
transform 1 0 5980 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_51
timestamp 1606120353
transform 1 0 5796 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_55
timestamp 1606120353
transform 1 0 6164 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__B
timestamp 1606120353
transform 1 0 8924 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__B1
timestamp 1606120353
transform 1 0 8280 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_76
timestamp 1606120353
transform 1 0 8096 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_57_80
timestamp 1606120353
transform 1 0 8464 0 1 33184
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_57_84
timestamp 1606120353
transform 1 0 8832 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_57_87
timestamp 1606120353
transform 1 0 9108 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_98
timestamp 1606120353
transform 1 0 10120 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_93
timestamp 1606120353
transform 1 0 9660 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_57_91
timestamp 1606120353
transform 1 0 9476 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__A
timestamp 1606120353
transform 1 0 9292 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1606120353
transform 1 0 9568 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0548_
timestamp 1606120353
transform 1 0 9844 0 1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_57_102
timestamp 1606120353
transform 1 0 10488 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__C
timestamp 1606120353
transform 1 0 10672 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0548__A
timestamp 1606120353
transform 1 0 10304 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_57_106
timestamp 1606120353
transform 1 0 10856 0 1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_57_118
timestamp 1606120353
transform 1 0 11960 0 1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_57_130
timestamp 1606120353
transform 1 0 13064 0 1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1606120353
transform 1 0 15180 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__A2
timestamp 1606120353
transform 1 0 14076 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__B1
timestamp 1606120353
transform 1 0 14444 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__A1
timestamp 1606120353
transform 1 0 14812 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_57_138
timestamp 1606120353
transform 1 0 13800 0 1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_57_143
timestamp 1606120353
transform 1 0 14260 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_147
timestamp 1606120353
transform 1 0 14628 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_151
timestamp 1606120353
transform 1 0 14996 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_154
timestamp 1606120353
transform 1 0 15272 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1103_
timestamp 1606120353
transform 1 0 16652 0 1 33184
box 0 -48 1196 592
use sky130_fd_sc_hd__buf_1  _1105_
timestamp 1606120353
transform 1 0 15640 0 1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__A1
timestamp 1606120353
transform 1 0 16468 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A1
timestamp 1606120353
transform 1 0 16100 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__A
timestamp 1606120353
transform 1 0 15456 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_161
timestamp 1606120353
transform 1 0 15916 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_165
timestamp 1606120353
transform 1 0 16284 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1606120353
transform -1 0 18860 0 1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__B1
timestamp 1606120353
transform 1 0 18032 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__A2
timestamp 1606120353
transform 1 0 18400 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_182
timestamp 1606120353
transform 1 0 17848 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_186
timestamp 1606120353
transform 1 0 18216 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1606120353
transform 1 0 1104 0 -1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1606120353
transform 1 0 1380 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_58_15
timestamp 1606120353
transform 1 0 2484 0 -1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1271_
timestamp 1606120353
transform 1 0 3220 0 -1 34272
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_8  FILLER_58_42
timestamp 1606120353
transform 1 0 4968 0 -1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__a21oi_4  _0751_
timestamp 1606120353
transform 1 0 6808 0 -1 34272
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1606120353
transform 1 0 6716 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__B1
timestamp 1606120353
transform 1 0 6256 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__B1
timestamp 1606120353
transform 1 0 5888 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_50
timestamp 1606120353
transform 1 0 5704 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_54
timestamp 1606120353
transform 1 0 6072 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_58_58
timestamp 1606120353
transform 1 0 6440 0 -1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_58_75
timestamp 1606120353
transform 1 0 8004 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_58_87
timestamp 1606120353
transform 1 0 9108 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__nand3_4  _0601_
timestamp 1606120353
transform 1 0 9292 0 -1 34272
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILLER_58_103
timestamp 1606120353
transform 1 0 10580 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1606120353
transform 1 0 12328 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_58_115
timestamp 1606120353
transform 1 0 11684 0 -1 34272
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_58_121
timestamp 1606120353
transform 1 0 12236 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_58_123
timestamp 1606120353
transform 1 0 12420 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__a21oi_4  _1107_
timestamp 1606120353
transform 1 0 14076 0 -1 34272
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_6  FILLER_58_135
timestamp 1606120353
transform 1 0 13524 0 -1 34272
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_58_154
timestamp 1606120353
transform 1 0 15272 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1113_
timestamp 1606120353
transform 1 0 16008 0 -1 34272
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__A2
timestamp 1606120353
transform 1 0 15824 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__B1
timestamp 1606120353
transform 1 0 15456 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_158
timestamp 1606120353
transform 1 0 15640 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_175
timestamp 1606120353
transform 1 0 17204 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1606120353
transform -1 0 18860 0 -1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1606120353
transform 1 0 17940 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__A1
timestamp 1606120353
transform 1 0 17388 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_58_179
timestamp 1606120353
transform 1 0 17572 0 -1 34272
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_58_184
timestamp 1606120353
transform 1 0 18032 0 -1 34272
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILLER_60_7
timestamp 1606120353
transform 1 0 1748 0 -1 35360
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1606120353
transform 1 0 1380 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_11
timestamp 1606120353
transform 1 0 2116 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_59_3
timestamp 1606120353
transform 1 0 1380 0 1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__D
timestamp 1606120353
transform 1 0 1564 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1606120353
transform 1 0 1104 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1606120353
transform 1 0 1104 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_59_19
timestamp 1606120353
transform 1 0 2852 0 1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_59_15
timestamp 1606120353
transform 1 0 2484 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__CLK
timestamp 1606120353
transform 1 0 2668 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__D
timestamp 1606120353
transform 1 0 2300 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1267_
timestamp 1606120353
transform 1 0 2300 0 -1 35360
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  FILLER_60_32
timestamp 1606120353
transform 1 0 4048 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_59_32
timestamp 1606120353
transform 1 0 4048 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_59_27
timestamp 1606120353
transform 1 0 3588 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A2
timestamp 1606120353
transform 1 0 3772 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1606120353
transform 1 0 3956 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_60_41
timestamp 1606120353
transform 1 0 4876 0 -1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_60_37
timestamp 1606120353
transform 1 0 4508 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__B1
timestamp 1606120353
transform 1 0 4692 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A1
timestamp 1606120353
transform 1 0 4324 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0834_
timestamp 1606120353
transform 1 0 4324 0 1 34272
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_60_54
timestamp 1606120353
transform 1 0 6072 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_60_49
timestamp 1606120353
transform 1 0 5612 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_59_52
timestamp 1606120353
transform 1 0 5888 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_48
timestamp 1606120353
transform 1 0 5520 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__A1_N
timestamp 1606120353
transform 1 0 5888 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A1
timestamp 1606120353
transform 1 0 5704 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__A2_N
timestamp 1606120353
transform 1 0 6072 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_60_58
timestamp 1606120353
transform 1 0 6440 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__B2
timestamp 1606120353
transform 1 0 6256 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1606120353
transform 1 0 6716 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__a2bb2oi_4  _0748_
timestamp 1606120353
transform 1 0 6256 0 1 34272
box 0 -48 1932 592
use sky130_fd_sc_hd__o21a_4  _0746_
timestamp 1606120353
transform 1 0 6808 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A2
timestamp 1606120353
transform 1 0 8372 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_77
timestamp 1606120353
transform 1 0 8188 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_59_81
timestamp 1606120353
transform 1 0 8556 0 1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_60_74
timestamp 1606120353
transform 1 0 7912 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_60_86
timestamp 1606120353
transform 1 0 9016 0 -1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_60_98
timestamp 1606120353
transform 1 0 10120 0 -1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_60_94
timestamp 1606120353
transform 1 0 9752 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_59_93
timestamp 1606120353
transform 1 0 9660 0 1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_59_89
timestamp 1606120353
transform 1 0 9292 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0518__A
timestamp 1606120353
transform 1 0 9936 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1606120353
transform 1 0 9568 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_60_102
timestamp 1606120353
transform 1 0 10488 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_59_101
timestamp 1606120353
transform 1 0 10396 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__A
timestamp 1606120353
transform 1 0 10580 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0537_
timestamp 1606120353
transform 1 0 10580 0 -1 35360
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILLER_59_105
timestamp 1606120353
transform 1 0 10764 0 1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1606120353
transform 1 0 12328 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_59_117
timestamp 1606120353
transform 1 0 11868 0 1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_59_129
timestamp 1606120353
transform 1 0 12972 0 1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_60_112
timestamp 1606120353
transform 1 0 11408 0 -1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_60_120
timestamp 1606120353
transform 1 0 12144 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_60_123
timestamp 1606120353
transform 1 0 12420 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_60_140
timestamp 1606120353
transform 1 0 13984 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_60_135
timestamp 1606120353
transform 1 0 13524 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_59_139
timestamp 1606120353
transform 1 0 13892 0 1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A
timestamp 1606120353
transform 1 0 13708 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1019_
timestamp 1606120353
transform 1 0 13708 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_60_144
timestamp 1606120353
transform 1 0 14352 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_59_147
timestamp 1606120353
transform 1 0 14628 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A
timestamp 1606120353
transform 1 0 14720 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A
timestamp 1606120353
transform 1 0 14168 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__B
timestamp 1606120353
transform 1 0 14536 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1045_
timestamp 1606120353
transform 1 0 14720 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_60_151
timestamp 1606120353
transform 1 0 14996 0 -1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_59_154
timestamp 1606120353
transform 1 0 15272 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_59_150
timestamp 1606120353
transform 1 0 14904 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1606120353
transform 1 0 15180 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_60_159
timestamp 1606120353
transform 1 0 15732 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_59_162
timestamp 1606120353
transform 1 0 16008 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_158
timestamp 1606120353
transform 1 0 15640 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__B1
timestamp 1606120353
transform 1 0 15824 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__A1
timestamp 1606120353
transform 1 0 16192 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A
timestamp 1606120353
transform 1 0 15824 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1054_
timestamp 1606120353
transform 1 0 15364 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_60_175
timestamp 1606120353
transform 1 0 17204 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_59_166
timestamp 1606120353
transform 1 0 16376 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _1116_
timestamp 1606120353
transform 1 0 16652 0 1 34272
box 0 -48 1196 592
use sky130_fd_sc_hd__o21ai_4  _1115_
timestamp 1606120353
transform 1 0 16008 0 -1 35360
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1606120353
transform -1 0 18860 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1606120353
transform -1 0 18860 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1606120353
transform 1 0 17940 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__A2
timestamp 1606120353
transform 1 0 17388 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__B1
timestamp 1606120353
transform 1 0 18032 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_182
timestamp 1606120353
transform 1 0 17848 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_59_186
timestamp 1606120353
transform 1 0 18216 0 1 34272
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_60_179
timestamp 1606120353
transform 1 0 17572 0 -1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_60_184
timestamp 1606120353
transform 1 0 18032 0 -1 35360
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1266_
timestamp 1606120353
transform 1 0 1472 0 1 35360
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1606120353
transform 1 0 1104 0 1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_61_3
timestamp 1606120353
transform 1 0 1380 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1606120353
transform 1 0 3956 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A
timestamp 1606120353
transform 1 0 4876 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_61_23
timestamp 1606120353
transform 1 0 3220 0 1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_61_32
timestamp 1606120353
transform 1 0 4048 0 1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_61_40
timestamp 1606120353
transform 1 0 4784 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_61_43
timestamp 1606120353
transform 1 0 5060 0 1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__inv_8  _0693_
timestamp 1606120353
transform 1 0 6072 0 1 35360
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B
timestamp 1606120353
transform 1 0 7084 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A
timestamp 1606120353
transform 1 0 5888 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_61_51
timestamp 1606120353
transform 1 0 5796 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_61_63
timestamp 1606120353
transform 1 0 6900 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_67
timestamp 1606120353
transform 1 0 7268 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A
timestamp 1606120353
transform 1 0 7452 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0758_
timestamp 1606120353
transform 1 0 7636 0 1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_61_74
timestamp 1606120353
transform 1 0 7912 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_78
timestamp 1606120353
transform 1 0 8280 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A
timestamp 1606120353
transform 1 0 8096 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__C
timestamp 1606120353
transform 1 0 8464 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_82
timestamp 1606120353
transform 1 0 8648 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A
timestamp 1606120353
transform 1 0 8832 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_86
timestamp 1606120353
transform 1 0 9016 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A1
timestamp 1606120353
transform 1 0 9200 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0518_
timestamp 1606120353
transform 1 0 9936 0 1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__nand2_4  _0529_
timestamp 1606120353
transform 1 0 10948 0 1 35360
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1606120353
transform 1 0 9568 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0529__B
timestamp 1606120353
transform 1 0 10764 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__A
timestamp 1606120353
transform 1 0 10396 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_90
timestamp 1606120353
transform 1 0 9384 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_61_93
timestamp 1606120353
transform 1 0 9660 0 1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_61_99
timestamp 1606120353
transform 1 0 10212 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_103
timestamp 1606120353
transform 1 0 10580 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0923_
timestamp 1606120353
transform 1 0 13156 0 1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A
timestamp 1606120353
transform 1 0 12972 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0529__A
timestamp 1606120353
transform 1 0 11960 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__CLK
timestamp 1606120353
transform 1 0 12512 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_116
timestamp 1606120353
transform 1 0 11776 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_61_120
timestamp 1606120353
transform 1 0 12144 0 1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_61_126
timestamp 1606120353
transform 1 0 12696 0 1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_61_134
timestamp 1606120353
transform 1 0 13432 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_138
timestamp 1606120353
transform 1 0 13800 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A
timestamp 1606120353
transform 1 0 13616 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A
timestamp 1606120353
transform 1 0 13984 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1038_
timestamp 1606120353
transform 1 0 14168 0 1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_61_145
timestamp 1606120353
transform 1 0 14444 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__C
timestamp 1606120353
transform 1 0 14628 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_149
timestamp 1606120353
transform 1 0 14812 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__D
timestamp 1606120353
transform 1 0 14996 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1606120353
transform 1 0 15180 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_61_154
timestamp 1606120353
transform 1 0 15272 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _1048_
timestamp 1606120353
transform 1 0 15364 0 1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _1124_
timestamp 1606120353
transform 1 0 16652 0 1 35360
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__A
timestamp 1606120353
transform 1 0 15824 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A
timestamp 1606120353
transform 1 0 16468 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_158
timestamp 1606120353
transform 1 0 15640 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_61_162
timestamp 1606120353
transform 1 0 16008 0 1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_61_166
timestamp 1606120353
transform 1 0 16376 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1606120353
transform -1 0 18860 0 1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__A2
timestamp 1606120353
transform 1 0 18032 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__B1
timestamp 1606120353
transform 1 0 18400 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_182
timestamp 1606120353
transform 1 0 17848 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_186
timestamp 1606120353
transform 1 0 18216 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1606120353
transform 1 0 1104 0 -1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__CLK
timestamp 1606120353
transform 1 0 1564 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1606120353
transform 1 0 1380 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_62_7
timestamp 1606120353
transform 1 0 1748 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_62_19
timestamp 1606120353
transform 1 0 2852 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__inv_8  _0804_
timestamp 1606120353
transform 1 0 4876 0 -1 36448
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__B2
timestamp 1606120353
transform 1 0 4692 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_62_31
timestamp 1606120353
transform 1 0 3956 0 -1 36448
box 0 -48 736 592
use sky130_fd_sc_hd__nand3_4  _0807_
timestamp 1606120353
transform 1 0 6808 0 -1 36448
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1606120353
transform 1 0 6716 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A1
timestamp 1606120353
transform 1 0 6532 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A2
timestamp 1606120353
transform 1 0 6164 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_62_50
timestamp 1606120353
transform 1 0 5704 0 -1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_62_54
timestamp 1606120353
transform 1 0 6072 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_62_57
timestamp 1606120353
transform 1 0 6348 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0732_
timestamp 1606120353
transform 1 0 8832 0 -1 36448
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__D1
timestamp 1606120353
transform 1 0 8464 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_62_76
timestamp 1606120353
transform 1 0 8096 0 -1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 1606120353
transform 1 0 8648 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0592_
timestamp 1606120353
transform 1 0 10764 0 -1 36448
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__A
timestamp 1606120353
transform 1 0 10580 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_62_93
timestamp 1606120353
transform 1 0 9660 0 -1 36448
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_62_101
timestamp 1606120353
transform 1 0 10396 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _1012_
timestamp 1606120353
transform 1 0 12972 0 -1 36448
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1606120353
transform 1 0 12328 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__C
timestamp 1606120353
transform 1 0 12144 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__C
timestamp 1606120353
transform 1 0 12604 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_62_114
timestamp 1606120353
transform 1 0 11592 0 -1 36448
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_62_123
timestamp 1606120353
transform 1 0 12420 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_127
timestamp 1606120353
transform 1 0 12788 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _1067_
timestamp 1606120353
transform 1 0 14536 0 -1 36448
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__C
timestamp 1606120353
transform 1 0 13984 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__A1
timestamp 1606120353
transform 1 0 14352 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_138
timestamp 1606120353
transform 1 0 13800 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_142
timestamp 1606120353
transform 1 0 14168 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1047_
timestamp 1606120353
transform 1 0 16836 0 -1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__A1
timestamp 1606120353
transform 1 0 16652 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__A2
timestamp 1606120353
transform 1 0 17296 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__B1
timestamp 1606120353
transform 1 0 16284 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_163
timestamp 1606120353
transform 1 0 16100 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_167
timestamp 1606120353
transform 1 0 16468 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_174
timestamp 1606120353
transform 1 0 17112 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1606120353
transform -1 0 18860 0 -1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1606120353
transform 1 0 17940 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_62_178
timestamp 1606120353
transform 1 0 17480 0 -1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_62_182
timestamp 1606120353
transform 1 0 17848 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_62_184
timestamp 1606120353
transform 1 0 18032 0 -1 36448
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1606120353
transform 1 0 1104 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__CLK
timestamp 1606120353
transform 1 0 1564 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1606120353
transform 1 0 1380 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_63_7
timestamp 1606120353
transform 1 0 1748 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_63_19
timestamp 1606120353
transform 1 0 2852 0 1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_63_32
timestamp 1606120353
transform 1 0 4048 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_63_29
timestamp 1606120353
transform 1 0 3772 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_25
timestamp 1606120353
transform 1 0 3404 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__CLK
timestamp 1606120353
transform 1 0 3220 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__D
timestamp 1606120353
transform 1 0 3588 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1606120353
transform 1 0 3956 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_63_37
timestamp 1606120353
transform 1 0 4508 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A1
timestamp 1606120353
transform 1 0 4324 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A2
timestamp 1606120353
transform 1 0 4692 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__a22oi_4  _0810_
timestamp 1606120353
transform 1 0 4876 0 1 36448
box 0 -48 1564 592
use sky130_fd_sc_hd__a21o_4  _0808_
timestamp 1606120353
transform 1 0 7176 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__B1
timestamp 1606120353
transform 1 0 6992 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__A
timestamp 1606120353
transform 1 0 6624 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_58
timestamp 1606120353
transform 1 0 6440 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_62
timestamp 1606120353
transform 1 0 6808 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A2
timestamp 1606120353
transform 1 0 8464 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B1
timestamp 1606120353
transform 1 0 8832 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__C1
timestamp 1606120353
transform 1 0 9200 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_78
timestamp 1606120353
transform 1 0 8280 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_82
timestamp 1606120353
transform 1 0 8648 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_86
timestamp 1606120353
transform 1 0 9016 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0596_
timestamp 1606120353
transform 1 0 10580 0 1 36448
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1606120353
transform 1 0 9568 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A
timestamp 1606120353
transform 1 0 9844 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__D
timestamp 1606120353
transform 1 0 10212 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_90
timestamp 1606120353
transform 1 0 9384 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_93
timestamp 1606120353
transform 1 0 9660 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_97
timestamp 1606120353
transform 1 0 10028 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_101
timestamp 1606120353
transform 1 0 10396 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_112
timestamp 1606120353
transform 1 0 11408 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_63_116
timestamp 1606120353
transform 1 0 11776 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0530__A
timestamp 1606120353
transform 1 0 11592 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A
timestamp 1606120353
transform 1 0 12052 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_121
timestamp 1606120353
transform 1 0 12236 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__B1
timestamp 1606120353
transform 1 0 12420 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1028_
timestamp 1606120353
transform 1 0 12604 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_63_128
timestamp 1606120353
transform 1 0 12880 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A
timestamp 1606120353
transform 1 0 13064 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_132
timestamp 1606120353
transform 1 0 13248 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1021_
timestamp 1606120353
transform 1 0 15272 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__and4_4  _1039_
timestamp 1606120353
transform 1 0 13616 0 1 36448
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1606120353
transform 1 0 15180 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__A
timestamp 1606120353
transform 1 0 13432 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__D
timestamp 1606120353
transform 1 0 14628 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__A2
timestamp 1606120353
transform 1 0 14996 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_145
timestamp 1606120353
transform 1 0 14444 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_149
timestamp 1606120353
transform 1 0 14812 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1120_
timestamp 1606120353
transform 1 0 16652 0 1 36448
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__A
timestamp 1606120353
transform 1 0 15732 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__A1
timestamp 1606120353
transform 1 0 16468 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__A1
timestamp 1606120353
transform 1 0 16100 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_157
timestamp 1606120353
transform 1 0 15548 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_161
timestamp 1606120353
transform 1 0 15916 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_165
timestamp 1606120353
transform 1 0 16284 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1606120353
transform -1 0 18860 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__A2
timestamp 1606120353
transform 1 0 18032 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_182
timestamp 1606120353
transform 1 0 17848 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_63_186
timestamp 1606120353
transform 1 0 18216 0 1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1606120353
transform 1 0 1104 0 -1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__D
timestamp 1606120353
transform 1 0 1564 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__D
timestamp 1606120353
transform 1 0 1932 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__CLK
timestamp 1606120353
transform 1 0 3036 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__CLK
timestamp 1606120353
transform 1 0 2300 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1606120353
transform 1 0 1380 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_7
timestamp 1606120353
transform 1 0 1748 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_11
timestamp 1606120353
transform 1 0 2116 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_64_15
timestamp 1606120353
transform 1 0 2484 0 -1 37536
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1150_
timestamp 1606120353
transform 1 0 3588 0 -1 37536
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__CLK
timestamp 1606120353
transform 1 0 3404 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_23
timestamp 1606120353
transform 1 0 3220 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_46
timestamp 1606120353
transform 1 0 5336 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__B1
timestamp 1606120353
transform 1 0 5520 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_64_50
timestamp 1606120353
transform 1 0 5704 0 -1 37536
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_64_54
timestamp 1606120353
transform 1 0 6072 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A1
timestamp 1606120353
transform 1 0 6164 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1606120353
transform 1 0 6348 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A2
timestamp 1606120353
transform 1 0 6532 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1606120353
transform 1 0 6716 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0692_
timestamp 1606120353
transform 1 0 6808 0 -1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_64_65
timestamp 1606120353
transform 1 0 7084 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__a2111oi_4  _0740_
timestamp 1606120353
transform 1 0 8464 0 -1 37536
box 0 -48 2024 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A
timestamp 1606120353
transform 1 0 8004 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__C
timestamp 1606120353
transform 1 0 7636 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__A
timestamp 1606120353
transform 1 0 7268 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_69
timestamp 1606120353
transform 1 0 7452 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_73
timestamp 1606120353
transform 1 0 7820 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_64_77
timestamp 1606120353
transform 1 0 8188 0 -1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0530_
timestamp 1606120353
transform 1 0 11224 0 -1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__B
timestamp 1606120353
transform 1 0 10672 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__D
timestamp 1606120353
transform 1 0 11040 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_102
timestamp 1606120353
transform 1 0 10488 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_106
timestamp 1606120353
transform 1 0 10856 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _1015_
timestamp 1606120353
transform 1 0 12512 0 -1 37536
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1606120353
transform 1 0 12328 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__B
timestamp 1606120353
transform 1 0 11960 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_64_113
timestamp 1606120353
transform 1 0 11500 0 -1 37536
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_64_117
timestamp 1606120353
transform 1 0 11868 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_64_120
timestamp 1606120353
transform 1 0 12144 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_64_123
timestamp 1606120353
transform 1 0 12420 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__o21ai_4  _1125_
timestamp 1606120353
transform 1 0 14076 0 -1 37536
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__B
timestamp 1606120353
transform 1 0 13616 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_64_133
timestamp 1606120353
transform 1 0 13340 0 -1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_64_138
timestamp 1606120353
transform 1 0 13800 0 -1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_64_154
timestamp 1606120353
transform 1 0 15272 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1122_
timestamp 1606120353
transform 1 0 16008 0 -1 37536
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__C
timestamp 1606120353
transform 1 0 15824 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__D
timestamp 1606120353
transform 1 0 15456 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_158
timestamp 1606120353
transform 1 0 15640 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_175
timestamp 1606120353
transform 1 0 17204 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1606120353
transform -1 0 18860 0 -1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1606120353
transform 1 0 17940 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__B1
timestamp 1606120353
transform 1 0 17388 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_64_179
timestamp 1606120353
transform 1 0 17572 0 -1 37536
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_64_184
timestamp 1606120353
transform 1 0 18032 0 -1 37536
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1269_
timestamp 1606120353
transform 1 0 1472 0 1 37536
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1606120353
transform 1 0 1104 0 1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_65_3
timestamp 1606120353
transform 1 0 1380 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1270_
timestamp 1606120353
transform 1 0 4048 0 1 37536
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1606120353
transform 1 0 3956 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__D
timestamp 1606120353
transform 1 0 3772 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__D
timestamp 1606120353
transform 1 0 3404 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_23
timestamp 1606120353
transform 1 0 3220 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_27
timestamp 1606120353
transform 1 0 3588 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0809_
timestamp 1606120353
transform 1 0 6532 0 1 37536
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__B1
timestamp 1606120353
transform 1 0 6348 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A
timestamp 1606120353
transform 1 0 5980 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_51
timestamp 1606120353
transform 1 0 5796 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_55
timestamp 1606120353
transform 1 0 6164 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0750_
timestamp 1606120353
transform 1 0 8464 0 1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__B
timestamp 1606120353
transform 1 0 8004 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__C
timestamp 1606120353
transform 1 0 9016 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_65_72
timestamp 1606120353
transform 1 0 7728 0 1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_65_77
timestamp 1606120353
transform 1 0 8188 0 1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_65_83
timestamp 1606120353
transform 1 0 8740 0 1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_65_88
timestamp 1606120353
transform 1 0 9200 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0734_
timestamp 1606120353
transform 1 0 9660 0 1 37536
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1606120353
transform 1 0 9568 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__A
timestamp 1606120353
transform 1 0 10764 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__B
timestamp 1606120353
transform 1 0 9384 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__B
timestamp 1606120353
transform 1 0 11132 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_65_102
timestamp 1606120353
transform 1 0 10488 0 1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_65_107
timestamp 1606120353
transform 1 0 10948 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__nand3_4  _0641_
timestamp 1606120353
transform 1 0 11960 0 1 37536
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__A
timestamp 1606120353
transform 1 0 11776 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_65_111
timestamp 1606120353
transform 1 0 11316 0 1 37536
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_65_115
timestamp 1606120353
transform 1 0 11684 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_65_132
timestamp 1606120353
transform 1 0 13248 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__C
timestamp 1606120353
transform 1 0 13432 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_136
timestamp 1606120353
transform 1 0 13616 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A
timestamp 1606120353
transform 1 0 13800 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_140
timestamp 1606120353
transform 1 0 13984 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1016_
timestamp 1606120353
transform 1 0 14168 0 1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_65_145
timestamp 1606120353
transform 1 0 14444 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A
timestamp 1606120353
transform 1 0 14628 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_149
timestamp 1606120353
transform 1 0 14812 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__B
timestamp 1606120353
transform 1 0 14996 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1606120353
transform 1 0 15180 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_65_154
timestamp 1606120353
transform 1 0 15272 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _1055_
timestamp 1606120353
transform 1 0 16008 0 1 37536
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__B
timestamp 1606120353
transform 1 0 15824 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__D
timestamp 1606120353
transform 1 0 15456 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_158
timestamp 1606120353
transform 1 0 15640 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1606120353
transform -1 0 18860 0 1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__A
timestamp 1606120353
transform 1 0 17756 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_179
timestamp 1606120353
transform 1 0 17572 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_65_183
timestamp 1606120353
transform 1 0 17940 0 1 37536
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_65_189
timestamp 1606120353
transform 1 0 18492 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_67_11
timestamp 1606120353
transform 1 0 2116 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_67_3
timestamp 1606120353
transform 1 0 1380 0 1 38624
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_66_3
timestamp 1606120353
transform 1 0 1380 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1606120353
transform 1 0 1104 0 1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1606120353
transform 1 0 1104 0 -1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_67_22
timestamp 1606120353
transform 1 0 3128 0 1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_67_18
timestamp 1606120353
transform 1 0 2760 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_14
timestamp 1606120353
transform 1 0 2392 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A
timestamp 1606120353
transform 1 0 2208 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__A
timestamp 1606120353
transform 1 0 2576 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__B
timestamp 1606120353
transform 1 0 2944 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1268_
timestamp 1606120353
transform 1 0 1472 0 -1 38624
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_2  FILLER_67_27
timestamp 1606120353
transform 1 0 3588 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_27
timestamp 1606120353
transform 1 0 3588 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_23
timestamp 1606120353
transform 1 0 3220 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A2
timestamp 1606120353
transform 1 0 3404 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A
timestamp 1606120353
transform 1 0 3772 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__B1_N
timestamp 1606120353
transform 1 0 3404 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A1
timestamp 1606120353
transform 1 0 3772 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1606120353
transform 1 0 3956 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1166_
timestamp 1606120353
transform 1 0 3956 0 -1 38624
box 0 -48 1748 592
use sky130_fd_sc_hd__a21bo_4  _0812_
timestamp 1606120353
transform 1 0 4048 0 1 38624
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_67_54
timestamp 1606120353
transform 1 0 6072 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_67_49
timestamp 1606120353
transform 1 0 5612 0 1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_67_45
timestamp 1606120353
transform 1 0 5244 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_66_54
timestamp 1606120353
transform 1 0 6072 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_66_50
timestamp 1606120353
transform 1 0 5704 0 -1 38624
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__C
timestamp 1606120353
transform 1 0 6164 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__B
timestamp 1606120353
transform 1 0 5428 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B
timestamp 1606120353
transform 1 0 5888 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_58
timestamp 1606120353
transform 1 0 6440 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_66_65
timestamp 1606120353
transform 1 0 7084 0 -1 38624
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_66_57
timestamp 1606120353
transform 1 0 6348 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__D
timestamp 1606120353
transform 1 0 6532 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A
timestamp 1606120353
transform 1 0 6256 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__B
timestamp 1606120353
transform 1 0 6624 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1606120353
transform 1 0 6716 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0749_
timestamp 1606120353
transform 1 0 6808 0 -1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__nand3_4  _0759_
timestamp 1606120353
transform 1 0 6808 0 1 38624
box 0 -48 1288 592
use sky130_fd_sc_hd__nand3_4  _0553_
timestamp 1606120353
transform 1 0 8280 0 1 38624
box 0 -48 1288 592
use sky130_fd_sc_hd__nand4_4  _0731_
timestamp 1606120353
transform 1 0 8004 0 -1 38624
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0553__B
timestamp 1606120353
transform 1 0 7820 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0553__C
timestamp 1606120353
transform 1 0 7452 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_71
timestamp 1606120353
transform 1 0 7636 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_76
timestamp 1606120353
transform 1 0 8096 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_67_93
timestamp 1606120353
transform 1 0 9660 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_66_96
timestamp 1606120353
transform 1 0 9936 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_92
timestamp 1606120353
transform 1 0 9568 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__C
timestamp 1606120353
transform 1 0 10120 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__A
timestamp 1606120353
transform 1 0 9752 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1606120353
transform 1 0 9568 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_66_104
timestamp 1606120353
transform 1 0 10672 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_66_100
timestamp 1606120353
transform 1 0 10304 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__B
timestamp 1606120353
transform 1 0 10488 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0597_
timestamp 1606120353
transform 1 0 10764 0 -1 38624
box 0 -48 828 592
use sky130_fd_sc_hd__nand4_4  _0710_
timestamp 1606120353
transform 1 0 9752 0 1 38624
box 0 -48 1564 592
use sky130_fd_sc_hd__fill_2  FILLER_67_116
timestamp 1606120353
transform 1 0 11776 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_67_111
timestamp 1606120353
transform 1 0 11316 0 1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_66_118
timestamp 1606120353
transform 1 0 11960 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_114
timestamp 1606120353
transform 1 0 11592 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__B
timestamp 1606120353
transform 1 0 11776 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__B
timestamp 1606120353
transform 1 0 11592 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__A
timestamp 1606120353
transform 1 0 12144 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__D
timestamp 1606120353
transform 1 0 11960 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_66_123
timestamp 1606120353
transform 1 0 12420 0 -1 38624
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__B
timestamp 1606120353
transform 1 0 12788 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1606120353
transform 1 0 12328 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__or3_4  _1127_
timestamp 1606120353
transform 1 0 12972 0 -1 38624
box 0 -48 828 592
use sky130_fd_sc_hd__nand3_4  _0642_
timestamp 1606120353
transform 1 0 12144 0 1 38624
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_67_138
timestamp 1606120353
transform 1 0 13800 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_134
timestamp 1606120353
transform 1 0 13432 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_142
timestamp 1606120353
transform 1 0 14168 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_138
timestamp 1606120353
transform 1 0 13800 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__B1
timestamp 1606120353
transform 1 0 13616 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__C
timestamp 1606120353
transform 1 0 13984 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A
timestamp 1606120353
transform 1 0 13984 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1013_
timestamp 1606120353
transform 1 0 14168 0 1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_67_154
timestamp 1606120353
transform 1 0 15272 0 1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_67_149
timestamp 1606120353
transform 1 0 14812 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_145
timestamp 1606120353
transform 1 0 14444 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__D
timestamp 1606120353
transform 1 0 14996 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__C
timestamp 1606120353
transform 1 0 14352 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A
timestamp 1606120353
transform 1 0 14628 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1606120353
transform 1 0 15180 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__nand4_4  _1071_
timestamp 1606120353
transform 1 0 14536 0 -1 38624
box 0 -48 1564 592
use sky130_fd_sc_hd__fill_2  FILLER_67_159
timestamp 1606120353
transform 1 0 15732 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_163
timestamp 1606120353
transform 1 0 16100 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__A
timestamp 1606120353
transform 1 0 16284 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A
timestamp 1606120353
transform 1 0 15548 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__C
timestamp 1606120353
transform 1 0 15916 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_174
timestamp 1606120353
transform 1 0 17112 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_167
timestamp 1606120353
transform 1 0 16468 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__D
timestamp 1606120353
transform 1 0 17296 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__A
timestamp 1606120353
transform 1 0 16652 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1046_
timestamp 1606120353
transform 1 0 16836 0 -1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__nand4_4  _1049_
timestamp 1606120353
transform 1 0 16100 0 1 38624
box 0 -48 1564 592
use sky130_fd_sc_hd__fill_2  FILLER_67_180
timestamp 1606120353
transform 1 0 17664 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_66_182
timestamp 1606120353
transform 1 0 17848 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_66_178
timestamp 1606120353
transform 1 0 17480 0 -1 38624
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__B
timestamp 1606120353
transform 1 0 17848 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_188
timestamp 1606120353
transform 1 0 18400 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_184
timestamp 1606120353
transform 1 0 18032 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_66_184
timestamp 1606120353
transform 1 0 18032 0 -1 38624
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__B
timestamp 1606120353
transform 1 0 18216 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1606120353
transform 1 0 17940 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1606120353
transform -1 0 18860 0 1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1606120353
transform -1 0 18860 0 -1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__nand2_4  _0811_
timestamp 1606120353
transform 1 0 2944 0 -1 39712
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1606120353
transform 1 0 1104 0 -1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1606120353
transform 1 0 1380 0 -1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_68_15
timestamp 1606120353
transform 1 0 2484 0 -1 39712
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_68_19
timestamp 1606120353
transform 1 0 2852 0 -1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__nor2_4  _0877_
timestamp 1606120353
transform 1 0 4508 0 -1 39712
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A1
timestamp 1606120353
transform 1 0 4232 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_68_29
timestamp 1606120353
transform 1 0 3772 0 -1 39712
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_68_33
timestamp 1606120353
transform 1 0 4140 0 -1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_68_36
timestamp 1606120353
transform 1 0 4416 0 -1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_68_50
timestamp 1606120353
transform 1 0 5704 0 -1 39712
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_68_46
timestamp 1606120353
transform 1 0 5336 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__A
timestamp 1606120353
transform 1 0 5520 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_68_62
timestamp 1606120353
transform 1 0 6808 0 -1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_68_57
timestamp 1606120353
transform 1 0 6348 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_68_54
timestamp 1606120353
transform 1 0 6072 0 -1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__B1
timestamp 1606120353
transform 1 0 6532 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A2
timestamp 1606120353
transform 1 0 6164 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1606120353
transform 1 0 6716 0 -1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__nor2_4  _0575_
timestamp 1606120353
transform 1 0 7084 0 -1 39712
box 0 -48 828 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 8740 0 -1 39712
box 0 -48 1840 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1606120353
transform 1 0 8556 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0553__A
timestamp 1606120353
transform 1 0 8188 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_68_74
timestamp 1606120353
transform 1 0 7912 0 -1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_68_79
timestamp 1606120353
transform 1 0 8372 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__nand2_4  _1031_
timestamp 1606120353
transform 1 0 10764 0 -1 39712
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_68_103
timestamp 1606120353
transform 1 0 10580 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1272_
timestamp 1606120353
transform 1 0 12512 0 -1 39712
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1606120353
transform 1 0 12328 0 -1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__C
timestamp 1606120353
transform 1 0 11868 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_68_114
timestamp 1606120353
transform 1 0 11592 0 -1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_68_119
timestamp 1606120353
transform 1 0 12052 0 -1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_68_123
timestamp 1606120353
transform 1 0 12420 0 -1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A1
timestamp 1606120353
transform 1 0 14444 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A4
timestamp 1606120353
transform 1 0 14812 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_68_143
timestamp 1606120353
transform 1 0 14260 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_68_147
timestamp 1606120353
transform 1 0 14628 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_68_151
timestamp 1606120353
transform 1 0 14996 0 -1 39712
box 0 -48 368 592
use sky130_fd_sc_hd__nand4_4  _1092_
timestamp 1606120353
transform 1 0 15548 0 -1 39712
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__B
timestamp 1606120353
transform 1 0 15364 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__D
timestamp 1606120353
transform 1 0 17296 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_68_174
timestamp 1606120353
transform 1 0 17112 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1606120353
transform -1 0 18860 0 -1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1606120353
transform 1 0 17940 0 -1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_68_178
timestamp 1606120353
transform 1 0 17480 0 -1 39712
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_68_182
timestamp 1606120353
transform 1 0 17848 0 -1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_68_184
timestamp 1606120353
transform 1 0 18032 0 -1 39712
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1606120353
transform 1 0 1104 0 1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1606120353
transform 1 0 1380 0 1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_69_15
timestamp 1606120353
transform 1 0 2484 0 1 39712
box 0 -48 736 592
use sky130_fd_sc_hd__a21oi_4  _0878_
timestamp 1606120353
transform 1 0 4232 0 1 39712
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1606120353
transform 1 0 3956 0 1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A2
timestamp 1606120353
transform 1 0 3772 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__B1
timestamp 1606120353
transform 1 0 3404 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_23
timestamp 1606120353
transform 1 0 3220 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_27
timestamp 1606120353
transform 1 0 3588 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_32
timestamp 1606120353
transform 1 0 4048 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__a41oi_4  _0761_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 6164 0 1 39712
box 0 -48 2024 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A1
timestamp 1606120353
transform 1 0 5980 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A4
timestamp 1606120353
transform 1 0 5612 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_47
timestamp 1606120353
transform 1 0 5428 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_51
timestamp 1606120353
transform 1 0 5796 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__A
timestamp 1606120353
transform 1 0 8372 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__B
timestamp 1606120353
transform 1 0 8740 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_77
timestamp 1606120353
transform 1 0 8188 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_81
timestamp 1606120353
transform 1 0 8556 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_69_85
timestamp 1606120353
transform 1 0 8924 0 1 39712
box 0 -48 368 592
use sky130_fd_sc_hd__nand2_4  _0757_
timestamp 1606120353
transform 1 0 9660 0 1 39712
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1606120353
transform 1 0 9568 0 1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A
timestamp 1606120353
transform 1 0 9384 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__C
timestamp 1606120353
transform 1 0 10764 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A
timestamp 1606120353
transform 1 0 11132 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_69_89
timestamp 1606120353
transform 1 0 9292 0 1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_69_102
timestamp 1606120353
transform 1 0 10488 0 1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_69_107
timestamp 1606120353
transform 1 0 10948 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__nand3_4  _0643_
timestamp 1606120353
transform 1 0 11868 0 1 39712
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__A
timestamp 1606120353
transform 1 0 11684 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_69_111
timestamp 1606120353
transform 1 0 11316 0 1 39712
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_69_131
timestamp 1606120353
transform 1 0 13156 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_135
timestamp 1606120353
transform 1 0 13524 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__B
timestamp 1606120353
transform 1 0 13340 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__A
timestamp 1606120353
transform 1 0 13708 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0598_
timestamp 1606120353
transform 1 0 13892 0 1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_69_142
timestamp 1606120353
transform 1 0 14168 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0598__A
timestamp 1606120353
transform 1 0 14352 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_146
timestamp 1606120353
transform 1 0 14536 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_69_150
timestamp 1606120353
transform 1 0 14904 0 1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A2
timestamp 1606120353
transform 1 0 14720 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1606120353
transform 1 0 15180 0 1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_69_154
timestamp 1606120353
transform 1 0 15272 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _1085_
timestamp 1606120353
transform 1 0 16008 0 1 39712
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__C
timestamp 1606120353
transform 1 0 15824 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A3
timestamp 1606120353
transform 1 0 15456 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_158
timestamp 1606120353
transform 1 0 15640 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1606120353
transform -1 0 18860 0 1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__A
timestamp 1606120353
transform 1 0 17756 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_179
timestamp 1606120353
transform 1 0 17572 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_69_183
timestamp 1606120353
transform 1 0 17940 0 1 39712
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_69_189
timestamp 1606120353
transform 1 0 18492 0 1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1606120353
transform 1 0 1104 0 -1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__D
timestamp 1606120353
transform 1 0 1564 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__CLK
timestamp 1606120353
transform 1 0 1932 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_3
timestamp 1606120353
transform 1 0 1380 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_7
timestamp 1606120353
transform 1 0 1748 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_70_11
timestamp 1606120353
transform 1 0 2116 0 -1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__inv_8  _0797_
timestamp 1606120353
transform 1 0 4784 0 -1 40800
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__B1
timestamp 1606120353
transform 1 0 4600 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__B1
timestamp 1606120353
transform 1 0 4232 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_70_23
timestamp 1606120353
transform 1 0 3220 0 -1 40800
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_70_31
timestamp 1606120353
transform 1 0 3956 0 -1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_70_36
timestamp 1606120353
transform 1 0 4416 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_49
timestamp 1606120353
transform 1 0 5612 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__D
timestamp 1606120353
transform 1 0 5796 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_53
timestamp 1606120353
transform 1 0 5980 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_57
timestamp 1606120353
transform 1 0 6348 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A3
timestamp 1606120353
transform 1 0 6164 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A
timestamp 1606120353
transform 1 0 6532 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1606120353
transform 1 0 6716 0 -1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_70_62
timestamp 1606120353
transform 1 0 6808 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A2
timestamp 1606120353
transform 1 0 6992 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_66
timestamp 1606120353
transform 1 0 7176 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _0551_
timestamp 1606120353
transform 1 0 8372 0 -1 40800
box 0 -48 1564 592
use sky130_fd_sc_hd__buf_1  _1082_
timestamp 1606120353
transform 1 0 7360 0 -1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__C
timestamp 1606120353
transform 1 0 8188 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__A
timestamp 1606120353
transform 1 0 7820 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_71
timestamp 1606120353
transform 1 0 7636 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_75
timestamp 1606120353
transform 1 0 8004 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__or3_4  _1109_
timestamp 1606120353
transform 1 0 10764 0 -1 40800
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0541__A
timestamp 1606120353
transform 1 0 10120 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0541__C
timestamp 1606120353
transform 1 0 10488 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_96
timestamp 1606120353
transform 1 0 9936 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_100
timestamp 1606120353
transform 1 0 10304 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_70_104
timestamp 1606120353
transform 1 0 10672 0 -1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__nor2_4  _1060_
timestamp 1606120353
transform 1 0 12512 0 -1 40800
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1606120353
transform 1 0 12328 0 -1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__A
timestamp 1606120353
transform 1 0 11960 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_70_114
timestamp 1606120353
transform 1 0 11592 0 -1 40800
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_70_120
timestamp 1606120353
transform 1 0 12144 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_70_123
timestamp 1606120353
transform 1 0 12420 0 -1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__a41oi_4  _1061_
timestamp 1606120353
transform 1 0 14076 0 -1 40800
box 0 -48 2024 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A
timestamp 1606120353
transform 1 0 13524 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__B
timestamp 1606120353
transform 1 0 13892 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_133
timestamp 1606120353
transform 1 0 13340 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_137
timestamp 1606120353
transform 1 0 13708 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1014_
timestamp 1606120353
transform 1 0 16836 0 -1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__A
timestamp 1606120353
transform 1 0 16284 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__A
timestamp 1606120353
transform 1 0 16652 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__D
timestamp 1606120353
transform 1 0 17296 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_163
timestamp 1606120353
transform 1 0 16100 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_167
timestamp 1606120353
transform 1 0 16468 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_174
timestamp 1606120353
transform 1 0 17112 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1606120353
transform -1 0 18860 0 -1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1606120353
transform 1 0 17940 0 -1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_70_178
timestamp 1606120353
transform 1 0 17480 0 -1 40800
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_70_182
timestamp 1606120353
transform 1 0 17848 0 -1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_70_184
timestamp 1606120353
transform 1 0 18032 0 -1 40800
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1274_
timestamp 1606120353
transform 1 0 1472 0 1 40800
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1606120353
transform 1 0 1104 0 1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_71_3
timestamp 1606120353
transform 1 0 1380 0 1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__o21ai_4  _0847_
timestamp 1606120353
transform 1 0 4692 0 1 40800
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1606120353
transform 1 0 3956 0 1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A1
timestamp 1606120353
transform 1 0 4508 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A2
timestamp 1606120353
transform 1 0 3772 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_71_23
timestamp 1606120353
transform 1 0 3220 0 1 40800
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILLER_71_32
timestamp 1606120353
transform 1 0 4048 0 1 40800
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_71_36
timestamp 1606120353
transform 1 0 4416 0 1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__o21ai_4  _0798_
timestamp 1606120353
transform 1 0 6624 0 1 40800
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__B1
timestamp 1606120353
transform 1 0 6440 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A2
timestamp 1606120353
transform 1 0 6072 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_52
timestamp 1606120353
transform 1 0 5888 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_56
timestamp 1606120353
transform 1 0 6256 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1075_
timestamp 1606120353
transform 1 0 8556 0 1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0552__C
timestamp 1606120353
transform 1 0 9016 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0552__A
timestamp 1606120353
transform 1 0 8372 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0552__B
timestamp 1606120353
transform 1 0 8004 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_73
timestamp 1606120353
transform 1 0 7820 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_77
timestamp 1606120353
transform 1 0 8188 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_84
timestamp 1606120353
transform 1 0 8832 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_88
timestamp 1606120353
transform 1 0 9200 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _0541_
timestamp 1606120353
transform 1 0 9660 0 1 40800
box 0 -48 1564 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1606120353
transform 1 0 9568 0 1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0541__D
timestamp 1606120353
transform 1 0 9384 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_110
timestamp 1606120353
transform 1 0 11224 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _0645_
timestamp 1606120353
transform 1 0 11960 0 1 40800
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__C
timestamp 1606120353
transform 1 0 11776 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__C
timestamp 1606120353
transform 1 0 11408 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_114
timestamp 1606120353
transform 1 0 11592 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_135
timestamp 1606120353
transform 1 0 13524 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_139
timestamp 1606120353
transform 1 0 13892 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__A
timestamp 1606120353
transform 1 0 13708 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_71_143
timestamp 1606120353
transform 1 0 14260 0 1 40800
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A
timestamp 1606120353
transform 1 0 14076 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__C
timestamp 1606120353
transform 1 0 14628 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_149
timestamp 1606120353
transform 1 0 14812 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__B
timestamp 1606120353
transform 1 0 14996 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_154
timestamp 1606120353
transform 1 0 15272 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1606120353
transform 1 0 15180 0 1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__nand4_4  _1088_
timestamp 1606120353
transform 1 0 15824 0 1 40800
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A
timestamp 1606120353
transform 1 0 15456 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_158
timestamp 1606120353
transform 1 0 15640 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1606120353
transform -1 0 18860 0 1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__B
timestamp 1606120353
transform 1 0 17572 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__B
timestamp 1606120353
transform 1 0 17940 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_177
timestamp 1606120353
transform 1 0 17388 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_181
timestamp 1606120353
transform 1 0 17756 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_71_185
timestamp 1606120353
transform 1 0 18124 0 1 40800
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_71_189
timestamp 1606120353
transform 1 0 18492 0 1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1275_
timestamp 1606120353
transform 1 0 1472 0 1 41888
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1606120353
transform 1 0 1104 0 -1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1606120353
transform 1 0 1104 0 1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__D
timestamp 1606120353
transform 1 0 1564 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__CLK
timestamp 1606120353
transform 1 0 1932 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_3
timestamp 1606120353
transform 1 0 1380 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_7
timestamp 1606120353
transform 1 0 1748 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_72_11
timestamp 1606120353
transform 1 0 2116 0 -1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_73_3
timestamp 1606120353
transform 1 0 1380 0 1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__D
timestamp 1606120353
transform 1 0 3404 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__CLK
timestamp 1606120353
transform 1 0 3404 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_23
timestamp 1606120353
transform 1 0 3220 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_73_23
timestamp 1606120353
transform 1 0 3220 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_73_27
timestamp 1606120353
transform 1 0 3588 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1606120353
transform 1 0 3956 0 1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__B1
timestamp 1606120353
transform 1 0 3772 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_72_33
timestamp 1606120353
transform 1 0 4140 0 -1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_73_32
timestamp 1606120353
transform 1 0 4048 0 1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_72_27
timestamp 1606120353
transform 1 0 3588 0 -1 41888
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_73_37
timestamp 1606120353
transform 1 0 4508 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_36
timestamp 1606120353
transform 1 0 4416 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__B2
timestamp 1606120353
transform 1 0 4232 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__A1
timestamp 1606120353
transform 1 0 4324 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A1
timestamp 1606120353
transform 1 0 4600 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__A2
timestamp 1606120353
transform 1 0 4692 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__a22oi_4  _0801_
timestamp 1606120353
transform 1 0 4876 0 1 41888
box 0 -48 1564 592
use sky130_fd_sc_hd__o21ai_4  _0799_
timestamp 1606120353
transform 1 0 4784 0 -1 41888
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1606120353
transform 1 0 6716 0 -1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__C1
timestamp 1606120353
transform 1 0 7084 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A1
timestamp 1606120353
transform 1 0 6716 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0552__D
timestamp 1606120353
transform 1 0 7176 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A1
timestamp 1606120353
transform 1 0 6532 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_72_53
timestamp 1606120353
transform 1 0 5980 0 -1 41888
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILLER_72_62
timestamp 1606120353
transform 1 0 6808 0 -1 41888
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_73_58
timestamp 1606120353
transform 1 0 6440 0 1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_73_63
timestamp 1606120353
transform 1 0 6900 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_73_67
timestamp 1606120353
transform 1 0 7268 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_76
timestamp 1606120353
transform 1 0 8096 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_72
timestamp 1606120353
transform 1 0 7728 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_68
timestamp 1606120353
transform 1 0 7360 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__A1
timestamp 1606120353
transform 1 0 7544 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__B1
timestamp 1606120353
transform 1 0 7912 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__A2
timestamp 1606120353
transform 1 0 7452 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_73_88
timestamp 1606120353
transform 1 0 9200 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_73_84
timestamp 1606120353
transform 1 0 8832 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A2
timestamp 1606120353
transform 1 0 9016 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__D1
timestamp 1606120353
transform 1 0 8280 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0676_
timestamp 1606120353
transform 1 0 7636 0 1 41888
box 0 -48 1196 592
use sky130_fd_sc_hd__nand4_4  _0552_
timestamp 1606120353
transform 1 0 8464 0 -1 41888
box 0 -48 1564 592
use sky130_fd_sc_hd__fill_2  FILLER_73_96
timestamp 1606120353
transform 1 0 9936 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_97
timestamp 1606120353
transform 1 0 10028 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__C
timestamp 1606120353
transform 1 0 9384 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__A
timestamp 1606120353
transform 1 0 10120 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0541__B
timestamp 1606120353
transform 1 0 10212 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1606120353
transform 1 0 9568 0 1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0584_
timestamp 1606120353
transform 1 0 9660 0 1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_73_100
timestamp 1606120353
transform 1 0 10304 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_101
timestamp 1606120353
transform 1 0 10396 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__A
timestamp 1606120353
transform 1 0 10580 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__A
timestamp 1606120353
transform 1 0 10488 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _1020_
timestamp 1606120353
transform 1 0 10764 0 -1 41888
box 0 -48 828 592
use sky130_fd_sc_hd__nand3_4  _0661_
timestamp 1606120353
transform 1 0 10672 0 1 41888
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_73_118
timestamp 1606120353
transform 1 0 11960 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_120
timestamp 1606120353
transform 1 0 12144 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_72_114
timestamp 1606120353
transform 1 0 11592 0 -1 41888
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__B
timestamp 1606120353
transform 1 0 11960 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__C
timestamp 1606120353
transform 1 0 12144 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_73_131
timestamp 1606120353
transform 1 0 13156 0 1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_73_126
timestamp 1606120353
transform 1 0 12696 0 1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_73_122
timestamp 1606120353
transform 1 0 12328 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__A1
timestamp 1606120353
transform 1 0 12972 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__D
timestamp 1606120353
transform 1 0 12512 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1606120353
transform 1 0 12328 0 -1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__o21ai_4  _1131_
timestamp 1606120353
transform 1 0 13248 0 1 41888
box 0 -48 1196 592
use sky130_fd_sc_hd__nand3_4  _0644_
timestamp 1606120353
transform 1 0 12420 0 -1 41888
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_72_141
timestamp 1606120353
transform 1 0 14076 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_137
timestamp 1606120353
transform 1 0 13708 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__B1
timestamp 1606120353
transform 1 0 14260 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A1
timestamp 1606120353
transform 1 0 13892 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A
timestamp 1606120353
transform 1 0 14628 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_145
timestamp 1606120353
transform 1 0 14444 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_73_145
timestamp 1606120353
transform 1 0 14444 0 1 41888
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__C
timestamp 1606120353
transform 1 0 14904 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__D
timestamp 1606120353
transform 1 0 14996 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_149
timestamp 1606120353
transform 1 0 14812 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_73_149
timestamp 1606120353
transform 1 0 14812 0 1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1606120353
transform 1 0 15180 0 1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_73_152
timestamp 1606120353
transform 1 0 15088 0 1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_73_154
timestamp 1606120353
transform 1 0 15272 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _1022_
timestamp 1606120353
transform 1 0 15180 0 -1 41888
box 0 -48 1564 592
use sky130_fd_sc_hd__nand4_4  _1083_
timestamp 1606120353
transform 1 0 15824 0 1 41888
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__D
timestamp 1606120353
transform 1 0 15456 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__A
timestamp 1606120353
transform 1 0 16928 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__C
timestamp 1606120353
transform 1 0 17296 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_170
timestamp 1606120353
transform 1 0 16744 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_174
timestamp 1606120353
transform 1 0 17112 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_73_158
timestamp 1606120353
transform 1 0 15640 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_73_181
timestamp 1606120353
transform 1 0 17756 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_73_177
timestamp 1606120353
transform 1 0 17388 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_72_182
timestamp 1606120353
transform 1 0 17848 0 -1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_72_178
timestamp 1606120353
transform 1 0 17480 0 -1 41888
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__B
timestamp 1606120353
transform 1 0 17572 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_73_185
timestamp 1606120353
transform 1 0 18124 0 1 41888
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_72_184
timestamp 1606120353
transform 1 0 18032 0 -1 41888
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__C
timestamp 1606120353
transform 1 0 17940 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1606120353
transform 1 0 17940 0 -1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_73_189
timestamp 1606120353
transform 1 0 18492 0 1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1606120353
transform -1 0 18860 0 1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1606120353
transform -1 0 18860 0 -1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1606120353
transform 1 0 1104 0 -1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__D
timestamp 1606120353
transform 1 0 1564 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__D
timestamp 1606120353
transform 1 0 1932 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__CLK
timestamp 1606120353
transform 1 0 2300 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_3
timestamp 1606120353
transform 1 0 1380 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_7
timestamp 1606120353
transform 1 0 1748 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_11
timestamp 1606120353
transform 1 0 2116 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_74_15
timestamp 1606120353
transform 1 0 2484 0 -1 42976
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1149_
timestamp 1606120353
transform 1 0 3404 0 -1 42976
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_2  FILLER_74_23
timestamp 1606120353
transform 1 0 3220 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_74_44
timestamp 1606120353
transform 1 0 5152 0 -1 42976
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_74_48
timestamp 1606120353
transform 1 0 5520 0 -1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_74_51
timestamp 1606120353
transform 1 0 5796 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__B
timestamp 1606120353
transform 1 0 5612 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_74_55
timestamp 1606120353
transform 1 0 6164 0 -1 42976
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__D
timestamp 1606120353
transform 1 0 5980 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__A
timestamp 1606120353
transform 1 0 6532 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_62
timestamp 1606120353
transform 1 0 6808 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A2
timestamp 1606120353
transform 1 0 6992 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1606120353
transform 1 0 6716 0 -1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_74_66
timestamp 1606120353
transform 1 0 7176 0 -1 42976
box 0 -48 368 592
use sky130_fd_sc_hd__a2111oi_4  _0562_
timestamp 1606120353
transform 1 0 7912 0 -1 42976
box 0 -48 2024 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__B1_N
timestamp 1606120353
transform 1 0 7636 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_74_70
timestamp 1606120353
transform 1 0 7544 0 -1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_74_73
timestamp 1606120353
transform 1 0 7820 0 -1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__and3_4  _0665_
timestamp 1606120353
transform 1 0 10764 0 -1 42976
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__B
timestamp 1606120353
transform 1 0 10580 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__C
timestamp 1606120353
transform 1 0 10212 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_74_96
timestamp 1606120353
transform 1 0 9936 0 -1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_74_101
timestamp 1606120353
transform 1 0 10396 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1130_
timestamp 1606120353
transform 1 0 12972 0 -1 42976
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1606120353
transform 1 0 12328 0 -1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A2
timestamp 1606120353
transform 1 0 12788 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__A2
timestamp 1606120353
transform 1 0 12144 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__B
timestamp 1606120353
transform 1 0 11776 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_114
timestamp 1606120353
transform 1 0 11592 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_118
timestamp 1606120353
transform 1 0 11960 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_74_123
timestamp 1606120353
transform 1 0 12420 0 -1 42976
box 0 -48 368 592
use sky130_fd_sc_hd__nand4_4  _1077_
timestamp 1606120353
transform 1 0 14904 0 -1 42976
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A
timestamp 1606120353
transform 1 0 14720 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__B
timestamp 1606120353
transform 1 0 14352 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_142
timestamp 1606120353
transform 1 0 14168 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_146
timestamp 1606120353
transform 1 0 14536 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__C
timestamp 1606120353
transform 1 0 16652 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__D
timestamp 1606120353
transform 1 0 17020 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_167
timestamp 1606120353
transform 1 0 16468 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_171
timestamp 1606120353
transform 1 0 16836 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_175
timestamp 1606120353
transform 1 0 17204 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1606120353
transform -1 0 18860 0 -1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1606120353
transform 1 0 17940 0 -1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__D
timestamp 1606120353
transform 1 0 17388 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_74_179
timestamp 1606120353
transform 1 0 17572 0 -1 42976
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_74_184
timestamp 1606120353
transform 1 0 18032 0 -1 42976
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1276_
timestamp 1606120353
transform 1 0 1472 0 1 42976
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1606120353
transform 1 0 1104 0 1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_75_3
timestamp 1606120353
transform 1 0 1380 0 1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__nand2_4  _0802_
timestamp 1606120353
transform 1 0 4048 0 1 42976
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1606120353
transform 1 0 3956 0 1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A1
timestamp 1606120353
transform 1 0 3772 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__B
timestamp 1606120353
transform 1 0 3404 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__B1_N
timestamp 1606120353
transform 1 0 5060 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_23
timestamp 1606120353
transform 1 0 3220 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_27
timestamp 1606120353
transform 1 0 3588 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_41
timestamp 1606120353
transform 1 0 4876 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _0837_
timestamp 1606120353
transform 1 0 5612 0 1 42976
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__C
timestamp 1606120353
transform 1 0 5428 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_45
timestamp 1606120353
transform 1 0 5244 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_66
timestamp 1606120353
transform 1 0 7176 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0670_
timestamp 1606120353
transform 1 0 8004 0 1 42976
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A1
timestamp 1606120353
transform 1 0 7360 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__B
timestamp 1606120353
transform 1 0 9016 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__B1
timestamp 1606120353
transform 1 0 7728 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_70
timestamp 1606120353
transform 1 0 7544 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_75_74
timestamp 1606120353
transform 1 0 7912 0 1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_75_84
timestamp 1606120353
transform 1 0 8832 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_88
timestamp 1606120353
transform 1 0 9200 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__nand3_4  _0675_
timestamp 1606120353
transform 1 0 9660 0 1 42976
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1606120353
transform 1 0 9568 0 1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__A
timestamp 1606120353
transform 1 0 9384 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__B
timestamp 1606120353
transform 1 0 11132 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_107
timestamp 1606120353
transform 1 0 10948 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0646_
timestamp 1606120353
transform 1 0 12420 0 1 42976
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__A
timestamp 1606120353
transform 1 0 12236 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__B
timestamp 1606120353
transform 1 0 11868 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__A
timestamp 1606120353
transform 1 0 11500 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_111
timestamp 1606120353
transform 1 0 11316 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_115
timestamp 1606120353
transform 1 0 11684 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_119
timestamp 1606120353
transform 1 0 12052 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_132
timestamp 1606120353
transform 1 0 13248 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_136
timestamp 1606120353
transform 1 0 13616 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__D
timestamp 1606120353
transform 1 0 13432 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__D
timestamp 1606120353
transform 1 0 13800 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0600_
timestamp 1606120353
transform 1 0 13984 0 1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_75_143
timestamp 1606120353
transform 1 0 14260 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_75_147
timestamp 1606120353
transform 1 0 14628 0 1 42976
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0600__A
timestamp 1606120353
transform 1 0 14444 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__C
timestamp 1606120353
transform 1 0 14996 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_75_154
timestamp 1606120353
transform 1 0 15272 0 1 42976
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1606120353
transform 1 0 15180 0 1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__nand4_4  _1074_
timestamp 1606120353
transform 1 0 16008 0 1 42976
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__B
timestamp 1606120353
transform 1 0 15640 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_160
timestamp 1606120353
transform 1 0 15824 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1606120353
transform -1 0 18860 0 1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__B
timestamp 1606120353
transform 1 0 17756 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_179
timestamp 1606120353
transform 1 0 17572 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_75_183
timestamp 1606120353
transform 1 0 17940 0 1 42976
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_75_189
timestamp 1606120353
transform 1 0 18492 0 1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1277_
timestamp 1606120353
transform 1 0 1472 0 -1 44064
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1606120353
transform 1 0 1104 0 -1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_76_3
timestamp 1606120353
transform 1 0 1380 0 -1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__a21bo_4  _0803_
timestamp 1606120353
transform 1 0 3956 0 -1 44064
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A2
timestamp 1606120353
transform 1 0 3772 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A
timestamp 1606120353
transform 1 0 3404 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_23
timestamp 1606120353
transform 1 0 3220 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_27
timestamp 1606120353
transform 1 0 3588 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_76_44
timestamp 1606120353
transform 1 0 5152 0 -1 44064
box 0 -48 368 592
use sky130_fd_sc_hd__o21ai_4  _0800_
timestamp 1606120353
transform 1 0 6900 0 -1 44064
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1606120353
transform 1 0 6716 0 -1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__B1
timestamp 1606120353
transform 1 0 6532 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A
timestamp 1606120353
transform 1 0 5612 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A2
timestamp 1606120353
transform 1 0 6164 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_76_48
timestamp 1606120353
transform 1 0 5520 0 -1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_76_51
timestamp 1606120353
transform 1 0 5796 0 -1 44064
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_76_57
timestamp 1606120353
transform 1 0 6348 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_76_62
timestamp 1606120353
transform 1 0 6808 0 -1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0531__B
timestamp 1606120353
transform 1 0 8740 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A1
timestamp 1606120353
transform 1 0 8280 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_76
timestamp 1606120353
transform 1 0 8096 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_76_80
timestamp 1606120353
transform 1 0 8464 0 -1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_76_85
timestamp 1606120353
transform 1 0 8924 0 -1 44064
box 0 -48 368 592
use sky130_fd_sc_hd__nand3_4  _0677_
timestamp 1606120353
transform 1 0 9936 0 -1 44064
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__A1
timestamp 1606120353
transform 1 0 9660 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__B
timestamp 1606120353
transform 1 0 9292 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_91
timestamp 1606120353
transform 1 0 9476 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_76_95
timestamp 1606120353
transform 1 0 9844 0 -1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_76_110
timestamp 1606120353
transform 1 0 11224 0 -1 44064
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_76_120
timestamp 1606120353
transform 1 0 12144 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_116
timestamp 1606120353
transform 1 0 11776 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__C
timestamp 1606120353
transform 1 0 11960 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__A
timestamp 1606120353
transform 1 0 11592 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_127
timestamp 1606120353
transform 1 0 12788 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_123
timestamp 1606120353
transform 1 0 12420 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__C
timestamp 1606120353
transform 1 0 12604 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__B1
timestamp 1606120353
transform 1 0 12972 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1606120353
transform 1 0 12328 0 -1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1178_
timestamp 1606120353
transform 1 0 13156 0 -1 44064
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1606120353
transform 1 0 15088 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_150
timestamp 1606120353
transform 1 0 14904 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_154
timestamp 1606120353
transform 1 0 15272 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _1065_
timestamp 1606120353
transform 1 0 15640 0 -1 44064
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__A
timestamp 1606120353
transform 1 0 15456 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_175
timestamp 1606120353
transform 1 0 17204 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1606120353
transform -1 0 18860 0 -1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1606120353
transform 1 0 17940 0 -1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__C
timestamp 1606120353
transform 1 0 17388 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_76_179
timestamp 1606120353
transform 1 0 17572 0 -1 44064
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_76_184
timestamp 1606120353
transform 1 0 18032 0 -1 44064
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1606120353
transform 1 0 1104 0 1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__CLK
timestamp 1606120353
transform 1 0 1564 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_3
timestamp 1606120353
transform 1 0 1380 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_77_7
timestamp 1606120353
transform 1 0 1748 0 1 44064
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_77_19
timestamp 1606120353
transform 1 0 2852 0 1 44064
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__B1
timestamp 1606120353
transform 1 0 3404 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_27
timestamp 1606120353
transform 1 0 3588 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A1
timestamp 1606120353
transform 1 0 3772 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_32
timestamp 1606120353
transform 1 0 4048 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A2
timestamp 1606120353
transform 1 0 4232 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1606120353
transform 1 0 3956 0 1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_77_36
timestamp 1606120353
transform 1 0 4416 0 1 44064
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_77_42
timestamp 1606120353
transform 1 0 4968 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A1
timestamp 1606120353
transform 1 0 4784 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A2
timestamp 1606120353
transform 1 0 5152 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0838_
timestamp 1606120353
transform 1 0 5336 0 1 44064
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A2
timestamp 1606120353
transform 1 0 7084 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__B1
timestamp 1606120353
transform 1 0 6716 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_59
timestamp 1606120353
transform 1 0 6532 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_63
timestamp 1606120353
transform 1 0 6900 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__a21oi_4  _0769_
timestamp 1606120353
transform 1 0 7268 0 1 44064
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0531__A
timestamp 1606120353
transform 1 0 8740 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_77_80
timestamp 1606120353
transform 1 0 8464 0 1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_77_85
timestamp 1606120353
transform 1 0 8924 0 1 44064
box 0 -48 368 592
use sky130_fd_sc_hd__o21a_4  _0561_
timestamp 1606120353
transform 1 0 9660 0 1 44064
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1606120353
transform 1 0 9568 0 1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__B1
timestamp 1606120353
transform 1 0 9384 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__A
timestamp 1606120353
transform 1 0 10948 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_77_89
timestamp 1606120353
transform 1 0 9292 0 1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_77_105
timestamp 1606120353
transform 1 0 10764 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_77_109
timestamp 1606120353
transform 1 0 11132 0 1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__nand3_4  _0658_
timestamp 1606120353
transform 1 0 11592 0 1 44064
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__D
timestamp 1606120353
transform 1 0 13156 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__C
timestamp 1606120353
transform 1 0 11408 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_77_128
timestamp 1606120353
transform 1 0 12880 0 1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__nand2_4  _0647_
timestamp 1606120353
transform 1 0 13616 0 1 44064
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1606120353
transform 1 0 15180 0 1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__A
timestamp 1606120353
transform 1 0 14628 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__B
timestamp 1606120353
transform 1 0 14996 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_77_133
timestamp 1606120353
transform 1 0 13340 0 1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_77_145
timestamp 1606120353
transform 1 0 14444 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_149
timestamp 1606120353
transform 1 0 14812 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_77_154
timestamp 1606120353
transform 1 0 15272 0 1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__nand4_4  _1059_
timestamp 1606120353
transform 1 0 16100 0 1 44064
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__C
timestamp 1606120353
transform 1 0 15916 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__B
timestamp 1606120353
transform 1 0 15548 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_159
timestamp 1606120353
transform 1 0 15732 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1606120353
transform -1 0 18860 0 1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__B
timestamp 1606120353
transform 1 0 17848 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_180
timestamp 1606120353
transform 1 0 17664 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_77_184
timestamp 1606120353
transform 1 0 18032 0 1 44064
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1606120353
transform 1 0 1104 0 -1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__D
timestamp 1606120353
transform 1 0 1564 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__CLK
timestamp 1606120353
transform 1 0 1932 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_3
timestamp 1606120353
transform 1 0 1380 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_7
timestamp 1606120353
transform 1 0 1748 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_78_11
timestamp 1606120353
transform 1 0 2116 0 -1 45152
box 0 -48 1104 592
use sky130_fd_sc_hd__a21oi_4  _0876_
timestamp 1606120353
transform 1 0 4140 0 -1 45152
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_8  FILLER_78_23
timestamp 1606120353
transform 1 0 3220 0 -1 45152
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_78_31
timestamp 1606120353
transform 1 0 3956 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0780_
timestamp 1606120353
transform 1 0 6808 0 -1 45152
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1606120353
transform 1 0 6716 0 -1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__B
timestamp 1606120353
transform 1 0 5520 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A1
timestamp 1606120353
transform 1 0 6532 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__B1
timestamp 1606120353
transform 1 0 5888 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_46
timestamp 1606120353
transform 1 0 5336 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_50
timestamp 1606120353
transform 1 0 5704 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_78_54
timestamp 1606120353
transform 1 0 6072 0 -1 45152
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_78_58
timestamp 1606120353
transform 1 0 6440 0 -1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__nor2_4  _0531_
timestamp 1606120353
transform 1 0 8740 0 -1 45152
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__C
timestamp 1606120353
transform 1 0 8096 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_74
timestamp 1606120353
transform 1 0 7912 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_78_78
timestamp 1606120353
transform 1 0 8280 0 -1 45152
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_78_82
timestamp 1606120353
transform 1 0 8648 0 -1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__nand3_4  _0656_
timestamp 1606120353
transform 1 0 10304 0 -1 45152
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__A2
timestamp 1606120353
transform 1 0 9752 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__A
timestamp 1606120353
transform 1 0 10120 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_92
timestamp 1606120353
transform 1 0 9568 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_96
timestamp 1606120353
transform 1 0 9936 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_118
timestamp 1606120353
transform 1 0 11960 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_114
timestamp 1606120353
transform 1 0 11592 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__B
timestamp 1606120353
transform 1 0 12144 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__A
timestamp 1606120353
transform 1 0 11776 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_127
timestamp 1606120353
transform 1 0 12788 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_123
timestamp 1606120353
transform 1 0 12420 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__D
timestamp 1606120353
transform 1 0 12972 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__C
timestamp 1606120353
transform 1 0 12604 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1606120353
transform 1 0 12328 0 -1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1179_
timestamp 1606120353
transform 1 0 13156 0 -1 45152
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__D
timestamp 1606120353
transform 1 0 15088 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_150
timestamp 1606120353
transform 1 0 14904 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_154
timestamp 1606120353
transform 1 0 15272 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _1090_
timestamp 1606120353
transform 1 0 15640 0 -1 45152
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__A
timestamp 1606120353
transform 1 0 15456 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_175
timestamp 1606120353
transform 1 0 17204 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1606120353
transform -1 0 18860 0 -1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1606120353
transform 1 0 17940 0 -1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A2
timestamp 1606120353
transform 1 0 17388 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_78_179
timestamp 1606120353
transform 1 0 17572 0 -1 45152
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_78_184
timestamp 1606120353
transform 1 0 18032 0 -1 45152
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1278_
timestamp 1606120353
transform 1 0 1472 0 1 45152
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1606120353
transform 1 0 1104 0 1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1606120353
transform 1 0 1104 0 -1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__D
timestamp 1606120353
transform 1 0 1564 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__CLK
timestamp 1606120353
transform 1 0 1932 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_79_3
timestamp 1606120353
transform 1 0 1380 0 1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1606120353
transform 1 0 1380 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_80_7
timestamp 1606120353
transform 1 0 1748 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_80_11
timestamp 1606120353
transform 1 0 2116 0 -1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_80_23
timestamp 1606120353
transform 1 0 3220 0 -1 46240
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_79_32
timestamp 1606120353
transform 1 0 4048 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_79_23
timestamp 1606120353
transform 1 0 3220 0 1 45152
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__D
timestamp 1606120353
transform 1 0 3772 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1606120353
transform 1 0 3956 0 1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_79_44
timestamp 1606120353
transform 1 0 5152 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_40
timestamp 1606120353
transform 1 0 4784 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_36
timestamp 1606120353
transform 1 0 4416 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__CLK
timestamp 1606120353
transform 1 0 4232 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__D
timestamp 1606120353
transform 1 0 4600 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A
timestamp 1606120353
transform 1 0 4968 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1165_
timestamp 1606120353
transform 1 0 3772 0 -1 46240
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_2  FILLER_80_52
timestamp 1606120353
transform 1 0 5888 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_80_48
timestamp 1606120353
transform 1 0 5520 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__D
timestamp 1606120353
transform 1 0 6072 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__A
timestamp 1606120353
transform 1 0 5704 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__C
timestamp 1606120353
transform 1 0 5336 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_80_65
timestamp 1606120353
transform 1 0 7084 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_80_60
timestamp 1606120353
transform 1 0 6624 0 -1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_80_56
timestamp 1606120353
transform 1 0 6256 0 -1 46240
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_79_65
timestamp 1606120353
transform 1 0 7084 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1606120353
transform 1 0 6716 0 -1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0745_
timestamp 1606120353
transform 1 0 6808 0 -1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__nand4_4  _0850_
timestamp 1606120353
transform 1 0 5520 0 1 45152
box 0 -48 1564 592
use sky130_fd_sc_hd__decap_4  FILLER_80_69
timestamp 1606120353
transform 1 0 7452 0 -1 46240
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_79_69
timestamp 1606120353
transform 1 0 7452 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__A
timestamp 1606120353
transform 1 0 7268 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__A
timestamp 1606120353
transform 1 0 7268 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__B
timestamp 1606120353
transform 1 0 7636 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0768_
timestamp 1606120353
transform 1 0 7820 0 1 45152
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILLER_80_86
timestamp 1606120353
transform 1 0 9016 0 -1 46240
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_79_86
timestamp 1606120353
transform 1 0 9016 0 1 45152
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_79_82
timestamp 1606120353
transform 1 0 8648 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__A
timestamp 1606120353
transform 1 0 8832 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__nor3_4  _0560_
timestamp 1606120353
transform 1 0 7820 0 -1 46240
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_80_96
timestamp 1606120353
transform 1 0 9936 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_93
timestamp 1606120353
transform 1 0 9660 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0582__B
timestamp 1606120353
transform 1 0 9752 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0582__A
timestamp 1606120353
transform 1 0 9384 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1606120353
transform 1 0 9568 0 1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__nor2_4  _0582_
timestamp 1606120353
transform 1 0 9844 0 1 45152
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_79_104
timestamp 1606120353
transform 1 0 10672 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__D
timestamp 1606120353
transform 1 0 10120 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__B
timestamp 1606120353
transform 1 0 10856 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0713_
timestamp 1606120353
transform 1 0 10304 0 -1 46240
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILLER_80_109
timestamp 1606120353
transform 1 0 11132 0 -1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_79_108
timestamp 1606120353
transform 1 0 11040 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__C
timestamp 1606120353
transform 1 0 11224 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_80_118
timestamp 1606120353
transform 1 0 11960 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_80_114
timestamp 1606120353
transform 1 0 11592 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__B
timestamp 1606120353
transform 1 0 12144 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__B
timestamp 1606120353
transform 1 0 11776 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__C
timestamp 1606120353
transform 1 0 11408 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_80_132
timestamp 1606120353
transform 1 0 13248 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_130
timestamp 1606120353
transform 1 0 13064 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_126
timestamp 1606120353
transform 1 0 12696 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__B
timestamp 1606120353
transform 1 0 13248 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__A
timestamp 1606120353
transform 1 0 12880 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1606120353
transform 1 0 12328 0 -1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0660_
timestamp 1606120353
transform 1 0 12420 0 -1 46240
box 0 -48 828 592
use sky130_fd_sc_hd__nand3_4  _0659_
timestamp 1606120353
transform 1 0 11408 0 1 45152
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_6  FILLER_80_140
timestamp 1606120353
transform 1 0 13984 0 -1 46240
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_80_136
timestamp 1606120353
transform 1 0 13616 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_138
timestamp 1606120353
transform 1 0 13800 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_134
timestamp 1606120353
transform 1 0 13432 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__CLK
timestamp 1606120353
transform 1 0 13800 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__CLK
timestamp 1606120353
transform 1 0 13432 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__CLK
timestamp 1606120353
transform 1 0 13616 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A
timestamp 1606120353
transform 1 0 13984 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_149
timestamp 1606120353
transform 1 0 14812 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_145
timestamp 1606120353
transform 1 0 14444 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__A
timestamp 1606120353
transform 1 0 14628 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1073_
timestamp 1606120353
transform 1 0 14168 0 1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _1017_
timestamp 1606120353
transform 1 0 14536 0 -1 46240
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_79_154
timestamp 1606120353
transform 1 0 15272 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__B1
timestamp 1606120353
transform 1 0 14996 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1606120353
transform 1 0 15180 0 1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_80_159
timestamp 1606120353
transform 1 0 15732 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_80_155
timestamp 1606120353
transform 1 0 15364 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_163
timestamp 1606120353
transform 1 0 16100 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_159
timestamp 1606120353
transform 1 0 15732 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__A1
timestamp 1606120353
transform 1 0 15548 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__A2
timestamp 1606120353
transform 1 0 15916 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__D
timestamp 1606120353
transform 1 0 16284 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__A
timestamp 1606120353
transform 1 0 15916 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1018_
timestamp 1606120353
transform 1 0 15456 0 1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_80_175
timestamp 1606120353
transform 1 0 17204 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_79_167
timestamp 1606120353
transform 1 0 16468 0 1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__o21a_4  _1114_
timestamp 1606120353
transform 1 0 16744 0 1 45152
box 0 -48 1104 592
use sky130_fd_sc_hd__o21a_4  _1111_
timestamp 1606120353
transform 1 0 16100 0 -1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1606120353
transform -1 0 18860 0 1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1606120353
transform -1 0 18860 0 -1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1606120353
transform 1 0 17940 0 -1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A1
timestamp 1606120353
transform 1 0 17388 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__B1
timestamp 1606120353
transform 1 0 18032 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_182
timestamp 1606120353
transform 1 0 17848 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_79_186
timestamp 1606120353
transform 1 0 18216 0 1 45152
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_80_179
timestamp 1606120353
transform 1 0 17572 0 -1 46240
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_80_184
timestamp 1606120353
transform 1 0 18032 0 -1 46240
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1279_
timestamp 1606120353
transform 1 0 1472 0 1 46240
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1606120353
transform 1 0 1104 0 1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_81_3
timestamp 1606120353
transform 1 0 1380 0 1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_81_23
timestamp 1606120353
transform 1 0 3220 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__B
timestamp 1606120353
transform 1 0 3404 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_27
timestamp 1606120353
transform 1 0 3588 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__A
timestamp 1606120353
transform 1 0 3772 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_32
timestamp 1606120353
transform 1 0 4048 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1606120353
transform 1 0 3956 0 1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__A1
timestamp 1606120353
transform 1 0 4232 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_36
timestamp 1606120353
transform 1 0 4416 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__A2
timestamp 1606120353
transform 1 0 4600 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_40
timestamp 1606120353
transform 1 0 4784 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__B
timestamp 1606120353
transform 1 0 4968 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_44
timestamp 1606120353
transform 1 0 5152 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _0841_
timestamp 1606120353
transform 1 0 5520 0 1 46240
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__C
timestamp 1606120353
transform 1 0 5336 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_81_65
timestamp 1606120353
transform 1 0 7084 0 1 46240
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__B
timestamp 1606120353
transform 1 0 8004 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A
timestamp 1606120353
transform 1 0 8372 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__C
timestamp 1606120353
transform 1 0 8740 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__D
timestamp 1606120353
transform 1 0 7636 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_73
timestamp 1606120353
transform 1 0 7820 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_77
timestamp 1606120353
transform 1 0 8188 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_81
timestamp 1606120353
transform 1 0 8556 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_81_85
timestamp 1606120353
transform 1 0 8924 0 1 46240
box 0 -48 552 592
use sky130_fd_sc_hd__buf_1  _0733_
timestamp 1606120353
transform 1 0 9660 0 1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1606120353
transform 1 0 9568 0 1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A
timestamp 1606120353
transform 1 0 10120 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A
timestamp 1606120353
transform 1 0 10488 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_81_91
timestamp 1606120353
transform 1 0 9476 0 1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_81_96
timestamp 1606120353
transform 1 0 9936 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_100
timestamp 1606120353
transform 1 0 10304 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_81_104
timestamp 1606120353
transform 1 0 10672 0 1 46240
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _0583_
timestamp 1606120353
transform 1 0 11408 0 1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1182_
timestamp 1606120353
transform 1 0 12696 0 1 46240
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__D
timestamp 1606120353
transform 1 0 12512 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__A
timestamp 1606120353
transform 1 0 11868 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_115
timestamp 1606120353
transform 1 0 11684 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_81_119
timestamp 1606120353
transform 1 0 12052 0 1 46240
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_81_123
timestamp 1606120353
transform 1 0 12420 0 1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1606120353
transform 1 0 15180 0 1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_81_145
timestamp 1606120353
transform 1 0 14444 0 1 46240
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_81_154
timestamp 1606120353
transform 1 0 15272 0 1 46240
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _1057_
timestamp 1606120353
transform 1 0 16008 0 1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _1106_
timestamp 1606120353
transform 1 0 17020 0 1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A
timestamp 1606120353
transform 1 0 16468 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A
timestamp 1606120353
transform 1 0 16836 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_165
timestamp 1606120353
transform 1 0 16284 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_169
timestamp 1606120353
transform 1 0 16652 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_176
timestamp 1606120353
transform 1 0 17296 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1606120353
transform -1 0 18860 0 1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A
timestamp 1606120353
transform 1 0 17480 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_81_180
timestamp 1606120353
transform 1 0 17664 0 1 46240
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_81_188
timestamp 1606120353
transform 1 0 18400 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1606120353
transform 1 0 1104 0 -1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__D
timestamp 1606120353
transform 1 0 1564 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__CLK
timestamp 1606120353
transform 1 0 1932 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_82_3
timestamp 1606120353
transform 1 0 1380 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_82_7
timestamp 1606120353
transform 1 0 1748 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_82_11
timestamp 1606120353
transform 1 0 2116 0 -1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__o21ai_4  _0842_
timestamp 1606120353
transform 1 0 4784 0 -1 47328
box 0 -48 1196 592
use sky130_fd_sc_hd__nor2_4  _0875_
timestamp 1606120353
transform 1 0 3220 0 -1 47328
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__B1
timestamp 1606120353
transform 1 0 4600 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_82_32
timestamp 1606120353
transform 1 0 4048 0 -1 47328
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1606120353
transform 1 0 6716 0 -1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__D
timestamp 1606120353
transform 1 0 6164 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_82_53
timestamp 1606120353
transform 1 0 5980 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_82_57
timestamp 1606120353
transform 1 0 6348 0 -1 47328
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_82_62
timestamp 1606120353
transform 1 0 6808 0 -1 47328
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_82_66
timestamp 1606120353
transform 1 0 7176 0 -1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__nand4_4  _0783_
timestamp 1606120353
transform 1 0 8004 0 -1 47328
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A1
timestamp 1606120353
transform 1 0 7268 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_82_69
timestamp 1606120353
transform 1 0 7452 0 -1 47328
box 0 -48 552 592
use sky130_fd_sc_hd__inv_8  _0779_
timestamp 1606120353
transform 1 0 10304 0 -1 47328
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__C
timestamp 1606120353
transform 1 0 10120 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__D
timestamp 1606120353
transform 1 0 9752 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_82_92
timestamp 1606120353
transform 1 0 9568 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_82_96
timestamp 1606120353
transform 1 0 9936 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_82_109
timestamp 1606120353
transform 1 0 11132 0 -1 47328
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1181_
timestamp 1606120353
transform 1 0 12972 0 -1 47328
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1606120353
transform 1 0 12328 0 -1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__D
timestamp 1606120353
transform 1 0 12696 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__A
timestamp 1606120353
transform 1 0 11592 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__CLK
timestamp 1606120353
transform 1 0 12144 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_82_113
timestamp 1606120353
transform 1 0 11500 0 -1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_82_116
timestamp 1606120353
transform 1 0 11776 0 -1 47328
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_82_123
timestamp 1606120353
transform 1 0 12420 0 -1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_82_128
timestamp 1606120353
transform 1 0 12880 0 -1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_82_148
timestamp 1606120353
transform 1 0 14720 0 -1 47328
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _1121_
timestamp 1606120353
transform 1 0 16928 0 -1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A
timestamp 1606120353
transform 1 0 15640 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__C
timestamp 1606120353
transform 1 0 16008 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__C
timestamp 1606120353
transform 1 0 16376 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_82_156
timestamp 1606120353
transform 1 0 15456 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_82_160
timestamp 1606120353
transform 1 0 15824 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_82_164
timestamp 1606120353
transform 1 0 16192 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_82_168
timestamp 1606120353
transform 1 0 16560 0 -1 47328
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_82_175
timestamp 1606120353
transform 1 0 17204 0 -1 47328
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1606120353
transform -1 0 18860 0 -1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1606120353
transform 1 0 17940 0 -1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_82_184
timestamp 1606120353
transform 1 0 18032 0 -1 47328
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1280_
timestamp 1606120353
transform 1 0 1472 0 1 47328
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1606120353
transform 1 0 1104 0 1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_83_3
timestamp 1606120353
transform 1 0 1380 0 1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1606120353
transform 1 0 3956 0 1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__B
timestamp 1606120353
transform 1 0 4968 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__A
timestamp 1606120353
transform 1 0 4600 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__A
timestamp 1606120353
transform 1 0 4232 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_83_23
timestamp 1606120353
transform 1 0 3220 0 1 47328
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_83_32
timestamp 1606120353
transform 1 0 4048 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_36
timestamp 1606120353
transform 1 0 4416 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_40
timestamp 1606120353
transform 1 0 4784 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_44
timestamp 1606120353
transform 1 0 5152 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _0859_
timestamp 1606120353
transform 1 0 5520 0 1 47328
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__C
timestamp 1606120353
transform 1 0 5336 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_65
timestamp 1606120353
transform 1 0 7084 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0784_
timestamp 1606120353
transform 1 0 8004 0 1 47328
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__A
timestamp 1606120353
transform 1 0 9016 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A2
timestamp 1606120353
transform 1 0 7268 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__B1
timestamp 1606120353
transform 1 0 7636 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_69
timestamp 1606120353
transform 1 0 7452 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_73
timestamp 1606120353
transform 1 0 7820 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_84
timestamp 1606120353
transform 1 0 8832 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_88
timestamp 1606120353
transform 1 0 9200 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0532_
timestamp 1606120353
transform 1 0 9660 0 1 47328
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1606120353
transform 1 0 9568 0 1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0532__A
timestamp 1606120353
transform 1 0 9384 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__B
timestamp 1606120353
transform 1 0 10672 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__A
timestamp 1606120353
transform 1 0 11040 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_102
timestamp 1606120353
transform 1 0 10488 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_106
timestamp 1606120353
transform 1 0 10856 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_110
timestamp 1606120353
transform 1 0 11224 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__nand3_4  _0657_
timestamp 1606120353
transform 1 0 11592 0 1 47328
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__D
timestamp 1606120353
transform 1 0 13064 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__B
timestamp 1606120353
transform 1 0 11408 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_128
timestamp 1606120353
transform 1 0 12880 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_132
timestamp 1606120353
transform 1 0 13248 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1606120353
transform 1 0 15180 0 1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__B
timestamp 1606120353
transform 1 0 14996 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__CLK
timestamp 1606120353
transform 1 0 13432 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__CLK
timestamp 1606120353
transform 1 0 13800 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_136
timestamp 1606120353
transform 1 0 13616 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_83_140
timestamp 1606120353
transform 1 0 13984 0 1 47328
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_83_148
timestamp 1606120353
transform 1 0 14720 0 1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_83_154
timestamp 1606120353
transform 1 0 15272 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _1110_
timestamp 1606120353
transform 1 0 15640 0 1 47328
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A
timestamp 1606120353
transform 1 0 15456 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__B
timestamp 1606120353
transform 1 0 16652 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_167
timestamp 1606120353
transform 1 0 16468 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_83_171
timestamp 1606120353
transform 1 0 16836 0 1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1606120353
transform -1 0 18860 0 1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_83_183
timestamp 1606120353
transform 1 0 17940 0 1 47328
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_83_189
timestamp 1606120353
transform 1 0 18492 0 1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1606120353
transform 1 0 1104 0 -1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1282__D
timestamp 1606120353
transform 1 0 1564 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_3
timestamp 1606120353
transform 1 0 1380 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_84_7
timestamp 1606120353
transform 1 0 1748 0 -1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_84_19
timestamp 1606120353
transform 1 0 2852 0 -1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__inv_8  _0559_
timestamp 1606120353
transform 1 0 5152 0 -1 48416
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__B
timestamp 1606120353
transform 1 0 4784 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_84_31
timestamp 1606120353
transform 1 0 3956 0 -1 48416
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_84_39
timestamp 1606120353
transform 1 0 4692 0 -1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_84_42
timestamp 1606120353
transform 1 0 4968 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1606120353
transform 1 0 6716 0 -1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__B1
timestamp 1606120353
transform 1 0 6992 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__C1
timestamp 1606120353
transform 1 0 6532 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__A1
timestamp 1606120353
transform 1 0 6164 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_53
timestamp 1606120353
transform 1 0 5980 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_57
timestamp 1606120353
transform 1 0 6348 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_62
timestamp 1606120353
transform 1 0 6808 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_84_66
timestamp 1606120353
transform 1 0 7176 0 -1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0521_
timestamp 1606120353
transform 1 0 9200 0 -1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__a21oi_4  _0789_
timestamp 1606120353
transform 1 0 7268 0 -1 48416
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__C
timestamp 1606120353
transform 1 0 9016 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A
timestamp 1606120353
transform 1 0 8648 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_80
timestamp 1606120353
transform 1 0 8464 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_84
timestamp 1606120353
transform 1 0 8832 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _0711_
timestamp 1606120353
transform 1 0 10304 0 -1 48416
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0532__B
timestamp 1606120353
transform 1 0 9660 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__B
timestamp 1606120353
transform 1 0 10120 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_91
timestamp 1606120353
transform 1 0 9476 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_84_95
timestamp 1606120353
transform 1 0 9844 0 -1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_84_109
timestamp 1606120353
transform 1 0 11132 0 -1 48416
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_84_120
timestamp 1606120353
transform 1 0 12144 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_116
timestamp 1606120353
transform 1 0 11776 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_84_113
timestamp 1606120353
transform 1 0 11500 0 -1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__D
timestamp 1606120353
transform 1 0 11960 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__C
timestamp 1606120353
transform 1 0 11592 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_127
timestamp 1606120353
transform 1 0 12788 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_123
timestamp 1606120353
transform 1 0 12420 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__C
timestamp 1606120353
transform 1 0 12604 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1606120353
transform 1 0 12328 0 -1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1183_
timestamp 1606120353
transform 1 0 12972 0 -1 48416
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_8  FILLER_84_148
timestamp 1606120353
transform 1 0 14720 0 -1 48416
box 0 -48 736 592
use sky130_fd_sc_hd__and3_4  _1137_
timestamp 1606120353
transform 1 0 15640 0 -1 48416
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__A1
timestamp 1606120353
transform 1 0 16652 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A1
timestamp 1606120353
transform 1 0 17020 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_156
timestamp 1606120353
transform 1 0 15456 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_167
timestamp 1606120353
transform 1 0 16468 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_171
timestamp 1606120353
transform 1 0 16836 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_175
timestamp 1606120353
transform 1 0 17204 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1606120353
transform -1 0 18860 0 -1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1606120353
transform 1 0 17940 0 -1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__B1
timestamp 1606120353
transform 1 0 17388 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_84_179
timestamp 1606120353
transform 1 0 17572 0 -1 48416
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_84_184
timestamp 1606120353
transform 1 0 18032 0 -1 48416
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILLER_86_7
timestamp 1606120353
transform 1 0 1748 0 -1 49504
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1606120353
transform 1 0 1380 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_85_3
timestamp 1606120353
transform 1 0 1380 0 1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1282__CLK
timestamp 1606120353
transform 1 0 1564 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1606120353
transform 1 0 1104 0 -1 49504
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1606120353
transform 1 0 1104 0 1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_86_16
timestamp 1606120353
transform 1 0 2576 0 -1 49504
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_86_13
timestamp 1606120353
transform 1 0 2300 0 -1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A1
timestamp 1606120353
transform 1 0 2944 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__B
timestamp 1606120353
transform 1 0 2392 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1282_
timestamp 1606120353
transform 1 0 1472 0 1 48416
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1147_
timestamp 1606120353
transform 1 0 3128 0 -1 49504
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_2  FILLER_85_27
timestamp 1606120353
transform 1 0 3588 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_23
timestamp 1606120353
transform 1 0 3220 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__CLK
timestamp 1606120353
transform 1 0 3772 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__D
timestamp 1606120353
transform 1 0 3404 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1606120353
transform 1 0 3956 0 1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_85_32
timestamp 1606120353
transform 1 0 4048 0 1 48416
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A
timestamp 1606120353
transform 1 0 4600 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__nand2_4  _0864_
timestamp 1606120353
transform 1 0 4784 0 1 48416
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_86_41
timestamp 1606120353
transform 1 0 4876 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__B2
timestamp 1606120353
transform 1 0 5060 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_86_45
timestamp 1606120353
transform 1 0 5244 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_clk_A
timestamp 1606120353
transform 1 0 5428 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_49
timestamp 1606120353
transform 1 0 5612 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_86_49
timestamp 1606120353
transform 1 0 5612 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__B1
timestamp 1606120353
transform 1 0 5796 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__A1
timestamp 1606120353
transform 1 0 5796 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_53
timestamp 1606120353
transform 1 0 5980 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_86_53
timestamp 1606120353
transform 1 0 5980 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__A2
timestamp 1606120353
transform 1 0 6164 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A4
timestamp 1606120353
transform 1 0 6164 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_86_57
timestamp 1606120353
transform 1 0 6348 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_57
timestamp 1606120353
transform 1 0 6348 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A3
timestamp 1606120353
transform 1 0 6532 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__A2
timestamp 1606120353
transform 1 0 6532 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1606120353
transform 1 0 6716 0 -1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__a211o_4  _0791_
timestamp 1606120353
transform 1 0 6808 0 -1 49504
box 0 -48 1288 592
use sky130_fd_sc_hd__a211o_4  _0771_
timestamp 1606120353
transform 1 0 6716 0 1 48416
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_86_76
timestamp 1606120353
transform 1 0 8096 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_75
timestamp 1606120353
transform 1 0 8004 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__C1
timestamp 1606120353
transform 1 0 8188 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__D
timestamp 1606120353
transform 1 0 8280 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_86_80
timestamp 1606120353
transform 1 0 8464 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_85_79
timestamp 1606120353
transform 1 0 8372 0 1 48416
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__C
timestamp 1606120353
transform 1 0 8648 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_85_86
timestamp 1606120353
transform 1 0 9016 0 1 48416
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_85_83
timestamp 1606120353
transform 1 0 8740 0 1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0533__A
timestamp 1606120353
transform 1 0 8832 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0533_
timestamp 1606120353
transform 1 0 8832 0 -1 49504
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_86_87
timestamp 1606120353
transform 1 0 9108 0 -1 49504
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_86_96
timestamp 1606120353
transform 1 0 9936 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_86_92
timestamp 1606120353
transform 1 0 9568 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_85_93
timestamp 1606120353
transform 1 0 9660 0 1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__C
timestamp 1606120353
transform 1 0 9384 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__B
timestamp 1606120353
transform 1 0 9752 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__A
timestamp 1606120353
transform 1 0 9384 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1606120353
transform 1 0 9568 0 1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0716_
timestamp 1606120353
transform 1 0 10120 0 -1 49504
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_86_107
timestamp 1606120353
transform 1 0 10948 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__B
timestamp 1606120353
transform 1 0 11132 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _0595_
timestamp 1606120353
transform 1 0 9752 0 1 48416
box 0 -48 1564 592
use sky130_fd_sc_hd__decap_3  FILLER_86_115
timestamp 1606120353
transform 1 0 11684 0 -1 49504
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_86_111
timestamp 1606120353
transform 1 0 11316 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_115
timestamp 1606120353
transform 1 0 11684 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_111
timestamp 1606120353
transform 1 0 11316 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__A2
timestamp 1606120353
transform 1 0 11500 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__A
timestamp 1606120353
transform 1 0 11960 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__D
timestamp 1606120353
transform 1 0 11868 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A
timestamp 1606120353
transform 1 0 11500 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0611_
timestamp 1606120353
transform 1 0 12052 0 1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_86_120
timestamp 1606120353
transform 1 0 12144 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_126
timestamp 1606120353
transform 1 0 12696 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_122
timestamp 1606120353
transform 1 0 12328 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__A
timestamp 1606120353
transform 1 0 12880 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A
timestamp 1606120353
transform 1 0 12512 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1606120353
transform 1 0 12328 0 -1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__and3_4  _0714_
timestamp 1606120353
transform 1 0 12420 0 -1 49504
box 0 -48 828 592
use sky130_fd_sc_hd__decap_4  FILLER_86_132
timestamp 1606120353
transform 1 0 13248 0 -1 49504
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_85_130
timestamp 1606120353
transform 1 0 13064 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__B
timestamp 1606120353
transform 1 0 13248 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_86_138
timestamp 1606120353
transform 1 0 13800 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_140
timestamp 1606120353
transform 1 0 13984 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_85_134
timestamp 1606120353
transform 1 0 13432 0 1 48416
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__C
timestamp 1606120353
transform 1 0 13800 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__C
timestamp 1606120353
transform 1 0 13984 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__B
timestamp 1606120353
transform 1 0 13616 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_86_142
timestamp 1606120353
transform 1 0 14168 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_85_148
timestamp 1606120353
transform 1 0 14720 0 1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_85_144
timestamp 1606120353
transform 1 0 14352 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_clk_A
timestamp 1606120353
transform 1 0 14352 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__B
timestamp 1606120353
transform 1 0 14168 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__A
timestamp 1606120353
transform 1 0 14536 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _1128_
timestamp 1606120353
transform 1 0 14536 0 -1 49504
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__B1
timestamp 1606120353
transform 1 0 14996 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1606120353
transform 1 0 15180 0 1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _1101_
timestamp 1606120353
transform 1 0 15272 0 1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_86_159
timestamp 1606120353
transform 1 0 15732 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_86_155
timestamp 1606120353
transform 1 0 15364 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_85_165
timestamp 1606120353
transform 1 0 16284 0 1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_85_161
timestamp 1606120353
transform 1 0 15916 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_157
timestamp 1606120353
transform 1 0 15548 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__D
timestamp 1606120353
transform 1 0 15916 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__A2
timestamp 1606120353
transform 1 0 16100 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__A
timestamp 1606120353
transform 1 0 15732 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__C
timestamp 1606120353
transform 1 0 15548 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_86_175
timestamp 1606120353
transform 1 0 17204 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A2
timestamp 1606120353
transform 1 0 16560 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _1123_
timestamp 1606120353
transform 1 0 16100 0 -1 49504
box 0 -48 1104 592
use sky130_fd_sc_hd__o21a_4  _1119_
timestamp 1606120353
transform 1 0 16744 0 1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1606120353
transform -1 0 18860 0 1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1606120353
transform -1 0 18860 0 -1 49504
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1606120353
transform 1 0 17940 0 -1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__B1
timestamp 1606120353
transform 1 0 17388 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_85_182
timestamp 1606120353
transform 1 0 17848 0 1 48416
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_86_179
timestamp 1606120353
transform 1 0 17572 0 -1 49504
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_86_184
timestamp 1606120353
transform 1 0 18032 0 -1 49504
box 0 -48 552 592
use sky130_fd_sc_hd__nand2_4  _0776_
timestamp 1606120353
transform 1 0 2392 0 1 49504
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1606120353
transform 1 0 1104 0 1 49504
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__A
timestamp 1606120353
transform 1 0 2208 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_87_3
timestamp 1606120353
transform 1 0 1380 0 1 49504
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_87_11
timestamp 1606120353
transform 1 0 2116 0 1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_87_32
timestamp 1606120353
transform 1 0 4048 0 1 49504
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_87_27
timestamp 1606120353
transform 1 0 3588 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_23
timestamp 1606120353
transform 1 0 3220 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__B1_N
timestamp 1606120353
transform 1 0 3772 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A2
timestamp 1606120353
transform 1 0 3404 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1606120353
transform 1 0 3956 0 1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_87_38
timestamp 1606120353
transform 1 0 4600 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__B1
timestamp 1606120353
transform 1 0 4416 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A2_N
timestamp 1606120353
transform 1 0 4784 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__a2bb2o_4  _0772_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 4968 0 1 49504
box 0 -48 1472 592
use sky130_fd_sc_hd__o41a_4  _0790_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 7176 0 1 49504
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A2
timestamp 1606120353
transform 1 0 6992 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A1
timestamp 1606120353
transform 1 0 6624 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_58
timestamp 1606120353
transform 1 0 6440 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_62
timestamp 1606120353
transform 1 0 6808 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__A1
timestamp 1606120353
transform 1 0 8924 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_83
timestamp 1606120353
transform 1 0 8740 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_87
timestamp 1606120353
transform 1 0 9108 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _0723_
timestamp 1606120353
transform 1 0 9660 0 1 49504
box 0 -48 1564 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1606120353
transform 1 0 9568 0 1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__B1
timestamp 1606120353
transform 1 0 9292 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_87_91
timestamp 1606120353
transform 1 0 9476 0 1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_87_110
timestamp 1606120353
transform 1 0 11224 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _0717_
timestamp 1606120353
transform 1 0 11960 0 1 49504
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__D
timestamp 1606120353
transform 1 0 13064 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__A
timestamp 1606120353
transform 1 0 11408 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__B
timestamp 1606120353
transform 1 0 11776 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_114
timestamp 1606120353
transform 1 0 11592 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_87_127
timestamp 1606120353
transform 1 0 12788 0 1 49504
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_87_132
timestamp 1606120353
transform 1 0 13248 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1076_
timestamp 1606120353
transform 1 0 15272 0 1 49504
box 0 -48 276 592
use sky130_fd_sc_hd__and3_4  _1118_
timestamp 1606120353
transform 1 0 13616 0 1 49504
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1606120353
transform 1 0 15180 0 1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__B
timestamp 1606120353
transform 1 0 14996 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__A
timestamp 1606120353
transform 1 0 13432 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__C
timestamp 1606120353
transform 1 0 14628 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_145
timestamp 1606120353
transform 1 0 14444 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_149
timestamp 1606120353
transform 1 0 14812 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1135_
timestamp 1606120353
transform 1 0 16652 0 1 49504
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__A
timestamp 1606120353
transform 1 0 15732 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A
timestamp 1606120353
transform 1 0 16100 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__A1
timestamp 1606120353
transform 1 0 16468 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_157
timestamp 1606120353
transform 1 0 15548 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_161
timestamp 1606120353
transform 1 0 15916 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_165
timestamp 1606120353
transform 1 0 16284 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1606120353
transform -1 0 18860 0 1 49504
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_87_182
timestamp 1606120353
transform 1 0 17848 0 1 49504
box 0 -48 736 592
use sky130_fd_sc_hd__a21bo_4  _0777_
timestamp 1606120353
transform 1 0 3128 0 -1 50592
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1606120353
transform 1 0 1104 0 -1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__D
timestamp 1606120353
transform 1 0 1564 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_3
timestamp 1606120353
transform 1 0 1380 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_88_7
timestamp 1606120353
transform 1 0 1748 0 -1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_88_19
timestamp 1606120353
transform 1 0 2852 0 -1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A1_N
timestamp 1606120353
transform 1 0 4968 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__D
timestamp 1606120353
transform 1 0 4600 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_88_35
timestamp 1606120353
transform 1 0 4324 0 -1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_88_40
timestamp 1606120353
transform 1 0 4784 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_88_44
timestamp 1606120353
transform 1 0 5152 0 -1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__A3
timestamp 1606120353
transform 1 0 5428 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_49
timestamp 1606120353
transform 1 0 5612 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__B2
timestamp 1606120353
transform 1 0 5796 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_53
timestamp 1606120353
transform 1 0 5980 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B1
timestamp 1606120353
transform 1 0 6164 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_57
timestamp 1606120353
transform 1 0 6348 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__A4
timestamp 1606120353
transform 1 0 6532 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_62
timestamp 1606120353
transform 1 0 6808 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1606120353
transform 1 0 6716 0 -1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__C
timestamp 1606120353
transform 1 0 6992 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_66
timestamp 1606120353
transform 1 0 7176 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__a2111o_4  _0739_
timestamp 1606120353
transform 1 0 8648 0 -1 50592
box 0 -48 1564 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk
timestamp 1606120353
transform 1 0 8372 0 -1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__C1
timestamp 1606120353
transform 1 0 8188 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__D1
timestamp 1606120353
transform 1 0 7820 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__A2
timestamp 1606120353
transform 1 0 7360 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_88_70
timestamp 1606120353
transform 1 0 7544 0 -1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_88_75
timestamp 1606120353
transform 1 0 8004 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__B
timestamp 1606120353
transform 1 0 10764 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__A
timestamp 1606120353
transform 1 0 11132 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__A
timestamp 1606120353
transform 1 0 10396 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_99
timestamp 1606120353
transform 1 0 10212 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_103
timestamp 1606120353
transform 1 0 10580 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_107
timestamp 1606120353
transform 1 0 10948 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_118
timestamp 1606120353
transform 1 0 11960 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_114
timestamp 1606120353
transform 1 0 11592 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__B1
timestamp 1606120353
transform 1 0 12144 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__C
timestamp 1606120353
transform 1 0 11776 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0593_
timestamp 1606120353
transform 1 0 11316 0 -1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_88_127
timestamp 1606120353
transform 1 0 12788 0 -1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_88_123
timestamp 1606120353
transform 1 0 12420 0 -1 50592
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__A1
timestamp 1606120353
transform 1 0 12880 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1606120353
transform 1 0 12328 0 -1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1187_
timestamp 1606120353
transform 1 0 13064 0 -1 50592
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__D
timestamp 1606120353
transform 1 0 14996 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_149
timestamp 1606120353
transform 1 0 14812 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_153
timestamp 1606120353
transform 1 0 15180 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _1108_
timestamp 1606120353
transform 1 0 15548 0 -1 50592
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__C
timestamp 1606120353
transform 1 0 15364 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__A2
timestamp 1606120353
transform 1 0 17296 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_174
timestamp 1606120353
transform 1 0 17112 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1606120353
transform -1 0 18860 0 -1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1606120353
transform 1 0 17940 0 -1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_88_178
timestamp 1606120353
transform 1 0 17480 0 -1 50592
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_88_182
timestamp 1606120353
transform 1 0 17848 0 -1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_88_184
timestamp 1606120353
transform 1 0 18032 0 -1 50592
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1281_
timestamp 1606120353
transform 1 0 1472 0 1 50592
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1606120353
transform 1 0 1104 0 1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_89_3
timestamp 1606120353
transform 1 0 1380 0 1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_89_23
timestamp 1606120353
transform 1 0 3220 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_clk_A
timestamp 1606120353
transform 1 0 3404 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_27
timestamp 1606120353
transform 1 0 3588 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A1
timestamp 1606120353
transform 1 0 3772 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1606120353
transform 1 0 3956 0 1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0704_
timestamp 1606120353
transform 1 0 4048 0 1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_89_35
timestamp 1606120353
transform 1 0 4324 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__A
timestamp 1606120353
transform 1 0 4508 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_39
timestamp 1606120353
transform 1 0 4692 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_89_43
timestamp 1606120353
transform 1 0 5060 0 1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A2
timestamp 1606120353
transform 1 0 4876 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_clk
timestamp 1606120353
transform 1 0 5152 0 1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1606120353
transform 1 0 6164 0 1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1606120353
transform 1 0 5796 0 1 50592
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_89_47
timestamp 1606120353
transform 1 0 5428 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__B1
timestamp 1606120353
transform 1 0 5612 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_62
timestamp 1606120353
transform 1 0 6808 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_58
timestamp 1606120353
transform 1 0 6440 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A
timestamp 1606120353
transform 1 0 6256 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__B
timestamp 1606120353
transform 1 0 6624 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__A1
timestamp 1606120353
transform 1 0 6992 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__o41a_4  _0770_
timestamp 1606120353
transform 1 0 7176 0 1 50592
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__B1
timestamp 1606120353
transform 1 0 8924 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_83
timestamp 1606120353
transform 1 0 8740 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_87
timestamp 1606120353
transform 1 0 9108 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__nor4_4  _0719_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 10212 0 1 50592
box 0 -48 1564 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1606120353
transform 1 0 9568 0 1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__C
timestamp 1606120353
transform 1 0 10028 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__A2
timestamp 1606120353
transform 1 0 9292 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_89_91
timestamp 1606120353
transform 1 0 9476 0 1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_89_93
timestamp 1606120353
transform 1 0 9660 0 1 50592
box 0 -48 368 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_clk
timestamp 1606120353
transform 1 0 12512 0 1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__D
timestamp 1606120353
transform 1 0 12972 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__B
timestamp 1606120353
transform 1 0 11960 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__B1
timestamp 1606120353
transform 1 0 12328 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_116
timestamp 1606120353
transform 1 0 11776 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_120
timestamp 1606120353
transform 1 0 12144 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_127
timestamp 1606120353
transform 1 0 12788 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_131
timestamp 1606120353
transform 1 0 13156 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1058_
timestamp 1606120353
transform 1 0 15272 0 1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__o21a_4  _1129_
timestamp 1606120353
transform 1 0 13340 0 1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1606120353
transform 1 0 15180 0 1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__B
timestamp 1606120353
transform 1 0 14996 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__A2
timestamp 1606120353
transform 1 0 14628 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_145
timestamp 1606120353
transform 1 0 14444 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_149
timestamp 1606120353
transform 1 0 14812 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1134_
timestamp 1606120353
transform 1 0 16652 0 1 50592
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__A
timestamp 1606120353
transform 1 0 15732 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A
timestamp 1606120353
transform 1 0 16100 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A1
timestamp 1606120353
transform 1 0 16468 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_157
timestamp 1606120353
transform 1 0 15548 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_161
timestamp 1606120353
transform 1 0 15916 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_165
timestamp 1606120353
transform 1 0 16284 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1606120353
transform -1 0 18860 0 1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__CLK
timestamp 1606120353
transform 1 0 18032 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_182
timestamp 1606120353
transform 1 0 17848 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_89_186
timestamp 1606120353
transform 1 0 18216 0 1 50592
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1606120353
transform 1 0 1104 0 -1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__CLK
timestamp 1606120353
transform 1 0 3128 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__CLK
timestamp 1606120353
transform 1 0 1564 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_3
timestamp 1606120353
transform 1 0 1380 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_90_7
timestamp 1606120353
transform 1 0 1748 0 -1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_90_19
timestamp 1606120353
transform 1 0 2852 0 -1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _0855_
timestamp 1606120353
transform 1 0 4692 0 -1 51680
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A2
timestamp 1606120353
transform 1 0 4048 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__B1
timestamp 1606120353
transform 1 0 4508 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_90_24
timestamp 1606120353
transform 1 0 3312 0 -1 51680
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_90_34
timestamp 1606120353
transform 1 0 4232 0 -1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__and4_4  _0712_
timestamp 1606120353
transform 1 0 6900 0 -1 51680
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1606120353
transform 1 0 6716 0 -1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__B1
timestamp 1606120353
transform 1 0 6532 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__B1
timestamp 1606120353
transform 1 0 6072 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_52
timestamp 1606120353
transform 1 0 5888 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_90_56
timestamp 1606120353
transform 1 0 6256 0 -1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_90_62
timestamp 1606120353
transform 1 0 6808 0 -1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__a32o_4  _0785_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 8464 0 -1 51680
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__A1
timestamp 1606120353
transform 1 0 8280 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__A3
timestamp 1606120353
transform 1 0 7912 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_72
timestamp 1606120353
transform 1 0 7728 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_76
timestamp 1606120353
transform 1 0 8096 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0718_
timestamp 1606120353
transform 1 0 10764 0 -1 51680
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A1
timestamp 1606120353
transform 1 0 10580 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__A
timestamp 1606120353
transform 1 0 10212 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_97
timestamp 1606120353
transform 1 0 10028 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_101
timestamp 1606120353
transform 1 0 10396 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1180_
timestamp 1606120353
transform 1 0 12880 0 -1 51680
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1606120353
transform 1 0 12328 0 -1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__D
timestamp 1606120353
transform 1 0 11776 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__B1
timestamp 1606120353
transform 1 0 12696 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A2
timestamp 1606120353
transform 1 0 12144 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_114
timestamp 1606120353
transform 1 0 11592 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_118
timestamp 1606120353
transform 1 0 11960 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_90_123
timestamp 1606120353
transform 1 0 12420 0 -1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__C
timestamp 1606120353
transform 1 0 14812 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__D
timestamp 1606120353
transform 1 0 15180 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_147
timestamp 1606120353
transform 1 0 14628 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_151
timestamp 1606120353
transform 1 0 14996 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _1117_
timestamp 1606120353
transform 1 0 15364 0 -1 51680
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A2
timestamp 1606120353
transform 1 0 17112 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_172
timestamp 1606120353
transform 1 0 16928 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_176
timestamp 1606120353
transform 1 0 17296 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1606120353
transform -1 0 18860 0 -1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1606120353
transform 1 0 17940 0 -1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__B1
timestamp 1606120353
transform 1 0 17480 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_90_180
timestamp 1606120353
transform 1 0 17664 0 -1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_90_184
timestamp 1606120353
transform 1 0 18032 0 -1 51680
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1606120353
transform 1 0 1104 0 1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__C
timestamp 1606120353
transform 1 0 3036 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__D
timestamp 1606120353
transform 1 0 2668 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_91_3
timestamp 1606120353
transform 1 0 1380 0 1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_91_15
timestamp 1606120353
transform 1 0 2484 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_19
timestamp 1606120353
transform 1 0 2852 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0867_
timestamp 1606120353
transform 1 0 4048 0 1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1606120353
transform 1 0 3956 0 1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A1
timestamp 1606120353
transform 1 0 3772 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__B1
timestamp 1606120353
transform 1 0 3404 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_23
timestamp 1606120353
transform 1 0 3220 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_27
timestamp 1606120353
transform 1 0 3588 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_44
timestamp 1606120353
transform 1 0 5152 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__a2bb2o_4  _0792_
timestamp 1606120353
transform 1 0 5888 0 1 51680
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__A2_N
timestamp 1606120353
transform 1 0 5704 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__A1_N
timestamp 1606120353
transform 1 0 5336 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_48
timestamp 1606120353
transform 1 0 5520 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_68
timestamp 1606120353
transform 1 0 7360 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_72
timestamp 1606120353
transform 1 0 7728 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A2_N
timestamp 1606120353
transform 1 0 7544 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__B2
timestamp 1606120353
transform 1 0 7912 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_76
timestamp 1606120353
transform 1 0 8096 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A1_N
timestamp 1606120353
transform 1 0 8280 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_91_80
timestamp 1606120353
transform 1 0 8464 0 1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0526_
timestamp 1606120353
transform 1 0 8556 0 1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_91_84
timestamp 1606120353
transform 1 0 8832 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0526__A
timestamp 1606120353
transform 1 0 9016 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_88
timestamp 1606120353
transform 1 0 9200 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__a2111oi_4  _0715_
timestamp 1606120353
transform 1 0 10580 0 1 51680
box 0 -48 2024 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1606120353
transform 1 0 9568 0 1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__B
timestamp 1606120353
transform 1 0 10304 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__A
timestamp 1606120353
transform 1 0 9936 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__C1
timestamp 1606120353
transform 1 0 9384 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_91_93
timestamp 1606120353
transform 1 0 9660 0 1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_91_98
timestamp 1606120353
transform 1 0 10120 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_91_102
timestamp 1606120353
transform 1 0 10488 0 1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__A1
timestamp 1606120353
transform 1 0 13156 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A1
timestamp 1606120353
transform 1 0 12788 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_125
timestamp 1606120353
transform 1 0 12604 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_129
timestamp 1606120353
transform 1 0 12972 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _1133_
timestamp 1606120353
transform 1 0 13340 0 1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1606120353
transform 1 0 15180 0 1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__B
timestamp 1606120353
transform 1 0 14628 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__A
timestamp 1606120353
transform 1 0 14996 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_145
timestamp 1606120353
transform 1 0 14444 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_149
timestamp 1606120353
transform 1 0 14812 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_154
timestamp 1606120353
transform 1 0 15272 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _1095_
timestamp 1606120353
transform 1 0 15456 0 1 51680
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__B
timestamp 1606120353
transform 1 0 17204 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_173
timestamp 1606120353
transform 1 0 17020 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1606120353
transform -1 0 18860 0 1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__A
timestamp 1606120353
transform 1 0 17572 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__C
timestamp 1606120353
transform 1 0 17940 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_177
timestamp 1606120353
transform 1 0 17388 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_181
timestamp 1606120353
transform 1 0 17756 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_91_185
timestamp 1606120353
transform 1 0 18124 0 1 51680
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_91_189
timestamp 1606120353
transform 1 0 18492 0 1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_93_3
timestamp 1606120353
transform 1 0 1380 0 1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_92_11
timestamp 1606120353
transform 1 0 2116 0 -1 52768
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_92_7
timestamp 1606120353
transform 1 0 1748 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_3
timestamp 1606120353
transform 1 0 1380 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__CLK
timestamp 1606120353
transform 1 0 1932 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__D
timestamp 1606120353
transform 1 0 1564 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1606120353
transform 1 0 1104 0 1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1606120353
transform 1 0 1104 0 -1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_92_21
timestamp 1606120353
transform 1 0 3036 0 -1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__B1
timestamp 1606120353
transform 1 0 2852 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1159_
timestamp 1606120353
transform 1 0 3128 0 -1 52768
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1148_
timestamp 1606120353
transform 1 0 1472 0 1 52768
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1162_
timestamp 1606120353
transform 1 0 4232 0 1 52768
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1606120353
transform 1 0 3956 0 1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__A1
timestamp 1606120353
transform 1 0 3404 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__B
timestamp 1606120353
transform 1 0 5060 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A
timestamp 1606120353
transform 1 0 3772 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_41
timestamp 1606120353
transform 1 0 4876 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_93_23
timestamp 1606120353
transform 1 0 3220 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_93_27
timestamp 1606120353
transform 1 0 3588 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_93_32
timestamp 1606120353
transform 1 0 4048 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_93_53
timestamp 1606120353
transform 1 0 5980 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_52
timestamp 1606120353
transform 1 0 5888 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_45
timestamp 1606120353
transform 1 0 5244 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__A
timestamp 1606120353
transform 1 0 5428 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__B2
timestamp 1606120353
transform 1 0 6072 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__B1
timestamp 1606120353
transform 1 0 6164 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0577_
timestamp 1606120353
transform 1 0 5612 0 -1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_93_57
timestamp 1606120353
transform 1 0 6348 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_92_56
timestamp 1606120353
transform 1 0 6256 0 -1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A1
timestamp 1606120353
transform 1 0 6532 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__A
timestamp 1606120353
transform 1 0 6532 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1606120353
transform 1 0 6716 0 -1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__a21oi_4  _0782_
timestamp 1606120353
transform 1 0 6716 0 1 52768
box 0 -48 1196 592
use sky130_fd_sc_hd__a2bb2oi_4  _0781_
timestamp 1606120353
transform 1 0 6808 0 -1 52768
box 0 -48 1932 592
use sky130_fd_sc_hd__fill_2  FILLER_93_74
timestamp 1606120353
transform 1 0 7912 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_93_78
timestamp 1606120353
transform 1 0 8280 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__A
timestamp 1606120353
transform 1 0 8096 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_93_82
timestamp 1606120353
transform 1 0 8648 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__C
timestamp 1606120353
transform 1 0 8464 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_93_86
timestamp 1606120353
transform 1 0 9016 0 1 52768
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_92_83
timestamp 1606120353
transform 1 0 8740 0 -1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__B1
timestamp 1606120353
transform 1 0 9016 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__B
timestamp 1606120353
transform 1 0 8832 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_88
timestamp 1606120353
transform 1 0 9200 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_93_93
timestamp 1606120353
transform 1 0 9660 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_96
timestamp 1606120353
transform 1 0 9936 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_92
timestamp 1606120353
transform 1 0 9568 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__A2
timestamp 1606120353
transform 1 0 9384 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__A1
timestamp 1606120353
transform 1 0 9384 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__A1
timestamp 1606120353
transform 1 0 9844 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__D1
timestamp 1606120353
transform 1 0 9752 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__B1
timestamp 1606120353
transform 1 0 10120 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1606120353
transform 1 0 9568 0 1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_93_110
timestamp 1606120353
transform 1 0 11224 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1143_
timestamp 1606120353
transform 1 0 10028 0 1 52768
box 0 -48 1196 592
use sky130_fd_sc_hd__nand3_4  _0636_
timestamp 1606120353
transform 1 0 10304 0 -1 52768
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_93_114
timestamp 1606120353
transform 1 0 11592 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_120
timestamp 1606120353
transform 1 0 12144 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_92_114
timestamp 1606120353
transform 1 0 11592 0 -1 52768
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__A2
timestamp 1606120353
transform 1 0 11408 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0624__C
timestamp 1606120353
transform 1 0 11960 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__B
timestamp 1606120353
transform 1 0 11776 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_93_132
timestamp 1606120353
transform 1 0 13248 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1606120353
transform 1 0 12328 0 -1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__o21ai_4  _1140_
timestamp 1606120353
transform 1 0 12420 0 -1 52768
box 0 -48 1196 592
use sky130_fd_sc_hd__nand3_4  _0624_
timestamp 1606120353
transform 1 0 11960 0 1 52768
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_93_143
timestamp 1606120353
transform 1 0 14260 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_93_136
timestamp 1606120353
transform 1 0 13616 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_140
timestamp 1606120353
transform 1 0 13984 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_136
timestamp 1606120353
transform 1 0 13616 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__D
timestamp 1606120353
transform 1 0 13800 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__A2
timestamp 1606120353
transform 1 0 13800 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__A
timestamp 1606120353
transform 1 0 14168 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__A
timestamp 1606120353
transform 1 0 13432 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0528_
timestamp 1606120353
transform 1 0 13984 0 1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_93_154
timestamp 1606120353
transform 1 0 15272 0 1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_93_147
timestamp 1606120353
transform 1 0 14628 0 1 52768
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__B
timestamp 1606120353
transform 1 0 14996 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0528__A
timestamp 1606120353
transform 1 0 14444 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1606120353
transform 1 0 15180 0 1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__nand4_4  _1126_
timestamp 1606120353
transform 1 0 14352 0 -1 52768
box 0 -48 1564 592
use sky130_fd_sc_hd__fill_2  FILLER_92_165
timestamp 1606120353
transform 1 0 16284 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_161
timestamp 1606120353
transform 1 0 15916 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__B
timestamp 1606120353
transform 1 0 16100 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_93_176
timestamp 1606120353
transform 1 0 17296 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_93_172
timestamp 1606120353
transform 1 0 16928 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_92_175
timestamp 1606120353
transform 1 0 17204 0 -1 52768
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_92_169
timestamp 1606120353
transform 1 0 16652 0 -1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__C
timestamp 1606120353
transform 1 0 16468 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__D
timestamp 1606120353
transform 1 0 17112 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1132_
timestamp 1606120353
transform 1 0 16928 0 -1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__nand4_4  _1097_
timestamp 1606120353
transform 1 0 15364 0 1 52768
box 0 -48 1564 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1606120353
transform -1 0 18860 0 -1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1606120353
transform -1 0 18860 0 1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1606120353
transform 1 0 17940 0 -1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__C
timestamp 1606120353
transform 1 0 17480 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__C
timestamp 1606120353
transform 1 0 17848 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_92_184
timestamp 1606120353
transform 1 0 18032 0 -1 52768
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_93_180
timestamp 1606120353
transform 1 0 17664 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_93_184
timestamp 1606120353
transform 1 0 18032 0 1 52768
box 0 -48 552 592
use sky130_fd_sc_hd__o21a_4  _0858_
timestamp 1606120353
transform 1 0 2852 0 -1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1606120353
transform 1 0 1104 0 -1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A2
timestamp 1606120353
transform 1 0 1564 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__B
timestamp 1606120353
transform 1 0 2208 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__A2
timestamp 1606120353
transform 1 0 2668 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_3
timestamp 1606120353
transform 1 0 1380 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_94_7
timestamp 1606120353
transform 1 0 1748 0 -1 53856
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_94_11
timestamp 1606120353
transform 1 0 2116 0 -1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_94_14
timestamp 1606120353
transform 1 0 2392 0 -1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__or2_4  _0866_
timestamp 1606120353
transform 1 0 4692 0 -1 53856
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__D
timestamp 1606120353
transform 1 0 4232 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_94_31
timestamp 1606120353
transform 1 0 3956 0 -1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_94_36
timestamp 1606120353
transform 1 0 4416 0 -1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_94_46
timestamp 1606120353
transform 1 0 5336 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_50
timestamp 1606120353
transform 1 0 5704 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_clk_A
timestamp 1606120353
transform 1 0 5520 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__D
timestamp 1606120353
transform 1 0 5888 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_clk
timestamp 1606120353
transform 1 0 6072 0 -1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_94_57
timestamp 1606120353
transform 1 0 6348 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A2
timestamp 1606120353
transform 1 0 6532 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_62
timestamp 1606120353
transform 1 0 6808 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1606120353
transform 1 0 6716 0 -1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0545_
timestamp 1606120353
transform 1 0 6992 0 -1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__nand4_4  _0764_
timestamp 1606120353
transform 1 0 8004 0 -1 53856
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__C
timestamp 1606120353
transform 1 0 7636 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_94_67
timestamp 1606120353
transform 1 0 7268 0 -1 53856
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_94_73
timestamp 1606120353
transform 1 0 7820 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1142_
timestamp 1606120353
transform 1 0 10396 0 -1 53856
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__A2
timestamp 1606120353
transform 1 0 9752 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__B1
timestamp 1606120353
transform 1 0 10120 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_92
timestamp 1606120353
transform 1 0 9568 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_96
timestamp 1606120353
transform 1 0 9936 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_94_100
timestamp 1606120353
transform 1 0 10304 0 -1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__nand3_4  _0635_
timestamp 1606120353
transform 1 0 12420 0 -1 53856
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1606120353
transform 1 0 12328 0 -1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0624__A
timestamp 1606120353
transform 1 0 11960 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_94_114
timestamp 1606120353
transform 1 0 11592 0 -1 53856
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_94_120
timestamp 1606120353
transform 1 0 12144 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _1102_
timestamp 1606120353
transform 1 0 15272 0 -1 53856
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__A
timestamp 1606120353
transform 1 0 15088 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__A
timestamp 1606120353
transform 1 0 14720 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__D
timestamp 1606120353
transform 1 0 14352 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A2
timestamp 1606120353
transform 1 0 13892 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_137
timestamp 1606120353
transform 1 0 13708 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_94_141
timestamp 1606120353
transform 1 0 14076 0 -1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_94_146
timestamp 1606120353
transform 1 0 14536 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_150
timestamp 1606120353
transform 1 0 14904 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0624__B
timestamp 1606120353
transform 1 0 17020 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_171
timestamp 1606120353
transform 1 0 16836 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_94_175
timestamp 1606120353
transform 1 0 17204 0 -1 53856
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1606120353
transform -1 0 18860 0 -1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1606120353
transform 1 0 17940 0 -1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_94_184
timestamp 1606120353
transform 1 0 18032 0 -1 53856
box 0 -48 552 592
use sky130_fd_sc_hd__a21bo_4  _0796_
timestamp 1606120353
transform 1 0 1380 0 1 53856
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1606120353
transform 1 0 1104 0 1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__A
timestamp 1606120353
transform 1 0 2760 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_16
timestamp 1606120353
transform 1 0 2576 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_95_20
timestamp 1606120353
transform 1 0 2944 0 1 53856
box 0 -48 736 592
use sky130_fd_sc_hd__or2_4  _0857_
timestamp 1606120353
transform 1 0 4048 0 1 53856
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1606120353
transform 1 0 3956 0 1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__B
timestamp 1606120353
transform 1 0 4876 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__A
timestamp 1606120353
transform 1 0 3772 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_95_28
timestamp 1606120353
transform 1 0 3680 0 1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_95_39
timestamp 1606120353
transform 1 0 4692 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_43
timestamp 1606120353
transform 1 0 5060 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_47
timestamp 1606120353
transform 1 0 5428 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__A
timestamp 1606120353
transform 1 0 5244 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_clk_A
timestamp 1606120353
transform 1 0 5612 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_51
timestamp 1606120353
transform 1 0 5796 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__C
timestamp 1606120353
transform 1 0 5980 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_clk
timestamp 1606120353
transform 1 0 6164 0 1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_95_58
timestamp 1606120353
transform 1 0 6440 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0525_
timestamp 1606120353
transform 1 0 6624 0 1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_95_63
timestamp 1606120353
transform 1 0 6900 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0525__A
timestamp 1606120353
transform 1 0 7084 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__nor3_4  _0763_
timestamp 1606120353
transform 1 0 7636 0 1 53856
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A
timestamp 1606120353
transform 1 0 7452 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A
timestamp 1606120353
transform 1 0 9016 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_67
timestamp 1606120353
transform 1 0 7268 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_84
timestamp 1606120353
transform 1 0 8832 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_88
timestamp 1606120353
transform 1 0 9200 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0765_
timestamp 1606120353
transform 1 0 9660 0 1 53856
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1606120353
transform 1 0 9568 0 1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__A1
timestamp 1606120353
transform 1 0 9384 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0581__A
timestamp 1606120353
transform 1 0 11040 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_106
timestamp 1606120353
transform 1 0 10856 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_110
timestamp 1606120353
transform 1 0 11224 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__nand3_4  _0640_
timestamp 1606120353
transform 1 0 12052 0 1 53856
box 0 -48 1288 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_clk
timestamp 1606120353
transform 1 0 11592 0 1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0581__B
timestamp 1606120353
transform 1 0 11408 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_117
timestamp 1606120353
transform 1 0 11868 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_137
timestamp 1606120353
transform 1 0 13708 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_133
timestamp 1606120353
transform 1 0 13340 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__D
timestamp 1606120353
transform 1 0 13892 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__D
timestamp 1606120353
transform 1 0 13524 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0550_
timestamp 1606120353
transform 1 0 14076 0 1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_95_148
timestamp 1606120353
transform 1 0 14720 0 1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_95_144
timestamp 1606120353
transform 1 0 14352 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__A
timestamp 1606120353
transform 1 0 14996 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0550__A
timestamp 1606120353
transform 1 0 14536 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1606120353
transform 1 0 15180 0 1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__nand4_4  _1136_
timestamp 1606120353
transform 1 0 15272 0 1 53856
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A1
timestamp 1606120353
transform 1 0 17020 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_171
timestamp 1606120353
transform 1 0 16836 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_175
timestamp 1606120353
transform 1 0 17204 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1606120353
transform -1 0 18860 0 1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A2
timestamp 1606120353
transform 1 0 17388 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__B1
timestamp 1606120353
transform 1 0 17756 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_179
timestamp 1606120353
transform 1 0 17572 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_95_183
timestamp 1606120353
transform 1 0 17940 0 1 53856
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_95_189
timestamp 1606120353
transform 1 0 18492 0 1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__nand2_4  _0795_
timestamp 1606120353
transform 1 0 2208 0 -1 54944
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1606120353
transform 1 0 1104 0 -1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__B1_N
timestamp 1606120353
transform 1 0 1564 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A1
timestamp 1606120353
transform 1 0 1932 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_3
timestamp 1606120353
transform 1 0 1380 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_7
timestamp 1606120353
transform 1 0 1748 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_96_11
timestamp 1606120353
transform 1 0 2116 0 -1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_96_21
timestamp 1606120353
transform 1 0 3036 0 -1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__inv_8  _0756_
timestamp 1606120353
transform 1 0 5152 0 -1 54944
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__B
timestamp 1606120353
transform 1 0 4600 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_clk_A
timestamp 1606120353
transform 1 0 4968 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__CLK
timestamp 1606120353
transform 1 0 4232 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_96_33
timestamp 1606120353
transform 1 0 4140 0 -1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_96_36
timestamp 1606120353
transform 1 0 4416 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_40
timestamp 1606120353
transform 1 0 4784 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1606120353
transform 1 0 6716 0 -1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A
timestamp 1606120353
transform 1 0 7084 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__B1
timestamp 1606120353
transform 1 0 6532 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A1
timestamp 1606120353
transform 1 0 6164 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_53
timestamp 1606120353
transform 1 0 5980 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_57
timestamp 1606120353
transform 1 0 6348 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_96_62
timestamp 1606120353
transform 1 0 6808 0 -1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__nand3_4  _0708_
timestamp 1606120353
transform 1 0 8832 0 -1 54944
box 0 -48 1288 592
use sky130_fd_sc_hd__inv_8  _0738_
timestamp 1606120353
transform 1 0 7268 0 -1 54944
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__B
timestamp 1606120353
transform 1 0 8648 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__B
timestamp 1606120353
transform 1 0 8280 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_76
timestamp 1606120353
transform 1 0 8096 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_80
timestamp 1606120353
transform 1 0 8464 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0581_
timestamp 1606120353
transform 1 0 10856 0 -1 54944
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__B1
timestamp 1606120353
transform 1 0 10396 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_96_98
timestamp 1606120353
transform 1 0 10120 0 -1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_96_103
timestamp 1606120353
transform 1 0 10580 0 -1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_96_121
timestamp 1606120353
transform 1 0 12236 0 -1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_96_117
timestamp 1606120353
transform 1 0 11868 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_113
timestamp 1606120353
transform 1 0 11500 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0640__C
timestamp 1606120353
transform 1 0 11684 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0640__A
timestamp 1606120353
transform 1 0 12052 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_96_127
timestamp 1606120353
transform 1 0 12788 0 -1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_96_123
timestamp 1606120353
transform 1 0 12420 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__B1
timestamp 1606120353
transform 1 0 13064 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0640__B
timestamp 1606120353
transform 1 0 12604 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1606120353
transform 1 0 12328 0 -1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1188_
timestamp 1606120353
transform 1 0 13248 0 -1 54944
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__B
timestamp 1606120353
transform 1 0 15272 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_96_151
timestamp 1606120353
transform 1 0 14996 0 -1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _1139_
timestamp 1606120353
transform 1 0 16008 0 -1 54944
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__C
timestamp 1606120353
transform 1 0 15640 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_156
timestamp 1606120353
transform 1 0 15456 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_160
timestamp 1606120353
transform 1 0 15824 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_96_175
timestamp 1606120353
transform 1 0 17204 0 -1 54944
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1606120353
transform -1 0 18860 0 -1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1606120353
transform 1 0 17940 0 -1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_96_184
timestamp 1606120353
transform 1 0 18032 0 -1 54944
box 0 -48 552 592
use sky130_fd_sc_hd__buf_1  _0794_
timestamp 1606120353
transform 1 0 2944 0 1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1606120353
transform 1 0 1104 0 1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__CLK
timestamp 1606120353
transform 1 0 1564 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_3
timestamp 1606120353
transform 1 0 1380 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_97_7
timestamp 1606120353
transform 1 0 1748 0 1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_97_19
timestamp 1606120353
transform 1 0 2852 0 1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_97_23
timestamp 1606120353
transform 1 0 3220 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A
timestamp 1606120353
transform 1 0 3404 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_27
timestamp 1606120353
transform 1 0 3588 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A
timestamp 1606120353
transform 1 0 3772 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_32
timestamp 1606120353
transform 1 0 4048 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1606120353
transform 1 0 3956 0 1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0874_
timestamp 1606120353
transform 1 0 4232 0 1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_97_37
timestamp 1606120353
transform 1 0 4508 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_97_41
timestamp 1606120353
transform 1 0 4876 0 1 54944
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A
timestamp 1606120353
transform 1 0 4692 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0851_
timestamp 1606120353
transform 1 0 5428 0 1 54944
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__A1
timestamp 1606120353
transform 1 0 7176 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A2
timestamp 1606120353
transform 1 0 6808 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A2
timestamp 1606120353
transform 1 0 5244 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_60
timestamp 1606120353
transform 1 0 6624 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_64
timestamp 1606120353
transform 1 0 6992 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0806_
timestamp 1606120353
transform 1 0 7360 0 1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__B1
timestamp 1606120353
transform 1 0 8648 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__B2
timestamp 1606120353
transform 1 0 9016 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_80
timestamp 1606120353
transform 1 0 8464 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_84
timestamp 1606120353
transform 1 0 8832 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_88
timestamp 1606120353
transform 1 0 9200 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_96
timestamp 1606120353
transform 1 0 9936 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__A
timestamp 1606120353
transform 1 0 9384 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A
timestamp 1606120353
transform 1 0 10120 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1606120353
transform 1 0 9568 0 1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0730_
timestamp 1606120353
transform 1 0 9660 0 1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_97_104
timestamp 1606120353
transform 1 0 10672 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_100
timestamp 1606120353
transform 1 0 10304 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A1
timestamp 1606120353
transform 1 0 10856 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__B
timestamp 1606120353
transform 1 0 10488 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__a22oi_4  _0674_
timestamp 1606120353
transform 1 0 11040 0 1 54944
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__D
timestamp 1606120353
transform 1 0 13156 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__A
timestamp 1606120353
transform 1 0 12788 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_125
timestamp 1606120353
transform 1 0 12604 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_129
timestamp 1606120353
transform 1 0 12972 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _1138_
timestamp 1606120353
transform 1 0 13340 0 1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1186_
timestamp 1606120353
transform 1 0 15272 0 1 54944
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1606120353
transform 1 0 15180 0 1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__D
timestamp 1606120353
transform 1 0 14996 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__A2
timestamp 1606120353
transform 1 0 14628 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_145
timestamp 1606120353
transform 1 0 14444 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_149
timestamp 1606120353
transform 1 0 14812 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__A1
timestamp 1606120353
transform 1 0 17204 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_173
timestamp 1606120353
transform 1 0 17020 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1606120353
transform -1 0 18860 0 1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__A2
timestamp 1606120353
transform 1 0 17572 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_177
timestamp 1606120353
transform 1 0 17388 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_97_181
timestamp 1606120353
transform 1 0 17756 0 1 54944
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_97_189
timestamp 1606120353
transform 1 0 18492 0 1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1606120353
transform 1 0 1104 0 -1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__B
timestamp 1606120353
transform 1 0 2208 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__D
timestamp 1606120353
transform 1 0 1564 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_3
timestamp 1606120353
transform 1 0 1380 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_98_7
timestamp 1606120353
transform 1 0 1748 0 -1 56032
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_98_11
timestamp 1606120353
transform 1 0 2116 0 -1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_98_14
timestamp 1606120353
transform 1 0 2392 0 -1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__nand2_4  _0868_
timestamp 1606120353
transform 1 0 4600 0 -1 56032
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__D
timestamp 1606120353
transform 1 0 4048 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A1
timestamp 1606120353
transform 1 0 4416 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__CLK
timestamp 1606120353
transform 1 0 3680 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_26
timestamp 1606120353
transform 1 0 3496 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_30
timestamp 1606120353
transform 1 0 3864 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_34
timestamp 1606120353
transform 1 0 4232 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0813_
timestamp 1606120353
transform 1 0 6808 0 -1 56032
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1606120353
transform 1 0 6716 0 -1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_clk
timestamp 1606120353
transform 1 0 6440 0 -1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A1
timestamp 1606120353
transform 1 0 5612 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__B1
timestamp 1606120353
transform 1 0 5980 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_47
timestamp 1606120353
transform 1 0 5428 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_51
timestamp 1606120353
transform 1 0 5796 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_98_55
timestamp 1606120353
transform 1 0 6164 0 -1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__B
timestamp 1606120353
transform 1 0 9200 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__A2
timestamp 1606120353
transform 1 0 8188 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__D
timestamp 1606120353
transform 1 0 8832 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_75
timestamp 1606120353
transform 1 0 8004 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_98_79
timestamp 1606120353
transform 1 0 8372 0 -1 56032
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1606120353
transform 1 0 8740 0 -1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_98_86
timestamp 1606120353
transform 1 0 9016 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__nand3_4  _0579_
timestamp 1606120353
transform 1 0 9660 0 -1 56032
box 0 -48 1288 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_clk
timestamp 1606120353
transform 1 0 9384 0 -1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__B1
timestamp 1606120353
transform 1 0 11132 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_107
timestamp 1606120353
transform 1 0 10948 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_111
timestamp 1606120353
transform 1 0 11316 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A2
timestamp 1606120353
transform 1 0 11500 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_115
timestamp 1606120353
transform 1 0 11684 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A2
timestamp 1606120353
transform 1 0 11868 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_clk
timestamp 1606120353
transform 1 0 12052 0 -1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1606120353
transform 1 0 12328 0 -1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0576_
timestamp 1606120353
transform 1 0 12420 0 -1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_98_126
timestamp 1606120353
transform 1 0 12696 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__C
timestamp 1606120353
transform 1 0 12880 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_98_130
timestamp 1606120353
transform 1 0 13064 0 -1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1193_
timestamp 1606120353
transform 1 0 13616 0 -1 56032
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__A1
timestamp 1606120353
transform 1 0 13340 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_98_135
timestamp 1606120353
transform 1 0 13524 0 -1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__o21a_4  _1141_
timestamp 1606120353
transform 1 0 16100 0 -1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__B1
timestamp 1606120353
transform 1 0 15916 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__CLK
timestamp 1606120353
transform 1 0 15548 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_155
timestamp 1606120353
transform 1 0 15364 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_159
timestamp 1606120353
transform 1 0 15732 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_98_175
timestamp 1606120353
transform 1 0 17204 0 -1 56032
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1606120353
transform -1 0 18860 0 -1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1606120353
transform 1 0 17940 0 -1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_98_184
timestamp 1606120353
transform 1 0 18032 0 -1 56032
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_100_3
timestamp 1606120353
transform 1 0 1380 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_99_7
timestamp 1606120353
transform 1 0 1748 0 1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_99_3
timestamp 1606120353
transform 1 0 1380 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__B1_N
timestamp 1606120353
transform 1 0 1564 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A
timestamp 1606120353
transform 1 0 2024 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1606120353
transform 1 0 1104 0 -1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1606120353
transform 1 0 1104 0 1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_99_21
timestamp 1606120353
transform 1 0 3036 0 1 56032
box 0 -48 368 592
use sky130_fd_sc_hd__nand2_4  _0817_
timestamp 1606120353
transform 1 0 2208 0 1 56032
box 0 -48 828 592
use sky130_fd_sc_hd__dfxtp_4  _1151_
timestamp 1606120353
transform 1 0 1564 0 -1 57120
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_1  FILLER_100_33
timestamp 1606120353
transform 1 0 4140 0 -1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_100_28
timestamp 1606120353
transform 1 0 3680 0 -1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_100_24
timestamp 1606120353
transform 1 0 3312 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_27
timestamp 1606120353
transform 1 0 3588 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__CLK
timestamp 1606120353
transform 1 0 3404 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A1
timestamp 1606120353
transform 1 0 3496 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__D
timestamp 1606120353
transform 1 0 3772 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A2
timestamp 1606120353
transform 1 0 3956 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1606120353
transform 1 0 3956 0 1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1163_
timestamp 1606120353
transform 1 0 4048 0 1 56032
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1161_
timestamp 1606120353
transform 1 0 4232 0 -1 57120
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_2  FILLER_100_53
timestamp 1606120353
transform 1 0 5980 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_55
timestamp 1606120353
transform 1 0 6164 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_51
timestamp 1606120353
transform 1 0 5796 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__B1
timestamp 1606120353
transform 1 0 6164 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A2
timestamp 1606120353
transform 1 0 5980 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_100_57
timestamp 1606120353
transform 1 0 6348 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A2
timestamp 1606120353
transform 1 0 6532 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__B1
timestamp 1606120353
transform 1 0 6348 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1606120353
transform 1 0 6716 0 -1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__o21ai_4  _0860_
timestamp 1606120353
transform 1 0 6808 0 -1 57120
box 0 -48 1196 592
use sky130_fd_sc_hd__o21ai_4  _0824_
timestamp 1606120353
transform 1 0 6532 0 1 56032
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_100_75
timestamp 1606120353
transform 1 0 8004 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_99_76
timestamp 1606120353
transform 1 0 8096 0 1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_99_72
timestamp 1606120353
transform 1 0 7728 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__B1
timestamp 1606120353
transform 1 0 8188 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A1
timestamp 1606120353
transform 1 0 7912 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_100_86
timestamp 1606120353
transform 1 0 9016 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1606120353
transform 1 0 8740 0 -1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_100_79
timestamp 1606120353
transform 1 0 8372 0 -1 57120
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_99_84
timestamp 1606120353
transform 1 0 8832 0 1 56032
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A2
timestamp 1606120353
transform 1 0 8832 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0536__A
timestamp 1606120353
transform 1 0 8372 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__C
timestamp 1606120353
transform 1 0 9200 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0536_
timestamp 1606120353
transform 1 0 8556 0 1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__nand4_4  _0737_
timestamp 1606120353
transform 1 0 9200 0 -1 57120
box 0 -48 1564 592
use sky130_fd_sc_hd__a21bo_4  _0709_
timestamp 1606120353
transform 1 0 10120 0 1 56032
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1606120353
transform 1 0 9568 0 1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__A
timestamp 1606120353
transform 1 0 9844 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__A
timestamp 1606120353
transform 1 0 11132 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_90
timestamp 1606120353
transform 1 0 9384 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_93
timestamp 1606120353
transform 1 0 9660 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_99_97
timestamp 1606120353
transform 1 0 10028 0 1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_100_105
timestamp 1606120353
transform 1 0 10764 0 -1 57120
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_100_116
timestamp 1606120353
transform 1 0 11776 0 -1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_100_111
timestamp 1606120353
transform 1 0 11316 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_115
timestamp 1606120353
transform 1 0 11684 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_111
timestamp 1606120353
transform 1 0 11316 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A
timestamp 1606120353
transform 1 0 12052 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A1
timestamp 1606120353
transform 1 0 11868 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__B1_N
timestamp 1606120353
transform 1 0 11500 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_clk
timestamp 1606120353
transform 1 0 11500 0 -1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _0805_
timestamp 1606120353
transform 1 0 12052 0 1 56032
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILLER_100_121
timestamp 1606120353
transform 1 0 12236 0 -1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_99_128
timestamp 1606120353
transform 1 0 12880 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1606120353
transform 1 0 12328 0 -1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _0762_
timestamp 1606120353
transform 1 0 12420 0 -1 57120
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_100_132
timestamp 1606120353
transform 1 0 13248 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_132
timestamp 1606120353
transform 1 0 13248 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__A
timestamp 1606120353
transform 1 0 13064 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_100_136
timestamp 1606120353
transform 1 0 13616 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_140
timestamp 1606120353
transform 1 0 13984 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_136
timestamp 1606120353
transform 1 0 13616 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__CLK
timestamp 1606120353
transform 1 0 13800 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__CLK
timestamp 1606120353
transform 1 0 14168 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_clk_A
timestamp 1606120353
transform 1 0 13432 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_clk_A
timestamp 1606120353
transform 1 0 13800 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_clk_A
timestamp 1606120353
transform 1 0 13432 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_100_152
timestamp 1606120353
transform 1 0 15088 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_154
timestamp 1606120353
transform 1 0 15272 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_149
timestamp 1606120353
transform 1 0 14812 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_99_144
timestamp 1606120353
transform 1 0 14352 0 1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__CLK
timestamp 1606120353
transform 1 0 14628 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__CLK
timestamp 1606120353
transform 1 0 14996 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1606120353
transform 1 0 15180 0 1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_100_140
timestamp 1606120353
transform 1 0 13984 0 -1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1185_
timestamp 1606120353
transform 1 0 15272 0 -1 57120
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1194_
timestamp 1606120353
transform 1 0 16100 0 1 56032
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__D
timestamp 1606120353
transform 1 0 15916 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__D
timestamp 1606120353
transform 1 0 15456 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_99_158
timestamp 1606120353
transform 1 0 15640 0 1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_100_173
timestamp 1606120353
transform 1 0 17020 0 -1 57120
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1606120353
transform -1 0 18860 0 1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1606120353
transform -1 0 18860 0 -1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1606120353
transform 1 0 17940 0 -1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_99_182
timestamp 1606120353
transform 1 0 17848 0 1 56032
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_100_181
timestamp 1606120353
transform 1 0 17756 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_100_184
timestamp 1606120353
transform 1 0 18032 0 -1 57120
box 0 -48 552 592
use sky130_fd_sc_hd__o21a_4  _0869_
timestamp 1606120353
transform 1 0 2116 0 1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1606120353
transform 1 0 1104 0 1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__A2
timestamp 1606120353
transform 1 0 1564 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A2
timestamp 1606120353
transform 1 0 1932 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_3
timestamp 1606120353
transform 1 0 1380 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_7
timestamp 1606120353
transform 1 0 1748 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_23
timestamp 1606120353
transform 1 0 3220 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__B1
timestamp 1606120353
transform 1 0 3404 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_27
timestamp 1606120353
transform 1 0 3588 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__B1
timestamp 1606120353
transform 1 0 3772 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_32
timestamp 1606120353
transform 1 0 4048 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A1
timestamp 1606120353
transform 1 0 4232 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1606120353
transform 1 0 3956 0 1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_101_36
timestamp 1606120353
transform 1 0 4416 0 1 57120
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_101_40
timestamp 1606120353
transform 1 0 4784 0 1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A2
timestamp 1606120353
transform 1 0 4876 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_43
timestamp 1606120353
transform 1 0 5060 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__a2bb2oi_4  _0816_
timestamp 1606120353
transform 1 0 5796 0 1 57120
box 0 -48 1932 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A2_N
timestamp 1606120353
transform 1 0 5612 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__B2
timestamp 1606120353
transform 1 0 5244 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_47
timestamp 1606120353
transform 1 0 5428 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__B2
timestamp 1606120353
transform 1 0 7912 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__B1
timestamp 1606120353
transform 1 0 8832 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A1
timestamp 1606120353
transform 1 0 8280 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A1
timestamp 1606120353
transform 1 0 9200 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_72
timestamp 1606120353
transform 1 0 7728 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_76
timestamp 1606120353
transform 1 0 8096 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_101_80
timestamp 1606120353
transform 1 0 8464 0 1 57120
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_101_86
timestamp 1606120353
transform 1 0 9016 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_101_93
timestamp 1606120353
transform 1 0 9660 0 1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_101_90
timestamp 1606120353
transform 1 0 9384 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A
timestamp 1606120353
transform 1 0 9936 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1606120353
transform 1 0 9568 0 1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0539_
timestamp 1606120353
transform 1 0 10120 0 1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_101_105
timestamp 1606120353
transform 1 0 10764 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_101
timestamp 1606120353
transform 1 0 10396 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0539__A
timestamp 1606120353
transform 1 0 10580 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__C
timestamp 1606120353
transform 1 0 10948 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__nand3_4  _0639_
timestamp 1606120353
transform 1 0 11132 0 1 57120
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__B
timestamp 1606120353
transform 1 0 12604 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__A
timestamp 1606120353
transform 1 0 12972 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_123
timestamp 1606120353
transform 1 0 12420 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_127
timestamp 1606120353
transform 1 0 12788 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_131
timestamp 1606120353
transform 1 0 13156 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1606120353
transform 1 0 15180 0 1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__C
timestamp 1606120353
transform 1 0 13340 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_101_135
timestamp 1606120353
transform 1 0 13524 0 1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_101_147
timestamp 1606120353
transform 1 0 14628 0 1 57120
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILLER_101_154
timestamp 1606120353
transform 1 0 15272 0 1 57120
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1195_
timestamp 1606120353
transform 1 0 15916 0 1 57120
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__D
timestamp 1606120353
transform 1 0 15732 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_101_158
timestamp 1606120353
transform 1 0 15640 0 1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1606120353
transform -1 0 18860 0 1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_101_180
timestamp 1606120353
transform 1 0 17664 0 1 57120
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_101_188
timestamp 1606120353
transform 1 0 18400 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0818_
timestamp 1606120353
transform 1 0 1380 0 -1 58208
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1606120353
transform 1 0 1104 0 -1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A1
timestamp 1606120353
transform 1 0 2760 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A2
timestamp 1606120353
transform 1 0 3128 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_102_16
timestamp 1606120353
transform 1 0 2576 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_102_20
timestamp 1606120353
transform 1 0 2944 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0865_
timestamp 1606120353
transform 1 0 3956 0 -1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_clk_A
timestamp 1606120353
transform 1 0 3772 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_102_24
timestamp 1606120353
transform 1 0 3312 0 -1 58208
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_102_28
timestamp 1606120353
transform 1 0 3680 0 -1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_102_43
timestamp 1606120353
transform 1 0 5060 0 -1 58208
box 0 -48 368 592
use sky130_fd_sc_hd__o22a_4  _0821_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 6808 0 -1 58208
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1606120353
transform 1 0 6716 0 -1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_clk
timestamp 1606120353
transform 1 0 6440 0 -1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A1
timestamp 1606120353
transform 1 0 5428 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__B1
timestamp 1606120353
transform 1 0 5796 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A2
timestamp 1606120353
transform 1 0 6256 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_102_49
timestamp 1606120353
transform 1 0 5612 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_102_53
timestamp 1606120353
transform 1 0 5980 0 -1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__o21a_4  _0814_
timestamp 1606120353
transform 1 0 8832 0 -1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__C
timestamp 1606120353
transform 1 0 8464 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_102_76
timestamp 1606120353
transform 1 0 8096 0 -1 58208
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_102_82
timestamp 1606120353
transform 1 0 8648 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0819_
timestamp 1606120353
transform 1 0 10672 0 -1 58208
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A
timestamp 1606120353
transform 1 0 10120 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_clk_A
timestamp 1606120353
transform 1 0 10488 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_102_96
timestamp 1606120353
transform 1 0 9936 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_102_100
timestamp 1606120353
transform 1 0 10304 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__nand3_4  _0621_
timestamp 1606120353
transform 1 0 12420 0 -1 58208
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1606120353
transform 1 0 12328 0 -1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__B
timestamp 1606120353
transform 1 0 11684 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_102_113
timestamp 1606120353
transform 1 0 11500 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_102_117
timestamp 1606120353
transform 1 0 11868 0 -1 58208
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_102_121
timestamp 1606120353
transform 1 0 12236 0 -1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__D
timestamp 1606120353
transform 1 0 13892 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__CLK
timestamp 1606120353
transform 1 0 14260 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_102_137
timestamp 1606120353
transform 1 0 13708 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_102_141
timestamp 1606120353
transform 1 0 14076 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_102_145
timestamp 1606120353
transform 1 0 14444 0 -1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__CLK
timestamp 1606120353
transform 1 0 15916 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_102_157
timestamp 1606120353
transform 1 0 15548 0 -1 58208
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_102_163
timestamp 1606120353
transform 1 0 16100 0 -1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_102_175
timestamp 1606120353
transform 1 0 17204 0 -1 58208
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1606120353
transform -1 0 18860 0 -1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1606120353
transform 1 0 17940 0 -1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_102_184
timestamp 1606120353
transform 1 0 18032 0 -1 58208
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1152_
timestamp 1606120353
transform 1 0 1472 0 1 58208
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1606120353
transform 1 0 1104 0 1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_103_3
timestamp 1606120353
transform 1 0 1380 0 1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_103_23
timestamp 1606120353
transform 1 0 3220 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__A
timestamp 1606120353
transform 1 0 3404 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_103_27
timestamp 1606120353
transform 1 0 3588 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__B2
timestamp 1606120353
transform 1 0 3772 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1606120353
transform 1 0 3956 0 1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0705_
timestamp 1606120353
transform 1 0 4048 0 1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_103_35
timestamp 1606120353
transform 1 0 4324 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A
timestamp 1606120353
transform 1 0 4508 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_103_39
timestamp 1606120353
transform 1 0 4692 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_103_43
timestamp 1606120353
transform 1 0 5060 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__B1
timestamp 1606120353
transform 1 0 4876 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__a22oi_4  _0825_
timestamp 1606120353
transform 1 0 5428 0 1 58208
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A2
timestamp 1606120353
transform 1 0 7176 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A2
timestamp 1606120353
transform 1 0 5244 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_103_64
timestamp 1606120353
transform 1 0 6992 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0815_
timestamp 1606120353
transform 1 0 7728 0 1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__B
timestamp 1606120353
transform 1 0 9016 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A
timestamp 1606120353
transform 1 0 7544 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_103_68
timestamp 1606120353
transform 1 0 7360 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_103_84
timestamp 1606120353
transform 1 0 8832 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_103_88
timestamp 1606120353
transform 1 0 9200 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__nor3_4  _0729_
timestamp 1606120353
transform 1 0 9660 0 1 58208
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1606120353
transform 1 0 9568 0 1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0549__A
timestamp 1606120353
transform 1 0 11224 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__B
timestamp 1606120353
transform 1 0 9384 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_103_106
timestamp 1606120353
transform 1 0 10856 0 1 58208
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1184_
timestamp 1606120353
transform 1 0 12696 0 1 58208
box 0 -48 1748 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_clk
timestamp 1606120353
transform 1 0 12236 0 1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_clk_A
timestamp 1606120353
transform 1 0 12052 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__CLK
timestamp 1606120353
transform 1 0 11684 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_103_112
timestamp 1606120353
transform 1 0 11408 0 1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_103_117
timestamp 1606120353
transform 1 0 11868 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_103_124
timestamp 1606120353
transform 1 0 12512 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1606120353
transform 1 0 15180 0 1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_clk_A
timestamp 1606120353
transform 1 0 14628 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_103_145
timestamp 1606120353
transform 1 0 14444 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_103_149
timestamp 1606120353
transform 1 0 14812 0 1 58208
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_103_154
timestamp 1606120353
transform 1 0 15272 0 1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_103_166
timestamp 1606120353
transform 1 0 16376 0 1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1606120353
transform -1 0 18860 0 1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_103_178
timestamp 1606120353
transform 1 0 17480 0 1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__a21bo_4  _0827_
timestamp 1606120353
transform 1 0 1380 0 -1 59296
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1606120353
transform 1 0 1104 0 -1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__D
timestamp 1606120353
transform 1 0 2760 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__A1
timestamp 1606120353
transform 1 0 3128 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_104_16
timestamp 1606120353
transform 1 0 2576 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_104_20
timestamp 1606120353
transform 1 0 2944 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0703_
timestamp 1606120353
transform 1 0 3312 0 -1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__a21o_4  _0823_
timestamp 1606120353
transform 1 0 4876 0 -1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A1
timestamp 1606120353
transform 1 0 4692 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__CLK
timestamp 1606120353
transform 1 0 3772 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_104_27
timestamp 1606120353
transform 1 0 3588 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_104_31
timestamp 1606120353
transform 1 0 3956 0 -1 59296
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1606120353
transform 1 0 6716 0 -1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__B
timestamp 1606120353
transform 1 0 6992 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A1
timestamp 1606120353
transform 1 0 6532 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__B1
timestamp 1606120353
transform 1 0 6164 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_104_53
timestamp 1606120353
transform 1 0 5980 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_104_57
timestamp 1606120353
transform 1 0 6348 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_104_62
timestamp 1606120353
transform 1 0 6808 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_104_66
timestamp 1606120353
transform 1 0 7176 0 -1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__nand4_4  _0735_
timestamp 1606120353
transform 1 0 8464 0 -1 59296
box 0 -48 1564 592
use sky130_fd_sc_hd__buf_1  _0744_
timestamp 1606120353
transform 1 0 7452 0 -1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__A
timestamp 1606120353
transform 1 0 7912 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__B1
timestamp 1606120353
transform 1 0 8280 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_104_72
timestamp 1606120353
transform 1 0 7728 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_104_76
timestamp 1606120353
transform 1 0 8096 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0549_
timestamp 1606120353
transform 1 0 11224 0 -1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__C
timestamp 1606120353
transform 1 0 10212 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__A
timestamp 1606120353
transform 1 0 10764 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_104_97
timestamp 1606120353
transform 1 0 10028 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_104_101
timestamp 1606120353
transform 1 0 10396 0 -1 59296
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_104_107
timestamp 1606120353
transform 1 0 10948 0 -1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1606120353
transform 1 0 12328 0 -1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_clk
timestamp 1606120353
transform 1 0 13156 0 -1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__D
timestamp 1606120353
transform 1 0 12696 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__B
timestamp 1606120353
transform 1 0 12144 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__C
timestamp 1606120353
transform 1 0 11776 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_104_113
timestamp 1606120353
transform 1 0 11500 0 -1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_104_118
timestamp 1606120353
transform 1 0 11960 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_104_123
timestamp 1606120353
transform 1 0 12420 0 -1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_104_128
timestamp 1606120353
transform 1 0 12880 0 -1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1192_
timestamp 1606120353
transform 1 0 13432 0 -1 59296
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_8  FILLER_104_153
timestamp 1606120353
transform 1 0 15180 0 -1 59296
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__CLK
timestamp 1606120353
transform 1 0 16100 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_104_161
timestamp 1606120353
transform 1 0 15916 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_104_165
timestamp 1606120353
transform 1 0 16284 0 -1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1606120353
transform -1 0 18860 0 -1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1606120353
transform 1 0 17940 0 -1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_104_177
timestamp 1606120353
transform 1 0 17388 0 -1 59296
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILLER_104_184
timestamp 1606120353
transform 1 0 18032 0 -1 59296
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILLER_106_7
timestamp 1606120353
transform 1 0 1748 0 -1 60384
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_106_3
timestamp 1606120353
transform 1 0 1380 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_105_7
timestamp 1606120353
transform 1 0 1748 0 1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_105_3
timestamp 1606120353
transform 1 0 1380 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__D
timestamp 1606120353
transform 1 0 1564 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__B1_N
timestamp 1606120353
transform 1 0 1564 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1606120353
transform 1 0 1104 0 -1 60384
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1606120353
transform 1 0 1104 0 1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_106_17
timestamp 1606120353
transform 1 0 2668 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_106_13
timestamp 1606120353
transform 1 0 2300 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__B
timestamp 1606120353
transform 1 0 2484 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__B1
timestamp 1606120353
transform 1 0 2116 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__A
timestamp 1606120353
transform 1 0 2024 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__nand2_4  _0826_
timestamp 1606120353
transform 1 0 2208 0 1 59296
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_106_21
timestamp 1606120353
transform 1 0 3036 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_105_21
timestamp 1606120353
transform 1 0 3036 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A2
timestamp 1606120353
transform 1 0 2852 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_105_32
timestamp 1606120353
transform 1 0 4048 0 1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_105_29
timestamp 1606120353
transform 1 0 3772 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_105_25
timestamp 1606120353
transform 1 0 3404 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__CLK
timestamp 1606120353
transform 1 0 3588 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__D
timestamp 1606120353
transform 1 0 3220 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1606120353
transform 1 0 3956 0 1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_106_42
timestamp 1606120353
transform 1 0 4968 0 -1 60384
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_105_37
timestamp 1606120353
transform 1 0 4508 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_clk_A
timestamp 1606120353
transform 1 0 4324 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__A
timestamp 1606120353
transform 1 0 4692 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_clk
timestamp 1606120353
transform 1 0 4876 0 1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _0820_
timestamp 1606120353
transform 1 0 5152 0 1 59296
box 0 -48 828 592
use sky130_fd_sc_hd__dfxtp_4  _1154_
timestamp 1606120353
transform 1 0 3220 0 -1 60384
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  FILLER_106_50
timestamp 1606120353
transform 1 0 5704 0 -1 60384
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_105_53
timestamp 1606120353
transform 1 0 5980 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_clk_A
timestamp 1606120353
transform 1 0 5980 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A1_N
timestamp 1606120353
transform 1 0 6164 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_clk
timestamp 1606120353
transform 1 0 6164 0 -1 60384
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_106_66
timestamp 1606120353
transform 1 0 7176 0 -1 60384
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_106_62
timestamp 1606120353
transform 1 0 6808 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_106_58
timestamp 1606120353
transform 1 0 6440 0 -1 60384
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_105_61
timestamp 1606120353
transform 1 0 6716 0 1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_105_57
timestamp 1606120353
transform 1 0 6348 0 1 59296
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__C
timestamp 1606120353
transform 1 0 6992 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__A
timestamp 1606120353
transform 1 0 6808 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1606120353
transform 1 0 6716 0 -1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__nand3_4  _0822_
timestamp 1606120353
transform 1 0 6992 0 1 59296
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__A
timestamp 1606120353
transform 1 0 7912 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_106_80
timestamp 1606120353
transform 1 0 8464 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_106_76
timestamp 1606120353
transform 1 0 8096 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_105_84
timestamp 1606120353
transform 1 0 8832 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_105_78
timestamp 1606120353
transform 1 0 8280 0 1 59296
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0555__C
timestamp 1606120353
transform 1 0 8280 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A
timestamp 1606120353
transform 1 0 8648 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0736_
timestamp 1606120353
transform 1 0 8648 0 -1 60384
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_105_88
timestamp 1606120353
transform 1 0 9200 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__D
timestamp 1606120353
transform 1 0 9016 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_106_97
timestamp 1606120353
transform 1 0 10028 0 -1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_106_91
timestamp 1606120353
transform 1 0 9476 0 -1 60384
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILLER_105_93
timestamp 1606120353
transform 1 0 9660 0 1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__C
timestamp 1606120353
transform 1 0 9384 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__A
timestamp 1606120353
transform 1 0 10120 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__B
timestamp 1606120353
transform 1 0 9936 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1606120353
transform 1 0 9568 0 1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_106_104
timestamp 1606120353
transform 1 0 10672 0 -1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_106_100
timestamp 1606120353
transform 1 0 10304 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__B
timestamp 1606120353
transform 1 0 10488 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0638_
timestamp 1606120353
transform 1 0 10764 0 -1 60384
box 0 -48 828 592
use sky130_fd_sc_hd__nand3_4  _0580_
timestamp 1606120353
transform 1 0 10120 0 1 59296
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  FILLER_106_119
timestamp 1606120353
transform 1 0 12052 0 -1 60384
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_106_114
timestamp 1606120353
transform 1 0 11592 0 -1 60384
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_105_117
timestamp 1606120353
transform 1 0 11868 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_105_112
timestamp 1606120353
transform 1 0 11408 0 1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__A
timestamp 1606120353
transform 1 0 11868 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__A
timestamp 1606120353
transform 1 0 11684 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__A
timestamp 1606120353
transform 1 0 12052 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1606120353
transform 1 0 12328 0 -1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__nand4_4  _0626_
timestamp 1606120353
transform 1 0 12236 0 1 59296
box 0 -48 1564 592
use sky130_fd_sc_hd__nand3_4  _0623_
timestamp 1606120353
transform 1 0 12420 0 -1 60384
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_106_137
timestamp 1606120353
transform 1 0 13708 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_105_142
timestamp 1606120353
transform 1 0 14168 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_105_138
timestamp 1606120353
transform 1 0 13800 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__C
timestamp 1606120353
transform 1 0 13892 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__B
timestamp 1606120353
transform 1 0 13984 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_106_153
timestamp 1606120353
transform 1 0 15180 0 -1 60384
box 0 -48 736 592
use sky130_fd_sc_hd__decap_6  FILLER_105_154
timestamp 1606120353
transform 1 0 15272 0 1 59296
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_105_152
timestamp 1606120353
transform 1 0 15088 0 1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_105_146
timestamp 1606120353
transform 1 0 14536 0 1 59296
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__D
timestamp 1606120353
transform 1 0 14352 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1606120353
transform 1 0 15180 0 1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_106_141
timestamp 1606120353
transform 1 0 14076 0 -1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1198_
timestamp 1606120353
transform 1 0 16100 0 1 59296
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__D
timestamp 1606120353
transform 1 0 15916 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__CLK
timestamp 1606120353
transform 1 0 16100 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_105_160
timestamp 1606120353
transform 1 0 15824 0 1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_106_161
timestamp 1606120353
transform 1 0 15916 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_106_165
timestamp 1606120353
transform 1 0 16284 0 -1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1606120353
transform -1 0 18860 0 1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1606120353
transform -1 0 18860 0 -1 60384
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1606120353
transform 1 0 17940 0 -1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_105_182
timestamp 1606120353
transform 1 0 17848 0 1 59296
box 0 -48 736 592
use sky130_fd_sc_hd__decap_6  FILLER_106_177
timestamp 1606120353
transform 1 0 17388 0 -1 60384
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILLER_106_184
timestamp 1606120353
transform 1 0 18032 0 -1 60384
box 0 -48 552 592
use sky130_fd_sc_hd__o21a_4  _0836_
timestamp 1606120353
transform 1 0 2116 0 1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1606120353
transform 1 0 1104 0 1 60384
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A1
timestamp 1606120353
transform 1 0 1932 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__A1
timestamp 1606120353
transform 1 0 1564 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_107_3
timestamp 1606120353
transform 1 0 1380 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_107_7
timestamp 1606120353
transform 1 0 1748 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _0835_
timestamp 1606120353
transform 1 0 4048 0 1 60384
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1606120353
transform 1 0 3956 0 1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__B
timestamp 1606120353
transform 1 0 3772 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__B
timestamp 1606120353
transform 1 0 4876 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__A
timestamp 1606120353
transform 1 0 3404 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_107_23
timestamp 1606120353
transform 1 0 3220 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_107_27
timestamp 1606120353
transform 1 0 3588 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_107_39
timestamp 1606120353
transform 1 0 4692 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_107_43
timestamp 1606120353
transform 1 0 5060 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__A
timestamp 1606120353
transform 1 0 5244 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_107_47
timestamp 1606120353
transform 1 0 5428 0 1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_107_59
timestamp 1606120353
transform 1 0 6532 0 1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__inv_8  _0556_
timestamp 1606120353
transform 1 0 7912 0 1 60384
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0555__B
timestamp 1606120353
transform 1 0 8924 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0555__A
timestamp 1606120353
transform 1 0 7728 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_107_71
timestamp 1606120353
transform 1 0 7636 0 1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_107_83
timestamp 1606120353
transform 1 0 8740 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_107_87
timestamp 1606120353
transform 1 0 9108 0 1 60384
box 0 -48 276 592
use sky130_fd_sc_hd__nand2_4  _0637_
timestamp 1606120353
transform 1 0 10304 0 1 60384
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1606120353
transform 1 0 9568 0 1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__A
timestamp 1606120353
transform 1 0 10120 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__B
timestamp 1606120353
transform 1 0 9384 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_107_93
timestamp 1606120353
transform 1 0 9660 0 1 60384
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_107_97
timestamp 1606120353
transform 1 0 10028 0 1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_107_109
timestamp 1606120353
transform 1 0 11132 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__nand3_4  _0625_
timestamp 1606120353
transform 1 0 11868 0 1 60384
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__A
timestamp 1606120353
transform 1 0 11316 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__C
timestamp 1606120353
transform 1 0 11684 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_107_113
timestamp 1606120353
transform 1 0 11500 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_107_131
timestamp 1606120353
transform 1 0 13156 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1606120353
transform 1 0 15180 0 1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__D
timestamp 1606120353
transform 1 0 14720 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__A
timestamp 1606120353
transform 1 0 13340 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__B
timestamp 1606120353
transform 1 0 13708 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_107_135
timestamp 1606120353
transform 1 0 13524 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_107_139
timestamp 1606120353
transform 1 0 13892 0 1 60384
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_107_147
timestamp 1606120353
transform 1 0 14628 0 1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_107_150
timestamp 1606120353
transform 1 0 14904 0 1 60384
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_107_154
timestamp 1606120353
transform 1 0 15272 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1199_
timestamp 1606120353
transform 1 0 16100 0 1 60384
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__D
timestamp 1606120353
transform 1 0 15916 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__CLK
timestamp 1606120353
transform 1 0 15456 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_107_158
timestamp 1606120353
transform 1 0 15640 0 1 60384
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1606120353
transform -1 0 18860 0 1 60384
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_107_182
timestamp 1606120353
transform 1 0 17848 0 1 60384
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1153_
timestamp 1606120353
transform 1 0 1472 0 -1 61472
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1606120353
transform 1 0 1104 0 -1 61472
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_108_3
timestamp 1606120353
transform 1 0 1380 0 -1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _0848_
timestamp 1606120353
transform 1 0 3956 0 -1 61472
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A2
timestamp 1606120353
transform 1 0 3404 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__B
timestamp 1606120353
transform 1 0 3772 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__CLK
timestamp 1606120353
transform 1 0 4784 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_108_23
timestamp 1606120353
transform 1 0 3220 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_108_27
timestamp 1606120353
transform 1 0 3588 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_108_38
timestamp 1606120353
transform 1 0 4600 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_108_42
timestamp 1606120353
transform 1 0 4968 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1606120353
transform 1 0 6716 0 -1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_108_54
timestamp 1606120353
transform 1 0 6072 0 -1 61472
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_108_60
timestamp 1606120353
transform 1 0 6624 0 -1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_108_62
timestamp 1606120353
transform 1 0 6808 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__nand3_4  _0555_
timestamp 1606120353
transform 1 0 8188 0 -1 61472
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  FILLER_108_74
timestamp 1606120353
transform 1 0 7912 0 -1 61472
box 0 -48 276 592
use sky130_fd_sc_hd__nand2_4  _0616_
timestamp 1606120353
transform 1 0 10488 0 -1 61472
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__A
timestamp 1606120353
transform 1 0 9660 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__C
timestamp 1606120353
transform 1 0 10028 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_108_91
timestamp 1606120353
transform 1 0 9476 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_108_95
timestamp 1606120353
transform 1 0 9844 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_108_99
timestamp 1606120353
transform 1 0 10212 0 -1 61472
box 0 -48 276 592
use sky130_fd_sc_hd__nor2_4  _0634_
timestamp 1606120353
transform 1 0 12696 0 -1 61472
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1606120353
transform 1 0 12328 0 -1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__B
timestamp 1606120353
transform 1 0 11868 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_108_111
timestamp 1606120353
transform 1 0 11316 0 -1 61472
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILLER_108_119
timestamp 1606120353
transform 1 0 12052 0 -1 61472
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_108_123
timestamp 1606120353
transform 1 0 12420 0 -1 61472
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1189_
timestamp 1606120353
transform 1 0 14720 0 -1 61472
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_12  FILLER_108_135
timestamp 1606120353
transform 1 0 13524 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_108_147
timestamp 1606120353
transform 1 0 14628 0 -1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_108_167
timestamp 1606120353
transform 1 0 16468 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1606120353
transform -1 0 18860 0 -1 61472
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1606120353
transform 1 0 17940 0 -1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_108_179
timestamp 1606120353
transform 1 0 17572 0 -1 61472
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_108_184
timestamp 1606120353
transform 1 0 18032 0 -1 61472
box 0 -48 552 592
use sky130_fd_sc_hd__o21a_4  _0832_
timestamp 1606120353
transform 1 0 1472 0 1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1606120353
transform 1 0 1104 0 1 61472
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A1
timestamp 1606120353
transform 1 0 2944 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_109_3
timestamp 1606120353
transform 1 0 1380 0 1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_109_16
timestamp 1606120353
transform 1 0 2576 0 1 61472
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_109_22
timestamp 1606120353
transform 1 0 3128 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1157_
timestamp 1606120353
transform 1 0 4048 0 1 61472
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_608
timestamp 1606120353
transform 1 0 3956 0 1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__B1
timestamp 1606120353
transform 1 0 3312 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__A2
timestamp 1606120353
transform 1 0 3680 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_109_26
timestamp 1606120353
transform 1 0 3496 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_109_30
timestamp 1606120353
transform 1 0 3864 0 1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_109_51
timestamp 1606120353
transform 1 0 5796 0 1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_109_63
timestamp 1606120353
transform 1 0 6900 0 1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0554__A
timestamp 1606120353
transform 1 0 8740 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__A
timestamp 1606120353
transform 1 0 8372 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_109_75
timestamp 1606120353
transform 1 0 8004 0 1 61472
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_109_81
timestamp 1606120353
transform 1 0 8556 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_109_85
timestamp 1606120353
transform 1 0 8924 0 1 61472
box 0 -48 368 592
use sky130_fd_sc_hd__nor3_4  _0666_
timestamp 1606120353
transform 1 0 9660 0 1 61472
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_609
timestamp 1606120353
transform 1 0 9568 0 1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__B
timestamp 1606120353
transform 1 0 9384 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__A
timestamp 1606120353
transform 1 0 11040 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_109_89
timestamp 1606120353
transform 1 0 9292 0 1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_109_106
timestamp 1606120353
transform 1 0 10856 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_109_110
timestamp 1606120353
transform 1 0 11224 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__nand3_4  _0631_
timestamp 1606120353
transform 1 0 12328 0 1 61472
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__A
timestamp 1606120353
transform 1 0 12144 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__B
timestamp 1606120353
transform 1 0 11776 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__C
timestamp 1606120353
transform 1 0 11408 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_109_114
timestamp 1606120353
transform 1 0 11592 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_109_118
timestamp 1606120353
transform 1 0 11960 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_109_140
timestamp 1606120353
transform 1 0 13984 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_109_136
timestamp 1606120353
transform 1 0 13616 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__CLK
timestamp 1606120353
transform 1 0 14168 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__D
timestamp 1606120353
transform 1 0 13800 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_109_149
timestamp 1606120353
transform 1 0 14812 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_109_144
timestamp 1606120353
transform 1 0 14352 0 1 61472
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__CLK
timestamp 1606120353
transform 1 0 14628 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__D
timestamp 1606120353
transform 1 0 14996 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_610
timestamp 1606120353
transform 1 0 15180 0 1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1190_
timestamp 1606120353
transform 1 0 15272 0 1 61472
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_12  FILLER_109_173
timestamp 1606120353
transform 1 0 17020 0 1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1606120353
transform -1 0 18860 0 1 61472
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_109_185
timestamp 1606120353
transform 1 0 18124 0 1 61472
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_109_189
timestamp 1606120353
transform 1 0 18492 0 1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _0831_
timestamp 1606120353
transform 1 0 1564 0 -1 62560
box 0 -48 644 592
use sky130_fd_sc_hd__o21a_4  _0849_
timestamp 1606120353
transform 1 0 2944 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1606120353
transform 1 0 1104 0 -1 62560
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__A
timestamp 1606120353
transform 1 0 2392 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__B1
timestamp 1606120353
transform 1 0 2760 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_110_3
timestamp 1606120353
transform 1 0 1380 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_110_12
timestamp 1606120353
transform 1 0 2208 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_110_16
timestamp 1606120353
transform 1 0 2576 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__D
timestamp 1606120353
transform 1 0 4232 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__CLK
timestamp 1606120353
transform 1 0 4600 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_110_32
timestamp 1606120353
transform 1 0 4048 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_110_36
timestamp 1606120353
transform 1 0 4416 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_110_40
timestamp 1606120353
transform 1 0 4784 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_611
timestamp 1606120353
transform 1 0 6716 0 -1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_110_52
timestamp 1606120353
transform 1 0 5888 0 -1 62560
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_110_60
timestamp 1606120353
transform 1 0 6624 0 -1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_110_62
timestamp 1606120353
transform 1 0 6808 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__buf_1  _0554_
timestamp 1606120353
transform 1 0 8740 0 -1 62560
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__B1
timestamp 1606120353
transform 1 0 9200 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_110_74
timestamp 1606120353
transform 1 0 7912 0 -1 62560
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_110_82
timestamp 1606120353
transform 1 0 8648 0 -1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_110_86
timestamp 1606120353
transform 1 0 9016 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0587_
timestamp 1606120353
transform 1 0 9752 0 -1 62560
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _0622_
timestamp 1606120353
transform 1 0 10764 0 -1 62560
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__B
timestamp 1606120353
transform 1 0 10212 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__A
timestamp 1606120353
transform 1 0 10580 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__D1
timestamp 1606120353
transform 1 0 9568 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_110_90
timestamp 1606120353
transform 1 0 9384 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_110_97
timestamp 1606120353
transform 1 0 10028 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_110_101
timestamp 1606120353
transform 1 0 10396 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0534_
timestamp 1606120353
transform 1 0 12420 0 -1 62560
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_612
timestamp 1606120353
transform 1 0 12328 0 -1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0534__A
timestamp 1606120353
transform 1 0 12880 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_110_114
timestamp 1606120353
transform 1 0 11592 0 -1 62560
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_110_126
timestamp 1606120353
transform 1 0 12696 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_110_130
timestamp 1606120353
transform 1 0 13064 0 -1 62560
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1200_
timestamp 1606120353
transform 1 0 13708 0 -1 62560
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__D
timestamp 1606120353
transform 1 0 13524 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_110_134
timestamp 1606120353
transform 1 0 13432 0 -1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__A
timestamp 1606120353
transform 1 0 16008 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_110_156
timestamp 1606120353
transform 1 0 15456 0 -1 62560
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_110_164
timestamp 1606120353
transform 1 0 16192 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_110_176
timestamp 1606120353
transform 1 0 17296 0 -1 62560
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1606120353
transform -1 0 18860 0 -1 62560
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_613
timestamp 1606120353
transform 1 0 17940 0 -1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_110_182
timestamp 1606120353
transform 1 0 17848 0 -1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_110_184
timestamp 1606120353
transform 1 0 18032 0 -1 62560
box 0 -48 552 592
use sky130_fd_sc_hd__o21a_4  _0840_
timestamp 1606120353
transform 1 0 1472 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1606120353
transform 1 0 1104 0 1 62560
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A1
timestamp 1606120353
transform 1 0 2760 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__B1
timestamp 1606120353
transform 1 0 3128 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_111_3
timestamp 1606120353
transform 1 0 1380 0 1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_111_16
timestamp 1606120353
transform 1 0 2576 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_111_20
timestamp 1606120353
transform 1 0 2944 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _0844_
timestamp 1606120353
transform 1 0 4048 0 1 62560
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_614
timestamp 1606120353
transform 1 0 3956 0 1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__A
timestamp 1606120353
transform 1 0 4876 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__D
timestamp 1606120353
transform 1 0 3772 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_111_24
timestamp 1606120353
transform 1 0 3312 0 1 62560
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_111_28
timestamp 1606120353
transform 1 0 3680 0 1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_111_39
timestamp 1606120353
transform 1 0 4692 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_111_43
timestamp 1606120353
transform 1 0 5060 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0778_
timestamp 1606120353
transform 1 0 6256 0 1 62560
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A
timestamp 1606120353
transform 1 0 6072 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__CLK
timestamp 1606120353
transform 1 0 5244 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_111_47
timestamp 1606120353
transform 1 0 5428 0 1 62560
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_111_53
timestamp 1606120353
transform 1 0 5980 0 1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_111_65
timestamp 1606120353
transform 1 0 7084 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_111_69
timestamp 1606120353
transform 1 0 7452 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__B2
timestamp 1606120353
transform 1 0 7268 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0662__A
timestamp 1606120353
transform 1 0 7636 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_111_73
timestamp 1606120353
transform 1 0 7820 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__C1
timestamp 1606120353
transform 1 0 8004 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_111_77
timestamp 1606120353
transform 1 0 8188 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A1
timestamp 1606120353
transform 1 0 8372 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0520_
timestamp 1606120353
transform 1 0 8556 0 1 62560
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_111_84
timestamp 1606120353
transform 1 0 8832 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0520__A
timestamp 1606120353
transform 1 0 9016 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_111_88
timestamp 1606120353
transform 1 0 9200 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__nand3_4  _0667_
timestamp 1606120353
transform 1 0 9844 0 1 62560
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_615
timestamp 1606120353
transform 1 0 9568 0 1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A2
timestamp 1606120353
transform 1 0 9384 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_111_93
timestamp 1606120353
transform 1 0 9660 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_111_109
timestamp 1606120353
transform 1 0 11132 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1191_
timestamp 1606120353
transform 1 0 12696 0 1 62560
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__D
timestamp 1606120353
transform 1 0 12512 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0519__A
timestamp 1606120353
transform 1 0 12144 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__C
timestamp 1606120353
transform 1 0 11316 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_111_113
timestamp 1606120353
transform 1 0 11500 0 1 62560
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_111_119
timestamp 1606120353
transform 1 0 12052 0 1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_111_122
timestamp 1606120353
transform 1 0 12328 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_616
timestamp 1606120353
transform 1 0 15180 0 1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__D
timestamp 1606120353
transform 1 0 14996 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__CLK
timestamp 1606120353
transform 1 0 14628 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_111_145
timestamp 1606120353
transform 1 0 14444 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_111_149
timestamp 1606120353
transform 1 0 14812 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_111_154
timestamp 1606120353
transform 1 0 15272 0 1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1225_
timestamp 1606120353
transform 1 0 15364 0 1 62560
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_12  FILLER_111_174
timestamp 1606120353
transform 1 0 17112 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1606120353
transform -1 0 18860 0 1 62560
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_111_186
timestamp 1606120353
transform 1 0 18216 0 1 62560
box 0 -48 368 592
use sky130_fd_sc_hd__o21a_4  _0845_
timestamp 1606120353
transform 1 0 2116 0 1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1155_
timestamp 1606120353
transform 1 0 1472 0 -1 63648
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1606120353
transform 1 0 1104 0 -1 63648
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1606120353
transform 1 0 1104 0 1 63648
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A1
timestamp 1606120353
transform 1 0 1932 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A2
timestamp 1606120353
transform 1 0 1564 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_112_3
timestamp 1606120353
transform 1 0 1380 0 -1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_113_3
timestamp 1606120353
transform 1 0 1380 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_113_7
timestamp 1606120353
transform 1 0 1748 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__D
timestamp 1606120353
transform 1 0 3404 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__CLK
timestamp 1606120353
transform 1 0 3404 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_112_23
timestamp 1606120353
transform 1 0 3220 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_113_23
timestamp 1606120353
transform 1 0 3220 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__D
timestamp 1606120353
transform 1 0 3772 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_112_27
timestamp 1606120353
transform 1 0 3588 0 -1 63648
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_113_27
timestamp 1606120353
transform 1 0 3588 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_620
timestamp 1606120353
transform 1 0 3956 0 1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__B
timestamp 1606120353
transform 1 0 4048 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_112_31
timestamp 1606120353
transform 1 0 3956 0 -1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_113_32
timestamp 1606120353
transform 1 0 4048 0 1 63648
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_113_38
timestamp 1606120353
transform 1 0 4600 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__A
timestamp 1606120353
transform 1 0 4416 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A
timestamp 1606120353
transform 1 0 4784 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0887_
timestamp 1606120353
transform 1 0 4968 0 1 63648
box 0 -48 828 592
use sky130_fd_sc_hd__dfxtp_4  _1171_
timestamp 1606120353
transform 1 0 4232 0 -1 63648
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_1  FILLER_113_55
timestamp 1606120353
transform 1 0 6164 0 1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_113_51
timestamp 1606120353
transform 1 0 5796 0 1 63648
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_112_53
timestamp 1606120353
transform 1 0 5980 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A4
timestamp 1606120353
transform 1 0 6164 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_113_58
timestamp 1606120353
transform 1 0 6440 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_112_57
timestamp 1606120353
transform 1 0 6348 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A2
timestamp 1606120353
transform 1 0 6532 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__A1_N
timestamp 1606120353
transform 1 0 6256 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A3
timestamp 1606120353
transform 1 0 6624 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_617
timestamp 1606120353
transform 1 0 6716 0 -1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _0662_
timestamp 1606120353
transform 1 0 6808 0 -1 63648
box 0 -48 828 592
use sky130_fd_sc_hd__o41ai_4  _0788_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 6808 0 1 63648
box 0 -48 2024 592
use sky130_fd_sc_hd__a2111oi_4  _0673_
timestamp 1606120353
transform 1 0 8924 0 -1 63648
box 0 -48 2024 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__A1
timestamp 1606120353
transform 1 0 9016 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__A2_N
timestamp 1606120353
transform 1 0 7820 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__B1
timestamp 1606120353
transform 1 0 8188 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_112_71
timestamp 1606120353
transform 1 0 7636 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_112_75
timestamp 1606120353
transform 1 0 8004 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_112_79
timestamp 1606120353
transform 1 0 8372 0 -1 63648
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_113_84
timestamp 1606120353
transform 1 0 8832 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_113_88
timestamp 1606120353
transform 1 0 9200 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__a21oi_4  _0669_
timestamp 1606120353
transform 1 0 9660 0 1 63648
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_621
timestamp 1606120353
transform 1 0 9568 0 1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__B
timestamp 1606120353
transform 1 0 9384 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__C
timestamp 1606120353
transform 1 0 11040 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A
timestamp 1606120353
transform 1 0 11132 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_112_107
timestamp 1606120353
transform 1 0 10948 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_113_106
timestamp 1606120353
transform 1 0 10856 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_113_110
timestamp 1606120353
transform 1 0 11224 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_112_116
timestamp 1606120353
transform 1 0 11776 0 -1 63648
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILLER_112_111
timestamp 1606120353
transform 1 0 11316 0 -1 63648
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__B
timestamp 1606120353
transform 1 0 11592 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__A
timestamp 1606120353
transform 1 0 11408 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_113_131
timestamp 1606120353
transform 1 0 13156 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_113_127
timestamp 1606120353
transform 1 0 12788 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_112_130
timestamp 1606120353
transform 1 0 13064 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_112_126
timestamp 1606120353
transform 1 0 12696 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__CLK
timestamp 1606120353
transform 1 0 13248 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__CLK
timestamp 1606120353
transform 1 0 12880 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__D
timestamp 1606120353
transform 1 0 12972 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_618
timestamp 1606120353
transform 1 0 12328 0 -1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0519_
timestamp 1606120353
transform 1 0 12420 0 -1 63648
box 0 -48 276 592
use sky130_fd_sc_hd__nor3_4  _0617_
timestamp 1606120353
transform 1 0 11592 0 1 63648
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_1  FILLER_112_134
timestamp 1606120353
transform 1 0 13432 0 -1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__A
timestamp 1606120353
transform 1 0 13340 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0599_
timestamp 1606120353
transform 1 0 13524 0 1 63648
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_113_154
timestamp 1606120353
transform 1 0 15272 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_113_148
timestamp 1606120353
transform 1 0 14720 0 1 63648
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_113_144
timestamp 1606120353
transform 1 0 14352 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_112_154
timestamp 1606120353
transform 1 0 15272 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__CLK
timestamp 1606120353
transform 1 0 14996 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__B
timestamp 1606120353
transform 1 0 14536 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_622
timestamp 1606120353
transform 1 0 15180 0 1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1202_
timestamp 1606120353
transform 1 0 13524 0 -1 63648
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  FILLER_113_158
timestamp 1606120353
transform 1 0 15640 0 1 63648
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_112_165
timestamp 1606120353
transform 1 0 16284 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_112_158
timestamp 1606120353
transform 1 0 15640 0 -1 63648
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__CLK
timestamp 1606120353
transform 1 0 15456 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__D
timestamp 1606120353
transform 1 0 15916 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__D
timestamp 1606120353
transform 1 0 15456 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0574_
timestamp 1606120353
transform 1 0 16008 0 -1 63648
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__CLK
timestamp 1606120353
transform 1 0 16468 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_112_169
timestamp 1606120353
transform 1 0 16652 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1203_
timestamp 1606120353
transform 1 0 16100 0 1 63648
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1606120353
transform -1 0 18860 0 -1 63648
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1606120353
transform -1 0 18860 0 1 63648
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_619
timestamp 1606120353
transform 1 0 17940 0 -1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_112_181
timestamp 1606120353
transform 1 0 17756 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_112_184
timestamp 1606120353
transform 1 0 18032 0 -1 63648
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_113_182
timestamp 1606120353
transform 1 0 17848 0 1 63648
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1156_
timestamp 1606120353
transform 1 0 2760 0 -1 64736
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1606120353
transform 1 0 1104 0 -1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__B1
timestamp 1606120353
transform 1 0 2116 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A2
timestamp 1606120353
transform 1 0 2484 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__D
timestamp 1606120353
transform 1 0 1564 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_114_3
timestamp 1606120353
transform 1 0 1380 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_114_7
timestamp 1606120353
transform 1 0 1748 0 -1 64736
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_114_13
timestamp 1606120353
transform 1 0 2300 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_114_17
timestamp 1606120353
transform 1 0 2668 0 -1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__B
timestamp 1606120353
transform 1 0 4968 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_114_37
timestamp 1606120353
transform 1 0 4508 0 -1 64736
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_114_41
timestamp 1606120353
transform 1 0 4876 0 -1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_114_44
timestamp 1606120353
transform 1 0 5152 0 -1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_114_52
timestamp 1606120353
transform 1 0 5888 0 -1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_114_48
timestamp 1606120353
transform 1 0 5520 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__D
timestamp 1606120353
transform 1 0 5704 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__B1
timestamp 1606120353
transform 1 0 6164 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0863_
timestamp 1606120353
transform 1 0 5244 0 -1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_114_62
timestamp 1606120353
transform 1 0 6808 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_114_57
timestamp 1606120353
transform 1 0 6348 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A2
timestamp 1606120353
transform 1 0 6532 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A1
timestamp 1606120353
transform 1 0 6992 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_623
timestamp 1606120353
transform 1 0 6716 0 -1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__a2bb2oi_4  _0787_
timestamp 1606120353
transform 1 0 7176 0 -1 64736
box 0 -48 1932 592
use sky130_fd_sc_hd__fill_2  FILLER_114_87
timestamp 1606120353
transform 1 0 9108 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__nor3_4  _0672_
timestamp 1606120353
transform 1 0 9844 0 -1 64736
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__B
timestamp 1606120353
transform 1 0 11224 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__B1
timestamp 1606120353
transform 1 0 9660 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__A2
timestamp 1606120353
transform 1 0 9292 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_114_91
timestamp 1606120353
transform 1 0 9476 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_114_108
timestamp 1606120353
transform 1 0 11040 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1204_
timestamp 1606120353
transform 1 0 12972 0 -1 64736
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_624
timestamp 1606120353
transform 1 0 12328 0 -1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__D
timestamp 1606120353
transform 1 0 11592 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_114_112
timestamp 1606120353
transform 1 0 11408 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_114_116
timestamp 1606120353
transform 1 0 11776 0 -1 64736
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILLER_114_123
timestamp 1606120353
transform 1 0 12420 0 -1 64736
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_114_148
timestamp 1606120353
transform 1 0 14720 0 -1 64736
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1197_
timestamp 1606120353
transform 1 0 15456 0 -1 64736
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_8  FILLER_114_175
timestamp 1606120353
transform 1 0 17204 0 -1 64736
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1606120353
transform -1 0 18860 0 -1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_625
timestamp 1606120353
transform 1 0 17940 0 -1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_114_184
timestamp 1606120353
transform 1 0 18032 0 -1 64736
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _0839_
timestamp 1606120353
transform 1 0 2208 0 1 64736
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1606120353
transform 1 0 1104 0 1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A
timestamp 1606120353
transform 1 0 3128 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__A
timestamp 1606120353
transform 1 0 2024 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__CLK
timestamp 1606120353
transform 1 0 1656 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_115_3
timestamp 1606120353
transform 1 0 1380 0 1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_115_8
timestamp 1606120353
transform 1 0 1840 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_115_19
timestamp 1606120353
transform 1 0 2852 0 1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__nor2_4  _0895_
timestamp 1606120353
transform 1 0 4048 0 1 64736
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_626
timestamp 1606120353
transform 1 0 3956 0 1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__B
timestamp 1606120353
transform 1 0 3772 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__B
timestamp 1606120353
transform 1 0 5152 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_115_24
timestamp 1606120353
transform 1 0 3312 0 1 64736
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_115_28
timestamp 1606120353
transform 1 0 3680 0 1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_115_41
timestamp 1606120353
transform 1 0 4876 0 1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1164_
timestamp 1606120353
transform 1 0 5612 0 1 64736
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  FILLER_115_46
timestamp 1606120353
transform 1 0 5336 0 1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_115_68
timestamp 1606120353
transform 1 0 7360 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_115_72
timestamp 1606120353
transform 1 0 7728 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A3
timestamp 1606120353
transform 1 0 7544 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A4
timestamp 1606120353
transform 1 0 7912 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_115_76
timestamp 1606120353
transform 1 0 8096 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A1
timestamp 1606120353
transform 1 0 8280 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_115_80
timestamp 1606120353
transform 1 0 8464 0 1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0682_
timestamp 1606120353
transform 1 0 8556 0 1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_115_84
timestamp 1606120353
transform 1 0 8832 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__A
timestamp 1606120353
transform 1 0 9016 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_115_88
timestamp 1606120353
transform 1 0 9200 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0573_
timestamp 1606120353
transform 1 0 10120 0 1 64736
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_627
timestamp 1606120353
transform 1 0 9568 0 1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__B
timestamp 1606120353
transform 1 0 9936 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__C
timestamp 1606120353
transform 1 0 11132 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__C
timestamp 1606120353
transform 1 0 9384 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_115_93
timestamp 1606120353
transform 1 0 9660 0 1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_115_107
timestamp 1606120353
transform 1 0 10948 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0542_
timestamp 1606120353
transform 1 0 11684 0 1 64736
box 0 -48 828 592
use sky130_fd_sc_hd__buf_1  _0543_
timestamp 1606120353
transform 1 0 13248 0 1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__A
timestamp 1606120353
transform 1 0 11500 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__CLK
timestamp 1606120353
transform 1 0 13064 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_115_111
timestamp 1606120353
transform 1 0 11316 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_115_124
timestamp 1606120353
transform 1 0 12512 0 1 64736
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_628
timestamp 1606120353
transform 1 0 15180 0 1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__D
timestamp 1606120353
transform 1 0 13708 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0543__A
timestamp 1606120353
transform 1 0 14076 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_115_135
timestamp 1606120353
transform 1 0 13524 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_115_139
timestamp 1606120353
transform 1 0 13892 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_115_143
timestamp 1606120353
transform 1 0 14260 0 1 64736
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_115_151
timestamp 1606120353
transform 1 0 14996 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_115_154
timestamp 1606120353
transform 1 0 15272 0 1 64736
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1206_
timestamp 1606120353
transform 1 0 16100 0 1 64736
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__D
timestamp 1606120353
transform 1 0 15916 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_115_160
timestamp 1606120353
transform 1 0 15824 0 1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1606120353
transform -1 0 18860 0 1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_115_182
timestamp 1606120353
transform 1 0 17848 0 1 64736
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _0856_
timestamp 1606120353
transform 1 0 3128 0 -1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1606120353
transform 1 0 1104 0 -1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__B
timestamp 1606120353
transform 1 0 2208 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__B
timestamp 1606120353
transform 1 0 2576 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__CLK
timestamp 1606120353
transform 1 0 2944 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_116_3
timestamp 1606120353
transform 1 0 1380 0 -1 65824
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_116_11
timestamp 1606120353
transform 1 0 2116 0 -1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_116_14
timestamp 1606120353
transform 1 0 2392 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_116_18
timestamp 1606120353
transform 1 0 2760 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1175_
timestamp 1606120353
transform 1 0 4140 0 -1 65824
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__B1
timestamp 1606120353
transform 1 0 3956 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__A
timestamp 1606120353
transform 1 0 3588 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_116_25
timestamp 1606120353
transform 1 0 3404 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_116_29
timestamp 1606120353
transform 1 0 3772 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_629
timestamp 1606120353
transform 1 0 6716 0 -1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__A2_N
timestamp 1606120353
transform 1 0 6992 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__B1
timestamp 1606120353
transform 1 0 6532 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__CLK
timestamp 1606120353
transform 1 0 6072 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_116_52
timestamp 1606120353
transform 1 0 5888 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_116_56
timestamp 1606120353
transform 1 0 6256 0 -1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_116_62
timestamp 1606120353
transform 1 0 6808 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_116_66
timestamp 1606120353
transform 1 0 7176 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__o41ai_4  _0767_
timestamp 1606120353
transform 1 0 7360 0 -1 65824
box 0 -48 2024 592
use sky130_fd_sc_hd__and4_4  _0603_
timestamp 1606120353
transform 1 0 10764 0 -1 65824
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__A
timestamp 1606120353
transform 1 0 10120 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A
timestamp 1606120353
transform 1 0 9568 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_116_90
timestamp 1606120353
transform 1 0 9384 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_116_94
timestamp 1606120353
transform 1 0 9752 0 -1 65824
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_116_100
timestamp 1606120353
transform 1 0 10304 0 -1 65824
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_116_104
timestamp 1606120353
transform 1 0 10672 0 -1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_630
timestamp 1606120353
transform 1 0 12328 0 -1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__A
timestamp 1606120353
transform 1 0 12604 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__B
timestamp 1606120353
transform 1 0 12972 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__A
timestamp 1606120353
transform 1 0 11776 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_116_114
timestamp 1606120353
transform 1 0 11592 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_116_118
timestamp 1606120353
transform 1 0 11960 0 -1 65824
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_116_123
timestamp 1606120353
transform 1 0 12420 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_116_127
timestamp 1606120353
transform 1 0 12788 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_116_131
timestamp 1606120353
transform 1 0 13156 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1205_
timestamp 1606120353
transform 1 0 13340 0 -1 65824
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__CLK
timestamp 1606120353
transform 1 0 15272 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_116_152
timestamp 1606120353
transform 1 0 15088 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__CLK
timestamp 1606120353
transform 1 0 16100 0 -1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_116_156
timestamp 1606120353
transform 1 0 15456 0 -1 65824
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_116_162
timestamp 1606120353
transform 1 0 16008 0 -1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_116_165
timestamp 1606120353
transform 1 0 16284 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1606120353
transform -1 0 18860 0 -1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_631
timestamp 1606120353
transform 1 0 17940 0 -1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_116_177
timestamp 1606120353
transform 1 0 17388 0 -1 65824
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILLER_116_184
timestamp 1606120353
transform 1 0 18032 0 -1 65824
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_117_3
timestamp 1606120353
transform 1 0 1380 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1606120353
transform 1 0 1104 0 1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0702_
timestamp 1606120353
transform 1 0 1564 0 1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_117_8
timestamp 1606120353
transform 1 0 1840 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_117_12
timestamp 1606120353
transform 1 0 2208 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A
timestamp 1606120353
transform 1 0 2024 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A
timestamp 1606120353
transform 1 0 2392 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_117_16
timestamp 1606120353
transform 1 0 2576 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A
timestamp 1606120353
transform 1 0 2760 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0843_
timestamp 1606120353
transform 1 0 2944 0 1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__a21oi_4  _0888_
timestamp 1606120353
transform 1 0 4876 0 1 65824
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_632
timestamp 1606120353
transform 1 0 3956 0 1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__A1
timestamp 1606120353
transform 1 0 4692 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A
timestamp 1606120353
transform 1 0 3588 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A
timestamp 1606120353
transform 1 0 4324 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_117_23
timestamp 1606120353
transform 1 0 3220 0 1 65824
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_117_29
timestamp 1606120353
transform 1 0 3772 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_117_32
timestamp 1606120353
transform 1 0 4048 0 1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_117_37
timestamp 1606120353
transform 1 0 4508 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__a2bb2oi_4  _0766_
timestamp 1606120353
transform 1 0 6900 0 1 65824
box 0 -48 1932 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__A
timestamp 1606120353
transform 1 0 6716 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__A1_N
timestamp 1606120353
transform 1 0 6348 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_117_54
timestamp 1606120353
transform 1 0 6072 0 1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_117_59
timestamp 1606120353
transform 1 0 6532 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0538__A
timestamp 1606120353
transform 1 0 9016 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_117_84
timestamp 1606120353
transform 1 0 8832 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_117_88
timestamp 1606120353
transform 1 0 9200 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__B
timestamp 1606120353
transform 1 0 9384 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_633
timestamp 1606120353
transform 1 0 9568 0 1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_117_93
timestamp 1606120353
transform 1 0 9660 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__C
timestamp 1606120353
transform 1 0 9844 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_117_97
timestamp 1606120353
transform 1 0 10028 0 1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0594_
timestamp 1606120353
transform 1 0 10120 0 1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_117_101
timestamp 1606120353
transform 1 0 10396 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__A
timestamp 1606120353
transform 1 0 10580 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_117_105
timestamp 1606120353
transform 1 0 10764 0 1 65824
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__A
timestamp 1606120353
transform 1 0 11132 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0605_
timestamp 1606120353
transform 1 0 11316 0 1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__nand2_4  _0629_
timestamp 1606120353
transform 1 0 12604 0 1 65824
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__B
timestamp 1606120353
transform 1 0 12420 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__A
timestamp 1606120353
transform 1 0 12052 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_117_114
timestamp 1606120353
transform 1 0 11592 0 1 65824
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_117_118
timestamp 1606120353
transform 1 0 11960 0 1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_117_121
timestamp 1606120353
transform 1 0 12236 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_117_142
timestamp 1606120353
transform 1 0 14168 0 1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_117_138
timestamp 1606120353
transform 1 0 13800 0 1 65824
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_117_134
timestamp 1606120353
transform 1 0 13432 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__CLK
timestamp 1606120353
transform 1 0 14260 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__C
timestamp 1606120353
transform 1 0 13616 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_117_149
timestamp 1606120353
transform 1 0 14812 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_117_145
timestamp 1606120353
transform 1 0 14444 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__D
timestamp 1606120353
transform 1 0 14628 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__D
timestamp 1606120353
transform 1 0 14996 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_634
timestamp 1606120353
transform 1 0 15180 0 1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1196_
timestamp 1606120353
transform 1 0 15272 0 1 65824
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_12  FILLER_117_173
timestamp 1606120353
transform 1 0 17020 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1606120353
transform -1 0 18860 0 1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_117_185
timestamp 1606120353
transform 1 0 18124 0 1 65824
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_117_189
timestamp 1606120353
transform 1 0 18492 0 1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_119_3
timestamp 1606120353
transform 1 0 1380 0 1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_118_7
timestamp 1606120353
transform 1 0 1748 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_118_3
timestamp 1606120353
transform 1 0 1380 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__B1
timestamp 1606120353
transform 1 0 1932 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A
timestamp 1606120353
transform 1 0 1564 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1606120353
transform 1 0 1104 0 1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1606120353
transform 1 0 1104 0 -1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _0773_
timestamp 1606120353
transform 1 0 1472 0 1 66912
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_119_17
timestamp 1606120353
transform 1 0 2668 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_119_13
timestamp 1606120353
transform 1 0 2300 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_118_11
timestamp 1606120353
transform 1 0 2116 0 -1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A1
timestamp 1606120353
transform 1 0 2484 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _0852_
timestamp 1606120353
transform 1 0 2208 0 -1 66912
box 0 -48 644 592
use sky130_fd_sc_hd__decap_6  FILLER_119_21
timestamp 1606120353
transform 1 0 3036 0 1 66912
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_118_19
timestamp 1606120353
transform 1 0 2852 0 -1 66912
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A2
timestamp 1606120353
transform 1 0 2852 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_119_29
timestamp 1606120353
transform 1 0 3772 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_118_30
timestamp 1606120353
transform 1 0 3864 0 -1 66912
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__A
timestamp 1606120353
transform 1 0 3588 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_638
timestamp 1606120353
transform 1 0 3956 0 1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0774_
timestamp 1606120353
transform 1 0 3588 0 -1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_119_37
timestamp 1606120353
transform 1 0 4508 0 1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_119_32
timestamp 1606120353
transform 1 0 4048 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_118_40
timestamp 1606120353
transform 1 0 4784 0 -1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_118_36
timestamp 1606120353
transform 1 0 4416 0 -1 66912
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__A
timestamp 1606120353
transform 1 0 4232 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A1
timestamp 1606120353
transform 1 0 4784 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0775_
timestamp 1606120353
transform 1 0 4232 0 1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_119_42
timestamp 1606120353
transform 1 0 4968 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_118_43
timestamp 1606120353
transform 1 0 5060 0 -1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__A2
timestamp 1606120353
transform 1 0 4876 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A2
timestamp 1606120353
transform 1 0 5152 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__nand2_4  _0872_
timestamp 1606120353
transform 1 0 5152 0 -1 66912
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_118_53
timestamp 1606120353
transform 1 0 5980 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__B1
timestamp 1606120353
transform 1 0 6164 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A1
timestamp 1606120353
transform 1 0 6624 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__B1
timestamp 1606120353
transform 1 0 6532 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_118_57
timestamp 1606120353
transform 1 0 6348 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_119_58
timestamp 1606120353
transform 1 0 6440 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_635
timestamp 1606120353
transform 1 0 6716 0 -1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A
timestamp 1606120353
transform 1 0 6992 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__B2
timestamp 1606120353
transform 1 0 6992 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_118_62
timestamp 1606120353
transform 1 0 6808 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_118_66
timestamp 1606120353
transform 1 0 7176 0 -1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_119_62
timestamp 1606120353
transform 1 0 6808 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__nand2_4  _0879_
timestamp 1606120353
transform 1 0 7176 0 1 66912
box 0 -48 828 592
use sky130_fd_sc_hd__o21a_4  _0873_
timestamp 1606120353
transform 1 0 5336 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_118_72
timestamp 1606120353
transform 1 0 7728 0 -1 66912
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _0558_
timestamp 1606120353
transform 1 0 7452 0 -1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_119_79
timestamp 1606120353
transform 1 0 8372 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_119_75
timestamp 1606120353
transform 1 0 8004 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__A
timestamp 1606120353
transform 1 0 8556 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__B
timestamp 1606120353
transform 1 0 8188 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0538_
timestamp 1606120353
transform 1 0 8464 0 -1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_119_88
timestamp 1606120353
transform 1 0 9200 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_119_83
timestamp 1606120353
transform 1 0 8740 0 1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_118_83
timestamp 1606120353
transform 1 0 8740 0 -1 66912
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0535__A
timestamp 1606120353
transform 1 0 9016 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__C
timestamp 1606120353
transform 1 0 9292 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__B
timestamp 1606120353
transform 1 0 9384 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_639
timestamp 1606120353
transform 1 0 9568 0 1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_119_107
timestamp 1606120353
transform 1 0 10948 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_118_109
timestamp 1606120353
transform 1 0 11132 0 -1 66912
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_118_105
timestamp 1606120353
transform 1 0 10764 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__C
timestamp 1606120353
transform 1 0 10948 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__A
timestamp 1606120353
transform 1 0 11132 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__nand3_4  _0671_
timestamp 1606120353
transform 1 0 9476 0 -1 66912
box 0 -48 1288 592
use sky130_fd_sc_hd__nand3_4  _0668_
timestamp 1606120353
transform 1 0 9660 0 1 66912
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  FILLER_119_115
timestamp 1606120353
transform 1 0 11684 0 1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_119_111
timestamp 1606120353
transform 1 0 11316 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_118_118
timestamp 1606120353
transform 1 0 11960 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_118_115
timestamp 1606120353
transform 1 0 11684 0 -1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0627__C
timestamp 1606120353
transform 1 0 11776 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__B
timestamp 1606120353
transform 1 0 11500 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0627__A
timestamp 1606120353
transform 1 0 12144 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0627__B
timestamp 1606120353
transform 1 0 11960 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_636
timestamp 1606120353
transform 1 0 12328 0 -1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__nand3_4  _0628_
timestamp 1606120353
transform 1 0 12420 0 -1 66912
box 0 -48 1288 592
use sky130_fd_sc_hd__nand3_4  _0627_
timestamp 1606120353
transform 1 0 12144 0 1 66912
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_119_138
timestamp 1606120353
transform 1 0 13800 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_119_134
timestamp 1606120353
transform 1 0 13432 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__B
timestamp 1606120353
transform 1 0 13984 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__A
timestamp 1606120353
transform 1 0 13616 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0557_
timestamp 1606120353
transform 1 0 14168 0 1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_119_154
timestamp 1606120353
transform 1 0 15272 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_119_149
timestamp 1606120353
transform 1 0 14812 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_119_145
timestamp 1606120353
transform 1 0 14444 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_118_149
timestamp 1606120353
transform 1 0 14812 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__CLK
timestamp 1606120353
transform 1 0 14996 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0557__A
timestamp 1606120353
transform 1 0 14628 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_640
timestamp 1606120353
transform 1 0 15180 0 1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_118_137
timestamp 1606120353
transform 1 0 13708 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1226_
timestamp 1606120353
transform 1 0 14996 0 -1 66912
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1207_
timestamp 1606120353
transform 1 0 16100 0 1 66912
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__D
timestamp 1606120353
transform 1 0 15916 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__D
timestamp 1606120353
transform 1 0 15456 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__CLK
timestamp 1606120353
transform 1 0 16928 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_118_170
timestamp 1606120353
transform 1 0 16744 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_118_174
timestamp 1606120353
transform 1 0 17112 0 -1 66912
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_119_158
timestamp 1606120353
transform 1 0 15640 0 1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1606120353
transform -1 0 18860 0 -1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1606120353
transform -1 0 18860 0 1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_637
timestamp 1606120353
transform 1 0 17940 0 -1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_118_182
timestamp 1606120353
transform 1 0 17848 0 -1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_118_184
timestamp 1606120353
transform 1 0 18032 0 -1 66912
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_119_182
timestamp 1606120353
transform 1 0 17848 0 1 66912
box 0 -48 736 592
use sky130_fd_sc_hd__o21a_4  _0853_
timestamp 1606120353
transform 1 0 1748 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1606120353
transform 1 0 1104 0 -1 68000
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__B1
timestamp 1606120353
transform 1 0 1564 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__CLK
timestamp 1606120353
transform 1 0 3036 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_120_3
timestamp 1606120353
transform 1 0 1380 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_120_19
timestamp 1606120353
transform 1 0 2852 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0793_
timestamp 1606120353
transform 1 0 3588 0 -1 68000
box 0 -48 276 592
use sky130_fd_sc_hd__a21oi_4  _0896_
timestamp 1606120353
transform 1 0 4784 0 -1 68000
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__B1
timestamp 1606120353
transform 1 0 4600 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__B1
timestamp 1606120353
transform 1 0 4048 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A2
timestamp 1606120353
transform 1 0 3404 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_120_23
timestamp 1606120353
transform 1 0 3220 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_120_30
timestamp 1606120353
transform 1 0 3864 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_120_34
timestamp 1606120353
transform 1 0 4232 0 -1 68000
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _0589_
timestamp 1606120353
transform 1 0 6808 0 -1 68000
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_641
timestamp 1606120353
transform 1 0 6716 0 -1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A2
timestamp 1606120353
transform 1 0 6164 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_120_53
timestamp 1606120353
transform 1 0 5980 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_120_57
timestamp 1606120353
transform 1 0 6348 0 -1 68000
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__A1
timestamp 1606120353
transform 1 0 7820 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__B1
timestamp 1606120353
transform 1 0 8188 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_120_71
timestamp 1606120353
transform 1 0 7636 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_120_75
timestamp 1606120353
transform 1 0 8004 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_120_79
timestamp 1606120353
transform 1 0 8372 0 -1 68000
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_120_87
timestamp 1606120353
transform 1 0 9108 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0535_
timestamp 1606120353
transform 1 0 9292 0 -1 68000
box 0 -48 276 592
use sky130_fd_sc_hd__nand3_4  _0632_
timestamp 1606120353
transform 1 0 10304 0 -1 68000
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A
timestamp 1606120353
transform 1 0 9752 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__D
timestamp 1606120353
transform 1 0 10120 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_120_92
timestamp 1606120353
transform 1 0 9568 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_120_96
timestamp 1606120353
transform 1 0 9936 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__nand3_4  _0633_
timestamp 1606120353
transform 1 0 12420 0 -1 68000
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_642
timestamp 1606120353
transform 1 0 12328 0 -1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__C
timestamp 1606120353
transform 1 0 12144 0 -1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_120_114
timestamp 1606120353
transform 1 0 11592 0 -1 68000
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_120_137
timestamp 1606120353
transform 1 0 13708 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_120_149
timestamp 1606120353
transform 1 0 14812 0 -1 68000
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1227_
timestamp 1606120353
transform 1 0 15456 0 -1 68000
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_1  FILLER_120_155
timestamp 1606120353
transform 1 0 15364 0 -1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_120_175
timestamp 1606120353
transform 1 0 17204 0 -1 68000
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1606120353
transform -1 0 18860 0 -1 68000
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_643
timestamp 1606120353
transform 1 0 17940 0 -1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_120_184
timestamp 1606120353
transform 1 0 18032 0 -1 68000
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1158_
timestamp 1606120353
transform 1 0 1472 0 1 68000
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1606120353
transform 1 0 1104 0 1 68000
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_121_3
timestamp 1606120353
transform 1 0 1380 0 1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1176_
timestamp 1606120353
transform 1 0 4048 0 1 68000
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_644
timestamp 1606120353
transform 1 0 3956 0 1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__A1
timestamp 1606120353
transform 1 0 3404 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A1
timestamp 1606120353
transform 1 0 3772 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_121_23
timestamp 1606120353
transform 1 0 3220 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_121_27
timestamp 1606120353
transform 1 0 3588 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0870_
timestamp 1606120353
transform 1 0 6532 0 1 68000
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__B2
timestamp 1606120353
transform 1 0 6992 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A
timestamp 1606120353
transform 1 0 5980 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A
timestamp 1606120353
transform 1 0 6348 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_121_51
timestamp 1606120353
transform 1 0 5796 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_121_55
timestamp 1606120353
transform 1 0 6164 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_121_62
timestamp 1606120353
transform 1 0 6808 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_121_66
timestamp 1606120353
transform 1 0 7176 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0663_
timestamp 1606120353
transform 1 0 7544 0 1 68000
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__B
timestamp 1606120353
transform 1 0 9016 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__A
timestamp 1606120353
transform 1 0 8648 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__A2
timestamp 1606120353
transform 1 0 7360 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_121_79
timestamp 1606120353
transform 1 0 8372 0 1 68000
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_121_84
timestamp 1606120353
transform 1 0 8832 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_121_88
timestamp 1606120353
transform 1 0 9200 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0524_
timestamp 1606120353
transform 1 0 9752 0 1 68000
box 0 -48 276 592
use sky130_fd_sc_hd__nand3_4  _0606_
timestamp 1606120353
transform 1 0 10764 0 1 68000
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_645
timestamp 1606120353
transform 1 0 9568 0 1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__C
timestamp 1606120353
transform 1 0 9384 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__A
timestamp 1606120353
transform 1 0 10212 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0606__A
timestamp 1606120353
transform 1 0 10580 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_121_93
timestamp 1606120353
transform 1 0 9660 0 1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_121_97
timestamp 1606120353
transform 1 0 10028 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_121_101
timestamp 1606120353
transform 1 0 10396 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__nand2_4  _0630_
timestamp 1606120353
transform 1 0 12788 0 1 68000
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__A
timestamp 1606120353
transform 1 0 12420 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_121_119
timestamp 1606120353
transform 1 0 12052 0 1 68000
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_121_125
timestamp 1606120353
transform 1 0 12604 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_646
timestamp 1606120353
transform 1 0 15180 0 1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__A
timestamp 1606120353
transform 1 0 13800 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__B
timestamp 1606120353
transform 1 0 14168 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_121_136
timestamp 1606120353
transform 1 0 13616 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_121_140
timestamp 1606120353
transform 1 0 13984 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_121_144
timestamp 1606120353
transform 1 0 14352 0 1 68000
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_121_152
timestamp 1606120353
transform 1 0 15088 0 1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_121_154
timestamp 1606120353
transform 1 0 15272 0 1 68000
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1208_
timestamp 1606120353
transform 1 0 16100 0 1 68000
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__D
timestamp 1606120353
transform 1 0 15916 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_121_160
timestamp 1606120353
transform 1 0 15824 0 1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1606120353
transform -1 0 18860 0 1 68000
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_121_182
timestamp 1606120353
transform 1 0 17848 0 1 68000
box 0 -48 736 592
use sky130_fd_sc_hd__o21a_4  _0862_
timestamp 1606120353
transform 1 0 1656 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1606120353
transform 1 0 1104 0 -1 69088
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__D
timestamp 1606120353
transform 1 0 2944 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_122_3
timestamp 1606120353
transform 1 0 1380 0 -1 69088
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_122_18
timestamp 1606120353
transform 1 0 2760 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_122_22
timestamp 1606120353
transform 1 0 3128 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0898_
timestamp 1606120353
transform 1 0 3496 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__D
timestamp 1606120353
transform 1 0 4784 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__CLK
timestamp 1606120353
transform 1 0 3312 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_122_38
timestamp 1606120353
transform 1 0 4600 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_122_42
timestamp 1606120353
transform 1 0 4968 0 -1 69088
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _0830_
timestamp 1606120353
transform 1 0 5336 0 -1 69088
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_122_49
timestamp 1606120353
transform 1 0 5612 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__B1
timestamp 1606120353
transform 1 0 5796 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_122_53
timestamp 1606120353
transform 1 0 5980 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__A2
timestamp 1606120353
transform 1 0 6164 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_122_57
timestamp 1606120353
transform 1 0 6348 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__CLK
timestamp 1606120353
transform 1 0 6532 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_122_62
timestamp 1606120353
transform 1 0 6808 0 -1 69088
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_647
timestamp 1606120353
transform 1 0 6716 0 -1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0663__A
timestamp 1606120353
transform 1 0 7176 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _0664_
timestamp 1606120353
transform 1 0 7360 0 -1 69088
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__B
timestamp 1606120353
transform 1 0 9200 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__D
timestamp 1606120353
transform 1 0 8832 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_122_82
timestamp 1606120353
transform 1 0 8648 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_122_86
timestamp 1606120353
transform 1 0 9016 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _0615_
timestamp 1606120353
transform 1 0 9384 0 -1 69088
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0606__B
timestamp 1606120353
transform 1 0 11132 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_122_107
timestamp 1606120353
transform 1 0 10948 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_122_111
timestamp 1606120353
transform 1 0 11316 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0606__C
timestamp 1606120353
transform 1 0 11500 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_122_115
timestamp 1606120353
transform 1 0 11684 0 -1 69088
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_122_121
timestamp 1606120353
transform 1 0 12236 0 -1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__B
timestamp 1606120353
transform 1 0 12052 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_648
timestamp 1606120353
transform 1 0 12328 0 -1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_122_126
timestamp 1606120353
transform 1 0 12696 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0544_
timestamp 1606120353
transform 1 0 12420 0 -1 69088
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_122_130
timestamp 1606120353
transform 1 0 13064 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0630__B
timestamp 1606120353
transform 1 0 12880 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0630__A
timestamp 1606120353
transform 1 0 13248 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _1144_
timestamp 1606120353
transform 1 0 13800 0 -1 69088
box 0 -48 644 592
use sky130_fd_sc_hd__decap_4  FILLER_122_134
timestamp 1606120353
transform 1 0 13432 0 -1 69088
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_122_145
timestamp 1606120353
transform 1 0 14444 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__CLK
timestamp 1606120353
transform 1 0 16100 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_122_157
timestamp 1606120353
transform 1 0 15548 0 -1 69088
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_122_165
timestamp 1606120353
transform 1 0 16284 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1606120353
transform -1 0 18860 0 -1 69088
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_649
timestamp 1606120353
transform 1 0 17940 0 -1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_122_177
timestamp 1606120353
transform 1 0 17388 0 -1 69088
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILLER_122_184
timestamp 1606120353
transform 1 0 18032 0 -1 69088
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _0861_
timestamp 1606120353
transform 1 0 2116 0 1 69088
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1606120353
transform 1 0 1104 0 1 69088
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A
timestamp 1606120353
transform 1 0 2944 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__A2
timestamp 1606120353
transform 1 0 1656 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_123_3
timestamp 1606120353
transform 1 0 1380 0 1 69088
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_123_8
timestamp 1606120353
transform 1 0 1840 0 1 69088
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_123_18
timestamp 1606120353
transform 1 0 2760 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_123_22
timestamp 1606120353
transform 1 0 3128 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__nand2_4  _0897_
timestamp 1606120353
transform 1 0 4048 0 1 69088
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_650
timestamp 1606120353
transform 1 0 3956 0 1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__B
timestamp 1606120353
transform 1 0 3772 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A
timestamp 1606120353
transform 1 0 5060 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__B
timestamp 1606120353
transform 1 0 3312 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_123_26
timestamp 1606120353
transform 1 0 3496 0 1 69088
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_123_41
timestamp 1606120353
transform 1 0 4876 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0880_
timestamp 1606120353
transform 1 0 5796 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__A1
timestamp 1606120353
transform 1 0 5612 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__D
timestamp 1606120353
transform 1 0 7084 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_123_45
timestamp 1606120353
transform 1 0 5244 0 1 69088
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_123_63
timestamp 1606120353
transform 1 0 6900 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0586_
timestamp 1606120353
transform 1 0 7636 0 1 69088
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__C
timestamp 1606120353
transform 1 0 9016 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__C
timestamp 1606120353
transform 1 0 8648 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__A
timestamp 1606120353
transform 1 0 7452 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_123_67
timestamp 1606120353
transform 1 0 7268 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_123_80
timestamp 1606120353
transform 1 0 8464 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_123_84
timestamp 1606120353
transform 1 0 8832 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_123_88
timestamp 1606120353
transform 1 0 9200 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _0588_
timestamp 1606120353
transform 1 0 9752 0 1 69088
box 0 -48 1564 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_651
timestamp 1606120353
transform 1 0 9568 0 1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__B
timestamp 1606120353
transform 1 0 9384 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_123_93
timestamp 1606120353
transform 1 0 9660 0 1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__nand3_4  _0609_
timestamp 1606120353
transform 1 0 12052 0 1 69088
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__A
timestamp 1606120353
transform 1 0 11868 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__A
timestamp 1606120353
transform 1 0 11500 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_123_111
timestamp 1606120353
transform 1 0 11316 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_123_115
timestamp 1606120353
transform 1 0 11684 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_652
timestamp 1606120353
transform 1 0 15180 0 1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_123_133
timestamp 1606120353
transform 1 0 13340 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_123_145
timestamp 1606120353
transform 1 0 14444 0 1 69088
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_123_154
timestamp 1606120353
transform 1 0 15272 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_123_166
timestamp 1606120353
transform 1 0 16376 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1606120353
transform -1 0 18860 0 1 69088
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_123_178
timestamp 1606120353
transform 1 0 17480 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1160_
timestamp 1606120353
transform 1 0 1472 0 -1 70176
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1606120353
transform 1 0 1104 0 -1 70176
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_124_3
timestamp 1606120353
transform 1 0 1380 0 -1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0871_
timestamp 1606120353
transform 1 0 5060 0 -1 70176
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A
timestamp 1606120353
transform 1 0 4048 0 -1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_124_23
timestamp 1606120353
transform 1 0 3220 0 -1 70176
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_124_31
timestamp 1606120353
transform 1 0 3956 0 -1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_124_34
timestamp 1606120353
transform 1 0 4232 0 -1 70176
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_124_42
timestamp 1606120353
transform 1 0 4968 0 -1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1167_
timestamp 1606120353
transform 1 0 6808 0 -1 70176
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_653
timestamp 1606120353
transform 1 0 6716 0 -1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__B
timestamp 1606120353
transform 1 0 5796 0 -1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__A
timestamp 1606120353
transform 1 0 6532 0 -1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_124_46
timestamp 1606120353
transform 1 0 5336 0 -1 70176
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_124_50
timestamp 1606120353
transform 1 0 5704 0 -1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_124_53
timestamp 1606120353
transform 1 0 5980 0 -1 70176
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__A
timestamp 1606120353
transform 1 0 9108 0 -1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__A
timestamp 1606120353
transform 1 0 8740 0 -1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_124_81
timestamp 1606120353
transform 1 0 8556 0 -1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_124_85
timestamp 1606120353
transform 1 0 8924 0 -1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__nand4_4  _0590_
timestamp 1606120353
transform 1 0 9292 0 -1 70176
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__D
timestamp 1606120353
transform 1 0 11040 0 -1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_124_106
timestamp 1606120353
transform 1 0 10856 0 -1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_124_110
timestamp 1606120353
transform 1 0 11224 0 -1 70176
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_654
timestamp 1606120353
transform 1 0 12328 0 -1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__B
timestamp 1606120353
transform 1 0 11776 0 -1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__C
timestamp 1606120353
transform 1 0 12144 0 -1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_124_118
timestamp 1606120353
transform 1 0 11960 0 -1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_124_123
timestamp 1606120353
transform 1 0 12420 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_135
timestamp 1606120353
transform 1 0 13524 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_147
timestamp 1606120353
transform 1 0 14628 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_159
timestamp 1606120353
transform 1 0 15732 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_171
timestamp 1606120353
transform 1 0 16836 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1606120353
transform -1 0 18860 0 -1 70176
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_655
timestamp 1606120353
transform 1 0 17940 0 -1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_124_184
timestamp 1606120353
transform 1 0 18032 0 -1 70176
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1606120353
transform 1 0 1104 0 1 70176
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1606120353
transform 1 0 1104 0 -1 71264
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__D
timestamp 1606120353
transform 1 0 1564 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__CLK
timestamp 1606120353
transform 1 0 1932 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_125_3
timestamp 1606120353
transform 1 0 1380 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_125_7
timestamp 1606120353
transform 1 0 1748 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_125_11
timestamp 1606120353
transform 1 0 2116 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_3
timestamp 1606120353
transform 1 0 1380 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_15
timestamp 1606120353
transform 1 0 2484 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_126_31
timestamp 1606120353
transform 1 0 3956 0 -1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_126_27
timestamp 1606120353
transform 1 0 3588 0 -1 71264
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_125_23
timestamp 1606120353
transform 1 0 3220 0 1 70176
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_656
timestamp 1606120353
transform 1 0 3956 0 1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_125_40
timestamp 1606120353
transform 1 0 4784 0 1 70176
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_125_36
timestamp 1606120353
transform 1 0 4416 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_125_32
timestamp 1606120353
transform 1 0 4048 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__B
timestamp 1606120353
transform 1 0 4600 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A
timestamp 1606120353
transform 1 0 4232 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__nand2_4  _0893_
timestamp 1606120353
transform 1 0 4048 0 -1 71264
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_126_41
timestamp 1606120353
transform 1 0 4876 0 -1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__D
timestamp 1606120353
transform 1 0 5060 0 -1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_126_45
timestamp 1606120353
transform 1 0 5244 0 -1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_125_48
timestamp 1606120353
transform 1 0 5520 0 1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__CLK
timestamp 1606120353
transform 1 0 5428 0 -1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__A
timestamp 1606120353
transform 1 0 5612 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__nand2_4  _0885_
timestamp 1606120353
transform 1 0 5796 0 1 70176
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_125_66
timestamp 1606120353
transform 1 0 7176 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_125_60
timestamp 1606120353
transform 1 0 6624 0 1 70176
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__A2
timestamp 1606120353
transform 1 0 6992 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_659
timestamp 1606120353
transform 1 0 6716 0 -1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _0747_
timestamp 1606120353
transform 1 0 6808 0 -1 71264
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILLER_126_49
timestamp 1606120353
transform 1 0 5612 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_126_75
timestamp 1606120353
transform 1 0 8004 0 -1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_126_71
timestamp 1606120353
transform 1 0 7636 0 -1 71264
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__A2_N
timestamp 1606120353
transform 1 0 8096 0 -1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__A1
timestamp 1606120353
transform 1 0 7360 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_126_82
timestamp 1606120353
transform 1 0 8648 0 -1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_126_78
timestamp 1606120353
transform 1 0 8280 0 -1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_125_88
timestamp 1606120353
transform 1 0 9200 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_125_84
timestamp 1606120353
transform 1 0 8832 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__B2
timestamp 1606120353
transform 1 0 8464 0 -1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__B1
timestamp 1606120353
transform 1 0 9016 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0722_
timestamp 1606120353
transform 1 0 8832 0 -1 71264
box 0 -48 828 592
use sky130_fd_sc_hd__o22a_4  _0591_
timestamp 1606120353
transform 1 0 7544 0 1 70176
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_126_97
timestamp 1606120353
transform 1 0 10028 0 -1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_126_93
timestamp 1606120353
transform 1 0 9660 0 -1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_125_93
timestamp 1606120353
transform 1 0 9660 0 1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__C
timestamp 1606120353
transform 1 0 10212 0 -1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__B
timestamp 1606120353
transform 1 0 9844 0 -1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__A
timestamp 1606120353
transform 1 0 9384 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_657
timestamp 1606120353
transform 1 0 9568 0 1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_126_109
timestamp 1606120353
transform 1 0 11132 0 -1 71264
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_126_105
timestamp 1606120353
transform 1 0 10764 0 -1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_126_101
timestamp 1606120353
transform 1 0 10396 0 -1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_125_108
timestamp 1606120353
transform 1 0 11040 0 1 70176
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__A4
timestamp 1606120353
transform 1 0 10948 0 -1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__A2
timestamp 1606120353
transform 1 0 10580 0 -1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__nand3_4  _0607_
timestamp 1606120353
transform 1 0 9752 0 1 70176
box 0 -48 1288 592
use sky130_fd_sc_hd__nand3_4  _0608_
timestamp 1606120353
transform 1 0 11776 0 1 70176
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_660
timestamp 1606120353
transform 1 0 12328 0 -1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__A
timestamp 1606120353
transform 1 0 11592 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__C
timestamp 1606120353
transform 1 0 11776 0 -1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_125_130
timestamp 1606120353
transform 1 0 13064 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_126_115
timestamp 1606120353
transform 1 0 11684 0 -1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_126_118
timestamp 1606120353
transform 1 0 11960 0 -1 71264
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_126_123
timestamp 1606120353
transform 1 0 12420 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_658
timestamp 1606120353
transform 1 0 15180 0 1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_125_142
timestamp 1606120353
transform 1 0 14168 0 1 70176
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_125_150
timestamp 1606120353
transform 1 0 14904 0 1 70176
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_125_154
timestamp 1606120353
transform 1 0 15272 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_135
timestamp 1606120353
transform 1 0 13524 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_147
timestamp 1606120353
transform 1 0 14628 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__CLK
timestamp 1606120353
transform 1 0 16100 0 -1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_125_166
timestamp 1606120353
transform 1 0 16376 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_126_159
timestamp 1606120353
transform 1 0 15732 0 -1 71264
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_126_165
timestamp 1606120353
transform 1 0 16284 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1606120353
transform -1 0 18860 0 1 70176
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1606120353
transform -1 0 18860 0 -1 71264
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_661
timestamp 1606120353
transform 1 0 17940 0 -1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_125_178
timestamp 1606120353
transform 1 0 17480 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_126_177
timestamp 1606120353
transform 1 0 17388 0 -1 71264
box 0 -48 552 592
use sky130_fd_sc_hd__decap_6  FILLER_126_184
timestamp 1606120353
transform 1 0 18032 0 -1 71264
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1606120353
transform 1 0 1104 0 1 71264
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_127_3
timestamp 1606120353
transform 1 0 1380 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_127_15
timestamp 1606120353
transform 1 0 2484 0 1 71264
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_127_32
timestamp 1606120353
transform 1 0 4048 0 1 71264
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_127_29
timestamp 1606120353
transform 1 0 3772 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_127_25
timestamp 1606120353
transform 1 0 3404 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__CLK
timestamp 1606120353
transform 1 0 3220 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__D
timestamp 1606120353
transform 1 0 3588 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_662
timestamp 1606120353
transform 1 0 3956 0 1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_127_39
timestamp 1606120353
transform 1 0 4692 0 1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_127_36
timestamp 1606120353
transform 1 0 4416 0 1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A2
timestamp 1606120353
transform 1 0 4508 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1170_
timestamp 1606120353
transform 1 0 4784 0 1 71264
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__B1
timestamp 1606120353
transform 1 0 7084 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__A
timestamp 1606120353
transform 1 0 6716 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_127_59
timestamp 1606120353
transform 1 0 6532 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_127_63
timestamp 1606120353
transform 1 0 6900 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0721_
timestamp 1606120353
transform 1 0 7636 0 1 71264
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A1
timestamp 1606120353
transform 1 0 7452 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__A1_N
timestamp 1606120353
transform 1 0 9016 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_127_67
timestamp 1606120353
transform 1 0 7268 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_127_84
timestamp 1606120353
transform 1 0 8832 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_127_88
timestamp 1606120353
transform 1 0 9200 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__a41o_4  _0613_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 10580 0 1 71264
box 0 -48 1564 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_663
timestamp 1606120353
transform 1 0 9568 0 1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__A1
timestamp 1606120353
transform 1 0 10396 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__A3
timestamp 1606120353
transform 1 0 10028 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__B2
timestamp 1606120353
transform 1 0 9384 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_127_93
timestamp 1606120353
transform 1 0 9660 0 1 71264
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_127_99
timestamp 1606120353
transform 1 0 10212 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0612_
timestamp 1606120353
transform 1 0 12880 0 1 71264
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__A
timestamp 1606120353
transform 1 0 12696 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_127_120
timestamp 1606120353
transform 1 0 12144 0 1 71264
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_664
timestamp 1606120353
transform 1 0 15180 0 1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_127_137
timestamp 1606120353
transform 1 0 13708 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_127_149
timestamp 1606120353
transform 1 0 14812 0 1 71264
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_127_154
timestamp 1606120353
transform 1 0 15272 0 1 71264
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1201_
timestamp 1606120353
transform 1 0 16100 0 1 71264
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__D
timestamp 1606120353
transform 1 0 15916 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_127_160
timestamp 1606120353
transform 1 0 15824 0 1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1606120353
transform -1 0 18860 0 1 71264
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_127_182
timestamp 1606120353
transform 1 0 17848 0 1 71264
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1606120353
transform 1 0 1104 0 -1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_128_3
timestamp 1606120353
transform 1 0 1380 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_15
timestamp 1606120353
transform 1 0 2484 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1174_
timestamp 1606120353
transform 1 0 3588 0 -1 72352
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_2  FILLER_128_46
timestamp 1606120353
transform 1 0 5336 0 -1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__B1
timestamp 1606120353
transform 1 0 5520 0 -1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_128_50
timestamp 1606120353
transform 1 0 5704 0 -1 72352
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_128_54
timestamp 1606120353
transform 1 0 6072 0 -1 72352
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__CLK
timestamp 1606120353
transform 1 0 6164 0 -1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_128_57
timestamp 1606120353
transform 1 0 6348 0 -1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__B
timestamp 1606120353
transform 1 0 6532 0 -1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_128_62
timestamp 1606120353
transform 1 0 6808 0 -1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_665
timestamp 1606120353
transform 1 0 6716 0 -1 72352
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0540_
timestamp 1606120353
transform 1 0 7084 0 -1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__a2bb2oi_4  _0720_
timestamp 1606120353
transform 1 0 8096 0 -1 72352
box 0 -48 1932 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A2
timestamp 1606120353
transform 1 0 7636 0 -1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_128_68
timestamp 1606120353
transform 1 0 7360 0 -1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_128_73
timestamp 1606120353
transform 1 0 7820 0 -1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__A2
timestamp 1606120353
transform 1 0 10764 0 -1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__B1
timestamp 1606120353
transform 1 0 11132 0 -1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_128_97
timestamp 1606120353
transform 1 0 10028 0 -1 72352
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_128_107
timestamp 1606120353
transform 1 0 10948 0 -1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_666
timestamp 1606120353
transform 1 0 12328 0 -1 72352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_128_111
timestamp 1606120353
transform 1 0 11316 0 -1 72352
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_128_119
timestamp 1606120353
transform 1 0 12052 0 -1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_128_123
timestamp 1606120353
transform 1 0 12420 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_135
timestamp 1606120353
transform 1 0 13524 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_147
timestamp 1606120353
transform 1 0 14628 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_159
timestamp 1606120353
transform 1 0 15732 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_171
timestamp 1606120353
transform 1 0 16836 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1606120353
transform -1 0 18860 0 -1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_667
timestamp 1606120353
transform 1 0 17940 0 -1 72352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_128_184
timestamp 1606120353
transform 1 0 18032 0 -1 72352
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1606120353
transform 1 0 1104 0 1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A1
timestamp 1606120353
transform 1 0 2944 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A2
timestamp 1606120353
transform 1 0 2576 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_129_3
timestamp 1606120353
transform 1 0 1380 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_129_15
timestamp 1606120353
transform 1 0 2484 0 1 72352
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_129_18
timestamp 1606120353
transform 1 0 2760 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_129_22
timestamp 1606120353
transform 1 0 3128 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0886_
timestamp 1606120353
transform 1 0 4508 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_668
timestamp 1606120353
transform 1 0 3956 0 1 72352
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A1
timestamp 1606120353
transform 1 0 4324 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__B1
timestamp 1606120353
transform 1 0 3312 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__A2
timestamp 1606120353
transform 1 0 3772 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_129_26
timestamp 1606120353
transform 1 0 3496 0 1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_129_32
timestamp 1606120353
transform 1 0 4048 0 1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1168_
timestamp 1606120353
transform 1 0 6348 0 1 72352
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__A
timestamp 1606120353
transform 1 0 6164 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__A1
timestamp 1606120353
transform 1 0 5796 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_129_49
timestamp 1606120353
transform 1 0 5612 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_129_53
timestamp 1606120353
transform 1 0 5980 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__A1_N
timestamp 1606120353
transform 1 0 8372 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__A2_N
timestamp 1606120353
transform 1 0 8740 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__B2
timestamp 1606120353
transform 1 0 9108 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_129_76
timestamp 1606120353
transform 1 0 8096 0 1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_129_81
timestamp 1606120353
transform 1 0 8556 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_129_85
timestamp 1606120353
transform 1 0 8924 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__a32oi_4  _0604_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 10764 0 1 72352
box 0 -48 2024 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_669
timestamp 1606120353
transform 1 0 9568 0 1 72352
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__A3
timestamp 1606120353
transform 1 0 10580 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__A1
timestamp 1606120353
transform 1 0 10212 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__B1
timestamp 1606120353
transform 1 0 9844 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_129_89
timestamp 1606120353
transform 1 0 9292 0 1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_129_93
timestamp 1606120353
transform 1 0 9660 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_129_97
timestamp 1606120353
transform 1 0 10028 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_129_101
timestamp 1606120353
transform 1 0 10396 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_129_127
timestamp 1606120353
transform 1 0 12788 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_670
timestamp 1606120353
transform 1 0 15180 0 1 72352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_129_139
timestamp 1606120353
transform 1 0 13892 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_129_151
timestamp 1606120353
transform 1 0 14996 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_129_154
timestamp 1606120353
transform 1 0 15272 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_129_166
timestamp 1606120353
transform 1 0 16376 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1606120353
transform -1 0 18860 0 1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_129_178
timestamp 1606120353
transform 1 0 17480 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__o21a_4  _0894_
timestamp 1606120353
transform 1 0 2944 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1606120353
transform 1 0 1104 0 -1 73440
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__A
timestamp 1606120353
transform 1 0 2576 0 -1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_130_3
timestamp 1606120353
transform 1 0 1380 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_130_15
timestamp 1606120353
transform 1 0 2484 0 -1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_130_18
timestamp 1606120353
transform 1 0 2760 0 -1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0884_
timestamp 1606120353
transform 1 0 4784 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__B1
timestamp 1606120353
transform 1 0 4232 0 -1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__B1
timestamp 1606120353
transform 1 0 4600 0 -1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_130_32
timestamp 1606120353
transform 1 0 4048 0 -1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_130_36
timestamp 1606120353
transform 1 0 4416 0 -1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__nand2_4  _0881_
timestamp 1606120353
transform 1 0 6808 0 -1 73440
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_671
timestamp 1606120353
transform 1 0 6716 0 -1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__D
timestamp 1606120353
transform 1 0 6348 0 -1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_130_52
timestamp 1606120353
transform 1 0 5888 0 -1 73440
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_130_56
timestamp 1606120353
transform 1 0 6256 0 -1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_130_59
timestamp 1606120353
transform 1 0 6532 0 -1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__a2bb2oi_4  _0618_
timestamp 1606120353
transform 1 0 8372 0 -1 73440
box 0 -48 1932 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__B1
timestamp 1606120353
transform 1 0 8096 0 -1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_130_71
timestamp 1606120353
transform 1 0 7636 0 -1 73440
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_130_75
timestamp 1606120353
transform 1 0 8004 0 -1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_130_78
timestamp 1606120353
transform 1 0 8280 0 -1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__B1
timestamp 1606120353
transform 1 0 10764 0 -1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__B2
timestamp 1606120353
transform 1 0 11132 0 -1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_130_100
timestamp 1606120353
transform 1 0 10304 0 -1 73440
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_130_104
timestamp 1606120353
transform 1 0 10672 0 -1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_130_107
timestamp 1606120353
transform 1 0 10948 0 -1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_672
timestamp 1606120353
transform 1 0 12328 0 -1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_130_111
timestamp 1606120353
transform 1 0 11316 0 -1 73440
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_130_119
timestamp 1606120353
transform 1 0 12052 0 -1 73440
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_130_123
timestamp 1606120353
transform 1 0 12420 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_130_135
timestamp 1606120353
transform 1 0 13524 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_130_147
timestamp 1606120353
transform 1 0 14628 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_130_159
timestamp 1606120353
transform 1 0 15732 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_130_171
timestamp 1606120353
transform 1 0 16836 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1606120353
transform -1 0 18860 0 -1 73440
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_673
timestamp 1606120353
transform 1 0 17940 0 -1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_130_184
timestamp 1606120353
transform 1 0 18032 0 -1 73440
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _0891_
timestamp 1606120353
transform 1 0 2576 0 1 73440
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1606120353
transform 1 0 1104 0 1 73440
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__D
timestamp 1606120353
transform 1 0 2392 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__CLK
timestamp 1606120353
transform 1 0 2024 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_131_3
timestamp 1606120353
transform 1 0 1380 0 1 73440
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_131_9
timestamp 1606120353
transform 1 0 1932 0 1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_131_12
timestamp 1606120353
transform 1 0 2208 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0882_
timestamp 1606120353
transform 1 0 4232 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_674
timestamp 1606120353
transform 1 0 3956 0 1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__B
timestamp 1606120353
transform 1 0 3404 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A1
timestamp 1606120353
transform 1 0 3772 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_131_23
timestamp 1606120353
transform 1 0 3220 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_131_27
timestamp 1606120353
transform 1 0 3588 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_131_32
timestamp 1606120353
transform 1 0 4048 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1169_
timestamp 1606120353
transform 1 0 6072 0 1 73440
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__A
timestamp 1606120353
transform 1 0 5520 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__B
timestamp 1606120353
transform 1 0 5888 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_131_46
timestamp 1606120353
transform 1 0 5336 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_131_50
timestamp 1606120353
transform 1 0 5704 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0614__A
timestamp 1606120353
transform 1 0 8004 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_131_73
timestamp 1606120353
transform 1 0 7820 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_131_77
timestamp 1606120353
transform 1 0 8188 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__nand3_4  _0619_
timestamp 1606120353
transform 1 0 10028 0 1 73440
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_675
timestamp 1606120353
transform 1 0 9568 0 1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__A
timestamp 1606120353
transform 1 0 9844 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__C
timestamp 1606120353
transform 1 0 9384 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_131_89
timestamp 1606120353
transform 1 0 9292 0 1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_131_93
timestamp 1606120353
transform 1 0 9660 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_131_111
timestamp 1606120353
transform 1 0 11316 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_131_123
timestamp 1606120353
transform 1 0 12420 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_676
timestamp 1606120353
transform 1 0 15180 0 1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_131_135
timestamp 1606120353
transform 1 0 13524 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_131_147
timestamp 1606120353
transform 1 0 14628 0 1 73440
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_131_154
timestamp 1606120353
transform 1 0 15272 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_131_166
timestamp 1606120353
transform 1 0 16376 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1606120353
transform -1 0 18860 0 1 73440
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_131_178
timestamp 1606120353
transform 1 0 17480 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__o21a_4  _0892_
timestamp 1606120353
transform 1 0 2116 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1173_
timestamp 1606120353
transform 1 0 2668 0 -1 74528
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1606120353
transform 1 0 1104 0 -1 74528
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1606120353
transform 1 0 1104 0 1 74528
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__A1
timestamp 1606120353
transform 1 0 1932 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__B1
timestamp 1606120353
transform 1 0 2116 0 -1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_132_3
timestamp 1606120353
transform 1 0 1380 0 -1 74528
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_132_13
timestamp 1606120353
transform 1 0 2300 0 -1 74528
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_133_3
timestamp 1606120353
transform 1 0 1380 0 1 74528
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_133_32
timestamp 1606120353
transform 1 0 4048 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_133_27
timestamp 1606120353
transform 1 0 3588 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_133_23
timestamp 1606120353
transform 1 0 3220 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__A2
timestamp 1606120353
transform 1 0 3404 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__B1
timestamp 1606120353
transform 1 0 3772 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_680
timestamp 1606120353
transform 1 0 3956 0 1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_132_40
timestamp 1606120353
transform 1 0 4784 0 -1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_132_36
timestamp 1606120353
transform 1 0 4416 0 -1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__D
timestamp 1606120353
transform 1 0 4968 0 -1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A2
timestamp 1606120353
transform 1 0 4600 0 -1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__A1
timestamp 1606120353
transform 1 0 4232 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _0883_
timestamp 1606120353
transform 1 0 5152 0 -1 74528
box 0 -48 644 592
use sky130_fd_sc_hd__dfxtp_4  _1172_
timestamp 1606120353
transform 1 0 4416 0 1 74528
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  FILLER_132_51
timestamp 1606120353
transform 1 0 5796 0 -1 74528
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__D
timestamp 1606120353
transform 1 0 6072 0 -1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_133_55
timestamp 1606120353
transform 1 0 6164 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__B
timestamp 1606120353
transform 1 0 6348 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_132_56
timestamp 1606120353
transform 1 0 6256 0 -1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__CLK
timestamp 1606120353
transform 1 0 6440 0 -1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_133_59
timestamp 1606120353
transform 1 0 6532 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_677
timestamp 1606120353
transform 1 0 6716 0 -1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A
timestamp 1606120353
transform 1 0 6716 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_132_60
timestamp 1606120353
transform 1 0 6624 0 -1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_132_62
timestamp 1606120353
transform 1 0 6808 0 -1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_132_66
timestamp 1606120353
transform 1 0 7176 0 -1 74528
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__A
timestamp 1606120353
transform 1 0 6992 0 -1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__nand2_4  _0889_
timestamp 1606120353
transform 1 0 6900 0 1 74528
box 0 -48 828 592
use sky130_fd_sc_hd__inv_8  _0614_
timestamp 1606120353
transform 1 0 7636 0 -1 74528
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILLER_132_70
timestamp 1606120353
transform 1 0 7544 0 -1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_132_80
timestamp 1606120353
transform 1 0 8464 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_72
timestamp 1606120353
transform 1 0 7728 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_133_84
timestamp 1606120353
transform 1 0 8832 0 1 74528
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_681
timestamp 1606120353
transform 1 0 9568 0 1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__B
timestamp 1606120353
transform 1 0 10028 0 -1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_132_92
timestamp 1606120353
transform 1 0 9568 0 -1 74528
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_132_96
timestamp 1606120353
transform 1 0 9936 0 -1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_132_99
timestamp 1606120353
transform 1 0 10212 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_93
timestamp 1606120353
transform 1 0 9660 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_105
timestamp 1606120353
transform 1 0 10764 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_678
timestamp 1606120353
transform 1 0 12328 0 -1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_132_111
timestamp 1606120353
transform 1 0 11316 0 -1 74528
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_132_119
timestamp 1606120353
transform 1 0 12052 0 -1 74528
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_132_123
timestamp 1606120353
transform 1 0 12420 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_117
timestamp 1606120353
transform 1 0 11868 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_129
timestamp 1606120353
transform 1 0 12972 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_682
timestamp 1606120353
transform 1 0 15180 0 1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_132_135
timestamp 1606120353
transform 1 0 13524 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_132_147
timestamp 1606120353
transform 1 0 14628 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_141
timestamp 1606120353
transform 1 0 14076 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_154
timestamp 1606120353
transform 1 0 15272 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_132_159
timestamp 1606120353
transform 1 0 15732 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_132_171
timestamp 1606120353
transform 1 0 16836 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_166
timestamp 1606120353
transform 1 0 16376 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1606120353
transform -1 0 18860 0 -1 74528
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1606120353
transform -1 0 18860 0 1 74528
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_679
timestamp 1606120353
transform 1 0 17940 0 -1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_132_184
timestamp 1606120353
transform 1 0 18032 0 -1 74528
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_133_178
timestamp 1606120353
transform 1 0 17480 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1606120353
transform 1 0 1104 0 -1 75616
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__A2
timestamp 1606120353
transform 1 0 2116 0 -1 75616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_134_3
timestamp 1606120353
transform 1 0 1380 0 -1 75616
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_134_13
timestamp 1606120353
transform 1 0 2300 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__o21a_4  _0890_
timestamp 1606120353
transform 1 0 4324 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__CLK
timestamp 1606120353
transform 1 0 4140 0 -1 75616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_134_25
timestamp 1606120353
transform 1 0 3404 0 -1 75616
box 0 -48 736 592
use sky130_fd_sc_hd__inv_8  _0786_
timestamp 1606120353
transform 1 0 6992 0 -1 75616
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_683
timestamp 1606120353
transform 1 0 6716 0 -1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_134_47
timestamp 1606120353
transform 1 0 5428 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_134_59
timestamp 1606120353
transform 1 0 6532 0 -1 75616
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_134_62
timestamp 1606120353
transform 1 0 6808 0 -1 75616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_134_73
timestamp 1606120353
transform 1 0 7820 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_134_85
timestamp 1606120353
transform 1 0 8924 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_134_97
timestamp 1606120353
transform 1 0 10028 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_134_109
timestamp 1606120353
transform 1 0 11132 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_684
timestamp 1606120353
transform 1 0 12328 0 -1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_134_121
timestamp 1606120353
transform 1 0 12236 0 -1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_134_123
timestamp 1606120353
transform 1 0 12420 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_134_135
timestamp 1606120353
transform 1 0 13524 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_134_147
timestamp 1606120353
transform 1 0 14628 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_134_159
timestamp 1606120353
transform 1 0 15732 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_134_171
timestamp 1606120353
transform 1 0 16836 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1606120353
transform -1 0 18860 0 -1 75616
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_685
timestamp 1606120353
transform 1 0 17940 0 -1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_134_184
timestamp 1606120353
transform 1 0 18032 0 -1 75616
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1606120353
transform 1 0 1104 0 1 75616
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_135_3
timestamp 1606120353
transform 1 0 1380 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_15
timestamp 1606120353
transform 1 0 2484 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_686
timestamp 1606120353
transform 1 0 3956 0 1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_135_27
timestamp 1606120353
transform 1 0 3588 0 1 75616
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_135_32
timestamp 1606120353
transform 1 0 4048 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_44
timestamp 1606120353
transform 1 0 5152 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_56
timestamp 1606120353
transform 1 0 6256 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_68
timestamp 1606120353
transform 1 0 7360 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_80
timestamp 1606120353
transform 1 0 8464 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_687
timestamp 1606120353
transform 1 0 9568 0 1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_135_93
timestamp 1606120353
transform 1 0 9660 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_105
timestamp 1606120353
transform 1 0 10764 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_117
timestamp 1606120353
transform 1 0 11868 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_129
timestamp 1606120353
transform 1 0 12972 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_688
timestamp 1606120353
transform 1 0 15180 0 1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_135_141
timestamp 1606120353
transform 1 0 14076 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_154
timestamp 1606120353
transform 1 0 15272 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_166
timestamp 1606120353
transform 1 0 16376 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1606120353
transform -1 0 18860 0 1 75616
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_135_178
timestamp 1606120353
transform 1 0 17480 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1606120353
transform 1 0 1104 0 -1 76704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_136_3
timestamp 1606120353
transform 1 0 1380 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_15
timestamp 1606120353
transform 1 0 2484 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_27
timestamp 1606120353
transform 1 0 3588 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_39
timestamp 1606120353
transform 1 0 4692 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_689
timestamp 1606120353
transform 1 0 6716 0 -1 76704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_136_51
timestamp 1606120353
transform 1 0 5796 0 -1 76704
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_136_59
timestamp 1606120353
transform 1 0 6532 0 -1 76704
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_136_62
timestamp 1606120353
transform 1 0 6808 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_74
timestamp 1606120353
transform 1 0 7912 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_86
timestamp 1606120353
transform 1 0 9016 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_98
timestamp 1606120353
transform 1 0 10120 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_110
timestamp 1606120353
transform 1 0 11224 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_690
timestamp 1606120353
transform 1 0 12328 0 -1 76704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_136_123
timestamp 1606120353
transform 1 0 12420 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_135
timestamp 1606120353
transform 1 0 13524 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_147
timestamp 1606120353
transform 1 0 14628 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_159
timestamp 1606120353
transform 1 0 15732 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_171
timestamp 1606120353
transform 1 0 16836 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1606120353
transform -1 0 18860 0 -1 76704
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_691
timestamp 1606120353
transform 1 0 17940 0 -1 76704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_136_184
timestamp 1606120353
transform 1 0 18032 0 -1 76704
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1606120353
transform 1 0 1104 0 1 76704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_137_3
timestamp 1606120353
transform 1 0 1380 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_15
timestamp 1606120353
transform 1 0 2484 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_692
timestamp 1606120353
transform 1 0 3956 0 1 76704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_137_27
timestamp 1606120353
transform 1 0 3588 0 1 76704
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_137_32
timestamp 1606120353
transform 1 0 4048 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_44
timestamp 1606120353
transform 1 0 5152 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_56
timestamp 1606120353
transform 1 0 6256 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_68
timestamp 1606120353
transform 1 0 7360 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_80
timestamp 1606120353
transform 1 0 8464 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_693
timestamp 1606120353
transform 1 0 9568 0 1 76704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_137_93
timestamp 1606120353
transform 1 0 9660 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_105
timestamp 1606120353
transform 1 0 10764 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_117
timestamp 1606120353
transform 1 0 11868 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_129
timestamp 1606120353
transform 1 0 12972 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_694
timestamp 1606120353
transform 1 0 15180 0 1 76704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_137_141
timestamp 1606120353
transform 1 0 14076 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_154
timestamp 1606120353
transform 1 0 15272 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_166
timestamp 1606120353
transform 1 0 16376 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1606120353
transform -1 0 18860 0 1 76704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_137_178
timestamp 1606120353
transform 1 0 17480 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1606120353
transform 1 0 1104 0 -1 77792
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_138_3
timestamp 1606120353
transform 1 0 1380 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_138_15
timestamp 1606120353
transform 1 0 2484 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_695
timestamp 1606120353
transform 1 0 3956 0 -1 77792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_138_27
timestamp 1606120353
transform 1 0 3588 0 -1 77792
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_138_32
timestamp 1606120353
transform 1 0 4048 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_138_44
timestamp 1606120353
transform 1 0 5152 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_696
timestamp 1606120353
transform 1 0 6808 0 -1 77792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_138_56
timestamp 1606120353
transform 1 0 6256 0 -1 77792
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_138_63
timestamp 1606120353
transform 1 0 6900 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_138_75
timestamp 1606120353
transform 1 0 8004 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_138_87
timestamp 1606120353
transform 1 0 9108 0 -1 77792
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_697
timestamp 1606120353
transform 1 0 9660 0 -1 77792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_138_94
timestamp 1606120353
transform 1 0 9752 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_138_106
timestamp 1606120353
transform 1 0 10856 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_698
timestamp 1606120353
transform 1 0 12512 0 -1 77792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_138_118
timestamp 1606120353
transform 1 0 11960 0 -1 77792
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_138_125
timestamp 1606120353
transform 1 0 12604 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_138_137
timestamp 1606120353
transform 1 0 13708 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_138_149
timestamp 1606120353
transform 1 0 14812 0 -1 77792
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_699
timestamp 1606120353
transform 1 0 15364 0 -1 77792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_138_156
timestamp 1606120353
transform 1 0 15456 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_138_168
timestamp 1606120353
transform 1 0 16560 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1606120353
transform -1 0 18860 0 -1 77792
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_700
timestamp 1606120353
transform 1 0 18216 0 -1 77792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_138_180
timestamp 1606120353
transform 1 0 17664 0 -1 77792
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILLER_138_187
timestamp 1606120353
transform 1 0 18308 0 -1 77792
box 0 -48 276 592
<< labels >>
rlabel metal3 s 0 40264 480 40384 6 addr_r[0]
port 0 nsew default input
rlabel metal3 s 0 48152 480 48272 6 addr_r[10]
port 1 nsew default input
rlabel metal3 s 0 48968 480 49088 6 addr_r[11]
port 2 nsew default input
rlabel metal3 s 0 49784 480 49904 6 addr_r[12]
port 3 nsew default input
rlabel metal3 s 0 50600 480 50720 6 addr_r[13]
port 4 nsew default input
rlabel metal3 s 0 40944 480 41064 6 addr_r[1]
port 5 nsew default input
rlabel metal3 s 0 41760 480 41880 6 addr_r[2]
port 6 nsew default input
rlabel metal3 s 0 42576 480 42696 6 addr_r[3]
port 7 nsew default input
rlabel metal3 s 0 43392 480 43512 6 addr_r[4]
port 8 nsew default input
rlabel metal3 s 0 44208 480 44328 6 addr_r[5]
port 9 nsew default input
rlabel metal3 s 0 45024 480 45144 6 addr_r[6]
port 10 nsew default input
rlabel metal3 s 0 45840 480 45960 6 addr_r[7]
port 11 nsew default input
rlabel metal3 s 0 46656 480 46776 6 addr_r[8]
port 12 nsew default input
rlabel metal3 s 0 47336 480 47456 6 addr_r[9]
port 13 nsew default input
rlabel metal3 s 0 28976 480 29096 6 addr_w[0]
port 14 nsew default input
rlabel metal3 s 0 37000 480 37120 6 addr_w[10]
port 15 nsew default input
rlabel metal3 s 0 37816 480 37936 6 addr_w[11]
port 16 nsew default input
rlabel metal3 s 0 38632 480 38752 6 addr_w[12]
port 17 nsew default input
rlabel metal3 s 0 39448 480 39568 6 addr_w[13]
port 18 nsew default input
rlabel metal3 s 0 29792 480 29912 6 addr_w[1]
port 19 nsew default input
rlabel metal3 s 0 30608 480 30728 6 addr_w[2]
port 20 nsew default input
rlabel metal3 s 0 31424 480 31544 6 addr_w[3]
port 21 nsew default input
rlabel metal3 s 0 32240 480 32360 6 addr_w[4]
port 22 nsew default input
rlabel metal3 s 0 33056 480 33176 6 addr_w[5]
port 23 nsew default input
rlabel metal3 s 0 33736 480 33856 6 addr_w[6]
port 24 nsew default input
rlabel metal3 s 0 34552 480 34672 6 addr_w[7]
port 25 nsew default input
rlabel metal3 s 0 35368 480 35488 6 addr_w[8]
port 26 nsew default input
rlabel metal3 s 0 36184 480 36304 6 addr_w[9]
port 27 nsew default input
rlabel metal3 s 19520 73992 20000 74112 6 baseaddr_r_sync[0]
port 28 nsew default tristate
rlabel metal3 s 19520 74672 20000 74792 6 baseaddr_r_sync[1]
port 29 nsew default tristate
rlabel metal3 s 19520 75352 20000 75472 6 baseaddr_r_sync[2]
port 30 nsew default tristate
rlabel metal3 s 19520 76032 20000 76152 6 baseaddr_r_sync[3]
port 31 nsew default tristate
rlabel metal3 s 19520 76712 20000 76832 6 baseaddr_r_sync[4]
port 32 nsew default tristate
rlabel metal3 s 19520 77392 20000 77512 6 baseaddr_r_sync[5]
port 33 nsew default tristate
rlabel metal3 s 19520 78072 20000 78192 6 baseaddr_r_sync[6]
port 34 nsew default tristate
rlabel metal3 s 19520 78752 20000 78872 6 baseaddr_r_sync[7]
port 35 nsew default tristate
rlabel metal3 s 19520 79432 20000 79552 6 baseaddr_r_sync[8]
port 36 nsew default tristate
rlabel metal3 s 19520 67872 20000 67992 6 baseaddr_w_sync[0]
port 37 nsew default tristate
rlabel metal3 s 19520 68552 20000 68672 6 baseaddr_w_sync[1]
port 38 nsew default tristate
rlabel metal3 s 19520 69232 20000 69352 6 baseaddr_w_sync[2]
port 39 nsew default tristate
rlabel metal3 s 19520 69912 20000 70032 6 baseaddr_w_sync[3]
port 40 nsew default tristate
rlabel metal3 s 19520 70592 20000 70712 6 baseaddr_w_sync[4]
port 41 nsew default tristate
rlabel metal3 s 19520 71272 20000 71392 6 baseaddr_w_sync[5]
port 42 nsew default tristate
rlabel metal3 s 19520 71952 20000 72072 6 baseaddr_w_sync[6]
port 43 nsew default tristate
rlabel metal3 s 19520 72632 20000 72752 6 baseaddr_w_sync[7]
port 44 nsew default tristate
rlabel metal3 s 19520 73312 20000 73432 6 baseaddr_w_sync[8]
port 45 nsew default tristate
rlabel metal3 s 0 280 480 400 6 clk
port 46 nsew default input
rlabel metal3 s 0 51416 480 51536 6 conf[0]
port 47 nsew default input
rlabel metal3 s 0 52232 480 52352 6 conf[1]
port 48 nsew default input
rlabel metal3 s 0 53048 480 53168 6 conf[2]
port 49 nsew default input
rlabel metal3 s 0 26664 480 26784 6 csb
port 50 nsew default input
rlabel metal3 s 19520 65832 20000 65952 6 csb0_sync
port 51 nsew default tristate
rlabel metal3 s 19520 67192 20000 67312 6 csb1_sync
port 52 nsew default tristate
rlabel metal3 s 0 960 480 1080 6 d_fabric_in[0]
port 53 nsew default input
rlabel metal3 s 0 8984 480 9104 6 d_fabric_in[10]
port 54 nsew default input
rlabel metal3 s 0 9800 480 9920 6 d_fabric_in[11]
port 55 nsew default input
rlabel metal3 s 0 10616 480 10736 6 d_fabric_in[12]
port 56 nsew default input
rlabel metal3 s 0 11432 480 11552 6 d_fabric_in[13]
port 57 nsew default input
rlabel metal3 s 0 12248 480 12368 6 d_fabric_in[14]
port 58 nsew default input
rlabel metal3 s 0 13064 480 13184 6 d_fabric_in[15]
port 59 nsew default input
rlabel metal3 s 0 13744 480 13864 6 d_fabric_in[16]
port 60 nsew default input
rlabel metal3 s 0 14560 480 14680 6 d_fabric_in[17]
port 61 nsew default input
rlabel metal3 s 0 15376 480 15496 6 d_fabric_in[18]
port 62 nsew default input
rlabel metal3 s 0 16192 480 16312 6 d_fabric_in[19]
port 63 nsew default input
rlabel metal3 s 0 1776 480 1896 6 d_fabric_in[1]
port 64 nsew default input
rlabel metal3 s 0 17008 480 17128 6 d_fabric_in[20]
port 65 nsew default input
rlabel metal3 s 0 17824 480 17944 6 d_fabric_in[21]
port 66 nsew default input
rlabel metal3 s 0 18640 480 18760 6 d_fabric_in[22]
port 67 nsew default input
rlabel metal3 s 0 19456 480 19576 6 d_fabric_in[23]
port 68 nsew default input
rlabel metal3 s 0 20272 480 20392 6 d_fabric_in[24]
port 69 nsew default input
rlabel metal3 s 0 20952 480 21072 6 d_fabric_in[25]
port 70 nsew default input
rlabel metal3 s 0 21768 480 21888 6 d_fabric_in[26]
port 71 nsew default input
rlabel metal3 s 0 22584 480 22704 6 d_fabric_in[27]
port 72 nsew default input
rlabel metal3 s 0 23400 480 23520 6 d_fabric_in[28]
port 73 nsew default input
rlabel metal3 s 0 24216 480 24336 6 d_fabric_in[29]
port 74 nsew default input
rlabel metal3 s 0 2592 480 2712 6 d_fabric_in[2]
port 75 nsew default input
rlabel metal3 s 0 25032 480 25152 6 d_fabric_in[30]
port 76 nsew default input
rlabel metal3 s 0 25848 480 25968 6 d_fabric_in[31]
port 77 nsew default input
rlabel metal3 s 0 3408 480 3528 6 d_fabric_in[3]
port 78 nsew default input
rlabel metal3 s 0 4224 480 4344 6 d_fabric_in[4]
port 79 nsew default input
rlabel metal3 s 0 5040 480 5160 6 d_fabric_in[5]
port 80 nsew default input
rlabel metal3 s 0 5856 480 5976 6 d_fabric_in[6]
port 81 nsew default input
rlabel metal3 s 0 6672 480 6792 6 d_fabric_in[7]
port 82 nsew default input
rlabel metal3 s 0 7352 480 7472 6 d_fabric_in[8]
port 83 nsew default input
rlabel metal3 s 0 8168 480 8288 6 d_fabric_in[9]
port 84 nsew default input
rlabel metal3 s 0 54544 480 54664 6 d_fabric_out[0]
port 85 nsew default tristate
rlabel metal3 s 0 62568 480 62688 6 d_fabric_out[10]
port 86 nsew default tristate
rlabel metal3 s 0 63384 480 63504 6 d_fabric_out[11]
port 87 nsew default tristate
rlabel metal3 s 0 64200 480 64320 6 d_fabric_out[12]
port 88 nsew default tristate
rlabel metal3 s 0 65016 480 65136 6 d_fabric_out[13]
port 89 nsew default tristate
rlabel metal3 s 0 65832 480 65952 6 d_fabric_out[14]
port 90 nsew default tristate
rlabel metal3 s 0 66648 480 66768 6 d_fabric_out[15]
port 91 nsew default tristate
rlabel metal3 s 0 67328 480 67448 6 d_fabric_out[16]
port 92 nsew default tristate
rlabel metal3 s 0 68144 480 68264 6 d_fabric_out[17]
port 93 nsew default tristate
rlabel metal3 s 0 68960 480 69080 6 d_fabric_out[18]
port 94 nsew default tristate
rlabel metal3 s 0 69776 480 69896 6 d_fabric_out[19]
port 95 nsew default tristate
rlabel metal3 s 0 55360 480 55480 6 d_fabric_out[1]
port 96 nsew default tristate
rlabel metal3 s 0 70592 480 70712 6 d_fabric_out[20]
port 97 nsew default tristate
rlabel metal3 s 0 71408 480 71528 6 d_fabric_out[21]
port 98 nsew default tristate
rlabel metal3 s 0 72224 480 72344 6 d_fabric_out[22]
port 99 nsew default tristate
rlabel metal3 s 0 73040 480 73160 6 d_fabric_out[23]
port 100 nsew default tristate
rlabel metal3 s 0 73720 480 73840 6 d_fabric_out[24]
port 101 nsew default tristate
rlabel metal3 s 0 74536 480 74656 6 d_fabric_out[25]
port 102 nsew default tristate
rlabel metal3 s 0 75352 480 75472 6 d_fabric_out[26]
port 103 nsew default tristate
rlabel metal3 s 0 76168 480 76288 6 d_fabric_out[27]
port 104 nsew default tristate
rlabel metal3 s 0 76984 480 77104 6 d_fabric_out[28]
port 105 nsew default tristate
rlabel metal3 s 0 77800 480 77920 6 d_fabric_out[29]
port 106 nsew default tristate
rlabel metal3 s 0 56176 480 56296 6 d_fabric_out[2]
port 107 nsew default tristate
rlabel metal3 s 0 78616 480 78736 6 d_fabric_out[30]
port 108 nsew default tristate
rlabel metal3 s 0 79432 480 79552 6 d_fabric_out[31]
port 109 nsew default tristate
rlabel metal3 s 0 56992 480 57112 6 d_fabric_out[3]
port 110 nsew default tristate
rlabel metal3 s 0 57808 480 57928 6 d_fabric_out[4]
port 111 nsew default tristate
rlabel metal3 s 0 58624 480 58744 6 d_fabric_out[5]
port 112 nsew default tristate
rlabel metal3 s 0 59440 480 59560 6 d_fabric_out[6]
port 113 nsew default tristate
rlabel metal3 s 0 60256 480 60376 6 d_fabric_out[7]
port 114 nsew default tristate
rlabel metal3 s 0 60936 480 61056 6 d_fabric_out[8]
port 115 nsew default tristate
rlabel metal3 s 0 61752 480 61872 6 d_fabric_out[9]
port 116 nsew default tristate
rlabel metal3 s 19520 280 20000 400 6 d_sram_in[0]
port 117 nsew default tristate
rlabel metal3 s 19520 7080 20000 7200 6 d_sram_in[10]
port 118 nsew default tristate
rlabel metal3 s 19520 7760 20000 7880 6 d_sram_in[11]
port 119 nsew default tristate
rlabel metal3 s 19520 8440 20000 8560 6 d_sram_in[12]
port 120 nsew default tristate
rlabel metal3 s 19520 9120 20000 9240 6 d_sram_in[13]
port 121 nsew default tristate
rlabel metal3 s 19520 9800 20000 9920 6 d_sram_in[14]
port 122 nsew default tristate
rlabel metal3 s 19520 10480 20000 10600 6 d_sram_in[15]
port 123 nsew default tristate
rlabel metal3 s 19520 11160 20000 11280 6 d_sram_in[16]
port 124 nsew default tristate
rlabel metal3 s 19520 11840 20000 11960 6 d_sram_in[17]
port 125 nsew default tristate
rlabel metal3 s 19520 12520 20000 12640 6 d_sram_in[18]
port 126 nsew default tristate
rlabel metal3 s 19520 13200 20000 13320 6 d_sram_in[19]
port 127 nsew default tristate
rlabel metal3 s 19520 960 20000 1080 6 d_sram_in[1]
port 128 nsew default tristate
rlabel metal3 s 19520 13880 20000 14000 6 d_sram_in[20]
port 129 nsew default tristate
rlabel metal3 s 19520 14560 20000 14680 6 d_sram_in[21]
port 130 nsew default tristate
rlabel metal3 s 19520 15240 20000 15360 6 d_sram_in[22]
port 131 nsew default tristate
rlabel metal3 s 19520 15920 20000 16040 6 d_sram_in[23]
port 132 nsew default tristate
rlabel metal3 s 19520 16600 20000 16720 6 d_sram_in[24]
port 133 nsew default tristate
rlabel metal3 s 19520 17280 20000 17400 6 d_sram_in[25]
port 134 nsew default tristate
rlabel metal3 s 19520 17960 20000 18080 6 d_sram_in[26]
port 135 nsew default tristate
rlabel metal3 s 19520 18640 20000 18760 6 d_sram_in[27]
port 136 nsew default tristate
rlabel metal3 s 19520 19320 20000 19440 6 d_sram_in[28]
port 137 nsew default tristate
rlabel metal3 s 19520 20000 20000 20120 6 d_sram_in[29]
port 138 nsew default tristate
rlabel metal3 s 19520 1640 20000 1760 6 d_sram_in[2]
port 139 nsew default tristate
rlabel metal3 s 19520 20680 20000 20800 6 d_sram_in[30]
port 140 nsew default tristate
rlabel metal3 s 19520 21360 20000 21480 6 d_sram_in[31]
port 141 nsew default tristate
rlabel metal3 s 19520 2320 20000 2440 6 d_sram_in[3]
port 142 nsew default tristate
rlabel metal3 s 19520 3000 20000 3120 6 d_sram_in[4]
port 143 nsew default tristate
rlabel metal3 s 19520 3680 20000 3800 6 d_sram_in[5]
port 144 nsew default tristate
rlabel metal3 s 19520 4360 20000 4480 6 d_sram_in[6]
port 145 nsew default tristate
rlabel metal3 s 19520 5040 20000 5160 6 d_sram_in[7]
port 146 nsew default tristate
rlabel metal3 s 19520 5720 20000 5840 6 d_sram_in[8]
port 147 nsew default tristate
rlabel metal3 s 19520 6400 20000 6520 6 d_sram_in[9]
port 148 nsew default tristate
rlabel metal3 s 19520 43936 20000 44056 6 d_sram_out[0]
port 149 nsew default input
rlabel metal3 s 19520 50736 20000 50856 6 d_sram_out[10]
port 150 nsew default input
rlabel metal3 s 19520 51416 20000 51536 6 d_sram_out[11]
port 151 nsew default input
rlabel metal3 s 19520 52096 20000 52216 6 d_sram_out[12]
port 152 nsew default input
rlabel metal3 s 19520 52776 20000 52896 6 d_sram_out[13]
port 153 nsew default input
rlabel metal3 s 19520 53592 20000 53712 6 d_sram_out[14]
port 154 nsew default input
rlabel metal3 s 19520 54272 20000 54392 6 d_sram_out[15]
port 155 nsew default input
rlabel metal3 s 19520 54952 20000 55072 6 d_sram_out[16]
port 156 nsew default input
rlabel metal3 s 19520 55632 20000 55752 6 d_sram_out[17]
port 157 nsew default input
rlabel metal3 s 19520 56312 20000 56432 6 d_sram_out[18]
port 158 nsew default input
rlabel metal3 s 19520 56992 20000 57112 6 d_sram_out[19]
port 159 nsew default input
rlabel metal3 s 19520 44616 20000 44736 6 d_sram_out[1]
port 160 nsew default input
rlabel metal3 s 19520 57672 20000 57792 6 d_sram_out[20]
port 161 nsew default input
rlabel metal3 s 19520 58352 20000 58472 6 d_sram_out[21]
port 162 nsew default input
rlabel metal3 s 19520 59032 20000 59152 6 d_sram_out[22]
port 163 nsew default input
rlabel metal3 s 19520 59712 20000 59832 6 d_sram_out[23]
port 164 nsew default input
rlabel metal3 s 19520 60392 20000 60512 6 d_sram_out[24]
port 165 nsew default input
rlabel metal3 s 19520 61072 20000 61192 6 d_sram_out[25]
port 166 nsew default input
rlabel metal3 s 19520 61752 20000 61872 6 d_sram_out[26]
port 167 nsew default input
rlabel metal3 s 19520 62432 20000 62552 6 d_sram_out[27]
port 168 nsew default input
rlabel metal3 s 19520 63112 20000 63232 6 d_sram_out[28]
port 169 nsew default input
rlabel metal3 s 19520 63792 20000 63912 6 d_sram_out[29]
port 170 nsew default input
rlabel metal3 s 19520 45296 20000 45416 6 d_sram_out[2]
port 171 nsew default input
rlabel metal3 s 19520 64472 20000 64592 6 d_sram_out[30]
port 172 nsew default input
rlabel metal3 s 19520 65152 20000 65272 6 d_sram_out[31]
port 173 nsew default input
rlabel metal3 s 19520 45976 20000 46096 6 d_sram_out[3]
port 174 nsew default input
rlabel metal3 s 19520 46656 20000 46776 6 d_sram_out[4]
port 175 nsew default input
rlabel metal3 s 19520 47336 20000 47456 6 d_sram_out[5]
port 176 nsew default input
rlabel metal3 s 19520 48016 20000 48136 6 d_sram_out[6]
port 177 nsew default input
rlabel metal3 s 19520 48696 20000 48816 6 d_sram_out[7]
port 178 nsew default input
rlabel metal3 s 19520 49376 20000 49496 6 d_sram_out[8]
port 179 nsew default input
rlabel metal3 s 19520 50056 20000 50176 6 d_sram_out[9]
port 180 nsew default input
rlabel metal3 s 0 53728 480 53848 6 out_reg
port 181 nsew default input
rlabel metal3 s 0 28160 480 28280 6 reb
port 182 nsew default input
rlabel metal3 s 19520 22040 20000 22160 6 w_mask[0]
port 183 nsew default tristate
rlabel metal3 s 19520 28976 20000 29096 6 w_mask[10]
port 184 nsew default tristate
rlabel metal3 s 19520 29656 20000 29776 6 w_mask[11]
port 185 nsew default tristate
rlabel metal3 s 19520 30336 20000 30456 6 w_mask[12]
port 186 nsew default tristate
rlabel metal3 s 19520 31016 20000 31136 6 w_mask[13]
port 187 nsew default tristate
rlabel metal3 s 19520 31696 20000 31816 6 w_mask[14]
port 188 nsew default tristate
rlabel metal3 s 19520 32376 20000 32496 6 w_mask[15]
port 189 nsew default tristate
rlabel metal3 s 19520 33056 20000 33176 6 w_mask[16]
port 190 nsew default tristate
rlabel metal3 s 19520 33736 20000 33856 6 w_mask[17]
port 191 nsew default tristate
rlabel metal3 s 19520 34416 20000 34536 6 w_mask[18]
port 192 nsew default tristate
rlabel metal3 s 19520 35096 20000 35216 6 w_mask[19]
port 193 nsew default tristate
rlabel metal3 s 19520 22720 20000 22840 6 w_mask[1]
port 194 nsew default tristate
rlabel metal3 s 19520 35776 20000 35896 6 w_mask[20]
port 195 nsew default tristate
rlabel metal3 s 19520 36456 20000 36576 6 w_mask[21]
port 196 nsew default tristate
rlabel metal3 s 19520 37136 20000 37256 6 w_mask[22]
port 197 nsew default tristate
rlabel metal3 s 19520 37816 20000 37936 6 w_mask[23]
port 198 nsew default tristate
rlabel metal3 s 19520 38496 20000 38616 6 w_mask[24]
port 199 nsew default tristate
rlabel metal3 s 19520 39176 20000 39296 6 w_mask[25]
port 200 nsew default tristate
rlabel metal3 s 19520 39856 20000 39976 6 w_mask[26]
port 201 nsew default tristate
rlabel metal3 s 19520 40536 20000 40656 6 w_mask[27]
port 202 nsew default tristate
rlabel metal3 s 19520 41216 20000 41336 6 w_mask[28]
port 203 nsew default tristate
rlabel metal3 s 19520 41896 20000 42016 6 w_mask[29]
port 204 nsew default tristate
rlabel metal3 s 19520 23400 20000 23520 6 w_mask[2]
port 205 nsew default tristate
rlabel metal3 s 19520 42576 20000 42696 6 w_mask[30]
port 206 nsew default tristate
rlabel metal3 s 19520 43256 20000 43376 6 w_mask[31]
port 207 nsew default tristate
rlabel metal3 s 19520 24080 20000 24200 6 w_mask[3]
port 208 nsew default tristate
rlabel metal3 s 19520 24760 20000 24880 6 w_mask[4]
port 209 nsew default tristate
rlabel metal3 s 19520 25440 20000 25560 6 w_mask[5]
port 210 nsew default tristate
rlabel metal3 s 19520 26120 20000 26240 6 w_mask[6]
port 211 nsew default tristate
rlabel metal3 s 19520 26936 20000 27056 6 w_mask[7]
port 212 nsew default tristate
rlabel metal3 s 19520 27616 20000 27736 6 w_mask[8]
port 213 nsew default tristate
rlabel metal3 s 19520 28296 20000 28416 6 w_mask[9]
port 214 nsew default tristate
rlabel metal3 s 0 27344 480 27464 6 web
port 215 nsew default input
rlabel metal3 s 19520 66512 20000 66632 6 web0_sync
port 216 nsew default tristate
rlabel metal5 s 1104 15301 18860 15621 6 VPWR
port 217 nsew default input
rlabel metal5 s 1104 28635 18860 28955 6 VGND
port 218 nsew default input
<< end >>
