VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sram_ifc
  CLASS BLOCK ;
  FOREIGN sram_ifc ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 400.000 ;
  PIN addr_r[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 17.040 200.000 17.640 ;
    END
  END addr_r[0]
  PIN addr_r[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 357.040 200.000 357.640 ;
    END
  END addr_r[10]
  PIN addr_r[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 176.840 200.000 177.440 ;
    END
  END addr_r[11]
  PIN addr_r[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.090 396.000 92.370 400.000 ;
    END
  END addr_r[12]
  PIN addr_r[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 306.040 200.000 306.640 ;
    END
  END addr_r[13]
  PIN addr_r[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END addr_r[1]
  PIN addr_r[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 82.890 396.000 83.170 400.000 ;
    END
  END addr_r[2]
  PIN addr_r[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END addr_r[3]
  PIN addr_r[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END addr_r[4]
  PIN addr_r[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END addr_r[5]
  PIN addr_r[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END addr_r[6]
  PIN addr_r[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END addr_r[7]
  PIN addr_r[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END addr_r[8]
  PIN addr_r[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END addr_r[9]
  PIN addr_w[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END addr_w[0]
  PIN addr_w[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END addr_w[10]
  PIN addr_w[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END addr_w[11]
  PIN addr_w[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 3.440 200.000 4.040 ;
    END
  END addr_w[12]
  PIN addr_w[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END addr_w[13]
  PIN addr_w[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END addr_w[1]
  PIN addr_w[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 146.240 200.000 146.840 ;
    END
  END addr_w[2]
  PIN addr_w[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END addr_w[3]
  PIN addr_w[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 44.240 200.000 44.840 ;
    END
  END addr_w[4]
  PIN addr_w[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END addr_w[5]
  PIN addr_w[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END addr_w[6]
  PIN addr_w[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END addr_w[7]
  PIN addr_w[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END addr_w[8]
  PIN addr_w[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END addr_w[9]
  PIN baseaddr_r_sync[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 227.840 200.000 228.440 ;
    END
  END baseaddr_r_sync[0]
  PIN baseaddr_r_sync[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.090 396.000 115.370 400.000 ;
    END
  END baseaddr_r_sync[1]
  PIN baseaddr_r_sync[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 74.840 200.000 75.440 ;
    END
  END baseaddr_r_sync[2]
  PIN baseaddr_r_sync[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END baseaddr_r_sync[3]
  PIN baseaddr_r_sync[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 125.840 200.000 126.440 ;
    END
  END baseaddr_r_sync[4]
  PIN baseaddr_r_sync[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END baseaddr_r_sync[5]
  PIN baseaddr_r_sync[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 102.040 200.000 102.640 ;
    END
  END baseaddr_r_sync[6]
  PIN baseaddr_r_sync[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END baseaddr_r_sync[7]
  PIN baseaddr_r_sync[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.990 396.000 122.270 400.000 ;
    END
  END baseaddr_r_sync[8]
  PIN baseaddr_w_sync[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.490 396.000 18.770 400.000 ;
    END
  END baseaddr_w_sync[0]
  PIN baseaddr_w_sync[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 363.840 200.000 364.440 ;
    END
  END baseaddr_w_sync[1]
  PIN baseaddr_w_sync[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END baseaddr_w_sync[2]
  PIN baseaddr_w_sync[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END baseaddr_w_sync[3]
  PIN baseaddr_w_sync[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.890 396.000 37.170 400.000 ;
    END
  END baseaddr_w_sync[4]
  PIN baseaddr_w_sync[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 161.090 396.000 161.370 400.000 ;
    END
  END baseaddr_w_sync[5]
  PIN baseaddr_w_sync[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END baseaddr_w_sync[6]
  PIN baseaddr_w_sync[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END baseaddr_w_sync[7]
  PIN baseaddr_w_sync[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 23.840 200.000 24.440 ;
    END
  END baseaddr_w_sync[8]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END clk
  PIN conf[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.490 396.000 110.770 400.000 ;
    END
  END conf[0]
  PIN conf[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END conf[1]
  PIN conf[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 210.840 200.000 211.440 ;
    END
  END conf[2]
  PIN csb
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 61.240 200.000 61.840 ;
    END
  END csb
  PIN csb0_sync
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 184.090 396.000 184.370 400.000 ;
    END
  END csb0_sync
  PIN csb1_sync
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END csb1_sync
  PIN d_fabric_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 30.640 200.000 31.240 ;
    END
  END d_fabric_in[0]
  PIN d_fabric_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END d_fabric_in[10]
  PIN d_fabric_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.490 396.000 87.770 400.000 ;
    END
  END d_fabric_in[11]
  PIN d_fabric_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 391.040 200.000 391.640 ;
    END
  END d_fabric_in[12]
  PIN d_fabric_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END d_fabric_in[13]
  PIN d_fabric_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END d_fabric_in[14]
  PIN d_fabric_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END d_fabric_in[15]
  PIN d_fabric_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.590 396.000 126.870 400.000 ;
    END
  END d_fabric_in[16]
  PIN d_fabric_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 384.240 200.000 384.840 ;
    END
  END d_fabric_in[17]
  PIN d_fabric_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 326.440 200.000 327.040 ;
    END
  END d_fabric_in[18]
  PIN d_fabric_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 188.690 396.000 188.970 400.000 ;
    END
  END d_fabric_in[19]
  PIN d_fabric_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END d_fabric_in[1]
  PIN d_fabric_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END d_fabric_in[20]
  PIN d_fabric_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 312.840 200.000 313.440 ;
    END
  END d_fabric_in[21]
  PIN d_fabric_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 37.440 200.000 38.040 ;
    END
  END d_fabric_in[22]
  PIN d_fabric_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 268.640 200.000 269.240 ;
    END
  END d_fabric_in[23]
  PIN d_fabric_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END d_fabric_in[24]
  PIN d_fabric_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 144.990 396.000 145.270 400.000 ;
    END
  END d_fabric_in[25]
  PIN d_fabric_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 396.000 2.670 400.000 ;
    END
  END d_fabric_in[26]
  PIN d_fabric_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END d_fabric_in[27]
  PIN d_fabric_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 248.240 200.000 248.840 ;
    END
  END d_fabric_in[28]
  PIN d_fabric_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 285.640 200.000 286.240 ;
    END
  END d_fabric_in[29]
  PIN d_fabric_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END d_fabric_in[2]
  PIN d_fabric_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 68.040 200.000 68.640 ;
    END
  END d_fabric_in[30]
  PIN d_fabric_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END d_fabric_in[31]
  PIN d_fabric_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END d_fabric_in[3]
  PIN d_fabric_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 131.190 396.000 131.470 400.000 ;
    END
  END d_fabric_in[4]
  PIN d_fabric_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.890 396.000 106.170 400.000 ;
    END
  END d_fabric_in[5]
  PIN d_fabric_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END d_fabric_in[6]
  PIN d_fabric_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 397.840 200.000 398.440 ;
    END
  END d_fabric_in[7]
  PIN d_fabric_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END d_fabric_in[8]
  PIN d_fabric_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END d_fabric_in[9]
  PIN d_fabric_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END d_fabric_out[0]
  PIN d_fabric_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END d_fabric_out[10]
  PIN d_fabric_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END d_fabric_out[11]
  PIN d_fabric_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 343.440 200.000 344.040 ;
    END
  END d_fabric_out[12]
  PIN d_fabric_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END d_fabric_out[13]
  PIN d_fabric_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END d_fabric_out[14]
  PIN d_fabric_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.490 396.000 41.770 400.000 ;
    END
  END d_fabric_out[15]
  PIN d_fabric_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 282.240 200.000 282.840 ;
    END
  END d_fabric_out[16]
  PIN d_fabric_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 396.000 101.570 400.000 ;
    END
  END d_fabric_out[17]
  PIN d_fabric_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END d_fabric_out[18]
  PIN d_fabric_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 132.640 200.000 133.240 ;
    END
  END d_fabric_out[19]
  PIN d_fabric_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END d_fabric_out[1]
  PIN d_fabric_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END d_fabric_out[20]
  PIN d_fabric_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END d_fabric_out[21]
  PIN d_fabric_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END d_fabric_out[22]
  PIN d_fabric_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END d_fabric_out[23]
  PIN d_fabric_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 217.640 200.000 218.240 ;
    END
  END d_fabric_out[24]
  PIN d_fabric_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END d_fabric_out[25]
  PIN d_fabric_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END d_fabric_out[26]
  PIN d_fabric_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END d_fabric_out[27]
  PIN d_fabric_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.790 396.000 44.070 400.000 ;
    END
  END d_fabric_out[28]
  PIN d_fabric_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END d_fabric_out[29]
  PIN d_fabric_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 23.090 396.000 23.370 400.000 ;
    END
  END d_fabric_out[2]
  PIN d_fabric_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 62.190 396.000 62.470 400.000 ;
    END
  END d_fabric_out[30]
  PIN d_fabric_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 197.890 396.000 198.170 400.000 ;
    END
  END d_fabric_out[31]
  PIN d_fabric_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.590 396.000 149.870 400.000 ;
    END
  END d_fabric_out[3]
  PIN d_fabric_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END d_fabric_out[4]
  PIN d_fabric_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 340.040 200.000 340.640 ;
    END
  END d_fabric_out[5]
  PIN d_fabric_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 319.640 200.000 320.240 ;
    END
  END d_fabric_out[6]
  PIN d_fabric_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 255.040 200.000 255.640 ;
    END
  END d_fabric_out[7]
  PIN d_fabric_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END d_fabric_out[8]
  PIN d_fabric_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END d_fabric_out[9]
  PIN d_sram_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END d_sram_in[0]
  PIN d_sram_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 197.240 200.000 197.840 ;
    END
  END d_sram_in[10]
  PIN d_sram_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 190.440 200.000 191.040 ;
    END
  END d_sram_in[11]
  PIN d_sram_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 66.790 396.000 67.070 400.000 ;
    END
  END d_sram_in[12]
  PIN d_sram_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END d_sram_in[13]
  PIN d_sram_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END d_sram_in[14]
  PIN d_sram_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END d_sram_in[15]
  PIN d_sram_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 166.640 200.000 167.240 ;
    END
  END d_sram_in[16]
  PIN d_sram_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 112.240 200.000 112.840 ;
    END
  END d_sram_in[17]
  PIN d_sram_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END d_sram_in[18]
  PIN d_sram_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 370.640 200.000 371.240 ;
    END
  END d_sram_in[19]
  PIN d_sram_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.690 396.000 27.970 400.000 ;
    END
  END d_sram_in[1]
  PIN d_sram_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END d_sram_in[20]
  PIN d_sram_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 299.240 200.000 299.840 ;
    END
  END d_sram_in[21]
  PIN d_sram_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END d_sram_in[22]
  PIN d_sram_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END d_sram_in[23]
  PIN d_sram_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 81.640 200.000 82.240 ;
    END
  END d_sram_in[24]
  PIN d_sram_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 174.890 396.000 175.170 400.000 ;
    END
  END d_sram_in[25]
  PIN d_sram_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END d_sram_in[26]
  PIN d_sram_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.890 396.000 14.170 400.000 ;
    END
  END d_sram_in[27]
  PIN d_sram_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END d_sram_in[28]
  PIN d_sram_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 88.440 200.000 89.040 ;
    END
  END d_sram_in[29]
  PIN d_sram_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END d_sram_in[2]
  PIN d_sram_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.390 396.000 71.670 400.000 ;
    END
  END d_sram_in[30]
  PIN d_sram_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 153.040 200.000 153.640 ;
    END
  END d_sram_in[31]
  PIN d_sram_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END d_sram_in[3]
  PIN d_sram_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 48.390 396.000 48.670 400.000 ;
    END
  END d_sram_in[4]
  PIN d_sram_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 183.640 200.000 184.240 ;
    END
  END d_sram_in[5]
  PIN d_sram_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END d_sram_in[6]
  PIN d_sram_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END d_sram_in[7]
  PIN d_sram_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END d_sram_in[8]
  PIN d_sram_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 204.040 200.000 204.640 ;
    END
  END d_sram_in[9]
  PIN d_sram_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END d_sram_out[0]
  PIN d_sram_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END d_sram_out[10]
  PIN d_sram_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END d_sram_out[11]
  PIN d_sram_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END d_sram_out[12]
  PIN d_sram_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.590 396.000 80.870 400.000 ;
    END
  END d_sram_out[13]
  PIN d_sram_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END d_sram_out[14]
  PIN d_sram_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 165.690 396.000 165.970 400.000 ;
    END
  END d_sram_out[15]
  PIN d_sram_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END d_sram_out[16]
  PIN d_sram_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 377.440 200.000 378.040 ;
    END
  END d_sram_out[17]
  PIN d_sram_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END d_sram_out[18]
  PIN d_sram_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 154.190 396.000 154.470 400.000 ;
    END
  END d_sram_out[19]
  PIN d_sram_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 292.440 200.000 293.040 ;
    END
  END d_sram_out[1]
  PIN d_sram_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 108.840 200.000 109.440 ;
    END
  END d_sram_out[20]
  PIN d_sram_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END d_sram_out[21]
  PIN d_sram_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END d_sram_out[22]
  PIN d_sram_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 158.790 396.000 159.070 400.000 ;
    END
  END d_sram_out[23]
  PIN d_sram_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 51.040 200.000 51.640 ;
    END
  END d_sram_out[24]
  PIN d_sram_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END d_sram_out[25]
  PIN d_sram_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.290 396.000 170.570 400.000 ;
    END
  END d_sram_out[26]
  PIN d_sram_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 95.240 200.000 95.840 ;
    END
  END d_sram_out[27]
  PIN d_sram_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END d_sram_out[28]
  PIN d_sram_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END d_sram_out[29]
  PIN d_sram_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 350.240 200.000 350.840 ;
    END
  END d_sram_out[2]
  PIN d_sram_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END d_sram_out[30]
  PIN d_sram_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END d_sram_out[31]
  PIN d_sram_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 170.040 200.000 170.640 ;
    END
  END d_sram_out[3]
  PIN d_sram_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END d_sram_out[4]
  PIN d_sram_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END d_sram_out[5]
  PIN d_sram_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 196.000 261.840 200.000 262.440 ;
    END
  END d_sram_out[6]
  PIN d_sram_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END d_sram_out[7]
  PIN d_sram_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END d_sram_out[8]
  PIN d_sram_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END d_sram_out[9]
  PIN out_reg
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.790 396.000 136.070 400.000 ;
    END
  END out_reg
  PIN reb
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END reb
  PIN w_mask[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 54.440 200.000 55.040 ;
    END
  END w_mask[0]
  PIN w_mask[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 57.590 396.000 57.870 400.000 ;
    END
  END w_mask[10]
  PIN w_mask[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 333.240 200.000 333.840 ;
    END
  END w_mask[11]
  PIN w_mask[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END w_mask[12]
  PIN w_mask[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END w_mask[13]
  PIN w_mask[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END w_mask[14]
  PIN w_mask[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END w_mask[15]
  PIN w_mask[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 140.390 396.000 140.670 400.000 ;
    END
  END w_mask[16]
  PIN w_mask[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 193.290 396.000 193.570 400.000 ;
    END
  END w_mask[17]
  PIN w_mask[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 275.440 200.000 276.040 ;
    END
  END w_mask[18]
  PIN w_mask[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END w_mask[19]
  PIN w_mask[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 10.240 200.000 10.840 ;
    END
  END w_mask[1]
  PIN w_mask[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 9.290 396.000 9.570 400.000 ;
    END
  END w_mask[20]
  PIN w_mask[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END w_mask[21]
  PIN w_mask[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 119.690 396.000 119.970 400.000 ;
    END
  END w_mask[22]
  PIN w_mask[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END w_mask[23]
  PIN w_mask[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END w_mask[24]
  PIN w_mask[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END w_mask[25]
  PIN w_mask[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 96.690 396.000 96.970 400.000 ;
    END
  END w_mask[26]
  PIN w_mask[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4.690 396.000 4.970 400.000 ;
    END
  END w_mask[27]
  PIN w_mask[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.990 396.000 76.270 400.000 ;
    END
  END w_mask[28]
  PIN w_mask[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 179.490 396.000 179.770 400.000 ;
    END
  END w_mask[29]
  PIN w_mask[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 32.290 396.000 32.570 400.000 ;
    END
  END w_mask[2]
  PIN w_mask[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END w_mask[30]
  PIN w_mask[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END w_mask[31]
  PIN w_mask[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 241.440 200.000 242.040 ;
    END
  END w_mask[3]
  PIN w_mask[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 224.440 200.000 225.040 ;
    END
  END w_mask[4]
  PIN w_mask[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 52.990 396.000 53.270 400.000 ;
    END
  END w_mask[5]
  PIN w_mask[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 159.840 200.000 160.440 ;
    END
  END w_mask[6]
  PIN w_mask[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 119.040 200.000 119.640 ;
    END
  END w_mask[7]
  PIN w_mask[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 234.640 200.000 235.240 ;
    END
  END w_mask[8]
  PIN w_mask[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 196.000 139.440 200.000 140.040 ;
    END
  END w_mask[9]
  PIN web
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END web
  PIN web0_sync
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END web0_sync
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 194.120 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 194.120 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 389.045 ;
      LAYER met1 ;
        RECT 0.070 4.460 198.190 389.600 ;
      LAYER met2 ;
        RECT 0.100 395.720 2.110 398.325 ;
        RECT 2.950 395.720 4.410 398.325 ;
        RECT 5.250 395.720 9.010 398.325 ;
        RECT 9.850 395.720 13.610 398.325 ;
        RECT 14.450 395.720 18.210 398.325 ;
        RECT 19.050 395.720 22.810 398.325 ;
        RECT 23.650 395.720 27.410 398.325 ;
        RECT 28.250 395.720 32.010 398.325 ;
        RECT 32.850 395.720 36.610 398.325 ;
        RECT 37.450 395.720 41.210 398.325 ;
        RECT 42.050 395.720 43.510 398.325 ;
        RECT 44.350 395.720 48.110 398.325 ;
        RECT 48.950 395.720 52.710 398.325 ;
        RECT 53.550 395.720 57.310 398.325 ;
        RECT 58.150 395.720 61.910 398.325 ;
        RECT 62.750 395.720 66.510 398.325 ;
        RECT 67.350 395.720 71.110 398.325 ;
        RECT 71.950 395.720 75.710 398.325 ;
        RECT 76.550 395.720 80.310 398.325 ;
        RECT 81.150 395.720 82.610 398.325 ;
        RECT 83.450 395.720 87.210 398.325 ;
        RECT 88.050 395.720 91.810 398.325 ;
        RECT 92.650 395.720 96.410 398.325 ;
        RECT 97.250 395.720 101.010 398.325 ;
        RECT 101.850 395.720 105.610 398.325 ;
        RECT 106.450 395.720 110.210 398.325 ;
        RECT 111.050 395.720 114.810 398.325 ;
        RECT 115.650 395.720 119.410 398.325 ;
        RECT 120.250 395.720 121.710 398.325 ;
        RECT 122.550 395.720 126.310 398.325 ;
        RECT 127.150 395.720 130.910 398.325 ;
        RECT 131.750 395.720 135.510 398.325 ;
        RECT 136.350 395.720 140.110 398.325 ;
        RECT 140.950 395.720 144.710 398.325 ;
        RECT 145.550 395.720 149.310 398.325 ;
        RECT 150.150 395.720 153.910 398.325 ;
        RECT 154.750 395.720 158.510 398.325 ;
        RECT 159.350 395.720 160.810 398.325 ;
        RECT 161.650 395.720 165.410 398.325 ;
        RECT 166.250 395.720 170.010 398.325 ;
        RECT 170.850 395.720 174.610 398.325 ;
        RECT 175.450 395.720 179.210 398.325 ;
        RECT 180.050 395.720 183.810 398.325 ;
        RECT 184.650 395.720 188.410 398.325 ;
        RECT 189.250 395.720 193.010 398.325 ;
        RECT 193.850 395.720 197.610 398.325 ;
        RECT 0.100 4.280 198.170 395.720 ;
        RECT 0.650 0.835 2.110 4.280 ;
        RECT 2.950 0.835 6.710 4.280 ;
        RECT 7.550 0.835 11.310 4.280 ;
        RECT 12.150 0.835 15.910 4.280 ;
        RECT 16.750 0.835 20.510 4.280 ;
        RECT 21.350 0.835 25.110 4.280 ;
        RECT 25.950 0.835 29.710 4.280 ;
        RECT 30.550 0.835 34.310 4.280 ;
        RECT 35.150 0.835 38.910 4.280 ;
        RECT 39.750 0.835 41.210 4.280 ;
        RECT 42.050 0.835 45.810 4.280 ;
        RECT 46.650 0.835 50.410 4.280 ;
        RECT 51.250 0.835 55.010 4.280 ;
        RECT 55.850 0.835 59.610 4.280 ;
        RECT 60.450 0.835 64.210 4.280 ;
        RECT 65.050 0.835 68.810 4.280 ;
        RECT 69.650 0.835 73.410 4.280 ;
        RECT 74.250 0.835 78.010 4.280 ;
        RECT 78.850 0.835 80.310 4.280 ;
        RECT 81.150 0.835 84.910 4.280 ;
        RECT 85.750 0.835 89.510 4.280 ;
        RECT 90.350 0.835 94.110 4.280 ;
        RECT 94.950 0.835 98.710 4.280 ;
        RECT 99.550 0.835 103.310 4.280 ;
        RECT 104.150 0.835 107.910 4.280 ;
        RECT 108.750 0.835 112.510 4.280 ;
        RECT 113.350 0.835 117.110 4.280 ;
        RECT 117.950 0.835 119.410 4.280 ;
        RECT 120.250 0.835 124.010 4.280 ;
        RECT 124.850 0.835 128.610 4.280 ;
        RECT 129.450 0.835 133.210 4.280 ;
        RECT 134.050 0.835 137.810 4.280 ;
        RECT 138.650 0.835 142.410 4.280 ;
        RECT 143.250 0.835 147.010 4.280 ;
        RECT 147.850 0.835 151.610 4.280 ;
        RECT 152.450 0.835 156.210 4.280 ;
        RECT 157.050 0.835 158.510 4.280 ;
        RECT 159.350 0.835 163.110 4.280 ;
        RECT 163.950 0.835 167.710 4.280 ;
        RECT 168.550 0.835 172.310 4.280 ;
        RECT 173.150 0.835 176.910 4.280 ;
        RECT 177.750 0.835 181.510 4.280 ;
        RECT 182.350 0.835 186.110 4.280 ;
        RECT 186.950 0.835 190.710 4.280 ;
        RECT 191.550 0.835 195.310 4.280 ;
        RECT 196.150 0.835 197.610 4.280 ;
      LAYER met3 ;
        RECT 4.400 397.440 195.600 398.305 ;
        RECT 0.525 392.040 198.195 397.440 ;
        RECT 4.400 390.640 195.600 392.040 ;
        RECT 0.525 385.240 198.195 390.640 ;
        RECT 4.400 383.840 195.600 385.240 ;
        RECT 0.525 378.440 198.195 383.840 ;
        RECT 4.400 377.040 195.600 378.440 ;
        RECT 0.525 371.640 198.195 377.040 ;
        RECT 4.400 370.240 195.600 371.640 ;
        RECT 0.525 364.840 198.195 370.240 ;
        RECT 4.400 363.440 195.600 364.840 ;
        RECT 0.525 358.040 198.195 363.440 ;
        RECT 4.400 356.640 195.600 358.040 ;
        RECT 0.525 351.240 198.195 356.640 ;
        RECT 4.400 349.840 195.600 351.240 ;
        RECT 0.525 347.840 198.195 349.840 ;
        RECT 4.400 346.440 198.195 347.840 ;
        RECT 0.525 344.440 198.195 346.440 ;
        RECT 0.525 343.040 195.600 344.440 ;
        RECT 0.525 341.040 198.195 343.040 ;
        RECT 4.400 339.640 195.600 341.040 ;
        RECT 0.525 334.240 198.195 339.640 ;
        RECT 4.400 332.840 195.600 334.240 ;
        RECT 0.525 327.440 198.195 332.840 ;
        RECT 4.400 326.040 195.600 327.440 ;
        RECT 0.525 320.640 198.195 326.040 ;
        RECT 4.400 319.240 195.600 320.640 ;
        RECT 0.525 313.840 198.195 319.240 ;
        RECT 4.400 312.440 195.600 313.840 ;
        RECT 0.525 307.040 198.195 312.440 ;
        RECT 4.400 305.640 195.600 307.040 ;
        RECT 0.525 300.240 198.195 305.640 ;
        RECT 4.400 298.840 195.600 300.240 ;
        RECT 0.525 293.440 198.195 298.840 ;
        RECT 4.400 292.040 195.600 293.440 ;
        RECT 0.525 290.040 198.195 292.040 ;
        RECT 4.400 288.640 198.195 290.040 ;
        RECT 0.525 286.640 198.195 288.640 ;
        RECT 0.525 285.240 195.600 286.640 ;
        RECT 0.525 283.240 198.195 285.240 ;
        RECT 4.400 281.840 195.600 283.240 ;
        RECT 0.525 276.440 198.195 281.840 ;
        RECT 4.400 275.040 195.600 276.440 ;
        RECT 0.525 269.640 198.195 275.040 ;
        RECT 4.400 268.240 195.600 269.640 ;
        RECT 0.525 262.840 198.195 268.240 ;
        RECT 4.400 261.440 195.600 262.840 ;
        RECT 0.525 256.040 198.195 261.440 ;
        RECT 4.400 254.640 195.600 256.040 ;
        RECT 0.525 249.240 198.195 254.640 ;
        RECT 4.400 247.840 195.600 249.240 ;
        RECT 0.525 242.440 198.195 247.840 ;
        RECT 4.400 241.040 195.600 242.440 ;
        RECT 0.525 235.640 198.195 241.040 ;
        RECT 4.400 234.240 195.600 235.640 ;
        RECT 0.525 232.240 198.195 234.240 ;
        RECT 4.400 230.840 198.195 232.240 ;
        RECT 0.525 228.840 198.195 230.840 ;
        RECT 0.525 227.440 195.600 228.840 ;
        RECT 0.525 225.440 198.195 227.440 ;
        RECT 4.400 224.040 195.600 225.440 ;
        RECT 0.525 218.640 198.195 224.040 ;
        RECT 4.400 217.240 195.600 218.640 ;
        RECT 0.525 211.840 198.195 217.240 ;
        RECT 4.400 210.440 195.600 211.840 ;
        RECT 0.525 205.040 198.195 210.440 ;
        RECT 4.400 203.640 195.600 205.040 ;
        RECT 0.525 198.240 198.195 203.640 ;
        RECT 4.400 196.840 195.600 198.240 ;
        RECT 0.525 191.440 198.195 196.840 ;
        RECT 4.400 190.040 195.600 191.440 ;
        RECT 0.525 184.640 198.195 190.040 ;
        RECT 4.400 183.240 195.600 184.640 ;
        RECT 0.525 177.840 198.195 183.240 ;
        RECT 4.400 176.440 195.600 177.840 ;
        RECT 0.525 174.440 198.195 176.440 ;
        RECT 4.400 173.040 198.195 174.440 ;
        RECT 0.525 171.040 198.195 173.040 ;
        RECT 0.525 169.640 195.600 171.040 ;
        RECT 0.525 167.640 198.195 169.640 ;
        RECT 4.400 166.240 195.600 167.640 ;
        RECT 0.525 160.840 198.195 166.240 ;
        RECT 4.400 159.440 195.600 160.840 ;
        RECT 0.525 154.040 198.195 159.440 ;
        RECT 4.400 152.640 195.600 154.040 ;
        RECT 0.525 147.240 198.195 152.640 ;
        RECT 4.400 145.840 195.600 147.240 ;
        RECT 0.525 140.440 198.195 145.840 ;
        RECT 4.400 139.040 195.600 140.440 ;
        RECT 0.525 133.640 198.195 139.040 ;
        RECT 4.400 132.240 195.600 133.640 ;
        RECT 0.525 126.840 198.195 132.240 ;
        RECT 4.400 125.440 195.600 126.840 ;
        RECT 0.525 120.040 198.195 125.440 ;
        RECT 4.400 118.640 195.600 120.040 ;
        RECT 0.525 116.640 198.195 118.640 ;
        RECT 4.400 115.240 198.195 116.640 ;
        RECT 0.525 113.240 198.195 115.240 ;
        RECT 0.525 111.840 195.600 113.240 ;
        RECT 0.525 109.840 198.195 111.840 ;
        RECT 4.400 108.440 195.600 109.840 ;
        RECT 0.525 103.040 198.195 108.440 ;
        RECT 4.400 101.640 195.600 103.040 ;
        RECT 0.525 96.240 198.195 101.640 ;
        RECT 4.400 94.840 195.600 96.240 ;
        RECT 0.525 89.440 198.195 94.840 ;
        RECT 4.400 88.040 195.600 89.440 ;
        RECT 0.525 82.640 198.195 88.040 ;
        RECT 4.400 81.240 195.600 82.640 ;
        RECT 0.525 75.840 198.195 81.240 ;
        RECT 4.400 74.440 195.600 75.840 ;
        RECT 0.525 69.040 198.195 74.440 ;
        RECT 4.400 67.640 195.600 69.040 ;
        RECT 0.525 62.240 198.195 67.640 ;
        RECT 4.400 60.840 195.600 62.240 ;
        RECT 0.525 58.840 198.195 60.840 ;
        RECT 4.400 57.440 198.195 58.840 ;
        RECT 0.525 55.440 198.195 57.440 ;
        RECT 0.525 54.040 195.600 55.440 ;
        RECT 0.525 52.040 198.195 54.040 ;
        RECT 4.400 50.640 195.600 52.040 ;
        RECT 0.525 45.240 198.195 50.640 ;
        RECT 4.400 43.840 195.600 45.240 ;
        RECT 0.525 38.440 198.195 43.840 ;
        RECT 4.400 37.040 195.600 38.440 ;
        RECT 0.525 31.640 198.195 37.040 ;
        RECT 4.400 30.240 195.600 31.640 ;
        RECT 0.525 24.840 198.195 30.240 ;
        RECT 4.400 23.440 195.600 24.840 ;
        RECT 0.525 18.040 198.195 23.440 ;
        RECT 4.400 16.640 195.600 18.040 ;
        RECT 0.525 11.240 198.195 16.640 ;
        RECT 4.400 9.840 195.600 11.240 ;
        RECT 0.525 4.440 198.195 9.840 ;
        RECT 4.400 3.040 195.600 4.440 ;
        RECT 0.525 0.855 198.195 3.040 ;
      LAYER met4 ;
        RECT 21.040 4.255 178.610 389.200 ;
      LAYER met5 ;
        RECT 5.520 106.300 194.120 334.450 ;
  END
END sram_ifc
END LIBRARY

