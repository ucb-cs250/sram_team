* NGSPICE file created from sram_ifc.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 D Q CLK VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D Y VGND VPWR
.ends

.subckt sram_ifc addr_r[0] addr_r[10] addr_r[11] addr_r[12] addr_r[13] addr_r[1] addr_r[2]
+ addr_r[3] addr_r[4] addr_r[5] addr_r[6] addr_r[7] addr_r[8] addr_r[9] addr_w[0]
+ addr_w[10] addr_w[11] addr_w[12] addr_w[13] addr_w[1] addr_w[2] addr_w[3] addr_w[4]
+ addr_w[5] addr_w[6] addr_w[7] addr_w[8] addr_w[9] baseaddr_r_sync[0] baseaddr_r_sync[1]
+ baseaddr_r_sync[2] baseaddr_r_sync[3] baseaddr_r_sync[4] baseaddr_r_sync[5] baseaddr_r_sync[6]
+ baseaddr_r_sync[7] baseaddr_r_sync[8] baseaddr_w_sync[0] baseaddr_w_sync[1] baseaddr_w_sync[2]
+ baseaddr_w_sync[3] baseaddr_w_sync[4] baseaddr_w_sync[5] baseaddr_w_sync[6] baseaddr_w_sync[7]
+ baseaddr_w_sync[8] clk conf[0] conf[1] conf[2] csb csb0_sync csb1_sync d_fabric_in[0]
+ d_fabric_in[10] d_fabric_in[11] d_fabric_in[12] d_fabric_in[13] d_fabric_in[14]
+ d_fabric_in[15] d_fabric_in[16] d_fabric_in[17] d_fabric_in[18] d_fabric_in[19]
+ d_fabric_in[1] d_fabric_in[20] d_fabric_in[21] d_fabric_in[22] d_fabric_in[23] d_fabric_in[24]
+ d_fabric_in[25] d_fabric_in[26] d_fabric_in[27] d_fabric_in[28] d_fabric_in[29]
+ d_fabric_in[2] d_fabric_in[30] d_fabric_in[31] d_fabric_in[3] d_fabric_in[4] d_fabric_in[5]
+ d_fabric_in[6] d_fabric_in[7] d_fabric_in[8] d_fabric_in[9] d_fabric_out[0] d_fabric_out[10]
+ d_fabric_out[11] d_fabric_out[12] d_fabric_out[13] d_fabric_out[14] d_fabric_out[15]
+ d_fabric_out[16] d_fabric_out[17] d_fabric_out[18] d_fabric_out[19] d_fabric_out[1]
+ d_fabric_out[20] d_fabric_out[21] d_fabric_out[22] d_fabric_out[23] d_fabric_out[24]
+ d_fabric_out[25] d_fabric_out[26] d_fabric_out[27] d_fabric_out[28] d_fabric_out[29]
+ d_fabric_out[2] d_fabric_out[30] d_fabric_out[31] d_fabric_out[3] d_fabric_out[4]
+ d_fabric_out[5] d_fabric_out[6] d_fabric_out[7] d_fabric_out[8] d_fabric_out[9]
+ d_sram_in[0] d_sram_in[10] d_sram_in[11] d_sram_in[12] d_sram_in[13] d_sram_in[14]
+ d_sram_in[15] d_sram_in[16] d_sram_in[17] d_sram_in[18] d_sram_in[19] d_sram_in[1]
+ d_sram_in[20] d_sram_in[21] d_sram_in[22] d_sram_in[23] d_sram_in[24] d_sram_in[25]
+ d_sram_in[26] d_sram_in[27] d_sram_in[28] d_sram_in[29] d_sram_in[2] d_sram_in[30]
+ d_sram_in[31] d_sram_in[3] d_sram_in[4] d_sram_in[5] d_sram_in[6] d_sram_in[7] d_sram_in[8]
+ d_sram_in[9] d_sram_out[0] d_sram_out[10] d_sram_out[11] d_sram_out[12] d_sram_out[13]
+ d_sram_out[14] d_sram_out[15] d_sram_out[16] d_sram_out[17] d_sram_out[18] d_sram_out[19]
+ d_sram_out[1] d_sram_out[20] d_sram_out[21] d_sram_out[22] d_sram_out[23] d_sram_out[24]
+ d_sram_out[25] d_sram_out[26] d_sram_out[27] d_sram_out[28] d_sram_out[29] d_sram_out[2]
+ d_sram_out[30] d_sram_out[31] d_sram_out[3] d_sram_out[4] d_sram_out[5] d_sram_out[6]
+ d_sram_out[7] d_sram_out[8] d_sram_out[9] out_reg reb w_mask[0] w_mask[10] w_mask[11]
+ w_mask[12] w_mask[13] w_mask[14] w_mask[15] w_mask[16] w_mask[17] w_mask[18] w_mask[19]
+ w_mask[1] w_mask[20] w_mask[21] w_mask[22] w_mask[23] w_mask[24] w_mask[25] w_mask[26]
+ w_mask[27] w_mask[28] w_mask[29] w_mask[2] w_mask[30] w_mask[31] w_mask[3] w_mask[4]
+ w_mask[5] w_mask[6] w_mask[7] w_mask[8] w_mask[9] web web0_sync VPWR VGND
XFILLER_100_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0703__A _0703_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_188 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_98 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_206 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_291 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_51 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0613__A _0697_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_282 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0708__B1 _0707_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1104__CLK _1197_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_263 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0765__A2_N _0529_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_217 VGND VPWR sky130_fd_sc_hd__fill_2
X_0985_ _0985_/A _0985_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0523__A _0570_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_39 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_250 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0650__A2 _0623_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1127__CLK _1150_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_106 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_128 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0608__A _0542_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_228 VGND VPWR sky130_fd_sc_hd__decap_3
X_0770_ _0762_/X _1089_/D _0769_/X d_fabric_out[6] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_5_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_139 VGND VPWR sky130_fd_sc_hd__decap_4
X_1184_ d_fabric_in[18] _1184_/Q _1223_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0518__A _0517_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_150 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_239 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0632__A2 _0627_/Y VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_12_0_clk clkbuf_3_6_0_clk/X _1162_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0968_ _0968_/A _0968_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0899_ _0899_/A _0899_/B _0903_/C _1177_/Q _0899_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0700__B _0700_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_277 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_228 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0871__A2 _0833_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0623__A2 _0620_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_35 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_132 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1144__D d_sram_out[29] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0847__C1 _0846_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0862__A2 _0839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_60 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_194 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_93 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_119 VGND VPWR sky130_fd_sc_hd__decap_3
X_0822_ d_sram_in[0] _0880_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0753_ _0642_/D _0496_/A _0709_/X _0753_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_127_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0801__A _0776_/A VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_1_0_clk clkbuf_3_1_0_clk/A clkbuf_4_3_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_50_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_0684_ _0675_/X _0684_/B _0684_/C _0683_/X _0684_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_96_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_191 VGND VPWR sky130_fd_sc_hd__fill_2
X_1167_ d_fabric_in[1] _0827_/A _1188_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1098_ _1098_/D _1098_/Q _1126_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0853__A2 _0946_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0711__A _0659_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1030__A2 _1025_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_97 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_52 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_96 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_163 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1139__D d_sram_out[24] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0978__D _0991_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0780__A1 _0779_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0780__B2 _1091_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_71 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0994__C _0953_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_234 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_245 VGND VPWR sky130_fd_sc_hd__decap_4
X_1021_ _0973_/A _1021_/B _1017_/C _1017_/D _1022_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_46_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_70 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_81 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_153 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_197 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0930__B1_N _0873_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0805_ _0799_/X _1102_/Q _0742_/D _0801_/X d_fabric_out[19] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1012__A2 _0983_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0531__A _0580_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0736_ _0668_/X _0737_/A _0501_/X _0735_/X _0736_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_115_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_125 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_188 VGND VPWR sky130_fd_sc_hd__decap_12
X_0667_ _0493_/X _0750_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1065__C _0952_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0598_ _0569_/X _0701_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_29_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_139 VGND VPWR sky130_fd_sc_hd__decap_4
X_1219_ addr_r[7] baseaddr_r_sync[7] _1128_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1079__A2 _1040_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_172 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0826__A2 _0834_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_175 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_278 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_289 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0817__A2 _1110_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_62 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_153 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0616__A _0510_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_56 VGND VPWR sky130_fd_sc_hd__decap_12
X_0521_ _0521_/A _0740_/B _0738_/C _1127_/Q _0546_/B VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0753__A1 _0642_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_1004_ _1031_/D _1017_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0526__A _0525_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_197 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_217 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1160__CLK _1223_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0899__C _0903_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0719_ _0651_/Y _0719_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_106_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_201 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_142 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_87 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_86 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0602__C _0702_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0735__A1 _0521_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0735__B2 _0655_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1152__D _1160_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_120 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0991__D _0991_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_292 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0671__B1 _0681_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_93 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_170 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1183__CLK _1162_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_181 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_209 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_101 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_134 VGND VPWR sky130_fd_sc_hd__fill_2
X_0504_ _0504_/A _0533_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_100_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_212 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_226 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0703__B _0703_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_123 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_127 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_149 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_41 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0613__B _0701_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0708__A1 _0705_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1147__D _1155_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0892__B1 _0891_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_0984_ _1044_/A _0985_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_105_209 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_281 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0714__A _0713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_22 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0938__A1 _1196_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1060__B1 _1057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_85 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0608__B _0524_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0874__B1 _0873_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0624__A _0580_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0929__A1 _1188_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1051__B1 _1049_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1221__CLK _1221_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_1183_ d_fabric_in[17] _1183_/Q _1162_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_94_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0865__B1 _0844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_251 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0534__A _0533_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0967_ _0945_/Y _0966_/Y _0946_/X _0960_/X w_mask[1] VGND VPWR sky130_fd_sc_hd__a211o_4
X_0898_ _0895_/D _0877_/X _0897_/Y d_sram_in[10] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0700__C _0717_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_137 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_289 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0709__A _0501_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0856__B1 _0855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_27 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_47 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1033__B1 _1029_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_144 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_51 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0619__A _0619_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0847__B1 _0844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1160__D _1223_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_173 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_83 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_251 VGND VPWR sky130_fd_sc_hd__decap_12
X_0821_ _0662_/X _1114_/Q _0616_/C _0779_/X d_fabric_out[31] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_80_93 VGND VPWR sky130_fd_sc_hd__decap_12
X_0752_ _0532_/X _0751_/X _0719_/X _0752_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0683_ _0509_/B _0679_/X _0681_/X _0682_/X _0683_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_43_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_118 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0529__A _0529_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1117__CLK _1162_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1166_ d_fabric_in[0] d_sram_in[0] _1188_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_195 VGND VPWR sky130_fd_sc_hd__fill_2
X_1097_ _0795_/X _1097_/Q _1089_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_60_19 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_143 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_154 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_232 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0780__A2 _0778_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_210 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1155__D _1226_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_243 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0994__D _0972_/A VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_clk clkbuf_3_5_0_clk/X _1226_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1020_ _0998_/X _1018_/X _1019_/X w_mask[10] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_46_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_70 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_92 VGND VPWR sky130_fd_sc_hd__decap_8
X_0804_ _0799_/X _1101_/Q _0725_/D _0801_/X d_fabric_out[18] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_115_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_0735_ _0521_/A _0669_/X _0739_/D _0742_/D _0655_/B _0735_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_115_145 VGND VPWR sky130_fd_sc_hd__fill_2
X_0666_ _0663_/X _0660_/X _0665_/X d_fabric_out[0] VGND VPWR sky130_fd_sc_hd__a21o_4
X_0597_ _0725_/C _0597_/B _0597_/C _0619_/A VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_29_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_265 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0781__A1_N _0674_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_224 VGND VPWR sky130_fd_sc_hd__fill_2
X_1218_ addr_r[6] baseaddr_r_sync[6] _1109_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_151 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_132 VGND VPWR sky130_fd_sc_hd__fill_2
X_1149_ _1149_/D _0499_/A _1162_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_4_206 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0722__A _0722_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_195 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_0_0_clk clkbuf_3_1_0_clk/A clkbuf_4_0_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0616__B _0513_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_68 VGND VPWR sky130_fd_sc_hd__decap_12
X_0520_ _0540_/C _0738_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0753__A2 _0496_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_202 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_70 VGND VPWR sky130_fd_sc_hd__decap_12
X_1003_ _0972_/A _1031_/D VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_19_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_121 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_154 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0542__A _0542_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_270 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0899__D _1177_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0718_ _0718_/A _0716_/X _0501_/X _0717_/X _0718_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_0649_ _0626_/Y _0632_/X _0636_/Y _0647_/X _0648_/Y _0649_/X VGND VPWR sky130_fd_sc_hd__o41a_4
XFILLER_122_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0717__A _0722_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_99 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0602__D _0602_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0735__A2 _0669_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_192 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_84 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_227 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0627__A _0562_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_113 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0671__A1 _0521_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_135 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0671__B2 _0655_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_83 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_179 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_171 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VPWR sky130_fd_sc_hd__decap_3
X_0503_ _1150_/Q _0513_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_100_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_271 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0703__C _0701_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_87 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_146 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_135 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_97 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0613__C _0594_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0910__A _0866_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0708__A2 _0706_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1163__D _1163_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0892__A1 _0827_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1150__CLK _1150_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0983_ _0982_/X _0983_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0898__B1_N _0897_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_160 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_293 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0714__B _0714_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_105 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_127 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_296 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0938__A2 _0922_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1060__A1 _0992_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_160 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1173__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0874__A1 _0872_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_41 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0905__A _0861_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0929__A2 _0926_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1051__A1 _0965_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1158__D _1158_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_153 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_164 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0640__A _0580_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_7 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_93 VGND VPWR sky130_fd_sc_hd__decap_12
X_1182_ d_fabric_in[16] _1182_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_83_108 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0865__A1 _0827_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_174 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_293 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0815__A out_reg VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_296 VGND VPWR sky130_fd_sc_hd__decap_3
X_0966_ _0965_/X _0966_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0550__A _0549_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0897_ _0897_/A _0896_/X _0897_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_99_241 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0700__D _1130_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1196__CLK _1223_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_19 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_171 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0856__A1 _0851_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0725__A _0576_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_66 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1033__A1 _0945_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0619__B _0619_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_182 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0847__A1 _0880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0635__A _0526_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_296 VGND VPWR sky130_fd_sc_hd__decap_3
X_0820_ _0662_/X _1113_/Q _1145_/Q _0815_/X d_fabric_out[30] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_127_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_0751_ _0668_/X _1127_/Q _0635_/C _0751_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_0682_ _0722_/A _0738_/B _0540_/C _1128_/Q _0682_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_36_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_1165_ _1165_/D csb1_sync _1197_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1096_ _0793_/X _1096_/Q _1089_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_163 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0545__A _0540_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_0949_ _0949_/A _0955_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_118_187 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0774__B1 _0709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0829__A1 _0880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1211__CLK _1132_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_65 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_87 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_110 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_154 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0765__B1 _0668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_190 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_95 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1171__D d_fabric_in[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_185 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_166 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_177 VGND VPWR sky130_fd_sc_hd__decap_4
X_0803_ _0799_/X _1100_/Q _0681_/D _0801_/X d_fabric_out[17] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__0756__B1 _0755_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0734_ _0663_/X _1085_/D _0733_/X d_fabric_out[2] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_115_135 VGND VPWR sky130_fd_sc_hd__decap_8
X_0665_ _1083_/Q _0776_/A _0665_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_130_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_0596_ _1134_/Q _0580_/C _0718_/A _0526_/X _0595_/X _0597_/C VGND VPWR sky130_fd_sc_hd__a2111oi_4
XFILLER_69_233 VGND VPWR sky130_fd_sc_hd__decap_4
X_1217_ addr_r[5] baseaddr_r_sync[5] _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_1148_ _1148_/D _0498_/A _1162_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_111_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_1079_ _0985_/A _1040_/X _1075_/Y _1079_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0778__A2_N _0496_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_249 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0722__B _0492_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0747__B1 _0742_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_56 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_78 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_31 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_291 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_239 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_86 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0616__C _0616_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_188 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1107__CLK _1132_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_293 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1166__D d_fabric_in[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_82 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_130 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_247 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_93 VGND VPWR sky130_fd_sc_hd__decap_6
X_1002_ _0998_/X _1001_/X _0996_/X w_mask[7] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_19_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0823__A _1226_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_208 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0542__B _0513_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0717_ _0722_/D _0717_/B _0717_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0648_ _0509_/A _0703_/A _0622_/Y _0648_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_0579_ _0533_/X _0580_/C _0569_/X _1130_/Q _0579_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_111_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_269 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_206 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0717__B _0717_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_291 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_261 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_177 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_125 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_147 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0733__A _0733_/A VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_10_0_clk clkbuf_3_5_0_clk/X _1128_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_119_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0735__A3 _0739_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_210 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_225 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_298 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_206 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0908__A _0903_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0671__A2 _0669_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_150 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0643__A _0533_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0959__B1 _0958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_172 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_241 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0795__A1_N _0575_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0502_ _0502_/A _0509_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_39_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_147 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0553__A _0524_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0703__D _0702_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_103 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0728__A _0721_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_44 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_10 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_32 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0613__D _1141_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0910__B _0910_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0638__A _0722_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_239 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0892__A2 _0890_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_209 VGND VPWR sky130_fd_sc_hd__fill_2
X_0982_ _0982_/A _0982_/B _0991_/C _0991_/D _0982_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_66_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_211 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_106 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0548__A _0547_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_194 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1060__A2 _1059_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_233 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_239 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0874__A2 _0875_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0905__B _0904_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_86 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1051__A2 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_110 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_176 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1174__D d_fabric_in[8] VGND VPWR sky130_fd_sc_hd__diode_2
X_1181_ d_fabric_in[15] _1181_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_76_172 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0865__A2 _0859_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_93 VGND VPWR sky130_fd_sc_hd__decap_12
X_0965_ _0964_/X _0965_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0831__A _1226_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0896_ _0846_/A _0890_/X _0895_/X _0896_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1084__D _0712_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_109 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0856__A2 _0833_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_186 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_220 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0725__B _0544_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0741__A _0510_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1033__A2 _1032_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1140__CLK _1197_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_64 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_97 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0619__C _0619_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_153 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0847__A2 _0946_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_52 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0916__A _0903_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0635__B _0633_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1169__D d_fabric_in[3] VGND VPWR sky130_fd_sc_hd__diode_2
X_0750_ _0750_/A _0750_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0651__A _0500_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0681_ _0542_/A _0492_/C _0722_/C _0681_/D _0681_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_89_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_289 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_161 VGND VPWR sky130_fd_sc_hd__fill_2
X_1164_ web web0_sync _1197_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1095_ _1095_/D _1095_/Q _1089_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0545__B _0542_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0561__A _0517_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1163__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0948_ _0969_/A _0949_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_118_166 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0774__A1 _1122_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0879_ _0952_/C _1046_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_133_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0829__A2 _0826_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_153 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_134 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_44 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_189 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_245 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_177 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0765__B2 _0724_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_289 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_62 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_73 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0646__A _0642_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1186__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0802_ _0799_/X _1099_/Q _0655_/A _0801_/X d_fabric_out[16] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__0756__A1 _0663_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0733_ _0733_/A _1085_/Q _0733_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0664_ out_reg _0776_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_130_117 VGND VPWR sky130_fd_sc_hd__decap_8
X_0595_ _1132_/Q _0582_/X _0595_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_37_120 VGND VPWR sky130_fd_sc_hd__fill_2
X_1216_ addr_r[4] baseaddr_r_sync[4] _1197_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_84_248 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_259 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_92 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_164 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0556__A _0581_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1147_ _1155_/Q _1147_/Q _1150_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_111_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_1078_ _1032_/X _1070_/X _1076_/X w_mask[29] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_52_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_167 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0722__C _0722_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0747__A1 _0750_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0747__B2 _0496_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_106 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_229 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0616__D _0533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_20 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_42 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_117 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1182__D d_fabric_in[16] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_259 VGND VPWR sky130_fd_sc_hd__decap_12
X_1001_ _1000_/X _1001_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_19_153 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1000__A _0973_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0542__C _0544_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0716_ _0668_/A _0720_/A _0716_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1201__CLK _1128_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0647_ _0647_/A _0639_/X _0641_/X _0646_/X _0647_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_0578_ _0559_/X _0568_/Y _0574_/Y _0578_/D _0578_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XANTENNA__1092__D _0781_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_259 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_251 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0733__B _1085_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_264 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_215 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_237 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_42 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0908__B _0903_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_148 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0671__A3 _0676_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_140 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_151 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0643__B _0565_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_162 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0959__A1 _1055_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_173 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1081__B1 _1079_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1177__D d_fabric_in[11] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1224__CLK _1128_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_7 VGND VPWR sky130_fd_sc_hd__decap_12
X_0501_ _0500_/X _0501_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_11_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_281 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0834__A _0834_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1072__B1 _1071_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1087__D _0754_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_207 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0728__B _0722_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_23 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0744__A _0738_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_22 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1063__B1 _1061_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0810__B1 _0723_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_231 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_286 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_275 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_74 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0638__B _0558_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_251 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0654__A _0690_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0981_ _1031_/A _0982_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1054__B1 _1052_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_118 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0868__B1 _0867_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_140 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_240 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0564__A _0564_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0739__A _0722_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_107 VGND VPWR sky130_fd_sc_hd__fill_2
X_1180_ d_fabric_in[14] _0912_/D _1089_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1190__D d_fabric_in[24] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_162 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_276 VGND VPWR sky130_fd_sc_hd__decap_12
X_0964_ _1031_/A _1021_/B _0977_/A _0972_/A _0964_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0831__B _0841_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0895_ _0899_/A _0899_/B _0903_/C _0895_/D _0895_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_59_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_237 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1092__CLK _1126_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_232 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0725__C _0725_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_112 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0741__B _0513_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_165 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0916__B _0903_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_198 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0635__C _0635_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0932__A _0875_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_0680_ _0544_/C _0722_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1185__D d_fabric_in[19] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_143 VGND VPWR sky130_fd_sc_hd__fill_2
X_1163_ _1163_/D csb0_sync _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1094_ _0788_/X _1094_/Q _1089_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0545__C _0544_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1003__A _0972_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_202 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0842__A _0841_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0561__B _0564_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0947_ _0962_/A _0969_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_109_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0774__A2 _0659_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0878_ _0838_/A _0952_/C VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_133_159 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1095__D _1095_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_202 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_213 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_23 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_56 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_31 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_42 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_154 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0646__B _0643_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_113 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_62 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0662__A _0662_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0801_ _0776_/A _0801_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0756__A2 _0754_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0732_ out_reg _0733_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0663_ _0662_/X _0663_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0610__D1 _0609_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_0594_ _0725_/D _0594_/B _0718_/A VGND VPWR sky130_fd_sc_hd__and2_4
X_1215_ addr_r[3] baseaddr_r_sync[3] _1188_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0837__A _0943_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0556__B _0556_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1146_ d_sram_out[31] _0616_/C _1197_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_113 VGND VPWR sky130_fd_sc_hd__fill_1
X_1077_ _1025_/X _1070_/X _1076_/X w_mask[28] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_111_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1130__CLK _1223_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0572__A _0571_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_218 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0722__D _0722_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0747__A2 _0736_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_143 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_157 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_83 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_32 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_80 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1153__CLK _1226_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1000_ _0973_/A _0991_/B _1000_/C _0991_/D _1000_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_19_165 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_102 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_271 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_clk_A clk VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1000__B _0991_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0542__D _0542_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0715_ _0663_/X _0712_/X _0714_/X d_fabric_out[1] VGND VPWR sky130_fd_sc_hd__a21o_4
X_0646_ _0642_/X _0643_/X _0646_/C _0646_/D _0646_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA_clkbuf_4_9_0_clk_A clkbuf_4_9_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0577_ _0575_/Y _0576_/X _0518_/X _0701_/C _0578_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0567__A _0645_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_249 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_1129_ d_sram_out[14] _0724_/D _1214_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1176__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_32 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0908__C _0908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_102 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_271 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_241 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_105 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_130 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0643__C _0643_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_163 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0959__A2 _0838_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_174 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1081__A1 _1040_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0940__A _0962_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_221 VGND VPWR sky130_fd_sc_hd__decap_12
X_0500_ _0499_/X _0500_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1193__D d_fabric_in[27] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_296 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1011__A _1009_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1072__A1 _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_182 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1199__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_0629_ _0629_/A _0703_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_133_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0728__C _0723_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_219 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_241 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_79 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0744__B _0744_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1063__A1 _1001_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_171 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0810__B2 _0808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0810__A1 _0806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_298 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_182 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_74 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_96 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_296 VGND VPWR sky130_fd_sc_hd__decap_3
X_0980_ _0968_/X _0979_/X _0975_/Y w_mask[3] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__1054__A1 _0979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1188__D d_fabric_in[22] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_7 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0670__A _0602_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_193 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0868__A1 _0864_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1006__A _1005_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_208 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0845__A _0835_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1098__D _1098_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0580__A _0533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0739__B _0492_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_clk_A clkbuf_3_7_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0755__A _0733_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1214__CLK _1214_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_296 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0490__A _0556_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0795__B1 _1145_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0665__A _1083_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_288 VGND VPWR sky130_fd_sc_hd__decap_8
X_0963_ _0963_/A _1021_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0786__B1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0831__C _1042_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0894_ _0891_/D _0877_/X _0893_/Y d_sram_in[9] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_99_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_249 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0575__A _0724_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0710__B1 _0709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_27 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0725__D _0725_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0777__B1 _0776_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0741__C _0724_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_22 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_44 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0916__C _0908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_188 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0768__B1 _0766_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_51 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_269 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_192 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_122 VGND VPWR sky130_fd_sc_hd__fill_2
X_1162_ _1225_/Q _1162_/Q _1162_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1093_ _0784_/X _1093_/Q _1109_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_269 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0759__B1 _0719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0561__C _0510_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0946_ _0946_/A _0942_/Y _0946_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_9_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_0877_ _0922_/B _0877_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_126_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_258 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_269 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_169 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_56 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_3_0_clk_A clkbuf_2_2_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0646__C _0646_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0943__A _0943_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0989__B1 _0988_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0800_ _0713_/X _1098_/D _0799_/X _1098_/Q d_fabric_out[15] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1196__D d_fabric_in[30] VGND VPWR sky130_fd_sc_hd__diode_2
X_0731_ _0750_/A _0718_/X _0730_/X _0725_/D _0711_/X _1085_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_6_251 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0610__C1 _0608_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_149 VGND VPWR sky130_fd_sc_hd__fill_2
X_0662_ _0662_/A _0662_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0593_ _0587_/C _0594_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_123_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0913__B1 _0912_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_228 VGND VPWR sky130_fd_sc_hd__fill_2
X_1214_ addr_r[2] baseaddr_r_sync[2] _1214_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_111 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_291 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0837__B _0834_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1145_ d_sram_out[30] _1145_/Q _1197_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_92_250 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0556__C _0504_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1014__A _0982_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_136 VGND VPWR sky130_fd_sc_hd__fill_2
X_1076_ _0985_/A _1035_/X _1075_/Y _1076_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA_clkbuf_4_5_0_clk_A clkbuf_3_2_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_180 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_0929_ _1188_/Q _0926_/X _0870_/X d_sram_in[22] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0747__A3 _0746_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0904__B1 _0903_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_261 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0763__A _0733_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_62 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_95 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_206 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_291 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_239 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_177 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0673__A _0583_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1000__C _1000_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_274 VGND VPWR sky130_fd_sc_hd__fill_1
X_0714_ _0713_/X _0714_/B _0714_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0645_ _0645_/A _0565_/X _0643_/C _1121_/Q _0646_/D VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1009__A _1007_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0576_ _0517_/X _0565_/A _0576_/C _0513_/A _0576_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_57_217 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0848__A _0897_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0567__B _0580_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1128_ d_sram_out[13] _1128_/Q _1128_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1059_ _1043_/A _1059_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_15_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0583__A _0645_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_139 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_213 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_206 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0908__D _1179_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0493__A _0492_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_139 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_180 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_120 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0643__D _0724_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_87 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_153 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1081__A2 _1043_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_186 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0940__B _0970_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_233 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1120__CLK _1214_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0668__A _0668_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_1_0_0_clk_A clkbuf_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0577__A1_N _0575_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_139 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_180 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1011__B _1028_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1072__A2 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_128 VGND VPWR sky130_fd_sc_hd__fill_2
X_0628_ _0580_/B _0701_/C _0629_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_131_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0578__A _0559_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0559_ _0554_/Y _0557_/X _1128_/Q _0558_/X _0559_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0728__D _0728_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_264 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0744__C _0740_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_clk_A clkbuf_3_3_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1063__A2 _1059_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0810__A2 _1105_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1143__CLK _1089_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_3 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0488__A _1147_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13_0_clk_A clkbuf_3_6_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1054__A2 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0951__A _0963_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_132 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_7 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0868__A2 _0833_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_19 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0845__B _0834_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1022__A _1022_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0861__A _0861_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1166__CLK _1188_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0580__B _0580_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_109 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0739__C _0722_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0755__B _1087_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_23 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_45 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_67 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0771__A _0740_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0795__B2 _0711_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_239 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0946__A _0946_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0665__B _0776_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_201 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1189__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1199__D addr_w[1] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0681__A _0542_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0962_ _0962_/A _1031_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0786__B2 _1093_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0786__A1 _0779_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0893_ _0866_/A _0893_/B _0893_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_99_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_109 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1017__A _0973_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0710__A1 _0685_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_167 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0591__A _0591_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0777__A1 _0762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0741__D _1130_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_56 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_131 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_22 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_44 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0916__D _1181_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_178 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0768__B2 _0767_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0768__A1 _0723_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_171 VGND VPWR sky130_fd_sc_hd__decap_12
X_1161_ _1224_/Q _1161_/Q _1226_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0676__A _0521_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_101 VGND VPWR sky130_fd_sc_hd__decap_4
X_1092_ _0781_/X _1092_/Q _1126_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_237 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_215 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0759__A1 _0757_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0561__D _1150_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0945_ _0945_/A _0945_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_9_293 VGND VPWR sky130_fd_sc_hd__decap_6
X_0876_ _0875_/Y _0922_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1204__CLK _1188_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_1_0_clk_A clkbuf_4_0_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0931__A1 _1190_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0586__A _0517_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_126 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_69 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_180 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_22 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_194 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0496__A _0496_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0646__D _0646_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0989__A1 _0985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0943__B _0834_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_91 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1227__CLK _1188_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0730_ _1117_/Q _0549_/A _0719_/X _0729_/X _0730_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__0610__B1 _0607_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_296 VGND VPWR sky130_fd_sc_hd__decap_3
X_0661_ out_reg _0662_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_0592_ _0569_/X _0597_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_237 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0913__A1 _1172_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1213_ addr_r[1] baseaddr_r_sync[1] _1226_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0837__C _1042_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1144_ d_sram_out[29] _1112_/D _1188_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_1_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_156 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1014__B _1021_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0556__D _0564_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1075_ _1066_/B _1074_/X _1056_/C _1075_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_0928_ _1187_/Q _0926_/X _0867_/X d_sram_in[21] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_106_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_0859_ _0955_/D _0946_/A _0859_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_136_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0904__A1 _1170_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_270 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_35 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_41 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0763__B _1088_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0605__A2_N _0562_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_134 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_115 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0954__A _0953_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1000__D _0991_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0713_ out_reg _0713_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0644_ _0533_/X _0565_/X _0584_/C _0720_/A _0646_/C VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1009__B _1045_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_19 VGND VPWR sky130_fd_sc_hd__decap_12
X_0575_ _0724_/D _0575_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_111_153 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_164 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0567__C _0643_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1025__A _1024_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_240 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0864__A _1171_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1127_ d_sram_out[12] _1127_/Q _1150_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_80_210 VGND VPWR sky130_fd_sc_hd__fill_2
X_1058_ _0983_/X _1043_/X _1057_/X w_mask[20] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_15_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_107 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0583__B _0569_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_265 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_118 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_110 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_298 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_99 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0940__C _0977_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0949__A _0949_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0559__A2_N _0557_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0684__A _0675_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_210 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1057__B1 _1056_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_118 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_192 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0804__B1 _0725_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1011__C _0960_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_118 VGND VPWR sky130_fd_sc_hd__fill_2
X_0627_ _0562_/X _0627_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0859__A _0955_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0578__B _0568_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0558_ _0533_/A _1153_/Q _0576_/C _0513_/A _0558_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_133_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1095__CLK _1089_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0489_ _1150_/Q _0556_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_38_251 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0594__A _0725_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0744__D _0743_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_201 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_278 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0769__A _0733_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_99 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_3_0_clk clkbuf_2_2_0_clk/A clkbuf_3_7_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_44_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0679__A _0722_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_162 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_198 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0845__C _0841_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0580__C _0580_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_204 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0589__A _0579_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0961__C1 _0960_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0739__D _0739_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_110 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_35 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1110__CLK _1214_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_57 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0771__B _0655_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0894__B1_N _0893_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0499__A _0499_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_154 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_176 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0946__B _0942_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_146 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_91 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_179 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0962__A _0962_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0681__B _0492_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0961_ _0942_/Y _0945_/Y _0946_/X _0960_/X w_mask[0] VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__0786__A2 _0784_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0892_ _0827_/A _0890_/X _0891_/X _0893_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_57_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_257 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1017__B _0982_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_132 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0710__A2 _0708_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1133__CLK _1223_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0872__A _1173_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0591__B _0591_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0777__A2 _0775_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_68 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_56 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0768__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_110 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0957__A _0956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0676__B _0492_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1160_ _1223_/Q _1160_/Q _1223_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1156__CLK _1162_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1091_ _0778_/X _1091_/Q _1126_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0692__A _0739_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_249 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0759__A2 _0758_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0944_ _0968_/A _0945_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0875_ _0875_/A _0875_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_133_107 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1028__A _1028_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0931__A2 _0926_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_238 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0586__B _0565_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_179 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_129 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1179__CLK _1221_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_45 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_89 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_271 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_146 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0989__A2 _0974_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0943__C _0908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_76 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0610__A1 _0675_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0660_ _0681_/D _0496_/X _0659_/X _0660_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_108_192 VGND VPWR sky130_fd_sc_hd__fill_2
X_0591_ _0591_/A _0591_/B _0591_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_123_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0687__A _0675_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0913__A2 _1046_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1212_ addr_r[0] baseaddr_r_sync[0] _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_77_260 VGND VPWR sky130_fd_sc_hd__fill_2
X_1143_ d_sram_out[28] _0532_/A _1089_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_1_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1014__C _1017_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_116 VGND VPWR sky130_fd_sc_hd__fill_2
X_1074_ _1007_/X _1055_/B _0973_/C _1045_/D _1074_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_92_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_296 VGND VPWR sky130_fd_sc_hd__decap_3
X_0927_ _1186_/Q _0926_/X _0862_/X d_sram_in[20] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_106_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_0858_ _0852_/B _0955_/D VGND VPWR sky130_fd_sc_hd__buf_1
X_0789_ _0779_/X _0788_/X _0785_/X _1094_/Q d_fabric_out[11] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__0597__A _0725_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0904__A2 _0890_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_230 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_168 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_53 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_24 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_35 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_79 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_241 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_182 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0970__A _0970_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_276 VGND VPWR sky130_fd_sc_hd__decap_12
X_0712_ _0750_/A _0672_/X _0710_/Y _0681_/D _0711_/X _0712_/X VGND VPWR sky130_fd_sc_hd__a32o_4
X_0643_ _0533_/A _0565_/X _0643_/C _0724_/D _0643_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1009__C _0991_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_0574_ _0518_/X _0569_/X _0573_/Y _0574_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0898__A1 _0895_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_176 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0567__D _1118_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1126_ d_sram_out[11] _0737_/A _1126_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_116 VGND VPWR sky130_fd_sc_hd__decap_4
X_1057_ _1044_/X _1018_/X _1056_/Y _1057_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_15_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0583__C _0582_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_244 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0880__A _0880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_121 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0889__A1 _0887_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1217__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_149 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1101__D _0725_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_144 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0940__D _0972_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0577__B1 _0518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_93 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0965__A _0964_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0684__B _0684_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_244 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1057__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0804__A1 _0799_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk clk clkbuf_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_30_163 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0804__B2 _0801_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0568__B1 _0567_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_62 VGND VPWR sky130_fd_sc_hd__decap_12
X_0626_ _0540_/C _0702_/B _0626_/C _0626_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0859__B _0946_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_141 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_130 VGND VPWR sky130_fd_sc_hd__fill_2
X_0557_ _0556_/X _0557_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0578__C _0574_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1036__A _0960_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0875__A _0875_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0488_ _1147_/Q _0488_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_38_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_296 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0594__B _0594_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_222 VGND VPWR sky130_fd_sc_hd__fill_2
X_1109_ _1141_/Q _1109_/Q _1109_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_53_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_235 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0559__B1 _1128_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0769__B _1089_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_130 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0785__A _0662_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0731__B1 _0725_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_93 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_152 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0798__B1 _0797_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0679__B _0738_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_293 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0695__A _1134_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_200 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0789__B1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0580__D _1122_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0589__B _0580_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0961__B1 _0946_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0609_ _0723_/D _0594_/B _0609_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_37_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_11 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0499__B _1147_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_208 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_122 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_133 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_70 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0681__C _0722_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0960_ _0960_/A _0955_/X _0960_/C _0960_/X VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__1085__CLK _1150_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0891_ _0899_/A _0899_/B _0903_/C _0891_/D _0891_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_99_269 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_170 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_219 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1017__C _1017_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_166 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_39 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_clk clkbuf_2_2_0_clk/A clkbuf_3_5_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_100_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_54 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_98 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_144 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0676__C _0675_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1090_ _0775_/X _1090_/Q _1132_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_147 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0973__A _0973_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0692__B _0558_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_0943_ _0943_/A _0834_/A _0908_/C _1042_/D _0968_/A VGND VPWR sky130_fd_sc_hd__or4_4
X_0874_ _0872_/Y _0875_/A _0873_/X d_sram_in[7] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_133_119 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1028__B _1028_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_206 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1100__CLK _1132_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0586__C _0587_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1044__A _1044_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0883__A _0883_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_191 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_239 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_23 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1104__D _0675_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_11 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0943__D _1042_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0610__A2 _0582_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_70 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1123__CLK _1126_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0590_ _0540_/C _0701_/C _0509_/A _0578_/Y _0589_/Y _0591_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_41_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0968__A _0968_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0687__B _0690_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1211_ addr_w[13] _1042_/D _1132_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_103 VGND VPWR sky130_fd_sc_hd__fill_2
X_1142_ d_sram_out[27] _1142_/Q _1223_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1073_ _1022_/X _1070_/X _1071_/X w_mask[27] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_1_86 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1014__D _1017_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_150 VGND VPWR sky130_fd_sc_hd__fill_1
X_0926_ _0875_/Y _0926_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0857_ _1170_/Q _0857_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1039__A _0949_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0788_ _0554_/Y _0787_/X _0739_/D _0787_/X _0788_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_163 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_141 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0878__A _0838_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0597__B _0597_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_27 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1146__CLK _1197_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_209 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_99 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_92 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_194 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0711_ _0659_/A _0711_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_51_80 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_288 VGND VPWR sky130_fd_sc_hd__decap_8
X_0642_ _0517_/X _0565_/X _0587_/C _0642_/D _0642_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0573_ _0642_/D _0524_/X _1121_/Q _0587_/C _0573_/Y VGND VPWR sky130_fd_sc_hd__a22oi_4
XANTENNA__0698__A _0697_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1009__D _1045_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0898__A2 _0877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_1125_ d_sram_out[10] _0720_/A _1109_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0583__D _0583_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1056_ _1056_/A _1056_/B _1056_/C _1056_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__1169__CLK _1162_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0880__B _1046_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_0909_ _1171_/Q _0890_/X _0908_/X _0910_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_102_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_249 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0889__A2 _0877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_36 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_245 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_109 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_101 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_145 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_214 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0577__B2 _0701_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_72 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_269 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_98 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0684__C _0684_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1057__A2 _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0981__A _1031_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_172 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0804__A2 _1101_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_186 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_203 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0568__A1 _0560_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_74 VGND VPWR sky130_fd_sc_hd__decap_12
X_0625_ _0614_/Y _0529_/A _0603_/Y _0571_/X _0626_/C VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_97_120 VGND VPWR sky130_fd_sc_hd__fill_2
X_0556_ _0581_/A _0556_/B _0504_/A _0564_/A _0556_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_97_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0578__D _0578_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0487_ _1132_/Q _0681_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1036__B _1028_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_197 VGND VPWR sky130_fd_sc_hd__fill_2
X_1108_ _0602_/D _1108_/Q _1126_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1202__D addr_w[4] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0891__A _0899_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1039_ _0949_/A _1021_/B _1000_/C _1031_/D _1039_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_42_38 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0559__B2 _0558_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_269 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_120 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_24 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_220 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0731__B2 _0711_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0731__A1 _0750_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1112__D _1112_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0788__A2_N _0787_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_72 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0798__A1 _1130_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0679__C _0544_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_239 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_226 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0789__B2 _1094_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0789__A1 _0779_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1207__CLK _1150_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0589__C _0583_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0961__A1 _0942_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0608_ _0542_/D _0524_/X _0608_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0539_ _0576_/C _0542_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0886__A _0908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_49 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_127 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_149 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0499__C _0499_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1107__D _1107_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_145 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0681__D _0681_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0890_ _1046_/C _0890_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_138_180 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_237 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_182 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1017__D _1017_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_192 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0790__A1_N _0560_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_139 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_180 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0934__A1 _1192_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_270 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_178 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0870__B1 _0848_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0925__A1 _1185_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0676__D _0676_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_178 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_126 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0973__B _0982_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_181 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_281 VGND VPWR sky130_fd_sc_hd__decap_12
X_0942_ _0942_/A _0942_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_118_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_0873_ _0872_/Y _0838_/X _0854_/Y _0873_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_62_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_240 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0586__D _1117_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1210__D addr_w[12] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_197 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_35 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_23 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1120__D d_sram_out[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_83 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1020__B1 _1019_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_229 VGND VPWR sky130_fd_sc_hd__fill_2
X_1210_ addr_w[12] _0972_/A _1188_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_77_240 VGND VPWR sky130_fd_sc_hd__fill_2
X_1141_ d_sram_out[26] _1141_/Q _1223_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_77_295 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0984__A _1044_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_232 VGND VPWR sky130_fd_sc_hd__decap_3
X_1072_ _1018_/X _1070_/X _1071_/X w_mask[26] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_92_254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_276 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_clk clkbuf_1_0_0_clk/X clkbuf_3_3_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0925_ _1185_/Q _0907_/X _0855_/X d_sram_in[19] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0906__B1_N _0905_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1039__B _1021_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0856_ _0851_/Y _0833_/X _0855_/X d_sram_in[3] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0787_ _0496_/A _0787_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1098__CLK _1126_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_175 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0597__C _0597_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1055__A _0955_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_251 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_148 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1205__D addr_w[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_265 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1078__B1 _1076_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_170 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_118 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1002__B1 _0996_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_126 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1115__D d_sram_out[0] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1069__B1 _1067_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_107 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_287 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0816__B1 _0722_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_151 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_234 VGND VPWR sky130_fd_sc_hd__decap_12
X_0710_ _0685_/X _0708_/Y _0709_/X _0710_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0979__A _0979_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0641_ _0697_/A _0700_/B _0702_/C _1117_/Q _0641_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0572_ _0571_/X _0587_/C VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0698__B _0700_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_232 VGND VPWR sky130_fd_sc_hd__decap_8
X_1124_ d_sram_out[9] _0583_/D _1197_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_80_224 VGND VPWR sky130_fd_sc_hd__decap_3
X_1055_ _0955_/A _1055_/B _0973_/C _1045_/D _1056_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_33_151 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0807__B1 _0542_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_268 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_0908_ _0903_/A _0903_/B _0908_/C _1179_/Q _0908_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_134_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_0839_ _0838_/X _0839_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_206 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_15 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_265 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1113__CLK _1126_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_102 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0799__A _0662_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0684__D _0683_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_81 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_151 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_184 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_198 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0568__A2 _0562_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_86 VGND VPWR sky130_fd_sc_hd__decap_12
X_0624_ _0580_/B _0702_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0502__A _0502_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0555_ _1153_/Q _0564_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_97_154 VGND VPWR sky130_fd_sc_hd__fill_2
X_0486_ reb csb _1165_/D VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_38_210 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1136__CLK _1214_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_276 VGND VPWR sky130_fd_sc_hd__decap_12
X_1107_ _1107_/D _1107_/Q _1132_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0891__B _0899_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1038_ _0945_/A _1035_/X _1037_/X w_mask[14] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_21_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_36 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_165 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0731__A2 _0718_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_132 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0798__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_176 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0679__D _0679_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1159__CLK _1198_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_80 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0992__A _0991_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_238 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0789__A2 _0788_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0589__D _0588_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0961__A2 _0945_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0607_ _0740_/D _0643_/C _0607_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0538_ _0581_/A _0576_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_39 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_179 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1213__D addr_r[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_49 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1123__D d_sram_out[8] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_190 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_194 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0987__A _0955_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_293 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0934__A2 _0932_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0897__A _0897_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1208__D addr_w[10] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_127 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0870__A1 _0869_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_193 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0925__A2 _0907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0600__A _0645_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1118__D d_sram_out[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_93 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0973__C _0973_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_70 VGND VPWR sky130_fd_sc_hd__decap_3
X_0941_ _0940_/X _0942_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_13_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_0872_ _1173_/Q _0872_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_55_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0510__A _0510_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_171 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_219 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_47 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_35 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_110 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1020__A1 _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_162 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_208 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_70 VGND VPWR sky130_fd_sc_hd__fill_1
X_1140_ d_sram_out[25] _0602_/D _1197_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_211 VGND VPWR sky130_fd_sc_hd__decap_3
X_1071_ _0985_/A _1032_/X _1066_/Y _1071_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_92_266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_163 VGND VPWR sky130_fd_sc_hd__fill_2
X_0924_ _1184_/Q _0907_/X _0849_/X d_sram_in[18] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0505__A _0513_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0855_ _0851_/Y _0839_/X _0854_/Y _0855_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1039__C _1000_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0786_ _0779_/X _0784_/X _0785_/X _1093_/Q d_fabric_out[10] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_114_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_187 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0770__B1 _0769_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1055__B _1055_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_138 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_116 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_296 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1078__A1 _1032_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1221__D addr_r[9] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_12 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_182 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_141 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1002__A1 _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_97 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0761__B1 _0759_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_105 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1192__CLK _1221_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_116 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1069__A1 _1015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0816__A1 _0813_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_130 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0816__B2 _0815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1131__D d_sram_out[16] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_83 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_246 VGND VPWR sky130_fd_sc_hd__decap_12
X_0640_ _0580_/B _0700_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0571_ _0570_/X _0571_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0698__C _0594_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0752__B1 _0719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0995__A _0994_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_1123_ d_sram_out[8] _0502_/A _1126_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1054_ _0979_/X _1043_/X _1052_/X w_mask[19] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_25_108 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0807__A1 _0806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0807__B2 _0801_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_174 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_0907_ _0875_/Y _0907_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_119_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_0838_ _0838_/A _0838_/B _0838_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0769_ _0733_/A _1089_/Q _0769_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_0_218 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1066__A _1064_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1216__D addr_r[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_103 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0734__B1 _0733_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_0_0_clk clkbuf_1_0_0_clk/X clkbuf_3_1_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__1126__D d_sram_out[11] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_211 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_247 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1088__CLK _1089_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_122 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_98 VGND VPWR sky130_fd_sc_hd__decap_12
X_0623_ _1115_/Q _0620_/X _0622_/Y _0623_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_131_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_271 VGND VPWR sky130_fd_sc_hd__fill_1
X_0554_ _0737_/A _0554_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_97_144 VGND VPWR sky130_fd_sc_hd__fill_1
X_1106_ _0740_/D _1106_/Q _1126_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_38_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_203 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0891__C _0903_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1037_ _0985_/X _1001_/X _1036_/Y _1037_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_61_291 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_166 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_260 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_22 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_48 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_263 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0731__A3 _0730_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_188 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_148 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0603__A _0532_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_84 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_219 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0707__B1 _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0513__A _0513_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_208 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1103__CLK _1089_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0606_ _0645_/A _0724_/C VGND VPWR sky130_fd_sc_hd__buf_1
X_0537_ _0526_/X _0532_/X _0675_/C _0546_/C VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_112_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_239 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_62 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_239 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1126__CLK _1126_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0987__B _1055_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_80 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_117 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0508__A _0507_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0897__B _0896_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1074__A _1007_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_244 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_222 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1224__D addr_r[12] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_180 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_139 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_239 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0870__A2 _0839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1149__CLK _1162_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_272 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1134__D d_sram_out[19] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_139 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0973__D _0991_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_93 VGND VPWR sky130_fd_sc_hd__fill_1
X_0940_ _0962_/A _0970_/A _0977_/A _0972_/A _0940_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_9_232 VGND VPWR sky130_fd_sc_hd__decap_12
X_0871_ _0869_/Y _0833_/X _0870_/X d_sram_in[6] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_126_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0998__A _0968_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_209 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_220 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_180 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_191 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0660__B1_N _0659_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1219__D addr_r[7] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0701__A _0724_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_38 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_47 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_63 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1129__D d_sram_out[14] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0611__A _0724_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1020__A2 _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_220 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_264 VGND VPWR sky130_fd_sc_hd__fill_2
X_1070_ _1043_/A _1070_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_52_109 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_197 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0505__B _0533_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0923_ _1183_/Q _0922_/B _0844_/X _0922_/Y d_sram_in[17] VGND VPWR sky130_fd_sc_hd__a211o_4
X_0854_ _0854_/A _0854_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0785_ _0662_/X _0785_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0521__A _0521_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1039__D _1031_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0770__A1 _0762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_199 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1055__C _0973_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_234 VGND VPWR sky130_fd_sc_hd__fill_1
X_1199_ addr_w[1] baseaddr_w_sync[1] _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1078__A2 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_161 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1002__A2 _1001_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_155 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0761__A1 _0675_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_188 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0761__B2 _0760_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_231 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_264 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1069__A2 _1059_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_172 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0816__A2 _1109_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_62 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_95 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0606__A _0645_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_258 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_83 VGND VPWR sky130_fd_sc_hd__decap_3
X_0570_ _0570_/A _1150_/Q _0570_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0698__D _0584_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0752__A1 _0532_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_147 VGND VPWR sky130_fd_sc_hd__decap_6
X_1122_ d_sram_out[7] _1122_/Q _1126_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1053_ _0974_/X _1043_/X _1052_/X w_mask[18] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_80_248 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0807__A2 _1103_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0516__A _0504_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0906_ _1178_/Q _0877_/X _0905_/Y d_sram_in[12] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_119_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_0837_ _0943_/A _0834_/A _1042_/C _0838_/B VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_134_239 VGND VPWR sky130_fd_sc_hd__decap_6
X_0768_ _0723_/D _0750_/X _0766_/X _0767_/X _1089_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1066__B _1066_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0699_ _0694_/X _0699_/B _0699_/C _0699_/D _0699_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__1082__A csb VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_204 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_237 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_104 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_186 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_126 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_217 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0734__A1 _0663_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_201 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1142__D d_sram_out[27] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_131 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_259 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_101 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_71 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_178 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_93 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_291 VGND VPWR sky130_fd_sc_hd__decap_8
X_0622_ _0499_/A _0488_/Y _0499_/C _0622_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_0553_ _0524_/X _0701_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_1105_ _0723_/D _1105_/Q _1197_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_53_237 VGND VPWR sky130_fd_sc_hd__decap_4
X_1036_ _0960_/C _1028_/X _1036_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__0891__D _0891_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1182__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_239 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_9 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_272 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_34 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1227__D conf[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_145 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_112 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_74 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1137__D d_sram_out[22] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0707__A1 _0585_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_204 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_281 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_0605_ _0603_/Y _0562_/X _1142_/Q _0639_/B _0612_/C VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_0536_ _0725_/C _0675_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_26_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_170 VGND VPWR sky130_fd_sc_hd__fill_2
X_1019_ _0985_/X _0992_/X _1011_/Y _1019_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0704__A _0704_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0937__A1 _1195_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0919__B1_N _0918_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_126 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0873__B1 _0854_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_281 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0625__B1 _0603_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_62 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0614__A _1145_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_95 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1050__B1 _1049_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0928__A1 _1187_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_130 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_229 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0987__C _0991_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0524__A _0581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0919__A1 _1181_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1041__B1 _1037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1220__CLK _1226_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_262 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1074__B _1055_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_234 VGND VPWR sky130_fd_sc_hd__fill_1
X_0519_ _0518_/X _0540_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_100_256 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_140 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0855__B1 _0854_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_284 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_107 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0609__A _0723_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_73 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_84 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_170 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_162 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1150__D _1158_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0870_ _0869_/Y _0839_/X _0848_/Y _0870_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_70_93 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1023__B1 _1019_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_254 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0519__A _0518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_118 VGND VPWR sky130_fd_sc_hd__fill_2
X_0999_ _0953_/Y _1000_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0701__B _0701_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1116__CLK _1223_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0611__B _0597_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1145__D d_sram_out[30] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_107 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0819__B1 _0679_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_173 VGND VPWR sky130_fd_sc_hd__fill_2
X_0922_ _0922_/A _0922_/B _0922_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_0853_ _0827_/A _0946_/A _0844_/X _0852_/X _0854_/A VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_60_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_0784_ _0722_/D _0711_/X _0783_/X _0784_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0521__B _0740_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0770__A2 _1089_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1055__D _1045_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1139__CLK _1089_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_213 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_19 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_257 VGND VPWR sky130_fd_sc_hd__fill_2
X_1198_ addr_w[0] baseaddr_w_sync[0] _1198_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_198 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0746__C1 _0745_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_88 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0761__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_184 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_154 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0622__A _0499_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_270 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0752__A2 _0751_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1121_ d_sram_out[6] _1121_/Q _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1052_ _1044_/X _1015_/X _1048_/Y _1052_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_92_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_0905_ _0861_/A _0904_/X _0905_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__0532__A _0532_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0836_ _0835_/A _0943_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_127_281 VGND VPWR sky130_fd_sc_hd__decap_12
X_0767_ _1121_/Q _0659_/A _0709_/X _0767_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1066__C _1056_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0698_ _0697_/A _0700_/B _0594_/B _0584_/D _0699_/D VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_102_137 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1082__B web VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_249 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_105 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_154 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_127 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_198 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0967__C1 _0960_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_98 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_76 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_98 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0734__A2 _1085_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_7 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0617__A _0597_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_146 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_61 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0621_ _0591_/X _0619_/X _0620_/X _0621_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_124_251 VGND VPWR sky130_fd_sc_hd__decap_12
X_0552_ _1154_/Q _0591_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_97_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_1104_ _0675_/D _1104_/Q _1197_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0527__A _0581_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1035_ _1034_/X _1035_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_21_113 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_179 VGND VPWR sky130_fd_sc_hd__decap_4
X_0819_ _0813_/X _1112_/Q _0679_/D _0815_/X d_fabric_out[29] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_115_284 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_46 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_23 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_271 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_97 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0707__A2 _0622_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_105 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1153__D _1161_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_216 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_219 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_293 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0604_ _0557_/X _0639_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_0535_ _0535_/A _0725_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0615__A2_N _0576_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_227 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_193 VGND VPWR sky130_fd_sc_hd__decap_3
X_1018_ _1017_/X _1018_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0704__B _0704_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0937__A2 _0932_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0720__A _0720_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_105 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0873__A1 _0872_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0625__A1 _0614_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_293 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0625__B2 _0571_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_140 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1050__A1 _0942_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0928__A2 _0926_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1148__D _1148_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0630__A _0594_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0987__D _1045_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_93 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1172__CLK _1221_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0524__B _0544_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0919__A2 _0907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1041__A1 _0945_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0540__A _0542_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_274 VGND VPWR sky130_fd_sc_hd__fill_1
X_0518_ _0517_/X _0518_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1074__C _0973_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_268 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0855__A1 _0851_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0791__B1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1195__CLK _1198_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_52 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0609__B _0594_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1023__A1 _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0782__B1 _0762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_141 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0535__A _0535_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_0998_ _0968_/A _0998_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_117_176 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_165 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0773__B1 _0719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0701__C _0701_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_211 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_204 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_165 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_154 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_86 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_97 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0764__B1 _0763_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0611__C _0611_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_203 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0819__A1 _0813_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1161__D _1224_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0819__B2 _0815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1210__CLK _1188_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0921_ _0880_/A _0875_/A _0920_/X d_sram_in[16] VGND VPWR sky130_fd_sc_hd__a21o_4
X_0852_ _0851_/A _0852_/B _0852_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0783_ _0720_/A _0750_/A _0783_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_53_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_281 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0521__C _0738_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_233 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_152 VGND VPWR sky130_fd_sc_hd__fill_1
X_1197_ d_fabric_in[31] _1197_/Q _1197_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_83_269 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_174 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_100 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_144 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0746__B1 _0651_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_247 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_291 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_41 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0903__A _0903_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0622__B _0488_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1156__D _0841_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_251 VGND VPWR sky130_fd_sc_hd__decap_12
X_1120_ d_sram_out[5] _0584_/D _1214_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_76_93 VGND VPWR sky130_fd_sc_hd__decap_12
X_1051_ _0965_/X _1043_/X _1049_/X w_mask[17] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_65_258 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_291 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0813__A _0662_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0904_ _1170_/Q _0890_/X _0903_/X _0904_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0976__B1 _0975_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0835_ _0835_/A _0883_/A _1042_/C _0838_/A VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__0532__B _0717_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1106__CLK _1126_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_293 VGND VPWR sky130_fd_sc_hd__decap_6
X_0766_ _0609_/X _0765_/X _0719_/X _0766_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0697_ _0697_/A _0700_/B _0580_/C _1122_/Q _0699_/C VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_102_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_193 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_160 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0900__B1 _0899_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_122 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0723__A _0740_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0967__B1 _0946_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_208 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_63 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_85 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_111 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_8 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0617__B _0616_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_125 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1129__CLK _1214_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0633__A _0725_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_84 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0958__B1 _0875_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0620_ _0499_/A _1147_/Q _0499_/C _0620_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_0551_ _0509_/X _0546_/Y _0550_/X _0551_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_124_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_263 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_1103_ _0542_/D _1103_/Q _1089_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0808__A _0776_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1034_ _0949_/A _0956_/X _1000_/C _1031_/D _1034_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0527__B _0556_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0543__A _1107_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8_0_clk_A clkbuf_4_9_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0818_ _0813_/X _1111_/Q _0532_/A _0815_/X d_fabric_out[28] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_115_230 VGND VPWR sky130_fd_sc_hd__decap_12
X_0749_ _0663_/X _0747_/X _0748_/X d_fabric_out[3] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_115_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_35 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0718__A _0718_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_291 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_99 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_136 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_158 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_129 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_228 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0628__A _0580_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_0603_ _0532_/A _0603_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_98_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_0534_ _0533_/X _0535_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_117 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_139 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0538__A _0581_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1017_ _0973_/A _0982_/B _1017_/C _1017_/D _1017_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_34_250 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0704__C _0699_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0720__B _0737_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_233 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0873__A2 _0838_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_194 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_31 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0625__A2 _0529_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_53 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_152 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1050__A2 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1164__D web VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1041__A2 _1040_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0540__B _0738_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0517_ _0517_/A _0517_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1074__D _1045_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_172 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0855__A2 _0839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_111 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_5_0_clk_A clkbuf_3_5_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0791__A1 _0713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0791__B2 _1095_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_231 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_106 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_97 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_120 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_186 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_257 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1159__D _1222_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0641__A _0697_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1023__A2 _1022_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0782__A1 _0779_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0782__B2 _1092_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_289 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_175 VGND VPWR sky130_fd_sc_hd__fill_2
X_0997_ _0968_/X _0995_/X _0996_/X w_mask[6] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0773__A1 _0771_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0701__D _1132_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_161 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0726__A _0510_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1162__CLK _1162_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_188 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0764__A1 _0762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0819__A2 _1112_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_62 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0636__A _0675_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_123 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_167 VGND VPWR sky130_fd_sc_hd__fill_2
X_0920_ _1182_/Q _0875_/Y _0920_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0851_ _0851_/A _0851_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0782_ _0779_/X _0781_/X _0762_/X _1092_/Q d_fabric_out[9] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__0521__D _1127_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_158 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_237 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_142 VGND VPWR sky130_fd_sc_hd__fill_2
X_1196_ d_fabric_in[30] _1196_/Q _1223_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_36_186 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0546__A _0509_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_167 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1185__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_217 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_208 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0746__A1 _1118_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_201 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_204 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_77 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_237 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_101 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_270 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0903__B _0903_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_2_0_clk_A clkbuf_2_2_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0622__C _0499_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0902__B1_N _0901_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_204 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1172__D d_fabric_in[6] VGND VPWR sky130_fd_sc_hd__diode_2
X_1050_ _0942_/A _1043_/X _1049_/X w_mask[16] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_80_229 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_93 VGND VPWR sky130_fd_sc_hd__decap_8
X_0903_ _0903_/A _0903_/B _0903_/C _1178_/Q _0903_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0976__A1 _0968_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0834_ _0834_/A _0883_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_0765_ _0614_/Y _0529_/A _0668_/X _0724_/D _0765_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_0696_ _0518_/X _0701_/B _0702_/C _0742_/D _0699_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_102_117 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_4_0_clk_A clkbuf_3_2_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0900__A1 _0851_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_229 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_107 VGND VPWR sky130_fd_sc_hd__decap_3
X_1179_ d_fabric_in[13] _1179_/Q _1221_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_24_145 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_118 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0723__B _0740_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0967__A1 _0945_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_250 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_253 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1200__CLK _1126_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_123 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_262 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0914__A _0897_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0633__B _0702_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1080__B1 _1079_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0958__A1 _0883_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1167__D d_fabric_in[1] VGND VPWR sky130_fd_sc_hd__diode_2
X_0550_ _0549_/Y _0550_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_137 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_93 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_1102_ _1134_/Q _1102_/Q _1132_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_53_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_229 VGND VPWR sky130_fd_sc_hd__fill_2
X_1033_ _0945_/A _1032_/X _1029_/Y w_mask[13] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0824__A _0841_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1071__B1 _1066_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_209 VGND VPWR sky130_fd_sc_hd__fill_1
X_0817_ _0813_/X _1110_/Q _0739_/D _0815_/X d_fabric_out[27] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1223__CLK _1223_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_220 VGND VPWR sky130_fd_sc_hd__decap_3
X_0748_ _0733_/A _1086_/Q _0748_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0679_ _0722_/A _0738_/B _0544_/C _0679_/D _0679_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_88_126 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_47 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_207 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0718__B _0716_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_148 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1062__B1 _1061_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0628__B _0701_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0644__A _0533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1053__B1 _1052_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_170 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0800__B1 _0799_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_0602_ _0697_/A _0701_/B _0702_/C _0602_/D _0612_/B VGND VPWR sky130_fd_sc_hd__and4_4
X_0533_ _0533_/A _0533_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_256 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0867__B1 _0866_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_281 VGND VPWR sky130_fd_sc_hd__decap_12
X_1016_ _0998_/X _1015_/X _1012_/X w_mask[9] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0554__A _0737_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_262 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0704__D _0704_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0729__A _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1119__CLK _1109_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_clk_A clkbuf_3_1_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_22 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_12_0_clk_A clkbuf_3_6_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0639__A _0723_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0849__B1 _0848_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1180__D d_fabric_in[14] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_121 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_154 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_3 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0540__C _0540_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0516_ _0504_/A _0517_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_100_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0549__A _0549_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1090__D _0775_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_110 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_198 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_19 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_178 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0791__A2 _1095_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_114 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1091__CLK _1126_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_132 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_154 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_165 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_198 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0922__A _0922_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0641__B _0700_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0782__A2 _0781_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1175__D d_fabric_in[9] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_198 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0832__A _0831_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0996_ _0985_/X _0979_/X _0988_/Y _0996_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_117_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0773__A2 _0772_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1085__D _1085_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_246 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_173 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0726__B _0513_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_56 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0742__A _0576_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_66 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0764__A2 _1088_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_268 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_132 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0636__B _0702_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_146 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0652__A _0542_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0850_ _0830_/Y _0833_/X _0849_/X d_sram_in[2] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0781_ _0674_/A _0496_/X _0676_/D _0496_/X _0781_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_39_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_205 VGND VPWR sky130_fd_sc_hd__fill_2
X_1195_ d_fabric_in[29] _1195_/Q _1198_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0827__A _0827_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_165 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0546__B _0546_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_179 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0562__A _0561_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_229 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_0_0_clk_A clkbuf_4_0_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0979_ _0979_/A _0979_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0746__A2 _0549_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_235 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0737__A _0737_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_77 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_99 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_54 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0903__C _0903_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_76 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_84 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_121 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0647__A _0647_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_165 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_157 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_179 VGND VPWR sky130_fd_sc_hd__fill_2
X_0902_ _1177_/Q _0877_/X _0901_/Y d_sram_in[11] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0976__A2 _0974_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0833_ _0875_/A _0833_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0764_ _0762_/X _1088_/D _0763_/X d_fabric_out[5] VGND VPWR sky130_fd_sc_hd__a21o_4
X_0695_ _1134_/Q _0742_/D VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_110_173 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_205 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_238 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0900__A2 _0890_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0557__A _0556_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1152__CLK _1223_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_1178_ d_fabric_in[12] _1178_/Q _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_24_102 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_271 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_190 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0723__C _0722_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0967__A2 _0966_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_68 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_32 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_219 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_293 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_64 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0914__B _0913_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_296 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_138 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1080__A1 _1035_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0958__A2 _0841_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_127 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1183__D d_fabric_in[17] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1175__CLK _1221_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_1101_ _0725_/D _1101_/Q _1132_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0894__A1 _0891_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1032_ _1031_/X _1032_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_61_241 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_149 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1071__A1 _0985_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1001__A _1000_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0816_ _0813_/X _1109_/Q _0722_/D _0815_/X d_fabric_out[26] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__0840__A _1228_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0747_ _0750_/A _0736_/X _0746_/X _0742_/D _0496_/A _0747_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_130_202 VGND VPWR sky130_fd_sc_hd__decap_12
X_0678_ _1112_/D _0679_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1093__D _0784_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0718__C _0501_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_68 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_296 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1062__A1 _0995_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0750__A _0750_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1198__CLK _1198_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0573__B1 _1121_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_31 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_74 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0644__B _0565_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1053__A1 _0974_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1178__D d_fabric_in[12] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_160 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0800__B2 _1098_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0800__A1 _0713_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0601_ _0582_/X _0702_/C VGND VPWR sky130_fd_sc_hd__buf_1
X_0532_ _0532_/A _0717_/B _0532_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_98_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_268 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0867__A1 _0864_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_163 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_174 VGND VPWR sky130_fd_sc_hd__decap_3
X_1015_ _1014_/X _1015_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0835__A _0835_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_296 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1088__D _1088_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0570__A _0570_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_257 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0729__B _0720_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_34 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_208 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0745__A _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_99 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_187 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0794__B1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0639__B _0639_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0849__A1 _0830_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1213__CLK _1226_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0655__A _0655_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_132 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_3 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0540__D _0642_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_222 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0537__B1 _0675_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0515_ _0738_/B _0740_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0565__A _0565_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_44 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_144 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0922__B _0922_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0767__B1 _0709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0641__C _0702_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_236 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1191__D d_fabric_in[25] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_258 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_163 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1109__CLK _1109_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0995_ _0994_/X _0995_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_117_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0758__B1 _0687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_144 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_188 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0726__C _1145_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0742__B _0544_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0997__B1 _0996_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0749__B1 _0748_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_56 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_203 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0921__B1 _0920_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_75 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0636__C _0636_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_177 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_136 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_74 VGND VPWR sky130_fd_sc_hd__decap_12
X_0780_ _0779_/X _0778_/X _0762_/X _1091_/Q d_fabric_out[8] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1186__D d_fabric_in[20] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_7 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_203 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_247 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_258 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_217 VGND VPWR sky130_fd_sc_hd__fill_2
X_1194_ d_fabric_in[28] _1194_/Q _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1004__A _1031_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0546__C _0546_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_29 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0843__A _1044_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0978_ _0973_/A _0991_/B _1017_/C _0991_/D _0979_/A VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__1096__D _0793_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_133 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0737__B _0737_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_291 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_158 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_180 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_33 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0903__D _1178_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_193 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0647__B _0639_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_177 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_261 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0663__A _0662_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_191 VGND VPWR sky130_fd_sc_hd__decap_12
X_0901_ _0854_/A _0901_/B _0901_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_0832_ _0831_/X _0875_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_127_241 VGND VPWR sky130_fd_sc_hd__decap_3
X_0763_ _0733_/A _1088_/Q _0763_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0694_ _0535_/A _0700_/B _0582_/X _0737_/A _0694_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_51_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0838__A _0838_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_185 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_93 VGND VPWR sky130_fd_sc_hd__fill_2
X_1177_ d_fabric_in[11] _1177_/Q _1226_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_24_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_114 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_158 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_109 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0723__D _0723_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_7 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_277 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0748__A _0733_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_10 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_32 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1080__A2 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_51 VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_9_0_clk clkbuf_4_9_0_clk/A _1150_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_87_62 VGND VPWR sky130_fd_sc_hd__decap_4
X_1100_ _1132_/Q _1100_/Q _1132_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_38_239 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0894__A2 _0877_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1031_ _1031_/A _1021_/B _1000_/C _1031_/D _1031_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_46_261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_264 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1071__A2 _1032_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_200 VGND VPWR sky130_fd_sc_hd__decap_12
X_0815_ out_reg _0815_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0746_ _1118_/Q _0549_/A _0651_/Y _0745_/X _0746_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_0677_ _0668_/A _0669_/X _0738_/C _0584_/D _0684_/C VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0718__D _0717_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_242 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1062__A2 _1059_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_106 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0573__B2 _0587_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0573__A1 _0642_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_109 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_31 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0644__C _0584_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0941__A _0940_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1053__A2 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_143 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_165 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0800__A2 _1098_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1142__CLK _1223_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0600_ _0645_/A _0697_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0531_ _0580_/C _0717_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1194__D d_fabric_in[28] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0867__A2 _0839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_172 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_142 VGND VPWR sky130_fd_sc_hd__fill_2
X_1014_ _0982_/A _1021_/B _1017_/C _1017_/D _1014_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0835__B _0883_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0851__A _0851_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0570__B _1150_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_0729_ _0550_/X _0720_/X _0728_/X _0729_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_134_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_109 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_291 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0729__C _0728_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_46 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0745__B _0737_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_23 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_67 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1165__CLK _1197_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_199 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0794__B2 _1096_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0794__A1 _0713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0849__A2 _0839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_153 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_175 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0655__B _0655_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_145 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_212 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_270 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1189__D d_fabric_in[23] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_144 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0537__A1 _0526_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0514_ _0513_/X _0738_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_100_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1007__A _1031_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0915__B1_N _0914_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_186 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0846__A _0846_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1188__CLK _1188_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1099__D _0655_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0581__A _0581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0491__A _0544_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0767__A1 _1121_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0641__D _1117_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_98 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_182 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_0994_ _0949_/A _0956_/X _0953_/Y _0972_/A _0994_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0758__A1 _0668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_117 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_139 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0930__A1 _1189_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_259 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0576__A _0517_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_123 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0726__D _0725_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0997__A1 _0968_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0742__C _0725_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_125 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0749__A1 _0663_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1203__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_66 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0921__A1 _0880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0486__A reb VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_207 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0685__B1 _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_126 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_215 VGND VPWR sky130_fd_sc_hd__decap_4
X_1193_ d_fabric_in[27] _1193_/Q _1221_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_36_112 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0546__D _0546_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_137 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1226__CLK _1226_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0977_ _0977_/A _1017_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_10_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_69 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_123 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_178 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_126 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0647__C _0641_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_145 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0658__B1 _0651_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_189 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0944__A _0968_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__decap_3
X_0900_ _0851_/A _0890_/X _0899_/X _0901_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_41_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1197__D d_fabric_in[31] VGND VPWR sky130_fd_sc_hd__diode_2
X_0831_ _1226_/Q _0841_/B _1042_/C _0831_/X VGND VPWR sky130_fd_sc_hd__or3_4
X_0762_ _0662_/X _0762_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0693_ _0676_/D _0627_/Y _0692_/X _0704_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0838__B _0838_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1015__A _1014_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_281 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0649__B1 _0648_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1176_ d_fabric_in[10] _0895_/D _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0854__A _0854_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0821__B1 _0616_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_289 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_218 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0748__B _1086_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_197 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_240 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_276 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_88 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0812__B1 _0544_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_96 VGND VPWR sky130_fd_sc_hd__fill_2
X_1030_ _0945_/A _1025_/X _1029_/Y w_mask[12] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_46_273 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0674__A _0674_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0803__B1 _0681_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0814_ _0813_/X _1108_/Q _0676_/D _0808_/X d_fabric_out[25] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_115_212 VGND VPWR sky130_fd_sc_hd__decap_8
X_0745_ _0550_/X _0737_/X _0744_/X _0745_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_115_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_245 VGND VPWR sky130_fd_sc_hd__decap_8
X_0676_ _0521_/A _0492_/C _0675_/C _0676_/D _0684_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_130_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_195 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0781__A2_N _0496_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1228_ conf[2] _1228_/Q _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_16_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0584__A _0533_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1159_ _1222_/Q _1159_/Q _1198_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1047__B1 _0958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0573__A2 _0524_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1094__CLK _1089_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_184 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0730__C1 _0729_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_251 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0494__A _0493_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_43 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0644__D _0720_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1038__B1 _1037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_177 VGND VPWR sky130_fd_sc_hd__decap_6
X_0530_ _0643_/C _0580_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0669__A _0740_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1013_ _0998_/X _1006_/X _1012_/X w_mask[8] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_93_198 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0835__C _1042_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_93 VGND VPWR sky130_fd_sc_hd__decap_12
X_0728_ _0721_/X _0722_/X _0723_/X _0728_/D _0728_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_103_237 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_226 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0579__A _0533_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0659_ _0659_/A _0658_/Y _0659_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_134_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_154 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_232 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0745__C _0744_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_198 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_35 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_8_0_clk clkbuf_4_9_0_clk/A _1221_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_138_156 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0794__A2 _0793_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_158 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0489__A _1150_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_98 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_224 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0952__A _0955_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_260 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_271 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_123 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_156 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0537__A2 _0532_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_235 VGND VPWR sky130_fd_sc_hd__fill_2
X_0513_ _0513_/A _0513_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_100_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_176 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0846__B _0852_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0581__B _1150_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_235 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_132 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_23 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1132__CLK _1132_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0767__A2 _0659_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_92 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_216 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0947__A _0962_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_179 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0682__A _0722_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0993_ _0968_/X _0992_/X _0989_/X w_mask[5] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_74_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0758__A2 _1128_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_159 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1018__A _1017_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0930__A2 _0926_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_238 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0857__A _1170_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1155__CLK _1150_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0576__B _0565_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_15 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0592__A _0569_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0997__A2 _0995_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0742__D _0742_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0749__A2 _0747_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_151 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0921__A2 _0875_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_216 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0486__B csb VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0685__A1 _0674_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_94 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1178__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0929__B1_N _0870_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0677__A _0668_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1192_ d_fabric_in[26] _1192_/Q _1221_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_76_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_146 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_274 VGND VPWR sky130_fd_sc_hd__decap_12
X_0976_ _0968_/X _0974_/X _0975_/Y w_mask[2] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_59_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0587__A _0517_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_208 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_252 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_274 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_201 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_173 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0497__A _0497_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_102 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0647__D _0646_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_271 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0658__A1 _0501_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0658__B2 _0657_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_116 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_190 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_80 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_160 VGND VPWR sky130_fd_sc_hd__fill_2
X_0830_ _0846_/A _0830_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0960__A _0960_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_221 VGND VPWR sky130_fd_sc_hd__decap_12
X_0761_ _0675_/D _0750_/X _0759_/X _0760_/X _1088_/D VGND VPWR sky130_fd_sc_hd__o22a_4
X_0692_ _0739_/D _0558_/X _0692_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_37_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_154 VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0_clk clkbuf_0_clk/X clkbuf_2_2_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0649__A1 _0626_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_293 VGND VPWR sky130_fd_sc_hd__decap_6
X_1175_ d_fabric_in[9] _0891_/D _1221_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_296 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1031__A _1031_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0821__B2 _0779_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0821__A1 _0662_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_0959_ _1055_/B _0838_/B _0958_/X _0960_/C VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_118_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_165 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_127 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_266 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_288 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0812__A1 _0806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0812__B2 _0808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_108 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1216__CLK _1197_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0955__A _0955_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0674__B _0509_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_233 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0690__A _0544_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0803__A1 _0799_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0803__B2 _0801_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0813_ _0662_/A _0813_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0744_ _0738_/X _0744_/B _0740_/X _0743_/X _0744_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_0675_ _0740_/A _0669_/X _0675_/C _0675_/D _0675_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_130_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_208 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1026__A _0985_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1227_ conf[1] _0841_/B _1188_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1158_ _1158_/D _1158_/Q _1221_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0584__B _0565_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_222 VGND VPWR sky130_fd_sc_hd__fill_2
X_1089_ _1089_/D _1089_/Q _1089_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1047__A1 _1045_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_152 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0730__B1 _0719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_55 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_77 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1038__A1 _0945_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_174 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_1012_ _0985_/X _0983_/X _1011_/Y _1012_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_93_166 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0788__B1 _0739_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0727_ _0507_/Y _0724_/X _0727_/C _0726_/X _0728_/D VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0579__B _0580_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0658_ _0501_/X _0551_/Y _0650_/X _0651_/Y _0657_/X _0658_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
X_0589_ _0579_/X _0580_/X _0583_/X _0588_/X _0589_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XANTENNA__0712__B1 _0681_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0595__A _1132_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_168 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_126 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_92 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0952__B _0991_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_288 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_261 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_236 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_272 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_168 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_91 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0795__A2_N _0787_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0512_ _0722_/A _0521_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_66_111 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_136 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1084__CLK _1089_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_127 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_214 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_291 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_166 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_79 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_291 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_98 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0963__A _0963_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0682__B _0738_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0992_ _0991_/X _0992_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_8_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_62 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_7_0_clk clkbuf_4_7_0_clk/A _1223_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0576__C _0576_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1034__A _0949_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_188 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_180 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_163 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0685__A2 _0684_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_67 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0783__A _0720_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0677__B _0669_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1191_ d_fabric_in[25] _1191_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0765__A1_N _0614_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_209 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_286 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_191 VGND VPWR sky130_fd_sc_hd__fill_2
X_0975_ _0946_/A _0966_/Y _0960_/X _0975_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__1122__CLK _1126_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1029__A _0960_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_174 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0587__B _1153_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_141 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0658__A2 _0551_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_70 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_70 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0960__B _0955_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_233 VGND VPWR sky130_fd_sc_hd__decap_8
X_0760_ _0584_/D _0496_/A _0709_/X _0760_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1145__CLK _1197_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0691_ _1142_/Q _0739_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0688__A _0607_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_209 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0649__A2 _0632_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1174_ d_fabric_in[8] _0887_/D _1221_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1031__B _1021_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0821__A2 _1114_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_211 VGND VPWR sky130_fd_sc_hd__decap_3
X_0958_ _0883_/A _0841_/C _0875_/A _0958_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_21_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_214 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_288 VGND VPWR sky130_fd_sc_hd__decap_8
X_0889_ _0887_/D _0877_/X _0888_/Y d_sram_in[8] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_99_172 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0598__A _0569_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_201 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_139 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_234 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0928__B1_N _0867_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1168__CLK _1223_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_68 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0812__A2 _1107_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_87 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0955__B _0991_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_109 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_172 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0971__A _0977_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0690__B _0597_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0803__A2 _1100_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0812_ _0806_/X _1107_/Q _0544_/D _0808_/X d_fabric_out[24] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0743_ _0616_/X _0509_/B _0743_/C _0742_/X _0743_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_0674_ _0674_/A _0509_/B _0674_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_130_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_291 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1026__B _0995_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_175 VGND VPWR sky130_fd_sc_hd__decap_4
X_1226_ conf[0] _1226_/Q _1226_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1157_ _1228_/Q _1149_/D _1162_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0584__C _0584_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1042__A _0899_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1088_ _1088_/D _1088_/Q _1089_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0881__A _0835_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1047__A2 _0838_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_131 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_7 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_269 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_57 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0730__A1 _1117_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_74 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_245 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1102__D _1134_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1038__A2 _1035_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_131 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_135 VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0_clk clkbuf_0_clk/X clkbuf_1_0_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_22_93 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_239 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0966__A _0965_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_164 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_220 VGND VPWR sky130_fd_sc_hd__fill_2
X_1011_ _1009_/X _1028_/A _0960_/C _1011_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_97_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0788__B2 _0787_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0726_ _0510_/X _0513_/X _1145_/Q _0725_/C _0726_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_103_206 VGND VPWR sky130_fd_sc_hd__fill_2
X_0657_ _0668_/A _0502_/A _0655_/X _0656_/X _0657_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__0579__C _0569_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0588_ _0584_/X _0588_/B _0586_/X _0588_/D _0588_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_69_131 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0712__A1 _0750_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0876__A _0875_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0712__B2 _0711_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0595__B _0582_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_145 VGND VPWR sky130_fd_sc_hd__fill_2
X_1209_ addr_w[11] _0977_/A _1150_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_125 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_105 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1206__CLK _1221_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_104 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_251 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0952__C _0952_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_273 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_204 VGND VPWR sky130_fd_sc_hd__fill_2
X_0511_ _0510_/X _0722_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_3_171 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0696__A _0518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0933__A1 _1191_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0709_ _0501_/X _0709_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_36 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_192 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_117 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0621__B1 _0620_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_22 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0924__A1 _1184_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_270 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_137 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0682__C _0540_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0991_ _0982_/A _0991_/B _0991_/C _0991_/D _0991_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0860__B1 _0880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_296 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0915__A1 _0912_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_207 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_134 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0576__D _0513_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_251 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1034__B _0956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_284 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_148 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1200__D addr_w[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_117 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0906__A1 _1178_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_175 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_137 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0783__B _0750_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_170 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1110__D _1142_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_229 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0677__C _0738_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_91 VGND VPWR sky130_fd_sc_hd__decap_8
X_1190_ d_fabric_in[24] _1190_/Q _1197_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_76_240 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0974__A _0973_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_298 VGND VPWR sky130_fd_sc_hd__fill_1
X_0974_ _0973_/X _0974_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1029__B _1029_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0587__C _0587_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1045__A _0955_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0884__A _0903_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_107 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1077__B1 _1076_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_37 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_234 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1097__CLK _1089_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1105__D _0723_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0658__A3 _0650_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_265 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_22 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1068__B1 _1067_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_60 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_60 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_173 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_93 VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_6_0_clk clkbuf_4_7_0_clk/A _1132_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0960__C _0960_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_0690_ _0544_/C _0597_/B _0690_/C _0679_/D _0704_/A VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0969__A _0969_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0688__B _0687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_97 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0649__A3 _0636_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1173_ d_fabric_in[7] _1173_/Q _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_170 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1031__C _1000_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_162 VGND VPWR sky130_fd_sc_hd__fill_2
X_0957_ _0956_/X _1055_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0888_ _0888_/A _0887_/X _0861_/A _0888_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_133_226 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0879__A _0952_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_14 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0955__C _0991_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1112__CLK _1214_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_162 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_184 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0690__C _0690_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0811_ _0806_/X _1106_/Q _0740_/D _0808_/X d_fabric_out[23] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0742_ _0576_/C _0544_/B _0725_/C _0742_/D _0742_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_115_226 VGND VPWR sky130_fd_sc_hd__fill_2
X_0673_ _0583_/D _0674_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0699__A _0694_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_154 VGND VPWR sky130_fd_sc_hd__fill_2
X_1225_ addr_r[13] _1225_/Q _1198_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_243 VGND VPWR sky130_fd_sc_hd__fill_1
X_1156_ _0841_/B _1148_/D _1162_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0584__D _0584_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1042__B _0899_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1087_ _0754_/X _1087_/Q _1089_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_20_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0730__A2 _0549_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1135__CLK _1132_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_276 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_94 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_146 VGND VPWR sky130_fd_sc_hd__fill_2
X_1010_ _0949_/A _0956_/X _0952_/C _1028_/A VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_93_179 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0982__A _0982_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_180 VGND VPWR sky130_fd_sc_hd__decap_12
X_0725_ _0576_/C _0544_/B _0725_/C _0725_/D _0727_/C VGND VPWR sky130_fd_sc_hd__and4_4
X_0656_ _0544_/D _0717_/B _0656_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0579__D _1130_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0927__B1_N _0862_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1158__CLK _1221_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0587_ _0517_/X _1153_/Q _0587_/C _0720_/A _0588_/D VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_69_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_240 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0712__A2 _0672_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1208_ addr_w[10] _0962_/A _1150_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1203__D addr_w[5] VGND VPWR sky130_fd_sc_hd__diode_2
X_1139_ d_sram_out[24] _1107_/D _1089_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_137 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_179 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1113__D _1145_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_252 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_181 VGND VPWR sky130_fd_sc_hd__fill_2
X_0510_ _0510_/A _0510_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0977__A _0977_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0696__B _0701_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_205 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1048__A _1045_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0933__A2 _0932_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0708_ _0705_/X _0706_/Y _0707_/X _0708_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_89_205 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_238 VGND VPWR sky130_fd_sc_hd__fill_2
X_0639_ _0723_/D _0639_/B _0639_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0887__A _0899_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_113 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_146 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_171 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0621__A1 _0591_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_34 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0924__A2 _0907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1108__D _0602_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0797__A _0616_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_95 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_102 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_93 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0682__D _1128_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0990_ _0968_/X _0983_/X _0989_/X w_mask[4] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0860__A1 _0826_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0915__A2 _0907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0500__A _0499_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_113 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_168 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1034__C _1000_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_110 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0906__A2 _0877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_119 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_86 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_219 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1219__CLK _1128_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0677__D _0584_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_285 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_108 VGND VPWR sky130_fd_sc_hd__decap_3
X_0973_ _0973_/A _0982_/B _0973_/C _0991_/D _0973_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_72_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1029__C _1028_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0587__D _0720_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1045__B _1045_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_244 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_266 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1077__A1 _1025_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1211__D addr_w[13] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_27 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_246 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_154 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0760__B1 _0709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_68 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_296 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1068__A1 _1006_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_171 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_61 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1121__D d_sram_out[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_152 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_94 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_82 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0751__B1 _0635_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0985__A _0985_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1191__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1172_ d_fabric_in[6] _1172_/Q _1221_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0649__A4 _0647_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_244 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1031__D _1031_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0956_ _0970_/A _0956_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0887_ _0899_/A _0899_/B _0903_/C _0887_/D _0887_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_133_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_238 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0990__B1 _0989_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1056__A _1056_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0895__A _0899_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1206__D addr_w[8] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_26 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_258 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_163 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_74 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1116__D d_sram_out[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_200 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0955__D _0955_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0690__D _0679_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0810_ _0806_/X _1105_/Q _0723_/D _0808_/X d_fabric_out[22] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0741_ _0510_/X _0513_/X _0724_/C _1130_/Q _0743_/C VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0699__B _0699_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0672_ _0668_/X _0583_/D _0501_/X _0671_/X _0672_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_35_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_1224_ addr_r[12] _1224_/Q _1128_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1155_ _1226_/Q _1155_/Q _1150_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_203 VGND VPWR sky130_fd_sc_hd__fill_2
X_1086_ _0747_/X _1086_/Q _1162_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1042__C _1042_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_247 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1087__CLK _1089_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_166 VGND VPWR sky130_fd_sc_hd__decap_12
X_0939_ _1197_/Q _0922_/B _0918_/Y d_sram_in[31] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_121_208 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0715__B1 _0714_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_15 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_5_0_clk clkbuf_3_2_0_clk/X _1188_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_113_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_288 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_100 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_293 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0706__B1 _0622_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_122 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_177 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0982__B _0982_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0724_ _0510_/X _0513_/X _0724_/C _0724_/D _0724_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0503__A _1150_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_192 VGND VPWR sky130_fd_sc_hd__decap_12
X_0655_ _0655_/A _0655_/B _0655_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0586_ _0517_/A _0565_/A _0587_/C _1117_/Q _0586_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_69_177 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0712__A3 _0710_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_169 VGND VPWR sky130_fd_sc_hd__fill_2
X_1207_ addr_w[9] _0970_/A _1150_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_236 VGND VPWR sky130_fd_sc_hd__decap_8
X_1138_ d_sram_out[23] _0740_/D _1223_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1069_ _1015_/X _1059_/X _1067_/X w_mask[25] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_25_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_239 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0778__A1_N _0509_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1102__CLK _1132_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_169 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_180 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_239 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0696__C _0702_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0577__A2_N _0576_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_119 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1125__CLK _1109_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0707_ _0585_/D _0622_/Y _0550_/X _0707_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1048__B _1056_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0638_ _0722_/D _0558_/X _0647_/A VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0887__B _0899_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0569_ _1153_/Q _0569_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1064__A _1007_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1214__D addr_r[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_206 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0621__A2 _0619_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0909__B1 _0908_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_46 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0797__B _0659_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1124__D d_sram_out[9] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0911__B1_N _0910_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0860__A2 _0859_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1148__CLK _1162_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0988__A _0960_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_283 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1034__D _1031_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_128 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1059__A _1043_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1209__D addr_w[11] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_49 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1119__D d_sram_out[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_84 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0601__A _0582_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_220 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_234 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_183 VGND VPWR sky130_fd_sc_hd__fill_2
X_0972_ _0972_/A _0991_/D VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_65_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0511__A _0510_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1045__C _0973_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_201 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1077__A2 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_258 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_177 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0760__A1 _0584_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_234 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1068__A2 _1059_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_40 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_62 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_73 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_214 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0751__A1 _0668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_44 VGND VPWR sky130_fd_sc_hd__decap_12
X_1171_ d_fabric_in[5] _1171_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_267 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0506__A _0506_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_186 VGND VPWR sky130_fd_sc_hd__fill_2
X_0955_ _0955_/A _0991_/B _0991_/C _0955_/D _0955_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0886_ _0908_/C _0903_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0990__A1 _0968_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_142 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1056__B _1056_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_197 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0895__B _0899_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_169 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_245 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1222__D addr_r[10] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_215 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1209__CLK _1150_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_269 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1132__D d_sram_out[17] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_237 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_93 VGND VPWR sky130_fd_sc_hd__fill_2
X_0740_ _0740_/A _0740_/B _0722_/C _0740_/D _0740_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0671_ _0521_/A _0669_/X _0676_/D _0681_/D _0655_/B _0671_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__0699__C _0699_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_3 VGND VPWR sky130_fd_sc_hd__decap_4
X_1223_ addr_r[11] _1223_/Q _1223_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_96_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_1154_ _1162_/Q _1154_/Q _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_226 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1042__D _1042_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1085_ _1085_/D _1085_/Q _1150_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_259 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_112 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_270 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_178 VGND VPWR sky130_fd_sc_hd__decap_12
X_0938_ _1196_/Q _0922_/B _0914_/Y d_sram_in[30] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_106_206 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_228 VGND VPWR sky130_fd_sc_hd__decap_8
X_0869_ _1172_/Q _0869_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1217__D addr_r[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0715__A1 _0663_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_112 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_204 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_123 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1181__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_63 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1127__D d_sram_out[12] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0706__A1 _0674_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_71 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_159 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0982__C _0991_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_81 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_32 VGND VPWR sky130_fd_sc_hd__decap_12
X_0723_ _0740_/A _0740_/B _0722_/C _0723_/D _0723_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0654_ _0690_/C _0655_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_0585_ _0517_/A _0565_/A _0584_/C _0585_/D _0588_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_69_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_253 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_7_0_clk_A clkbuf_4_7_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1206_ addr_w[8] baseaddr_w_sync[8] _1221_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_1137_ d_sram_out[22] _0723_/D _1214_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1068_ _1006_/X _1059_/X _1067_/X w_mask[24] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_33_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_106 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0936__A1 _1194_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_231 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_74 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_210 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_96 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_243 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_128 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_95 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0604__A _0557_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0927__A1 _1186_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0696__D _0742_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_115 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_137 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0863__B1 _0862_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_80 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0615__B1 _1112_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_251 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_4_0_clk clkbuf_3_2_0_clk/X _1089_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0514__A _0513_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0706_ _0674_/A _0703_/A _0622_/Y _0706_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__1048__C _1056_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0637_ _1141_/Q _0722_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0887__C _0903_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_240 VGND VPWR sky130_fd_sc_hd__fill_2
X_0568_ _0560_/Y _0562_/X _0567_/Y _0568_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__1064__B _1045_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0499_ _0499_/A _1147_/Q _0499_/C _0499_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_54_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_192 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_218 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_120 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0909__A1 _1171_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_98 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_86 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_148 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1140__D d_sram_out[25] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0988__B _0988_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_262 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_232 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0509__A _0509_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_195 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1013__B1 _1012_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_175 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1075__A _1066_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_39 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1225__D addr_r[13] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_140 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_4_0_clk_A clkbuf_3_5_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_15_0_clk_A clkbuf_3_7_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1135__D d_sram_out[20] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_210 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0818__B1 _0532_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1115__CLK _1197_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_173 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_195 VGND VPWR sky130_fd_sc_hd__decap_12
X_0971_ _0977_/A _0973_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0999__A _0953_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1045__D _1045_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_140 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0809__B1 _0675_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_279 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_132 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0702__A _0724_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0760__A2 _0496_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0925__B1_N _0855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1138__CLK _1223_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_265 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_257 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_268 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_30 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_52 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_41 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_165 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_85 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_62 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0612__A _0599_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_281 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0736__C1 _0735_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0751__A2 _1127_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_210 VGND VPWR sky130_fd_sc_hd__fill_2
X_1170_ d_fabric_in[4] _1170_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_2_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_121 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_91 VGND VPWR sky130_fd_sc_hd__fill_1
X_0954_ _0953_/Y _0991_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_118_226 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_215 VGND VPWR sky130_fd_sc_hd__decap_8
X_0885_ _0841_/C _0908_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0522__A _0510_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_270 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0990__A2 _0983_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1056__C _1056_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_115 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0895__C _0903_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_159 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_24 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_238 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_192 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_73 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_216 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_84 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0607__A _0740_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1_0_clk_A clkbuf_1_0_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_154 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_50 VGND VPWR sky130_fd_sc_hd__fill_2
X_0670_ _0602_/D _0676_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0699__D _0699_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1222_ addr_r[10] _1222_/Q _1198_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_96_179 VGND VPWR sky130_fd_sc_hd__fill_1
X_1153_ _1161_/Q _1153_/Q _1226_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_1084_ _0712_/X _0714_/B _1089_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0517__A _0517_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0660__A1 _0681_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0937_ _1195_/Q _0932_/X _0910_/Y d_sram_in[29] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA_clkbuf_4_3_0_clk_A clkbuf_4_3_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0868_ _0864_/Y _0833_/X _0867_/X d_sram_in[5] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0799_ _0662_/A _0799_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_114_240 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0715__A2 _0712_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_216 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0706__A2 _0703_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_224 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1143__D d_sram_out[28] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_50 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_257 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0982__D _0991_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_227 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_44 VGND VPWR sky130_fd_sc_hd__decap_12
X_0722_ _0722_/A _0492_/C _0722_/C _0722_/D _0722_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0653_ _0740_/A _0668_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_40_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_0584_ _0533_/A _0565_/A _0584_/C _0584_/D _0584_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_69_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_232 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_265 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_1205_ addr_w[7] baseaddr_w_sync[7] _1197_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_84_149 VGND VPWR sky130_fd_sc_hd__fill_2
X_1136_ d_sram_out[21] _0675_/D _1214_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_227 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_182 VGND VPWR sky130_fd_sc_hd__fill_2
X_1067_ _1044_/X _1025_/X _1066_/Y _1067_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_33_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_118 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0936__A2 _0932_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1228__D conf[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_22 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_116 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_200 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_86 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0927__A2 _0926_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1138__D d_sram_out[23] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_208 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0620__A _0499_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_60 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0863__A1 _0857_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0615__B2 _0558_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_296 VGND VPWR sky130_fd_sc_hd__decap_3
X_0705_ _0705_/A _0686_/X _0705_/C _0705_/D _0705_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0530__A _0643_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0636_ _0675_/C _0702_/B _0636_/C _0636_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0887__D _0887_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0567_ _0645_/A _0580_/B _0643_/C _1118_/Q _0567_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_57_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_116 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0551__B1 _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1064__C _0973_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_138 VGND VPWR sky130_fd_sc_hd__fill_2
X_0498_ _0498_/A _0499_/C VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1171__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_182 VGND VPWR sky130_fd_sc_hd__fill_1
X_1119_ d_sram_out[4] _0642_/D _1109_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_110_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0705__A _0705_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_132 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0909__A2 _0890_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_clk_A clkbuf_3_1_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0790__B1 _0532_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_241 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_85 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_171 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_11_0_clk_A clkbuf_3_5_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_196 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_61 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0988__C _0960_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0781__B1 _0676_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_92 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_105 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1194__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_255 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0509__B _0509_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_141 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_163 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0525__A _0655_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1013__A1 _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0772__B1 _0668_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0619_ _0619_/A _0619_/B _0619_/C _0619_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__1075__B _1074_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_64 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_190 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_3_0_clk clkbuf_4_3_0_clk/A _1126_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_76_244 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0818__A1 _0813_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0818__B2 _0815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_72 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1151__D _1159_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_258 VGND VPWR sky130_fd_sc_hd__fill_2
X_0970_ _0970_/A _0982_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0754__B1 _0752_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_157 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0809__B2 _0808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0809__A1 _0806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_196 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0993__B1 _0989_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0702__B _0702_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_108 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_214 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_31 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_97 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_75 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_177 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0612__B _0612_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_293 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0736__B1 _0501_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_240 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1146__D d_sram_out[31] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_222 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_203 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_247 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_174 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0672__C1 _0671_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_166 VGND VPWR sky130_fd_sc_hd__fill_1
X_0953_ _0977_/A _0953_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_118_238 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_0884_ _0903_/B _0899_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0975__B1 _0960_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_133 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_177 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_155 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0895__D _0895_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_291 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_133 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0713__A out_reg VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_11 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1105__CLK _1197_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_171 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_225 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_52 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0607__B _0643_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_84 VGND VPWR sky130_fd_sc_hd__fill_2
X_1221_ addr_r[9] _1158_/D _1221_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_203 VGND VPWR sky130_fd_sc_hd__decap_12
X_1152_ _1160_/Q _0504_/A _1223_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1083_ _0660_/X _1083_/Q _1109_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_269 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0660__A2 _0496_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1128__CLK _1128_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_170 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0924__B1_N _0849_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0533__A _0533_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0936_ _1194_/Q _0932_/X _0905_/Y d_sram_in[28] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0867_ _0864_/Y _0839_/X _0866_/Y _0867_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0798_ _1130_/Q _0750_/X _0797_/X _1098_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0939__B1_N _0918_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_169 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_228 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_87 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_125 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_147 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_158 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0618__A _0591_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_56 VGND VPWR sky130_fd_sc_hd__decap_12
X_0721_ _0740_/A _0740_/B _0738_/C _1121_/Q _0721_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0652_ _0542_/A _0740_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0583_ _0645_/A _0569_/X _0582_/X _0583_/D _0583_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_33_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_117 VGND VPWR sky130_fd_sc_hd__decap_6
X_1204_ addr_w[6] baseaddr_w_sync[6] _1188_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0528__A _0527_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1135_ d_sram_out[20] _0542_/D _1132_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1066_ _1064_/X _1066_/B _1056_/C _1066_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_40_209 VGND VPWR sky130_fd_sc_hd__decap_4
X_0919_ _1181_/Q _0907_/X _0918_/Y d_sram_in[15] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_108_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_180 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_201 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_86 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0901__A _0854_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0620__B _1147_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_83 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1154__D _1162_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_180 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_150 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0863__A2 _0833_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_0704_ _0704_/A _0704_/B _0699_/X _0704_/D _0705_/D VGND VPWR sky130_fd_sc_hd__or4_4
X_0635_ _0526_/X _0633_/X _0635_/C _0636_/C VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_97_220 VGND VPWR sky130_fd_sc_hd__fill_2
X_0566_ _0565_/X _0580_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_264 VGND VPWR sky130_fd_sc_hd__decap_6
X_0497_ _0497_/A _0659_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0551__A1 _0509_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1064__D _0955_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1118_ d_sram_out[3] _1118_/Q _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1049_ _1044_/X _1006_/X _1048_/Y _1049_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_21_220 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0705__B _0686_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0721__A _0740_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0790__B2 _0787_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_99 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_168 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_97 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_194 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_131 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_175 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_202 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1149__D _1149_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0631__A _0535_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0781__B2 _0496_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_267 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0806__A _0662_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_186 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0525__B _0524_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1013__A2 _1006_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0541__A _0535_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0772__B2 _1130_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0772__A1 _0521_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0618_ _0591_/A _0618_/B _0618_/C _0705_/A _0619_/C VGND VPWR sky130_fd_sc_hd__nor4_4
XANTENNA__1075__C _1056_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0549_ _0549_/A _0549_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_85_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_150 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_183 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_153 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0716__A _0668_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_289 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0818__A2 _1111_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_62 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0626__A _0540_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_95 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_280 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1161__CLK _1226_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0754__A1 _0542_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_147 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0754__B2 _0753_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_245 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0809__A2 _1104_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_248 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0536__A _0725_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_167 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0790__A2_N _0787_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0993__A1 _0968_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0702__C _0702_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_191 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_120 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_21 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_76 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_156 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_87 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1184__CLK _1223_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_217 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0612__C _0612_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0736__A1 _0668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_215 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1162__D _1225_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0672__B1 _0501_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_93 VGND VPWR sky130_fd_sc_hd__decap_12
X_0952_ _0955_/A _0991_/B _0952_/C _0960_/A VGND VPWR sky130_fd_sc_hd__and3_4
X_0883_ _0883_/A _0903_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0975__A1 _0946_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_15 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_112 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_101 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_123 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_23 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_2_0_clk clkbuf_4_3_0_clk/A _1197_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_87_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_204 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_237 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_229 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1157__D _1228_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_1220_ addr_r[8] baseaddr_r_sync[8] _1226_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_1151_ _1159_/Q _0510_/A _1223_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_207 VGND VPWR sky130_fd_sc_hd__fill_2
X_1082_ csb web _1163_/D VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_45_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_218 VGND VPWR sky130_fd_sc_hd__fill_2
X_0935_ _1193_/Q _0932_/X _0901_/Y d_sram_in[27] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0866_ _0866_/A _0866_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_9_182 VGND VPWR sky130_fd_sc_hd__fill_1
X_0797_ _0616_/C _0659_/A _0797_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_114_264 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_19 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_148 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_170 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_104 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0724__A _0510_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_148 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0939__A1 _1197_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1061__B1 _1056_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_99 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_88 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1222__CLK _1198_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_137 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0618__B _0618_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_74 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_251 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0634__A _0542_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1052__B1 _1048_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_68 VGND VPWR sky130_fd_sc_hd__decap_12
X_0720_ _0720_/A _0737_/B _0720_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_0651_ _0500_/X _0651_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0582_ _0584_/C _0582_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_245 VGND VPWR sky130_fd_sc_hd__fill_2
X_1203_ addr_w[5] baseaddr_w_sync[5] _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_26_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_129 VGND VPWR sky130_fd_sc_hd__fill_2
X_1134_ d_sram_out[19] _1134_/Q _1132_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1065_ _1007_/X _1055_/B _0952_/C _1066_/B VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__0544__A _0510_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0918_ _0854_/A _0917_/X _0918_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_0849_ _0830_/Y _0839_/X _0848_/Y _0849_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_102_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0719__A _0651_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_184 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_224 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_251 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_268 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0901__B _0901_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0620__C _0499_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_107 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0605__A1_N _0603_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0629__A _0629_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1118__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1170__D d_fabric_in[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_83 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_240 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0938__B1_N _0914_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_210 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_93 VGND VPWR sky130_fd_sc_hd__decap_8
X_0703_ _0703_/A _0703_/B _0701_/X _0702_/X _0704_/D VGND VPWR sky130_fd_sc_hd__or4_4
X_0634_ _0542_/D _0690_/C _0635_/C VGND VPWR sky130_fd_sc_hd__and2_4
X_0565_ _0565_/A _0565_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0496_ _0496_/A _0496_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0551__A2 _0546_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0539__A _0576_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1117_ d_sram_out[2] _1117_/Q _1162_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_132 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_1048_ _1045_/X _1056_/A _1056_/C _1048_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_21_232 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0705__C _0705_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_19 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1016__B1 _1012_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0721__B _0740_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_10 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_76 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_143 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_64 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0912__A _0903_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0631__B _0690_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1165__D _1165_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_287 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_224 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1090__CLK _1132_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0559__A1_N _0554_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_121 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0822__A d_sram_in[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_167 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0772__A2 _0669_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0617_ _0597_/B _0616_/X _0705_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_105_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_0548_ _0547_/X _0549_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_235 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0716__B _0720_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0732__A out_reg VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_205 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0907__A _0875_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_165 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0626__B _0702_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0642__A _0517_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_292 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0754__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_205 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_260 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0552__A _1154_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0993__A2 _0992_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_281 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0702__D _1118_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0727__A _0507_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_238 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_22 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_44 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_44 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_135 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_88 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0612__D _0611_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0736__A2 _0737_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_257 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0637__A _1141_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_238 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_102 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0672__A1 _0668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_157 VGND VPWR sky130_fd_sc_hd__decap_3
X_0951_ _0963_/A _0991_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0882_ _0903_/A _0899_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0975__A2 _0966_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_107 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_249 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0547__A _0499_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_219 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_157 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_207 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_35 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_190 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1151__CLK _1223_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_97 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0920__A _1182_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_232 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0590__B1 _0578_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_7 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1173__D d_fabric_in[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_149 VGND VPWR sky130_fd_sc_hd__fill_2
X_1150_ _1158_/Q _1150_/Q _1150_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_1081_ _1040_/X _1043_/A _1079_/X w_mask[31] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_45_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_161 VGND VPWR sky130_fd_sc_hd__decap_6
X_0934_ _1192_/Q _0932_/X _0897_/Y d_sram_in[26] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0865_ _0827_/A _0859_/X _0844_/X _0866_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0830__A _0846_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0796_ _0713_/X _0795_/X _0785_/X _1097_/Q d_fabric_out[14] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_114_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1083__D _0660_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1174__CLK _1221_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_19 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_271 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_127 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0724__B _0513_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1061__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0939__A2 _0922_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_56 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0740__A _0740_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_105 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_216 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0618__C _0618_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_263 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0634__B _0690_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_296 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1052__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1168__D d_fabric_in[2] VGND VPWR sky130_fd_sc_hd__diode_2
X_0650_ _0621_/Y _0623_/X _0549_/Y _0649_/X _0650_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_0581_ _0581_/A _1150_/Q _0584_/C VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1197__CLK _1197_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_127 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_93 VGND VPWR sky130_fd_sc_hd__decap_8
X_1202_ addr_w[4] baseaddr_w_sync[4] _1214_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_19_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_171 VGND VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_1_0_clk clkbuf_4_0_0_clk/A _1109_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1133_ d_sram_out[18] _0725_/D _1223_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1064_ _1007_/X _1045_/B _0973_/C _0955_/D _1064_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_92_163 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0825__A _1228_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0544__B _0544_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0917_ _1173_/Q _1046_/C _0916_/X _0917_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0560__A _1127_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0848_ _0897_/A _0848_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0779_ _0776_/A _0779_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_68_19 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_235 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_208 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_152 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_225 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_263 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_258 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_11 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_269 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0793__B1 _0792_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_174 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0645__A _0645_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0784__B1 _0783_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0702_ _0724_/C _0702_/B _0702_/C _1118_/Q _0702_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0633_ _0725_/D _0702_/C _0633_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0564_ _0564_/A _0565_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0495_ _0497_/A _0496_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1116_ d_sram_out[1] _0585_/D _1223_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_196 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1212__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0555__A _1153_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_144 VGND VPWR sky130_fd_sc_hd__fill_1
X_1047_ _1045_/B _0838_/B _0958_/X _1056_/C VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_110_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_188 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0705__D _0705_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1016__A1 _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0775__B1 _0773_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0721__C _0738_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_22 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_32 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_155 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0912__B _0903_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0631__C _0702_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0766__B1 _0719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_222 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1181__D d_fabric_in[15] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_196 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_281 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0772__A3 _0616_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_127 VGND VPWR sky130_fd_sc_hd__decap_12
X_0616_ _0510_/A _0513_/A _0616_/C _0533_/X _0616_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_124_190 VGND VPWR sky130_fd_sc_hd__decap_12
X_0547_ _0499_/A _0488_/Y _0499_/C _0547_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_105_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_214 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1091__D _0778_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_258 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0996__B1 _0988_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1108__CLK _1126_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_56 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_179 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0937__B1_N _0910_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_31 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_239 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0626__C _0626_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0642__B _0565_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_96 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_7 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1176__D d_fabric_in[10] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_269 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_155 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0833__A _0875_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_293 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1086__D _0747_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0727__B _0724_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_12 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_56 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_67 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0743__A _0616_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_208 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_214 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_171 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_225 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0918__A _0854_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_74 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0657__C1 _0656_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_291 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_250 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_147 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0672__A2 _0583_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0653__A _0740_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0950_ _0970_/A _0963_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0829__B1_N _0922_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0881_ _0835_/A _0903_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_126_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0828__A _0827_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_209 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0547__B _0488_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_250 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0563__A _0517_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_219 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_191 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_47 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0738__A _0542_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_174 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_44 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0920__B _0875_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0590__B2 _0589_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0590__A1 _0540_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_117 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_239 VGND VPWR sky130_fd_sc_hd__decap_4
X_1080_ _1035_/X _1070_/X _1079_/X w_mask[30] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0933_ _1191_/Q _0932_/X _0893_/Y d_sram_in[25] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_13_180 VGND VPWR sky130_fd_sc_hd__decap_3
X_0864_ _1171_/Q _0864_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_9_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_211 VGND VPWR sky130_fd_sc_hd__decap_3
X_0795_ _0575_/Y _0787_/X _1145_/Q _0711_/X _0795_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0558__A _0533_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0724__C _0724_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1061__A2 _1022_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0740__B _0740_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_54 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_183 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_209 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0618__D _0705_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_97 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1052__A2 _1015_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0580_ _0533_/X _0580_/B _0580_/C _1122_/Q _0580_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1184__D d_fabric_in[18] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_117 VGND VPWR sky130_fd_sc_hd__fill_2
X_1201_ addr_w[3] baseaddr_w_sync[3] _1128_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_111_269 VGND VPWR sky130_fd_sc_hd__fill_1
X_1132_ d_sram_out[17] _1132_/Q _1132_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1063_ _1001_/X _1059_/X _1061_/X w_mask[23] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_33_220 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0544__C _0544_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0841__A _1226_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0916_ _0903_/A _0903_/B _0908_/C _1181_/Q _0916_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0847_ _0880_/A _0946_/A _0844_/X _0846_/X _0897_/A VGND VPWR sky130_fd_sc_hd__a211o_4
X_0778_ _0509_/A _0496_/X _0544_/D _0496_/X _0778_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1141__CLK _1223_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1094__D _0788_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_269 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_131 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_215 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_23 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0793__A1 _0679_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_113 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_172 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0926__A _0875_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_142 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0645__B _0565_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_80 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1179__D d_fabric_in[13] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0661__A out_reg VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1164__CLK _1197_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0701_ _0724_/C _0701_/B _0701_/C _1132_/Q _0701_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_128_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0784__A1 _0722_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0632_ _0544_/D _0627_/Y _0703_/A _0631_/X _0632_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_97_201 VGND VPWR sky130_fd_sc_hd__decap_3
X_0563_ _0517_/X _0645_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_31_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_245 VGND VPWR sky130_fd_sc_hd__fill_2
X_0494_ _0493_/X _0497_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_57_109 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_153 VGND VPWR sky130_fd_sc_hd__fill_2
X_1115_ d_sram_out[0] _1115_/Q _1197_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0836__A _0835_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_167 VGND VPWR sky130_fd_sc_hd__fill_2
X_1046_ _1007_/X _1045_/B _1046_/C _1056_/A VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_21_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1089__D _1089_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_111 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1016__A2 _1015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0571__A _0570_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0775__A1 _0740_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0775__B2 _0774_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0721__D _1121_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_22 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1187__CLK _1198_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_32 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0912__C _0908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0766__A1 _0609_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_147 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_0_0_clk clkbuf_4_0_0_clk/A _1214_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_5_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0631__D _1127_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_109 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0656__A _0544_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_167 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_139 VGND VPWR sky130_fd_sc_hd__decap_12
X_0615_ _0614_/Y _0576_/X _1112_/D _0558_/X _0618_/C VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_0546_ _0509_/B _0546_/B _0546_/C _0546_/D _0546_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_105_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_186 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0566__A _0565_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_270 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0693__B1 _0692_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_178 VGND VPWR sky130_fd_sc_hd__fill_2
X_1029_ _0960_/C _1029_/B _1028_/X _1029_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0996__A1 _0985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_66 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_112 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_76 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0788__A1_N _0554_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0642__C _0587_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_86 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_261 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1202__CLK _1214_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1192__D d_fabric_in[26] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0911__A1 _1179_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_115 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1010__A _0949_/A VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_7_0_clk clkbuf_3_7_0_clk/A clkbuf_3_7_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_104_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_194 VGND VPWR sky130_fd_sc_hd__decap_12
X_0529_ _0529_/A _0643_/C VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0902__A1 _1177_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_145 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0666__B1 _0665_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_13 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0727__C _0727_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_167 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_46 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_262 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_57 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0743__B _0509_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_23 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1225__CLK _1198_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_150 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_237 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0918__B _0917_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_112 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0657__B1 _0655_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_7 VGND VPWR sky130_fd_sc_hd__decap_12
X_0880_ _0880_/A _1046_/C _0888_/A VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1187__D d_fabric_in[21] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_159 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0828__B _0826_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0896__B1 _0895_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_18 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1005__A _0982_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0648__B1 _0622_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0547__C _0499_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_137 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0844__A d_sram_in[0] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0936__B1_N _0905_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1073__B1 _1071_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0820__B1 _1145_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1097__D _0795_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_181 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0738__B _0738_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_44 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_181 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0811__B1 _0740_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0590__A2 _0701_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0664__A out_reg VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_276 VGND VPWR sky130_fd_sc_hd__decap_12
X_0932_ _0875_/Y _0932_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0863_ _0857_/Y _0833_/X _0862_/X d_sram_in[4] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_9_174 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0802__B1 _0655_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_0794_ _0713_/X _0793_/X _0785_/X _1096_/Q d_fabric_out[13] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_87_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0839__A _0838_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0558__B _1153_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_207 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_251 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0574__A _0518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_221 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0724__D _0724_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0740__C _0722_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1037__B1 _1036_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_140 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_80 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0659__A _0659_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1200_ addr_w[2] baseaddr_w_sync[2] _1126_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1093__CLK _1109_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1131_ d_sram_out[16] _0655_/A _1109_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_77_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_121 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_132 VGND VPWR sky130_fd_sc_hd__fill_2
X_1062_ _0995_/X _1059_/X _1061_/X w_mask[22] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_18_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_243 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0544__D _0544_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0915_ _0912_/D _0907_/X _0914_/Y d_sram_in[14] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0841__B _0841_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0846_ _0846_/A _0852_/B _0846_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0777_ _0762_/X _0775_/X _0776_/X d_fabric_out[7] VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0569__A _1153_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_210 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_216 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1019__B1 _1011_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_35 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0793__A2 _0711_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_151 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_198 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0645__C _0643_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0942__A _0942_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0700_ _0535_/A _0700_/B _0717_/B _1130_/Q _0703_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_128_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0784__A2 _0711_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1195__D d_fabric_in[29] VGND VPWR sky130_fd_sc_hd__diode_2
X_0631_ _0535_/A _0690_/C _0702_/B _1127_/Q _0631_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0562_ _0561_/X _0562_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0493_ _0492_/X _0493_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_24_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_132 VGND VPWR sky130_fd_sc_hd__fill_2
X_1114_ _0616_/C _1114_/Q _1126_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_0_94 VGND VPWR sky130_fd_sc_hd__decap_6
X_1045_ _0955_/A _1045_/B _0973_/C _1045_/D _1045_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0852__A _0851_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0775__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_137 VGND VPWR sky130_fd_sc_hd__decap_12
X_0829_ _0880_/A _0826_/X _0922_/A d_sram_in[1] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_135_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_79 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_68 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_198 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_113 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0762__A _0662_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_239 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0912__D _0912_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0766__A2 _0765_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_192 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0923__C1 _0922_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_235 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_279 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_205 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_132 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0656__B _0717_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1131__CLK _1109_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0614_ _1145_/Q _0614_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_131_118 VGND VPWR sky130_fd_sc_hd__fill_2
X_0545_ _0540_/X _0542_/X _0544_/X _0546_/D VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__1008__A _0963_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_113 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_282 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_198 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0693__A1 _0676_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_157 VGND VPWR sky130_fd_sc_hd__fill_2
X_1028_ _1028_/A _1028_/B _1028_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_14_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0582__A _0584_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0996__A2 _0979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_170 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0757__A _0679_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_143 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1154__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_271 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0492__A _0499_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0642__D _0642_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_273 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0667__A _0493_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_238 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_249 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0911__A2 _0907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_293 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1010__B _0956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_129 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1177__CLK _1226_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0528_ _0527_/X _0529_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_58_205 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_249 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0902__A2 _0877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_271 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_124 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0666__A1 _0663_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0727__D _0726_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_47 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_105 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_58 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_285 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0743__C _0743_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_35 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_184 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0487__A _1132_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0657__A1 _0668_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_285 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0950__A _0970_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_90 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0896__A1 _0846_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_219 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1005__B _0982_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0648__A1 _0509_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0844__B _0826_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1021__A _0973_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1073__A1 _1022_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0820__A1 _0662_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0820__B2 _0815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_160 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0738__C _0738_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_208 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_219 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_230 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_160 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_193 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0811__A1 _0806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0811__B2 _0808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_257 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0590__A3 _0509_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_86 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_6_0_clk clkbuf_3_7_0_clk/A clkbuf_3_6_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0945__A _0945_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_288 VGND VPWR sky130_fd_sc_hd__decap_8
X_0931_ _1190_/Q _0926_/X _0888_/Y d_sram_in[24] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__1198__D addr_w[0] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0802__A1 _0799_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0680__A _0544_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0862_ _0857_/Y _0839_/X _0861_/Y _0862_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0802__B2 _0801_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0793_ _0679_/D _0711_/X _0792_/X _0793_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_54_3 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0558__C _0576_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1215__CLK _1188_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0574__B _0569_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_263 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_296 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0740__D _0740_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_208 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_67 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_62 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1037__A1 _0985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_152 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0796__B1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_145 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0659__B _0658_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_249 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0935__B1_N _0901_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_7 VGND VPWR sky130_fd_sc_hd__fill_2
X_1130_ d_sram_out[15] _1130_/Q _1223_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1061_ _1044_/X _1022_/X _1056_/Y _1061_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0675__A _0740_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_233 VGND VPWR sky130_fd_sc_hd__fill_2
X_0914_ _0897_/A _0913_/X _0914_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__0841__C _0841_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0845_ _0835_/A _0834_/A _0841_/C _0852_/B VGND VPWR sky130_fd_sc_hd__and3_4
X_0776_ _0776_/A _1090_/Q _0776_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_102_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_271 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0585__A _0517_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_59 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_206 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1019__A1 _0985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_47 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_135 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0778__B1 _0544_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_157 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0495__A _0497_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_166 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0645__D _1121_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_62 VGND VPWR sky130_fd_sc_hd__decap_12
X_0630_ _0594_/B _0690_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_136_190 VGND VPWR sky130_fd_sc_hd__decap_8
X_0561_ _0517_/A _0564_/A _0510_/A _1150_/Q _0561_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_97_236 VGND VPWR sky130_fd_sc_hd__fill_2
X_0492_ _0499_/A _0488_/Y _0492_/C _0498_/A _0492_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_17_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0889__B1_N _0888_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1113_ _1145_/Q _1113_/Q _1126_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_188 VGND VPWR sky130_fd_sc_hd__fill_2
X_1044_ _1044_/A _1044_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_80_147 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0852__B _0852_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_269 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_0828_ _0827_/Y _0826_/X _0922_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_134_149 VGND VPWR sky130_fd_sc_hd__decap_4
X_0759_ _0757_/X _0758_/X _0719_/X _0759_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_135_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_107 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_203 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_258 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_111 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_122 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1083__CLK _1109_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_171 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0923__B1 _0844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_100 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_80 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_125 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_147 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0953__A _0977_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_0613_ _0697_/A _0701_/B _0594_/B _1141_/Q _0618_/B VGND VPWR sky130_fd_sc_hd__and4_4
X_0544_ _0510_/X _0544_/B _0544_/C _0544_/D _0544_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_85_239 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1024__A _0982_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0693__A2 _0627_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_294 VGND VPWR sky130_fd_sc_hd__decap_4
X_1027_ _1031_/A _0956_/X _0953_/Y _0955_/D _1028_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_14_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_206 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0757__B _0717_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_89 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0492__B _0488_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_81 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0948__A _0969_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_250 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_209 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0683__A _0509_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1010__C _0952_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0596__D1 _0595_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_0527_ _0581_/A _0556_/B _0527_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0858__A _0852_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_228 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0666__A2 _0660_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0593__A _0587_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_15 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_37 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_139 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0743__D _0742_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_47 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_233 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1121__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_209 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0657__A2 _0502_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_147 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_76 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_70 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0678__A _1112_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0896__A2 _0890_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_261 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1005__C _1017_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0648__A2 _0703_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_231 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1073__A2 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1021__B _1021_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0820__A2 _1113_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1144__CLK _1188_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0588__A _0584_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0738__D _1122_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_117 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0811__A2 _1106_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_211 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_244 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_269 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0498__A _0498_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_201 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_234 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1167__CLK _1188_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_150 VGND VPWR sky130_fd_sc_hd__fill_1
X_0930_ _1189_/Q _0926_/X _0873_/X d_sram_in[23] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_13_194 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_110 VGND VPWR sky130_fd_sc_hd__fill_2
X_0861_ _0861_/A _0861_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0802__A2 _1099_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0792_ _1128_/Q _0493_/X _0792_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_47_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0558__D _0513_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_153 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_197 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0574__C _0573_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1032__A _1031_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_24 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_41 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_74 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1037__A2 _1001_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0796__A1 _0713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0796__B2 _1097_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_168 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_164 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0956__A _0970_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_101 VGND VPWR sky130_fd_sc_hd__fill_2
X_1060_ _0992_/X _1059_/X _1057_/X w_mask[21] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0675__B _0669_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_178 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0691__A _1142_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0913_ _1172_/Q _1046_/C _0912_/X _0913_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_0844_ d_sram_in[0] _0826_/X _0844_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_108_19 VGND VPWR sky130_fd_sc_hd__decap_12
X_0775_ _0740_/D _0750_/X _0773_/X _0774_/X _0775_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_102_206 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_239 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1027__A _1031_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_142 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0866__A _0866_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0585__B _0565_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1189_ d_fabric_in[23] _1189_/Q _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_207 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_229 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1019__A2 _0992_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0778__B2 _0496_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_169 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_5_0_clk clkbuf_3_5_0_clk/A clkbuf_3_5_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_58_56 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0776__A _0776_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_245 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1205__CLK _1197_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0560_ _1127_/Q _0560_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_97_215 VGND VPWR sky130_fd_sc_hd__decap_3
X_0491_ _0544_/B _0492_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0686__A _0675_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_101 VGND VPWR sky130_fd_sc_hd__fill_2
X_1112_ _1112_/D _1112_/Q _1214_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1043_ _1043_/A _1043_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_65_178 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_147 VGND VPWR sky130_fd_sc_hd__decap_12
X_0827_ _0827_/A _0827_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0758_ _0668_/X _1128_/Q _0687_/X _0758_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_135_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_0689_ _0738_/C _0597_/B _0689_/C _0705_/C VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_56_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_69 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0934__B1_N _0897_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1228__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0923__A1 _1183_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_178 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_137 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_0612_ _0599_/X _0612_/B _0612_/C _0611_/Y _0619_/B VGND VPWR sky130_fd_sc_hd__nor4_4
X_0543_ _1107_/D _0544_/D VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_167 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1024__B _0982_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1026_ _0985_/A _0995_/X _1029_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_61_170 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0850__B1 _0849_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1040__A _1039_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_178 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_35 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_137 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0492__C _0492_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_242 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1100__D _1132_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_183 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_240 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0964__A _1031_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_159 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0683__B _0679_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_192 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_220 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0596__C1 _0526_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0526_ _0525_/X _0526_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1035__A _1034_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_38 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1076__B1 _1075_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1009_ _1007_/X _1045_/B _0991_/C _1045_/D _1009_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_135_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_218 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_243 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1067__B1 _1066_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0814__B1 _0676_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_234 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1096__CLK _1089_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_280 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1005__D _1017_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_273 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0694__A _0535_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_221 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_254 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1058__B1 _1057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1021__C _1017_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0805__B1 _0742_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0869__A _1172_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0588__B _0588_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_134 VGND VPWR sky130_fd_sc_hd__fill_2
X_0509_ _0509_/A _0509_/B _0509_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_100_167 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_7_0_clk_A clkbuf_3_7_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1049__B1 _1048_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_256 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_289 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0779__A _0776_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_22 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_98 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_184 VGND VPWR sky130_fd_sc_hd__decap_8
X_0860_ _0826_/X _0859_/X _0880_/A _0861_/A VGND VPWR sky130_fd_sc_hd__o21a_4
X_0791_ _0713_/X _1095_/D _0785_/X _1095_/Q d_fabric_out[12] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_114_215 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0689__A _0738_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_110 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_213 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1111__CLK _1214_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_0989_ _0985_/X _0974_/X _0988_/Y _0989_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_105_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_204 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0599__A _0518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_110 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_36 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_154 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_53 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_57 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0796__A2 _0795_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_187 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_143 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0675__C _0675_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1134__CLK _1132_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0972__A _0972_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_0912_ _0903_/A _0903_/B _0908_/C _0912_/D _0912_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0843_ _1044_/A _0946_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_0774_ _1122_/Q _0659_/A _0709_/X _0774_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1027__B _0956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_176 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1043__A _1043_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0585__C _0584_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_135 VGND VPWR sky130_fd_sc_hd__fill_2
X_1188_ d_fabric_in[22] _1188_/Q _1188_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_17_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0882__A _0903_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_219 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_106 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1157__CLK _1162_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0776__B _1090_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_176 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1103__D _0542_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0792__A _1128_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_44 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_55 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_86 VGND VPWR sky130_fd_sc_hd__decap_12
X_0490_ _0556_/B _0544_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_249 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0686__B _0655_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1111_ _0532_/A _1111_/Q _1214_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_80_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_1042_ _0899_/A _0899_/B _1042_/C _1042_/D _1043_/A VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_0_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_159 VGND VPWR sky130_fd_sc_hd__decap_12
X_0826_ _0835_/A _0834_/A _1042_/C _0826_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0757_ _0679_/D _0717_/B _0757_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA_clkbuf_4_6_0_clk_A clkbuf_4_7_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0688_ _0607_/X _0687_/X _0689_/C VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0877__A _0922_/B VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_15_0_clk clkbuf_3_7_0_clk/X _1198_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_71_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_36 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_23 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_184 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0923__A2 _0922_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0787__A _0496_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_93 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_116 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_160 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_81 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_0611_ _0724_/C _0597_/B _0611_/C _0611_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_0542_ _0542_/A _0513_/X _0544_/C _0542_/D _0542_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0697__A _0697_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_146 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1024__C _1000_/C VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_4_0_clk clkbuf_3_5_0_clk/A clkbuf_4_9_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1025_ _1024_/X _1025_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_46_190 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0850__A1 _0830_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_193 VGND VPWR sky130_fd_sc_hd__fill_2
X_0809_ _0806_/X _1104_/Q _0675_/D _0808_/X d_fabric_out[21] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_115_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_263 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_116 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0492__D _0498_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_298 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_274 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_211 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0964__B _1021_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0683__C _0681_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_233 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_288 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_1_1_0_clk_A clkbuf_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_232 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0596__B1 _0718_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0525_ _0655_/A _0524_/X _0525_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0933__B1_N _0893_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0615__A1_N _0614_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1218__CLK _1109_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_149 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_28 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_277 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1076__A1 _0985_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1008_ _0963_/A _1045_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_34_193 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0890__A _1046_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1201__D addr_w[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_204 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_3_0_clk_A clkbuf_3_3_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_263 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_68 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_116 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_222 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1067__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1111__D _0532_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0814__B2 _0808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0814__A1 _0813_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_14_0_clk_A clkbuf_3_7_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_174 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_185 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_246 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_292 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_296 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0694__B _0700_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1058__A1 _0983_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_266 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1021__D _1017_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_152 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0805__A1 _0799_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0805__B2 _0801_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0588__C _0586_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0508_ _0507_/Y _0509_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1046__A _1007_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1190__CLK _1197_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0885__A _0841_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_244 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1049__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_163 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_268 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0980__B1 _0975_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_34 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_293 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1106__D _0740_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_93 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_258 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_167 VGND VPWR sky130_fd_sc_hd__fill_1
X_0790_ _0560_/Y _0787_/X _0532_/A _0787_/X _1095_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_7 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0689__B _0597_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_271 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_225 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_0988_ _0960_/A _0988_/B _0960_/C _0988_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_105_238 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0599__B _0701_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_199 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_98 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1086__CLK _1162_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_133 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_166 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0650__C1 _0649_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_208 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_0_0_clk_A clkbuf_1_0_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0675__D _0675_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_92 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_0911_ _1179_/Q _0907_/X _0910_/Y d_sram_in[13] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0842_ _0841_/X _1044_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0773_ _0771_/X _0772_/X _0719_/X _0773_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_52_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1027__C _0953_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_263 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_296 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0585__D _0585_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1187_ d_fabric_in[21] _1187_/Q _1198_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_83_169 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_2_0_clk_A clkbuf_4_3_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_209 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0632__C1 _0631_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_241 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_291 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0792__B _0493_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_180 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_269 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_67 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_105 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_98 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1101__CLK _1132_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1110_ _1142_/Q _1110_/Q _1214_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0686__C _0702_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0983__A _0982_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32 VGND VPWR sky130_fd_sc_hd__decap_12
X_1041_ _0945_/A _1040_/X _1037_/X w_mask[15] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_0_87 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_74 VGND VPWR sky130_fd_sc_hd__decap_12
X_0825_ _1228_/Q _1042_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_127_171 VGND VPWR sky130_fd_sc_hd__decap_12
X_0756_ _0663_/X _0754_/X _0755_/X d_fabric_out[4] VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0917__B1 _0916_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0687_ _0675_/D _0690_/C _0687_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_88_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_125 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_147 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1204__D addr_w[6] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0893__A _0866_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_38 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_180 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_191 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0853__C1 _0852_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_22 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_66 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_261 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1124__CLK _1197_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_35 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_239 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1114__D _0616_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_191 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_171 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_160 VGND VPWR sky130_fd_sc_hd__fill_1
X_0610_ _0675_/D _0582_/X _0607_/X _0608_/X _0609_/X _0611_/C VGND VPWR sky130_fd_sc_hd__a2111oi_4
XFILLER_124_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0978__A _0973_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0541_ _0535_/A _0544_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0697__B _0700_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1024__D _1017_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1024_ _0982_/A _0982_/B _1000_/C _1017_/D _1024_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0850__A2 _0833_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1147__CLK _1150_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0808_ _0776_/A _0808_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0888__A _0888_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0739_ _0722_/A _0492_/C _0722_/C _0739_/D _0744_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_39_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_15 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_180 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_211 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1109__D _1141_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_10_0_clk_A clkbuf_3_5_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_71 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_231 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0964__C _0977_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_109 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0683__D _0682_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_7 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_14_0_clk clkbuf_3_7_0_clk/X _1171_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0596__A1 _1134_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0524_ _0581_/A _0544_/B _0524_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0501__A _0500_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_209 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_128 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_29 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_109 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1076__A2 _1035_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1007_ _1031_/A _1007_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_135_214 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_216 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_177 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_139 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1067__A2 _1025_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_289 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_172 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_68 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_79 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_62 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0814__A2 _1108_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_197 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_258 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_3_0_clk clkbuf_3_3_0_clk/A clkbuf_4_7_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0694__C _0582_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_245 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1058__A2 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0991__A _0982_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_142 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0805__A2 _1102_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_225 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_291 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_164 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0588__D _0588_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0507_ _0737_/B _0507_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1046__B _1045_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_256 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1049__A2 _1006_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1212__D addr_r[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0980__A1 _0968_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_46 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_215 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1122__D d_sram_out[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_131 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1208__CLK _1150_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0689__C _0689_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0986__A _0955_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_98 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_201 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_237 VGND VPWR sky130_fd_sc_hd__decap_6
X_0987_ _0955_/A _1055_/B _0991_/C _1045_/D _0988_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_8_190 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0599__C _0701_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1207__D addr_w[9] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_245 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_105 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0650__B1 _0549_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_250 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1117__D d_sram_out[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_201 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_237 VGND VPWR sky130_fd_sc_hd__decap_6
X_0910_ _0866_/A _0910_/B _0910_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_41_281 VGND VPWR sky130_fd_sc_hd__decap_12
X_0841_ _1226_/Q _0841_/B _0841_/C _0841_/X VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__1180__CLK _1089_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0772_ _0521_/A _0669_/X _0616_/C _0668_/A _1130_/Q _0772_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_5_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1027__D _0955_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_148 VGND VPWR sky130_fd_sc_hd__fill_2
X_1186_ d_fabric_in[20] _1186_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_24_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0632__B1 _0703_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0935__A1 _1193_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_123 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_253 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_126 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0871__B1 _0870_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_79 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_117 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0623__B1 _0622_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_152 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0686__D _1128_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44 VGND VPWR sky130_fd_sc_hd__decap_12
X_1040_ _1039_/X _1040_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0862__B1 _0861_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0504__A _0504_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0824_ _0841_/B _0834_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0755_ _0733_/A _1087_/Q _0755_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0917__A1 _1173_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0686_ _0675_/C _0655_/B _0702_/B _1128_/Q _0686_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_88_207 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0893__B _0893_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1169_ d_fabric_in[3] _0851_/A _1162_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1070__A _1043_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0853__B1 _0844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1220__D addr_r[8] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_78 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_56 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0605__B1 _1142_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_183 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_47 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1030__B1 _1029_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_104 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_84 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_151 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1130__D d_sram_out[15] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_60 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_71 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0978__B _0991_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0540_ _0542_/A _0738_/B _0540_/C _0642_/D _0540_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1099__CLK _1132_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0697__C _0580_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0994__A _0949_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1023_ _0998_/X _1022_/X _1019_/X w_mask[11] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_53_107 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_298 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_173 VGND VPWR sky130_fd_sc_hd__fill_2
X_0807_ _0806_/X _1103_/Q _0542_/D _0801_/X d_fabric_out[20] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1012__B1 _1011_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0738_ _0542_/A _0738_/B _0738_/C _1122_/Q _0738_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0888__B _0887_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_0669_ _0740_/B _0669_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1065__A _1007_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_145 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_240 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1215__D addr_r[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_27 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1079__B1 _1075_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_140 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0826__B1 _1042_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_85 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_74 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1125__D d_sram_out[10] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_83 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0964__D _0972_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0817__B1 _0739_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_184 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0596__A2 _0580_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0523_ _0570_/A _0581_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_167 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_276 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1114__CLK _1126_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1006_ _1005_/X _1006_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_34_162 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0899__A _0899_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_228 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_221 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_268 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0602__A _0697_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_210 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1137__CLK _1214_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0694__D _0737_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_235 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0991__B _0991_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_173 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_80 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_3 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_190 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_215 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_237 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0512__A _0722_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_121 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_154 VGND VPWR sky130_fd_sc_hd__decap_3
X_0506_ _0506_/A _0737_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1046__C _1046_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_268 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_110 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_154 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0980__A2 _0979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_58 VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_13_0_clk clkbuf_3_6_0_clk/X _1185_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_133_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_73 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_110 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_176 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_114 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_213 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0507__A _0737_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0986_ _0955_/D _1045_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0599__D _1107_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_257 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1223__D addr_r[11] VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_2_0_clk clkbuf_3_3_0_clk/A clkbuf_3_2_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_42_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_49 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0650__A1 _0621_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_113 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_168 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1133__D d_sram_out[18] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_293 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_82 VGND VPWR sky130_fd_sc_hd__fill_2
X_0840_ _1228_/Q _0841_/C VGND VPWR sky130_fd_sc_hd__inv_8
X_0771_ _0740_/D _0655_/B _0771_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_38_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_146 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_127 VGND VPWR sky130_fd_sc_hd__fill_2
X_1185_ d_fabric_in[19] _1185_/Q _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_24_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0632__A1 _0544_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0969_ _0969_/A _0973_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0935__A2 _0932_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_109 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1218__D addr_r[6] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0700__A _0535_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_113 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_105 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0931__B1_N _0888_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_216 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0871__A1 _0869_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_293 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0623__A1 _1115_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_23 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1128__D d_sram_out[13] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_120 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_60 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_119 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0862__A1 _0857_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_98 VGND VPWR sky130_fd_sc_hd__decap_8
X_0823_ _1226_/Q _0835_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_80_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_0754_ _0542_/D _0750_/X _0752_/X _0753_/X _0754_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__0917__A2 _1046_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0685_ _0674_/X _0684_/Y _0550_/X _0685_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0520__A _0540_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_274 VGND VPWR sky130_fd_sc_hd__fill_1
X_1168_ d_fabric_in[2] _0846_/A _1223_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0853__A1 _0827_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1099_ _0655_/A _1099_/Q _1132_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0605__B2 _0639_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_296 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1030__A1 _0945_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1170__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_62 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_184 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0978__C _1017_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0780__B1 _0762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0697__D _1122_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_285 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0994__B _0956_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1022_ _1022_/A _1022_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0515__A _0738_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0806_ _0662_/A _0806_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_115_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1012__A1 _0985_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0737_ _0737_/A _0737_/B _0737_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_115_176 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0888__C _0861_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0668_ _0668_/A _0668_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1065__B _1055_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1193__CLK _1221_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0599_ _0518_/X _0701_/B _0701_/C _1107_/D _0599_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_37_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_119 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1079__A1 _0985_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0826__A1 _0835_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_165 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_64 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_187 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_62 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_203 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0817__A1 _0813_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0817__B2 _0815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1141__D d_sram_out[26] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_44 VGND VPWR sky130_fd_sc_hd__decap_12
X_0522_ _0510_/A _0570_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0753__B1 _0709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_179 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_214 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_225 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_236 VGND VPWR sky130_fd_sc_hd__fill_2
X_1005_ _0982_/A _0982_/B _1017_/C _1017_/D _1005_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_34_185 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0899__B _0899_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1226__D conf[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_146 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_135 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_255 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_247 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1089__CLK _1089_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_122 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0602__B _0701_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0735__B1 _0742_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1136__D d_sram_out[21] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_273 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_240 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0991__C _0991_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_280 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_180 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_0505_ _0513_/A _0533_/A _0506_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_100_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_200 VGND VPWR sky130_fd_sc_hd__decap_12
.ends

