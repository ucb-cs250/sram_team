* NGSPICE file created from sram_ifc.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 D Q CLK VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D Y VGND VPWR
.ends

.subckt sram_ifc addr_r[0] addr_r[10] addr_r[11] addr_r[12] addr_r[13] addr_r[1] addr_r[2]
+ addr_r[3] addr_r[4] addr_r[5] addr_r[6] addr_r[7] addr_r[8] addr_r[9] addr_w[0]
+ addr_w[10] addr_w[11] addr_w[12] addr_w[13] addr_w[1] addr_w[2] addr_w[3] addr_w[4]
+ addr_w[5] addr_w[6] addr_w[7] addr_w[8] addr_w[9] baseaddr_r_sync[0] baseaddr_r_sync[1]
+ baseaddr_r_sync[2] baseaddr_r_sync[3] baseaddr_r_sync[4] baseaddr_r_sync[5] baseaddr_r_sync[6]
+ baseaddr_r_sync[7] baseaddr_r_sync[8] baseaddr_w_sync[0] baseaddr_w_sync[1] baseaddr_w_sync[2]
+ baseaddr_w_sync[3] baseaddr_w_sync[4] baseaddr_w_sync[5] baseaddr_w_sync[6] baseaddr_w_sync[7]
+ baseaddr_w_sync[8] clk conf[0] conf[1] conf[2] csb csb0_sync csb1_sync d_fabric_in[0]
+ d_fabric_in[10] d_fabric_in[11] d_fabric_in[12] d_fabric_in[13] d_fabric_in[14]
+ d_fabric_in[15] d_fabric_in[16] d_fabric_in[17] d_fabric_in[18] d_fabric_in[19]
+ d_fabric_in[1] d_fabric_in[20] d_fabric_in[21] d_fabric_in[22] d_fabric_in[23] d_fabric_in[24]
+ d_fabric_in[25] d_fabric_in[26] d_fabric_in[27] d_fabric_in[28] d_fabric_in[29]
+ d_fabric_in[2] d_fabric_in[30] d_fabric_in[31] d_fabric_in[3] d_fabric_in[4] d_fabric_in[5]
+ d_fabric_in[6] d_fabric_in[7] d_fabric_in[8] d_fabric_in[9] d_fabric_out[0] d_fabric_out[10]
+ d_fabric_out[11] d_fabric_out[12] d_fabric_out[13] d_fabric_out[14] d_fabric_out[15]
+ d_fabric_out[16] d_fabric_out[17] d_fabric_out[18] d_fabric_out[19] d_fabric_out[1]
+ d_fabric_out[20] d_fabric_out[21] d_fabric_out[22] d_fabric_out[23] d_fabric_out[24]
+ d_fabric_out[25] d_fabric_out[26] d_fabric_out[27] d_fabric_out[28] d_fabric_out[29]
+ d_fabric_out[2] d_fabric_out[30] d_fabric_out[31] d_fabric_out[3] d_fabric_out[4]
+ d_fabric_out[5] d_fabric_out[6] d_fabric_out[7] d_fabric_out[8] d_fabric_out[9]
+ d_sram_in[0] d_sram_in[10] d_sram_in[11] d_sram_in[12] d_sram_in[13] d_sram_in[14]
+ d_sram_in[15] d_sram_in[16] d_sram_in[17] d_sram_in[18] d_sram_in[19] d_sram_in[1]
+ d_sram_in[20] d_sram_in[21] d_sram_in[22] d_sram_in[23] d_sram_in[24] d_sram_in[25]
+ d_sram_in[26] d_sram_in[27] d_sram_in[28] d_sram_in[29] d_sram_in[2] d_sram_in[30]
+ d_sram_in[31] d_sram_in[3] d_sram_in[4] d_sram_in[5] d_sram_in[6] d_sram_in[7] d_sram_in[8]
+ d_sram_in[9] d_sram_out[0] d_sram_out[10] d_sram_out[11] d_sram_out[12] d_sram_out[13]
+ d_sram_out[14] d_sram_out[15] d_sram_out[16] d_sram_out[17] d_sram_out[18] d_sram_out[19]
+ d_sram_out[1] d_sram_out[20] d_sram_out[21] d_sram_out[22] d_sram_out[23] d_sram_out[24]
+ d_sram_out[25] d_sram_out[26] d_sram_out[27] d_sram_out[28] d_sram_out[29] d_sram_out[2]
+ d_sram_out[30] d_sram_out[31] d_sram_out[3] d_sram_out[4] d_sram_out[5] d_sram_out[6]
+ d_sram_out[7] d_sram_out[8] d_sram_out[9] out_reg reb w_mask[0] w_mask[10] w_mask[11]
+ w_mask[12] w_mask[13] w_mask[14] w_mask[15] w_mask[16] w_mask[17] w_mask[18] w_mask[19]
+ w_mask[1] w_mask[20] w_mask[21] w_mask[22] w_mask[23] w_mask[24] w_mask[25] w_mask[26]
+ w_mask[27] w_mask[28] w_mask[29] w_mask[2] w_mask[30] w_mask[31] w_mask[3] w_mask[4]
+ w_mask[5] w_mask[6] w_mask[7] w_mask[8] w_mask[9] web web0_sync VPWR VGND
XFILLER_39_233 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_247 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_188 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0703__A _0703_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_63 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_85 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_239 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_188 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0613__A _0697_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_354 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1104__CLK _1104_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0708__B1 _0707_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0765__A2_N _0528_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0985_ _0984_/X _0985_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0523__A _0523_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_291 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0650__A2 _0623_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1127__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_368 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_225 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_62 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0608__A _0634_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0770_ _0762_/X _1089_/D _0769_/X d_fabric_out[6] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_5_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_353 VGND VPWR sky130_fd_sc_hd__fill_2
X_1184_ d_fabric_in[18] _1184_/Q _1184_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0518__A _0587_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_239 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0632__A2 _0627_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0968_ _0943_/X _0968_/X VGND VPWR sky130_fd_sc_hd__buf_1
Xclkbuf_4_12_0_clk clkbuf_3_6_0_clk/X _1196_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0899_ _0899_/A _0899_/B _0903_/C _1177_/Q _0899_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0700__B _0694_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_114 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0871__A2 _0833_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_294 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0623__A2 _0620_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_198 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1144__D d_sram_out[29] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_50 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0847__C1 _0846_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0862__A2 _0839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_367 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_261 VGND VPWR sky130_fd_sc_hd__decap_3
X_0822_ d_sram_in[0] _0880_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0753_ _0540_/D _0495_/X _0709_/X _0753_/X VGND VPWR sky130_fd_sc_hd__o21a_4
Xclkbuf_3_1_0_clk clkbuf_3_1_0_clk/A clkbuf_4_2_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0801__A _0665_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0684_ _0684_/A _0676_/X _0684_/C _0684_/D _0684_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_29_309 VGND VPWR sky130_fd_sc_hd__fill_2
X_1167_ d_fabric_in[1] _0827_/A _1152_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_44_19 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_312 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0853__A2 _0859_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1098_ _1098_/D _1098_/Q _1155_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1030__A2 _1025_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0711__A _0497_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_320 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_375 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_356 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_367 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_85 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_235 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1139__D d_sram_out[24] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0978__D _0982_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0780__A1 _0779_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0780__B2 _1091_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_82 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0994__C _0999_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1021_ _0973_/A _1021_/B _1021_/C _1021_/D _1021_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_34_334 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0930__B1_N _0873_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0805_ _0799_/X _1102_/Q _0695_/X _0801_/X d_fabric_out[19] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__0531__A _0530_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1012__A2 _0983_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0736_ _0668_/X _1126_/Q _0501_/X _0735_/X _0736_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_0667_ _0493_/X _0750_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1065__C _0878_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_19 VGND VPWR sky130_fd_sc_hd__fill_1
X_0598_ _0579_/C _0701_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_29_128 VGND VPWR sky130_fd_sc_hd__fill_2
X_1219_ addr_r[7] baseaddr_r_sync[7] _1108_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1079__A2 _1040_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_109 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_301 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0826__A2 _0845_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_120 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_348 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_65 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_400 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_40 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0817__A2 _1110_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_73 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0616__A _1151_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_315 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_95 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_56 VGND VPWR sky130_fd_sc_hd__decap_12
X_0521_ _0676_/A _0721_/B _0721_/C _1127_/Q _0521_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0753__A1 _0540_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_256 VGND VPWR sky130_fd_sc_hd__decap_12
X_1004_ _1031_/D _1021_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0526__A _0526_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_348 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1160__CLK _1152_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0899__C _0903_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0719_ _0651_/Y _0719_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_57_234 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_178 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_75 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0602__C _0633_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0735__B2 _0655_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0735__A1 _0676_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1152__D _1160_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_289 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_72 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0991__D _0982_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_134 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0671__B1 _0487_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1183__CLK _1191_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_385 VGND VPWR sky130_fd_sc_hd__decap_12
X_0504_ _1152_/Q _0584_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_39_201 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0703__B _0700_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_237 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_127 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0613__B _0701_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0708__A1 _0705_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1147__D _1155_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_215 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0892__B1 _0891_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_218 VGND VPWR sky130_fd_sc_hd__fill_2
X_0984_ _0843_/A _0984_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_67_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_259 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_229 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0714__A _0714_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_148 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_44 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0938__A1 _1196_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_88 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1060__B1 _1057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_204 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_30 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_373 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_52 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0608__B _0608_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0874__B1 _0873_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0624__A _0566_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0929__A1 _1188_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1051__B1 _1049_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1221__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_351 VGND VPWR sky130_fd_sc_hd__fill_2
X_1183_ d_fabric_in[17] _1183_/Q _1191_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0865__B1 _0844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_398 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0534__A _0616_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_284 VGND VPWR sky130_fd_sc_hd__decap_3
X_0967_ _0945_/Y _0966_/Y _0946_/X _0960_/X w_mask[1] VGND VPWR sky130_fd_sc_hd__a211o_4
X_0898_ _0895_/D _0877_/X _0897_/Y d_sram_in[10] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0700__C _0717_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0709__A _0501_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_365 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0856__B1 _0855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_262 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_98 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1033__B1 _1029_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0619__A _0597_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_170 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0847__B1 _0844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1160__D _1223_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_89 VGND VPWR sky130_fd_sc_hd__fill_1
X_0821_ _0663_/A _1114_/Q _1146_/Q _0779_/X d_fabric_out[31] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0752_ _0532_/X _0751_/X _0719_/X _0752_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0683_ _0674_/B _0679_/X _0681_/X _0683_/D _0684_/D VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0529__A _0528_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_170 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1117__CLK _1130_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_151 VGND VPWR sky130_fd_sc_hd__fill_2
X_1166_ d_fabric_in[0] d_sram_in[0] _1188_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_343 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_173 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_302 VGND VPWR sky130_fd_sc_hd__decap_4
X_1097_ _0795_/X _1097_/Q _1207_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_265 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_287 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_32 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_354 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_387 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_313 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_64 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_214 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0780__A2 _0778_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1155__D _1226_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_94 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0994__D _0972_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_343 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_365 VGND VPWR sky130_fd_sc_hd__fill_1
X_1020_ _0998_/X _1018_/X _1019_/X w_mask[10] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_46_140 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_11_0_clk clkbuf_3_5_0_clk/X _1130_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_34_324 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_184 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_165 VGND VPWR sky130_fd_sc_hd__fill_1
X_0804_ _0799_/X _1101_/Q _0594_/A _0801_/X d_fabric_out[18] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0735_ _0676_/A _0669_/X _0739_/D _0695_/X _0655_/B _0735_/X VGND VPWR sky130_fd_sc_hd__a32o_4
X_0666_ _0663_/X _0660_/X _0665_/X d_fabric_out[0] VGND VPWR sky130_fd_sc_hd__a21o_4
X_0597_ _0726_/D _0689_/B _0596_/Y _0597_/X VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__0781__A1_N _0674_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1218_ addr_r[6] baseaddr_r_sync[6] _1131_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_110 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_335 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_195 VGND VPWR sky130_fd_sc_hd__fill_2
X_1149_ _1149_/D _0620_/A _1196_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0722__A _0722_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_22 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_31 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_75 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_143 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_379 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_0_0_clk clkbuf_3_1_0_clk/A clkbuf_3_0_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0616__B _0616_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_338 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_68 VGND VPWR sky130_fd_sc_hd__decap_12
X_0520_ _0682_/C _0721_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_3_261 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0753__A2 _0495_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_235 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_268 VGND VPWR sky130_fd_sc_hd__decap_6
X_1003_ _0972_/A _1031_/D VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_19_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_165 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_187 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_371 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0542__A _0681_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0899__D _1177_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0718_ _0718_/A _0716_/X _0501_/X _0717_/X _0718_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_0649_ _0626_/Y _0632_/X _0636_/Y _0647_/X _0648_/Y _0649_/X VGND VPWR sky130_fd_sc_hd__o41a_4
XFILLER_25_132 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0717__A _0717_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_165 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_99 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0602__D _0602_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0735__A2 _0669_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_84 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0627__A _0562_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_143 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_198 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_187 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0671__A1 _0676_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_157 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0671__B2 _0655_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_179 VGND VPWR sky130_fd_sc_hd__fill_2
X_0503_ _1150_/Q _0616_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_39_257 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_113 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0703__C _0701_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_290 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_157 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_168 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_53 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_190 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_64 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0613__C _0594_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_97 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0708__A2 _0706_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0910__A _0910_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1163__D _1163_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_94 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0892__A1 _0827_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1150__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_293 VGND VPWR sky130_fd_sc_hd__fill_2
X_0983_ _0983_/A _0983_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0898__B1_N _0897_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_238 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0714__B _1084_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_23 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0938__A2 _0876_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1060__A1 _0992_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_304 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1173__CLK _1191_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_238 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0874__A1 _0872_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_219 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0905__A _0905_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0929__A2 _0926_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1051__A1 _0966_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1158__D _1158_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0640__A _0566_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_164 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_7 VGND VPWR sky130_fd_sc_hd__fill_2
X_1182_ d_fabric_in[16] _1182_/Q _1191_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_49_363 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0865__A1 _0827_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_282 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_219 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_293 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0815__A out_reg VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_263 VGND VPWR sky130_fd_sc_hd__fill_1
X_0966_ _0966_/A _0966_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0550__A _0549_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0897_ _0897_/A _0897_/B _0897_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__0700__D _1130_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1196__CLK _1196_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_333 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0856__A1 _0851_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0725__A _0725_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_403 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_44 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_77 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1033__A1 _0944_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_15 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0619__B _0612_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0847__A1 _0880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_344 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_355 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_366 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0635__A _0526_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0820_ _0663_/A _1113_/Q _1113_/D _0815_/X d_fabric_out[30] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0751_ _0668_/X _1127_/Q _0634_/X _0751_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_0682_ _0722_/A _0679_/B _0682_/C _1128_/Q _0683_/D VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_36_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_300 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_182 VGND VPWR sky130_fd_sc_hd__fill_1
X_1165_ _1165_/D csb1_sync _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_185 VGND VPWR sky130_fd_sc_hd__fill_2
X_1096_ _0793_/X _1096_/Q _1096_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0545__A _0540_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_391 VGND VPWR sky130_fd_sc_hd__decap_6
X_0949_ _1010_/A _1045_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0774__B1 _0709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_108 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0829__A1 _0880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1211__CLK _1133_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_336 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_32 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_226 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0765__B1 _0668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_108 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_322 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1171__D d_fabric_in[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_314 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_391 VGND VPWR sky130_fd_sc_hd__decap_6
X_0803_ _0799_/X _1100_/Q _0487_/X _0801_/X d_fabric_out[17] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_6_270 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0756__B1 _0755_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0734_ _0663_/X _1085_/D _0733_/X d_fabric_out[2] VGND VPWR sky130_fd_sc_hd__a21o_4
X_0665_ _1083_/Q _0665_/B _0665_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0596_ _1134_/Q _0530_/X _0718_/A _0526_/X _0595_/X _0596_/Y VGND VPWR sky130_fd_sc_hd__a2111oi_4
XFILLER_29_108 VGND VPWR sky130_fd_sc_hd__fill_2
X_1217_ addr_r[5] baseaddr_r_sync[5] _1096_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_325 VGND VPWR sky130_fd_sc_hd__fill_2
X_1148_ _1156_/Q _0498_/A _1155_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1079_ _0984_/X _1040_/X _1075_/Y _1079_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_40_306 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_317 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_177 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0778__A2_N _0496_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_328 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0722__B _0492_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0747__B1 _0695_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_141 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_20 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0616__C _1146_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1107__CLK _1104_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1166__D d_fabric_in[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_130 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_174 VGND VPWR sky130_fd_sc_hd__fill_2
X_1002_ _0998_/X _1001_/X _0996_/X w_mask[7] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_22_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0823__A _1226_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_383 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0542__B _0726_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0717_ _0717_/A _0717_/B _0717_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0648_ _0509_/A _0703_/A _0622_/Y _0648_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_0579_ _0616_/D _0530_/X _0579_/C _1130_/Q _0579_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_25_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_111 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0717__B _0717_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_23 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_155 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_56 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_45 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_78 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0733__A _0732_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_361 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_10_0_clk clkbuf_3_5_0_clk/X _1163_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0735__A3 _0739_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_210 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_247 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0908__A _0903_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_52 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_239 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_122 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_114 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0671__A2 _0669_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_361 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0643__A _0584_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0959__B1 _0958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_398 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0795__A1_N _0575_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0502_ _0502_/A _0509_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_39_225 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_239 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_125 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_147 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_158 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0553__A _0608_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0703__D _0702_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_90 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0728__A _0728_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_217 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_87 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0613__D _1141_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0910__B _0909_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_51 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0638__A _0717_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0892__A2 _0890_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0982_ _0982_/A _0982_/B _0982_/C _0982_/D _0983_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_8_162 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_3 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_217 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0548__A _0547_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_397 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_57 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1060__A2 _1059_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_316 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_76 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0874__A2 _0875_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_294 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_231 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0905__B _0904_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_286 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1051__A2 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_132 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_176 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1174__D d_fabric_in[8] VGND VPWR sky130_fd_sc_hd__diode_2
X_1181_ d_fabric_in[15] _1181_/Q _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_345 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0865__A2 _0859_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0965_ _0964_/X _0966_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0831__A _1226_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0896_ _0846_/A _0890_/X _0895_/X _0897_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1084__D _1084_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_106 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_117 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_80 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_139 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_183 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_312 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_345 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0856__A2 _0833_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0725__B _0491_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1033__A2 _1032_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0741__A _0510_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1140__CLK _1108_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_42 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0619__C _0618_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_312 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_97 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0847__A2 _0859_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_389 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0916__A _0903_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0635__B _0635_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_286 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1169__D d_fabric_in[3] VGND VPWR sky130_fd_sc_hd__diode_2
X_0750_ _0750_/A _0750_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0651__A _0500_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0681_ _0681_/A _0492_/C _0723_/C _0487_/X _0681_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_29_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_109 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_334 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_367 VGND VPWR sky130_fd_sc_hd__decap_8
X_1164_ web web0_sync _1145_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1095_ _1095_/D _1095_/Q _1207_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0545__B _0545_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1163__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0948_ _0969_/A _1010_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0561__A _0585_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0879_ _0878_/Y _0880_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0774__A1 _1122_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_312 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0829__A2 _0828_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_131 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0765__B2 _0724_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_301 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0646__A _0642_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_367 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_337 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1186__CLK _1130_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0802_ _0799_/X _1099_/Q _0655_/A _0801_/X d_fabric_out[16] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__0756__A1 _0663_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0733_ _0732_/X _1085_/Q _0733_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0664_ out_reg _0665_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0595_ _1132_/Q _0582_/X _0595_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_1216_ addr_r[4] baseaddr_r_sync[4] _1104_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0556__A _0581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_175 VGND VPWR sky130_fd_sc_hd__fill_2
X_1147_ _1155_/Q _1147_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_359 VGND VPWR sky130_fd_sc_hd__decap_6
X_1078_ _1032_/X _1070_/X _1076_/X w_mask[29] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_52_145 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0722__C _0723_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0747__A1 _0750_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0747__B2 _0495_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_54 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_167 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_370 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0616__D _0616_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_178 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1182__D d_fabric_in[16] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_153 VGND VPWR sky130_fd_sc_hd__fill_2
X_1001_ _1000_/X _1001_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_34_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_145 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1000__A _0973_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_395 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0542__C _0679_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0716_ _0668_/A _0716_/B _0716_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1201__CLK _1096_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0647_ _0647_/A _0647_/B _0647_/C _0646_/X _0647_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_0578_ _0559_/X _0578_/B _0574_/Y _0577_/X _0578_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XANTENNA__1092__D _0781_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_259 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_178 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_340 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0733__B _1085_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_204 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0908__B _0903_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_101 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_292 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0671__A3 _0676_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0643__B _0644_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0959__A1 _1065_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_333 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1081__B1 _1079_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1224__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1177__D d_fabric_in[11] VGND VPWR sky130_fd_sc_hd__diode_2
X_0501_ _0500_/X _0501_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_11_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_251 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0834__A _0845_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_273 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1072__B1 _1071_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1087__D _1087_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0728__B _0728_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_207 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_56 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_67 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0744__A _0738_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_262 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1063__B1 _1061_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_303 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0810__B1 _0723_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_63 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_85 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0638__B _0558_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_281 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0654__A _0654_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_251 VGND VPWR sky130_fd_sc_hd__fill_2
X_0981_ _1007_/A _0982_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_12_170 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1054__B1 _1052_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_380 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_354 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0868__B1 _0867_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_240 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0564__A _0555_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_295 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_328 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0739__A _0722_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_321 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_229 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_218 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_276 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_144 VGND VPWR sky130_fd_sc_hd__decap_12
X_1180_ d_fabric_in[14] _0912_/D _1145_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1190__D d_fabric_in[24] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_221 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_276 VGND VPWR sky130_fd_sc_hd__fill_2
X_0964_ _1007_/A _1021_/B _1209_/Q _0972_/A _0964_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0831__B _1156_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0895_ _0899_/A _0899_/B _0903_/C _0895_/D _0895_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1092__CLK _1145_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_357 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0725__C _0726_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0741__B _0726_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_32 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0916__B _0903_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0635__C _0634_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_276 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0932__A _0876_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0680_ _0679_/C _0723_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1185__D d_fabric_in[19] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_313 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_184 VGND VPWR sky130_fd_sc_hd__decap_6
X_1163_ _1163_/D csb0_sync _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1094_ _0788_/X _1094_/Q _1096_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_316 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_390 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1003__A _0972_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0545__C _0545_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_224 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0842__A _0841_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0947_ _0940_/A _0969_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0561__B _0555_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_279 VGND VPWR sky130_fd_sc_hd__fill_2
X_0878_ _0838_/A _0878_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0774__A2 _0497_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1095__D _1095_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_23 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_78 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_89 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_77 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_110 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0646__B _0643_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_168 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0662__A _0661_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0801_ _0665_/B _0801_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0756__A2 _1087_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0732_ out_reg _0732_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0610__D1 _0609_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0663_ _0663_/A _0663_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0594_ _0594_/A _0594_/B _0718_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_41_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_1215_ addr_r[3] baseaddr_r_sync[3] _1133_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_110 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0837__A _0836_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1146_ d_sram_out[31] _1146_/Q _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0556__B _0489_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_102 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1130__CLK _1130_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1077_ _1025_/X _1070_/X _1076_/X w_mask[28] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_33_360 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_371 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0572__A _0571_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0722__D _0717_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0747__A2 _0736_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_36 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_11 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_349 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_77 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_319 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_382 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_43 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_98 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_80 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_227 VGND VPWR sky130_fd_sc_hd__decap_8
X_1000_ _0973_/A _0952_/B _0999_/X _0982_/D _1000_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__1153__CLK _1130_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_157 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_clk_A clk VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1000__B _0952_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0542__D _0634_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0715_ _0663_/X _1084_/D _0714_/X d_fabric_out[1] VGND VPWR sky130_fd_sc_hd__a21o_4
X_0646_ _0642_/X _0643_/X _0644_/X _0645_/X _0646_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA_clkbuf_4_9_0_clk_A clkbuf_3_4_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0577_ _0575_/Y _0576_/X _0574_/A _0553_/X _0577_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_57_205 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0567__A _0606_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_249 VGND VPWR sky130_fd_sc_hd__fill_2
X_1129_ d_sram_out[14] _0724_/D _1104_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_40_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_79 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1176__CLK _1188_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0908__C _0908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_130 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_190 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_301 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0643__C _0529_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0959__A2 _0838_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_385 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1081__A1 _1040_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0940__A _0940_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0500_ _0499_/X _0500_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1193__D d_fabric_in[27] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_105 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1011__A _1009_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1072__A1 _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_70 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1199__CLK _1130_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0629_ _0628_/X _0703_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0728__C _0723_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_127 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0744__B _0739_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_296 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_160 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1063__A1 _1001_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_56 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0810__B2 _0808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0810__A1 _0806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_0980_ _0968_/X _0979_/X _0975_/Y w_mask[3] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__1188__D d_fabric_in[22] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1054__A1 _0979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0670__A _0602_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_182 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_392 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_311 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_366 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1006__A _1005_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0868__A1 _0864_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0845__A _0845_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_403 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_222 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_244 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1098__D _1098_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_288 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0580__A _0616_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0739__B _0492_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_clk_A clkbuf_3_7_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_12 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_34 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1214__CLK _1188_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0755__A _0732_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_285 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_255 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0490__A _0489_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0795__B1 _1113_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_322 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_355 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0665__A _1083_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0963_ _0950_/Y _1021_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0786__B1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0831__C _0831_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0894_ _0891_/D _0877_/X _0893_/Y d_sram_in[9] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_4_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_325 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0575__A _0724_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0710__B1 _0709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_200 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0725__D _0594_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_266 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0741__C _0741_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0777__B1 _0776_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_174 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0916__C _0908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0768__B1 _0766_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_163 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_347 VGND VPWR sky130_fd_sc_hd__decap_12
X_1162_ _1225_/Q _1162_/Q _1184_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1093_ _0784_/X _1093_/Q _1096_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_361 VGND VPWR sky130_fd_sc_hd__decap_12
X_0946_ _0859_/B _0946_/B _0946_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0561__C _1151_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_269 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0759__B1 _0719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_281 VGND VPWR sky130_fd_sc_hd__decap_12
X_0877_ _0876_/X _0877_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_18_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_391 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_57 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_269 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_56 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_314 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_3_0_clk_A clkbuf_2_2_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_347 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0646__C _0644_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_144 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_103 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0943__A _0836_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_147 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0989__B1 _0988_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0800_ _0714_/A _1098_/D _0799_/X _1098_/Q d_fabric_out[15] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0731_ _0750_/A _0718_/X _0730_/X _0594_/A _0711_/X _1085_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__1196__D d_fabric_in[30] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0610__C1 _0608_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0662_ _0661_/Y _0663_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0593_ _0586_/C _0594_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_34_3 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0913__B1 _0912_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_50 VGND VPWR sky130_fd_sc_hd__decap_8
X_1214_ addr_r[2] baseaddr_r_sync[2] _1188_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0837__B _0845_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_155 VGND VPWR sky130_fd_sc_hd__fill_2
X_1145_ d_sram_out[30] _1113_/D _1145_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0556__C _1152_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1014__A _0982_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_125 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_391 VGND VPWR sky130_fd_sc_hd__decap_6
X_1076_ _0984_/X _1035_/X _1075_/Y _1076_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA_clkbuf_4_5_0_clk_A clkbuf_4_5_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0929_ _1188_/Q _0926_/X _0870_/X d_sram_in[22] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0747__A3 _0746_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_59 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0904__B1 _0903_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_306 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_114 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_350 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0763__A _0732_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_394 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_191 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_287 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_188 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0673__A _0673_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_331 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1000__C _0999_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0714_ _0714_/A _1084_/Q _0714_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0645_ _0606_/A _0644_/B _0529_/Y _0721_/D _0645_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1009__A _1046_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0576_ _0587_/A _0584_/B _0725_/A _0616_/B _0576_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0848__A _0897_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0567__B _0566_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1128_ d_sram_out[13] _1128_/Q _1130_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_48 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0583__A _0606_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1059_ _1042_/Y _1059_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_31_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_213 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0908__D _0908_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_44 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_147 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0493__A _0493_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_131 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0643__D _0724_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_313 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1081__A2 _1042_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0940__B _1207_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1120__CLK _1131_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0668__A _0668_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_1_0_0_clk_A clkbuf_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0577__A1_N _0575_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_272 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_139 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1011__B _1011_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_172 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1072__A2 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_183 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_194 VGND VPWR sky130_fd_sc_hd__decap_8
X_0628_ _0566_/X _0553_/X _0628_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0578__A _0559_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0559_ _0554_/Y _0604_/A _1128_/Q _0558_/X _0559_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__0728__D _0727_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_294 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_275 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0744__C _0740_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_clk_A clkbuf_3_3_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1063__A2 _1059_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0810__A2 _1105_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1143__CLK _1096_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0488__A _1147_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_209 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_13_0_clk_A clkbuf_3_6_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_294 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_297 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_91 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0951__A _0950_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_121 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1054__A2 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_154 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_301 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0868__A2 _0833_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_209 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0845__B _0845_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1022__A _1021_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1166__CLK _1188_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0861__A _0905_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0580__B _0566_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0739__C _0723_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0755__B _1087_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_245 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0771__A _1138_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0795__B2 _0711_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_352 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_396 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_304 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0946__A _0859_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_367 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_389 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_264 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0665__B _0665_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_286 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1189__CLK _1184_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_256 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1199__D addr_w[1] VGND VPWR sky130_fd_sc_hd__diode_2
X_0962_ _0940_/A _1007_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_32_267 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0681__A _0681_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0786__B2 _1093_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0786__A1 _0779_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0893_ _0910_/A _0892_/X _0893_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_64_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1017__A _0973_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_175 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0710__A1 _0685_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_26 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0591__A _0552_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_48 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0741__D _1130_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0777__A1 _0762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_67 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_304 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_44 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0916__D _1181_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_223 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0768__B2 _0767_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0768__A1 _0723_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_182 VGND VPWR sky130_fd_sc_hd__fill_1
X_1161_ _1224_/Q _1161_/Q _1130_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0676__A _0676_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_112 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_326 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_359 VGND VPWR sky130_fd_sc_hd__decap_6
X_1092_ _0781_/X _1092_/Q _1145_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_60_373 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_237 VGND VPWR sky130_fd_sc_hd__fill_2
X_0945_ _0944_/X _0945_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0561__D _1150_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0759__A1 _0757_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_293 VGND VPWR sky130_fd_sc_hd__decap_12
X_0876_ _0876_/A _0876_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1204__CLK _1133_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1_0_clk_A clkbuf_3_0_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0931__A1 _1190_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0586__A _0585_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_36 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_351 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_403 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_66 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0496__A _0495_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_359 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0646__D _0645_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_115 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_159 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0989__A1 _0985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0943__B _0845_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1227__CLK _1133_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_91 VGND VPWR sky130_fd_sc_hd__fill_1
X_0730_ _1117_/Q _0548_/X _0719_/X _0729_/X _0730_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__0610__B1 _0688_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0661_ out_reg _0661_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_6_274 VGND VPWR sky130_fd_sc_hd__fill_1
X_0592_ _0579_/C _0689_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0913__A1 _1172_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1213_ addr_r[1] baseaddr_r_sync[1] _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_27_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0837__C _0831_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1144_ d_sram_out[29] _1112_/D _1207_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_1_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_370 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0556__D _0555_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1014__B _1021_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_329 VGND VPWR sky130_fd_sc_hd__decap_4
X_1075_ _1066_/B _1075_/B _1048_/C _1075_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_52_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_340 VGND VPWR sky130_fd_sc_hd__fill_2
X_0928_ _1187_/Q _0926_/X _0867_/X d_sram_in[21] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0859_ _0859_/A _0859_/B _0859_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0904__A1 _1170_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_46 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0763__B _0763_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_299 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0605__A2_N _0562_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_101 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0954__A _0999_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_178 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_181 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_343 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_398 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1000__D _0982_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0713_ out_reg _0714_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0644_ _0616_/D _0644_/B _0582_/A _0716_/B _0644_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1009__B _1046_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0575_ _0724_/D _0575_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0567__C _0529_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1025__A _1025_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1127_ d_sram_out[12] _1127_/Q _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_115 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0864__A _1171_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_27 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0583__B _0579_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_159 VGND VPWR sky130_fd_sc_hd__decap_3
X_1058_ _0983_/X _1043_/X _1057_/X w_mask[20] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_40_118 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_192 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_126 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_132 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_118 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_110 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_325 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0940__C _1209_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_398 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0949__A _1010_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_240 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0559__A2_N _0604_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0684__A _0684_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_210 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_265 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1057__B1 _1056_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0804__B1 _0594_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1011__C _0959_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_0627_ _0562_/X _0627_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0859__A _0859_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0578__B _0578_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0558_ _0584_/A _1153_/Q _0725_/A _0616_/B _0558_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1095__CLK _1207_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0489_ _1150_/Q _0489_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_26_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_251 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0594__A _0594_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_232 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0744__D _0744_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0769__A _0732_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_55 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_232 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_clk clkbuf_2_2_0_clk/A clkbuf_3_7_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_8_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_177 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_80 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0679__A _0722_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_335 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_232 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0845__C _0845_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_287 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_279 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0580__C _0530_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0589__A _0579_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0961__C1 _0960_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0739__D _0739_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_298 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1110__CLK _1108_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0771__B _0655_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_103 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0894__B1_N _0893_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0499__A _0620_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_316 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0946__B _0946_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0962__A _0940_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_235 VGND VPWR sky130_fd_sc_hd__decap_8
X_0961_ _0946_/B _0945_/Y _0946_/X _0960_/X w_mask[0] VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__0681__B _0492_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0786__A2 _0784_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0892_ _0827_/A _0890_/X _0891_/X _0892_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_57_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1017__B _0982_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_187 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0710__A2 _0708_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1133__CLK _1133_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_371 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_213 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0872__A _1173_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_279 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0591__B _0591_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0777__A2 _1090_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_213 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0768__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0957__A _1010_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_7 VGND VPWR sky130_fd_sc_hd__fill_2
X_1160_ _1223_/Q _1160_/Q _1152_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0676__B _0492_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1156__CLK _1155_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1091_ _0778_/X _1091_/Q _1145_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_308 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0692__A _0739_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0944_ _0943_/X _0944_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0759__A2 _0758_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0875_ _0875_/A _0876_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1028__A _1011_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0931__A2 _0926_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_305 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0586__B _0584_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_316 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_179 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_363 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_396 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1179__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_157 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_371 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0989__A2 _0974_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0943__C _0908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_70 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0610__A1 _0675_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0660_ _0487_/X _0496_/X _0659_/X _0660_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0591_ _0552_/Y _0591_/B _0591_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_40_91 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0687__A _0675_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0913__A2 _0880_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1212_ addr_r[0] baseaddr_r_sync[0] _1188_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_1_74 VGND VPWR sky130_fd_sc_hd__decap_4
X_1143_ d_sram_out[28] _0532_/A _1096_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1014__C _1021_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1074_ _1046_/A _1065_/B _1045_/C _1045_/D _1075_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_37_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_190 VGND VPWR sky130_fd_sc_hd__fill_2
X_0927_ _1186_/Q _0926_/X _0862_/X d_sram_in[20] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0858_ _0852_/B _0859_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0789_ _0779_/X _0788_/X _0785_/X _1094_/Q d_fabric_out[11] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__0597__A _0726_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0904__A2 _0890_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_69 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_127 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_311 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0970__A _1207_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0712_ _0750_/A _0672_/X _0710_/Y _0487_/X _0711_/X _1084_/D VGND VPWR sky130_fd_sc_hd__a32o_4
X_0643_ _0584_/A _0644_/B _0529_/Y _0724_/D _0643_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1009__C _0982_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0574_ _0574_/A _0579_/C _0573_/Y _0574_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0898__A1 _0895_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0567__D _0702_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1126_ d_sram_out[11] _1126_/Q _1145_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0583__C _0582_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1057_ _1044_/X _1018_/X _1056_/Y _1057_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_33_171 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0880__A _0880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_259 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_208 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0889__A1 _1174_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1217__CLK _1096_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_300 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_111 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1101__D _0594_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_182 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0940__D _0972_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0577__B1 _0574_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0965__A _0964_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0684__B _0676_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_296 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_160 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1057__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_288 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0804__A1 _0799_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk clk clkbuf_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XANTENNA__0804__B2 _0801_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0568__B1 _0567_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_62 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_51 VGND VPWR sky130_fd_sc_hd__decap_8
X_0626_ _0682_/C _0686_/C _0626_/C _0626_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0859__B _0859_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0578__C _0574_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0557_ _0556_/X _0604_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1036__A _0959_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_230 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0875__A _0875_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0488_ _1147_/Q _0488_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_38_263 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_27 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0594__B _0594_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_285 VGND VPWR sky130_fd_sc_hd__decap_3
X_1109_ _1141_/Q _1109_/Q _1096_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_13_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_163 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0559__B1 _1128_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0769__B _1089_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0785__A _0663_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0731__B1 _0594_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_274 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_244 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_255 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_141 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0798__B1 _0797_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0679__B _0679_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0695__A _1134_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_211 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_299 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0789__B1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_269 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0580__D _1122_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0961__B1 _0946_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0589__B _0589_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0609_ _0723_/D _0594_/B _0609_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_58_303 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_380 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_266 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_36 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_115 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0499__B _1147_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_255 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_0960_ _0988_/A _0955_/X _0959_/Y _0960_/X VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__0681__C _0723_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1085__CLK _1130_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0891_ _0899_/A _0899_/B _0903_/C _0891_/D _0891_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_67_122 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1017__C _1021_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_306 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_391 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_129 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_clk clkbuf_2_2_0_clk/A clkbuf_3_5_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_46_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_199 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_339 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0676__C _0676_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_199 VGND VPWR sky130_fd_sc_hd__fill_2
X_1090_ _1090_/D _1090_/Q _1155_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0973__A _0973_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0692__B _0558_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_320 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_228 VGND VPWR sky130_fd_sc_hd__fill_2
X_0943_ _0836_/Y _0845_/B _0908_/C _1042_/D _0943_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_0874_ _0872_/Y _0875_/A _0873_/X d_sram_in[7] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__1028__B _1028_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1100__CLK _1196_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0586__C _0586_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_328 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1044__A _0843_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_147 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0883__A _0883_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_331 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_26 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_306 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_339 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_125 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1104__D _0675_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_383 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_180 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0943__D _1042_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_191 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_375 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0610__A2 _0582_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1123__CLK _1145_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0590_ _0682_/C _0553_/X _0509_/A _0578_/Y _0589_/Y _0591_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__0968__A _0943_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0687__B _0654_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1211_ addr_w[13] _1042_/D _1133_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_1_31 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_114 VGND VPWR sky130_fd_sc_hd__fill_2
X_1142_ d_sram_out[27] _0691_/A _1096_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1014__D _1021_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1073_ _1022_/X _1070_/X _1071_/X w_mask[27] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_33_375 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_150 VGND VPWR sky130_fd_sc_hd__decap_3
X_0926_ _0876_/A _0926_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1039__A _1010_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0857_ _1170_/Q _0857_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0788_ _0554_/Y _0787_/X _0739_/D _0787_/X _0788_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__0878__A _0838_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0597__B _0689_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_139 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_47 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1146__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_257 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_84 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_294 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_150 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_323 VGND VPWR sky130_fd_sc_hd__fill_2
X_0711_ _0497_/X _0711_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0642_ _0587_/A _0644_/B _0586_/C _0540_/D _0642_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0698__A _0697_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0573_ _0540_/D _0608_/B _0721_/D _0586_/C _0573_/Y VGND VPWR sky130_fd_sc_hd__a22oi_4
XANTENNA__1009__D _1045_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0898__A2 _0877_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1125_ d_sram_out[10] _0716_/B _1131_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0583__D _0673_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1056_ _1048_/B _1055_/X _1048_/C _1056_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__1169__CLK _1188_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_323 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0880__B _0880_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_0909_ _1171_/Q _0890_/X _0908_/X _0909_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_0_249 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0889__A2 _0877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_242 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_134 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_161 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0577__B2 _0553_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0684__C _0684_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0981__A _1007_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_109 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1057__A2 _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0804__A2 _1101_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_131 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0568__A1 _0560_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_96 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_74 VGND VPWR sky130_fd_sc_hd__fill_2
X_0625_ _0614_/Y _0528_/X _0603_/Y _0571_/X _0626_/C VGND VPWR sky130_fd_sc_hd__o22a_4
X_0556_ _0581_/A _0489_/Y _1152_/Q _0555_/Y _0556_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0578__D _0577_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1036__B _1029_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0487_ _1132_/Q _0487_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_1108_ _0602_/D _1108_/Q _1108_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_13_109 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1202__D addr_w[4] VGND VPWR sky130_fd_sc_hd__diode_2
X_1039_ _1010_/A _1021_/B _0999_/X _1031_/D _1039_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0891__A _0899_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_49 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_175 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0559__B2 _0558_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0731__A1 _0750_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0731__B2 _0711_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_50 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1112__D _1112_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0788__A2_N _0787_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_289 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_72 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0798__A1 _1130_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_186 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_93 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0679__C _0679_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_215 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_226 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_248 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0789__B2 _1094_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0789__A1 _0779_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1207__CLK _1207_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0961__A1 _0946_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0589__C _0589_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0608_ _0634_/A _0608_/B _0608_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0539_ _0725_/A _0681_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0886__A _0908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_38 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_392 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_15 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_48 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_300 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0499__C _0620_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1107__D _0543_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_359 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_201 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_245 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_204 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_215 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0681__D _0487_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0890_ _0880_/B _0890_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_4_86 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1017__D _1021_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_329 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0790__A1_N _0560_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0934__A1 _1192_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_112 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_215 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0870__B1 _0848_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_40 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_62 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0925__A1 _1185_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_174 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_196 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_134 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0676__D _0676_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0973__B _0982_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_351 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_362 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_398 VGND VPWR sky130_fd_sc_hd__decap_6
X_0942_ _0942_/A _0946_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_13_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_281 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_230 VGND VPWR sky130_fd_sc_hd__decap_6
X_0873_ _0872_/Y _0839_/A _0854_/Y _0873_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_62_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0586__D _1117_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_362 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_207 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1210__D addr_w[12] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_318 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_362 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_395 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_332 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_398 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1120__D d_sram_out[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_240 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_288 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1020__B1 _1019_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1210_ addr_w[12] _0972_/A _1152_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1141_ d_sram_out[26] _1141_/Q _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0984__A _0843_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1072_ _1018_/X _1070_/X _1071_/X w_mask[26] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_37_159 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_1_0_clk clkbuf_1_0_0_clk/X clkbuf_3_3_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_33_387 VGND VPWR sky130_fd_sc_hd__decap_12
X_0925_ _1185_/Q _0907_/X _0855_/X d_sram_in[19] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0906__B1_N _0905_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1039__B _1021_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0856_ _0851_/Y _0833_/X _0855_/X d_sram_in[3] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0787_ _0495_/X _0787_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1098__CLK _1155_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1055__A _1045_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0597__C _0596_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_137 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_148 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1205__D addr_w[7] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1078__B1 _1076_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_321 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_181 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1002__B1 _0996_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_72 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_126 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1115__D d_sram_out[0] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1069__B1 _1067_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0816__B1 _0717_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_335 VGND VPWR sky130_fd_sc_hd__fill_1
X_0710_ _0685_/X _0708_/Y _0709_/X _0710_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0641_ _0697_/A _0694_/B _0633_/B _1117_/Q _0647_/C VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0979__A _0978_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0572_ _0571_/X _0586_/C VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0698__B _0694_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_280 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_243 VGND VPWR sky130_fd_sc_hd__fill_1
X_1124_ d_sram_out[9] _0673_/A _1104_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1055_ _1045_/A _1065_/B _1045_/C _1045_/D _1055_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0807__B1 _0634_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_357 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_0908_ _0903_/A _0903_/B _0908_/C _0908_/D _0908_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0839_ _0839_/A _0839_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_206 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_254 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1113__CLK _1130_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_102 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_324 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0799__A _0661_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_73 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_254 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0684__D _0684_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_4 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_184 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_173 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_110 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_187 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0568__A2 _0562_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0624_ _0566_/X _0686_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0502__A _0502_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0555_ _1153_/Q _0555_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0486_ reb csb _1165_/D VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1136__CLK _1104_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1107_ _0543_/A _1107_/Q _1104_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1038_ _0944_/X _1035_/X _1037_/X w_mask[14] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0891__B _0899_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_279 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_58 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_221 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0731__A2 _0718_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_298 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0798__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_331 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0679__D _0757_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1159__CLK _1191_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0992__A _0992_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_279 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0789__A2 _0788_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_191 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0961__A2 _0945_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0589__D _0589_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0607_ _1138_/Q _0529_/Y _0688_/A VGND VPWR sky130_fd_sc_hd__and2_4
X_0538_ _0581_/A _0725_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_58_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1213__D addr_r[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_367 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_213 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1123__D d_sram_out[8] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_268 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_271 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_293 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0987__A _1045_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_146 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_330 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1208__D addr_w[10] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0897__A _0897_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0934__A2 _0932_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_38 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_124 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_308 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_48 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_227 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_205 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_249 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0870__A1 _0869_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_293 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_85 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0925__A2 _0907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0600__A _0606_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1118__D d_sram_out[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_157 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0973__C _1045_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_300 VGND VPWR sky130_fd_sc_hd__decap_6
X_0941_ _0941_/A _0942_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0872_ _1173_/Q _0872_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_55_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0510__A _1151_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_308 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_374 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_193 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_219 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_344 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_355 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_252 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1020__A1 _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_70 VGND VPWR sky130_fd_sc_hd__fill_2
X_1140_ d_sram_out[25] _0602_/D _1108_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_1_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_99 VGND VPWR sky130_fd_sc_hd__fill_2
X_1071_ _0984_/X _1032_/X _1066_/Y _1071_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_33_344 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_130 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_399 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0505__A _0616_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0924_ _1184_/Q _0907_/X _0849_/X d_sram_in[18] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0855_ _0851_/Y _0839_/X _0854_/Y _0855_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1039__C _0999_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0786_ _0779_/X _0784_/X _0785_/X _1093_/Q d_fabric_out[10] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1055__B _1065_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0770__B1 _0769_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_127 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_17 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1078__A1 _1032_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1221__D addr_r[9] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_163 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1002__A1 _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0761__B1 _0759_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1192__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_62 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1069__A1 _1015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_119 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0816__A1 _0813_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0816__B2 _0815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1131__D d_sram_out[16] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_185 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_196 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_93 VGND VPWR sky130_fd_sc_hd__fill_1
X_0640_ _0566_/X _0694_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0571_ _0570_/X _0571_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0698__C _0594_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_292 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0995__A _0995_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0752__B1 _0719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_3 VGND VPWR sky130_fd_sc_hd__fill_1
X_1123_ d_sram_out[8] _0502_/A _1145_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_119 VGND VPWR sky130_fd_sc_hd__fill_1
X_1054_ _0979_/X _1043_/X _1052_/X w_mask[19] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0807__A1 _0806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0807__B2 _0801_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_336 VGND VPWR sky130_fd_sc_hd__fill_2
X_0907_ _0876_/A _0907_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0838_ _0838_/A _0838_/B _0839_/A VGND VPWR sky130_fd_sc_hd__and2_4
X_0769_ _0732_/X _1089_/Q _0769_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_0_218 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1066__A _1066_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1216__D addr_r[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_403 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_288 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_125 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0734__B1 _0733_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_0_0_clk clkbuf_1_0_0_clk/X clkbuf_3_1_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__1126__D d_sram_out[11] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_152 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_141 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_196 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1088__CLK _1155_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_0623_ _1115_/Q _0620_/X _0622_/Y _0623_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0554_ _1126_/Q _0554_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_38_200 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_222 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_19 VGND VPWR sky130_fd_sc_hd__fill_2
X_1106_ _1138_/Q _1106_/Q _1104_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1037_ _0985_/X _1001_/X _1036_/Y _1037_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0891__C _0903_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_280 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_15 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0731__A3 _0730_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_247 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_122 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_291 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_126 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_148 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0603__A _0532_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_398 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0707__B1 _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_92 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_258 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_206 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_291 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0513__A _0616_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1103__CLK _1133_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0606_ _0606_/A _0741_/C VGND VPWR sky130_fd_sc_hd__buf_1
X_0537_ _0526_/X _0532_/X _0676_/C _0537_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_49_339 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_291 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_261 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1126__CLK _1145_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0987__B _1065_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_114 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_372 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_342 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0508__A _0508_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_280 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0897__B _0897_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1074__A _1046_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_136 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1224__D addr_r[12] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0870__A2 _0839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_261 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1149__CLK _1196_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_97 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1134__D d_sram_out[19] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_309 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_139 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0973__D _0982_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_386 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_93 VGND VPWR sky130_fd_sc_hd__decap_12
X_0940_ _0940_/A _1207_/Q _1209_/Q _0972_/A _0941_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_13_272 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_243 VGND VPWR sky130_fd_sc_hd__fill_1
X_0871_ _0869_/Y _0833_/X _0870_/X d_sram_in[6] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0998__A _0943_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_3 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_172 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0660__B1_N _0659_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_323 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_367 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1219__D addr_r[7] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0701__A _0741_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_367 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_96 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_264 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1129__D d_sram_out[14] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_246 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0611__A _0741_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1020__A2 _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_34 VGND VPWR sky130_fd_sc_hd__fill_2
X_1070_ _1042_/Y _1070_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_45_150 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_323 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_194 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_186 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0505__B _0584_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0923_ _1183_/Q _0876_/X _0844_/X _0922_/Y d_sram_in[17] VGND VPWR sky130_fd_sc_hd__a211o_4
X_0854_ _0854_/A _0854_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0785_ _0663_/A _0785_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1039__D _1031_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0521__A _0676_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0770__A1 _0762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1055__C _1045_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_106 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1078__A2 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1199_ addr_w[1] baseaddr_w_sync[1] _1130_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_356 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1002__A2 _1001_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_87 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0761__A1 _0675_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0761__B2 _0760_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_41 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_52 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_301 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1069__A2 _1059_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_334 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_312 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0816__A2 _1109_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_142 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0606__A _0606_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_315 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_337 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_359 VGND VPWR sky130_fd_sc_hd__decap_12
X_0570_ _0523_/A _1150_/Q _0570_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0698__D _0677_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0752__A1 _0532_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1122_ d_sram_out[7] _1122_/Q _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_150 VGND VPWR sky130_fd_sc_hd__decap_3
X_1053_ _0974_/X _1043_/X _1052_/X w_mask[18] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_18_183 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0807__A2 _1103_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0516__A _1152_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_315 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_175 VGND VPWR sky130_fd_sc_hd__fill_2
X_0906_ _1178_/Q _0877_/X _0905_/Y d_sram_in[12] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0837_ _0836_/Y _0845_/B _0831_/C _0838_/B VGND VPWR sky130_fd_sc_hd__or3_4
X_0768_ _0723_/D _0750_/X _0766_/X _0767_/X _1089_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1066__B _1066_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0699_ _0694_/X _0696_/X _0699_/C _0698_/X _0699_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__1082__A csb VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_267 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_104 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_164 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_186 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_370 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0734__A1 _0663_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1142__D d_sram_out[27] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_278 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_215 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_6 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_60 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_330 VGND VPWR sky130_fd_sc_hd__decap_12
X_0622_ _0620_/A _0488_/Y _0620_/C _0622_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_0553_ _0608_/B _0553_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_1105_ _0723_/D _1105_/Q _1104_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_38_267 VGND VPWR sky130_fd_sc_hd__fill_2
X_1036_ _0959_/Y _1029_/C _1036_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__0891__D _0891_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_19 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_156 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1182__CLK _1191_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1227__D conf[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_234 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_278 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_63 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_85 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1137__D d_sram_out[22] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0707__A1 _1116_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_270 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_229 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0605_ _0603_/Y _0562_/X _0691_/A _0604_/Y _0612_/C VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_0536_ _0726_/D _0676_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_53_18 VGND VPWR sky130_fd_sc_hd__fill_2
X_1019_ _0985_/X _0992_/X _1011_/Y _1019_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0704__A _0690_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0937__A1 _1195_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_325 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0919__B1_N _0918_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_318 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_30 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_41 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0873__B1 _0854_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_270 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0625__B1 _0603_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_403 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0614__A _1113_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_95 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1050__B1 _1049_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0928__A1 _1187_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_152 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0987__C _0982_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_362 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_354 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_240 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0524__A _0581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1041__B1 _1037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0919__A1 _1181_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1220__CLK _1188_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1074__B _1065_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0519_ _0574_/A _0682_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_58_148 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_170 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0855__B1 _0854_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_104 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0609__A _0723_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_354 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1150__D _1150_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_240 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_200 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_0870_ _0869_/Y _0839_/X _0848_/Y _0870_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1023__B1 _1019_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0519__A _0574_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_151 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_184 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_398 VGND VPWR sky130_fd_sc_hd__decap_6
X_0999_ _0999_/A _0999_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0701__B _0701_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_343 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1116__CLK _1196_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_313 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_258 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_74 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0611__B _0689_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1145__D d_sram_out[30] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_321 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_376 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0819__B1 _0757_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_302 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_143 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_198 VGND VPWR sky130_fd_sc_hd__decap_12
X_0922_ _0828_/X _0876_/X _0922_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_0853_ _0827_/A _0859_/B _0844_/X _0852_/X _0854_/A VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_60_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_0784_ _0717_/A _0711_/X _0783_/X _0784_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0521__B _0721_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1055__D _1045_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0770__A2 _1089_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1139__CLK _1133_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1198_ addr_w[0] baseaddr_w_sync[0] _1133_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_36_162 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_346 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_143 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_239 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0746__C1 _0745_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0761__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_121 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_327 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0622__A _0620_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0752__A2 _0751_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_257 VGND VPWR sky130_fd_sc_hd__decap_8
X_1121_ d_sram_out[6] _0721_/D _1196_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1052_ _1044_/X _1015_/X _1048_/Y _1052_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_33_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_143 VGND VPWR sky130_fd_sc_hd__fill_2
X_0905_ _0905_/A _0904_/X _0905_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__0532__A _0532_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0836_ _0845_/A _0836_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0767_ _0721_/D _0497_/X _0709_/X _0767_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1066__C _1048_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0698_ _0697_/A _0694_/B _0594_/B _0677_/D _0698_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1082__B web VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_121 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_105 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_176 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0967__C1 _0960_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_382 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0734__A2 _1085_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_7 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0617__A _0689_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_72 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_78 VGND VPWR sky130_fd_sc_hd__decap_12
X_0621_ _0591_/X _0619_/X _0620_/X _0621_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0552_ _1154_/Q _0552_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_38_213 VGND VPWR sky130_fd_sc_hd__fill_1
X_1104_ _0675_/D _1104_/Q _1104_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1035_ _1034_/X _1035_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0527__A _0581_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0819_ _0813_/X _1112_/Q _0757_/A _0815_/X d_fabric_out[29] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_29_257 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_87 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_102 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_20 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_356 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0707__A2 _0622_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1153__D _1161_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_219 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_161 VGND VPWR sky130_fd_sc_hd__fill_2
X_0604_ _0604_/A _0604_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0535_ _0535_/A _0726_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0615__A2_N _0576_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_205 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_249 VGND VPWR sky130_fd_sc_hd__fill_2
X_1018_ _1018_/A _1018_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0704__B _0704_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0937__A2 _0932_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0720__A _0716_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0873__A1 _0872_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_400 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0625__A1 _0614_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0625__B2 _0571_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_74 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1050__A1 _0942_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0928__A2 _0926_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1148__D _1156_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0630__A _0594_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0987__D _1045_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_392 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1172__CLK _1130_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_388 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_219 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0524__B _0491_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1041__A1 _0944_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0919__A2 _0907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0540__A _0681_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0518_ _0587_/A _0574_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1074__C _1045_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_341 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_396 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0855__A1 _0851_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_44 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0791__B1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1195__CLK _1184_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_52 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0609__B _0594_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_96 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_311 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1023__A1 _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_7 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0782__B1 _0762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_108 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0535__A _0535_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0998_ _0943_/X _0998_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0701__C _0553_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0773__B1 _0719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_130 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_200 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_87 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_391 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0611__C _0610_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0764__B1 _0763_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0819__A1 _0813_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_58 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1161__D _1224_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0819__B2 _0815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_130 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1210__CLK _1152_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0921_ _0880_/A _0875_/A _0920_/X d_sram_in[16] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_60_166 VGND VPWR sky130_fd_sc_hd__decap_12
X_0852_ _0851_/A _0852_/B _0852_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0783_ _0716_/B _0750_/A _0783_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_53_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0521__C _0721_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_119 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_141 VGND VPWR sky130_fd_sc_hd__fill_2
X_1197_ d_fabric_in[31] _1197_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_24_325 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_155 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0746__B1 _0651_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_200 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_222 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_31 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_75 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_166 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_188 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_41 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0903__A _0903_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_74 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_85 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0622__B _0488_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1156__D _1156_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1120_ d_sram_out[5] _0677_/D _1131_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_269 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_130 VGND VPWR sky130_fd_sc_hd__fill_2
X_1051_ _0966_/A _1043_/X _1049_/X w_mask[17] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_18_163 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_188 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0813__A _0661_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0904_ _1170_/Q _0890_/X _0903_/X _0904_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0976__B1 _0975_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0835_ _0845_/A _0883_/A _0831_/C _0838_/A VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__1106__CLK _1104_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0532__B _0717_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0766_ _0609_/X _0765_/X _0719_/X _0766_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0697_ _0697_/A _0694_/B _0530_/X _1122_/Q _0699_/C VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0900__B1 _0899_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_280 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_100 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_350 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0723__A _0721_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0967__B1 _0946_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_77 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_258 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0617__B _0743_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_40 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1129__CLK _1104_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0633__A _0594_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_158 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_84 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0958__B1 _0875_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_354 VGND VPWR sky130_fd_sc_hd__decap_12
X_0620_ _0620_/A _1147_/Q _0620_/C _0620_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_0551_ _0509_/X _0546_/Y _0550_/X _0551_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_1103_ _0634_/A _1103_/Q _1133_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0808__A _0665_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1034_ _1010_/A _1010_/B _0999_/X _1031_/D _1034_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0527__B _0489_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0543__A _0543_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8_0_clk_A clkbuf_3_4_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0818_ _0813_/X _1111_/Q _0532_/A _0815_/X d_fabric_out[28] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0749_ _0663_/X _1086_/D _0748_/X d_fabric_out[3] VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0718__A _0718_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_22 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_291 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_191 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_368 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_309 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_95 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0628__A _0566_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_291 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_173 VGND VPWR sky130_fd_sc_hd__decap_8
X_0603_ _0532_/A _0603_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0534_ _0616_/D _0535_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0538__A _0581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_280 VGND VPWR sky130_fd_sc_hd__fill_2
X_1017_ _0973_/A _0982_/B _1021_/C _1021_/D _1018_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_34_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0704__C _0699_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0720__B _0720_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_331 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_217 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0873__A2 _0839_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_283 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0625__A2 _0528_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_231 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_253 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1050__A2 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1164__D web VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_250 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1041__A2 _1040_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0540__B _0679_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0517_ _0585_/A _0587_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1074__D _1045_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_320 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_353 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_194 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0855__A2 _0839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_264 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_5_0_clk_A clkbuf_3_5_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0791__A1 _0714_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0791__B2 _1095_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_135 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_150 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_194 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_257 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0641__A _0697_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1159__D _1222_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1023__A2 _1022_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0782__A1 _0779_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0782__B2 _1092_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_304 VGND VPWR sky130_fd_sc_hd__fill_1
X_0997_ _0968_/X _1026_/B _0996_/X w_mask[6] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0701__D _1132_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0773__A1 _0771_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_323 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0726__A _0510_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_370 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_32 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1162__CLK _1184_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_87 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0764__A1 _0762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_74 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_62 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0819__A2 _1112_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0636__A _0676_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_348 VGND VPWR sky130_fd_sc_hd__decap_12
X_0920_ _1182_/Q _0876_/A _0920_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_60_178 VGND VPWR sky130_fd_sc_hd__decap_6
X_0851_ _0851_/A _0851_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0782_ _0779_/X _0781_/X _0762_/X _1092_/Q d_fabric_out[9] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_5_271 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0521__D _1127_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1196_ d_fabric_in[30] _1196_/Q _1196_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_24_304 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0546__A _0674_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_197 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1185__CLK _1191_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_381 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0746__A1 _0702_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_234 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_77 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_307 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_53 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0903__B _0903_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0622__C _0620_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_2_0_clk_A clkbuf_2_2_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0902__B1_N _0901_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1172__D d_fabric_in[6] VGND VPWR sky130_fd_sc_hd__diode_2
X_1050_ _0942_/A _1043_/X _1049_/X w_mask[16] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_33_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_167 VGND VPWR sky130_fd_sc_hd__fill_2
X_0903_ _0903_/A _0903_/B _0903_/C _1178_/Q _0903_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0976__A1 _0968_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0834_ _0845_/B _0883_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_0765_ _0614_/Y _0528_/X _0668_/X _0724_/D _0765_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_0696_ _0574_/A _0701_/B _0633_/B _0695_/X _0696_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA_clkbuf_4_4_0_clk_A clkbuf_4_5_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_215 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0900__A1 _0851_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_292 VGND VPWR sky130_fd_sc_hd__decap_12
X_1179_ d_fabric_in[13] _0908_/D _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_107 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_145 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_118 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0723__B _0721_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0967__A1 _0945_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_89 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1200__CLK _1131_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_204 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_270 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_112 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_97 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_156 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0914__A _0897_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0633__B _0633_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_300 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1080__B1 _1079_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0958__A1 _0883_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1167__D d_fabric_in[1] VGND VPWR sky130_fd_sc_hd__diode_2
X_0550_ _0549_/Y _0550_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_1102_ _1134_/Q _1102_/Q _1207_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1033_ _0944_/X _1032_/X _1029_/Y w_mask[13] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0824__A _1156_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1071__B1 _1066_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1223__CLK _1152_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0817_ _0813_/X _1110_/Q _0739_/D _0815_/X d_fabric_out[27] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0748_ _0732_/X _1086_/Q _0748_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0679_ _0722_/A _0679_/B _0679_/C _0757_/A _0679_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0718__B _0716_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_270 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_295 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_11 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1062__B1 _1061_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0628__B _0553_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0644__A _0616_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_284 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_295 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1053__B1 _1052_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0800__B1 _0799_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0602_ _0697_/A _0701_/B _0633_/B _0602_/D _0612_/B VGND VPWR sky130_fd_sc_hd__and4_4
X_0533_ _0584_/A _0616_/D VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_3_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0867__B1 _0866_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_229 VGND VPWR sky130_fd_sc_hd__fill_2
X_1016_ _0998_/X _1015_/X _1012_/X w_mask[9] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0554__A _1126_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_284 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0704__D _0704_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0729__A _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_clk_A clkbuf_3_1_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1119__CLK _1131_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_343 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_88 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_210 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_276 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_12_0_clk_A clkbuf_3_6_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_129 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0639__A _0723_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_310 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0849__B1 _0848_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_376 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1180__D d_fabric_in[14] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_357 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_221 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_276 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0540__C _0682_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0516_ _1152_/Q _0585_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0549__A _0548_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_365 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1090__D _1090_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_287 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0791__A2 _1095_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_65 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1091__CLK _1145_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_335 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_236 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0922__A _0828_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0641__B _0694_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1175__D d_fabric_in[9] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0782__A2 _0781_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_313 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_173 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_327 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0832__A _0832_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0996_ _0985_/X _0979_/X _0988_/Y _0996_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0773__A2 _0772_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1085__D _1085_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_154 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0726__B _0726_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_165 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_45 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_213 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0742__A _0725_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_239 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_22 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0764__A2 _1088_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_38 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_313 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_302 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0636__B _0686_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_113 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0652__A _0681_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0850_ _0830_/Y _0833_/X _0849_/X d_sram_in[2] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0781_ _0674_/A _0496_/X _0676_/D _0496_/X _0781_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_5_261 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_283 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_121 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_132 VGND VPWR sky130_fd_sc_hd__decap_3
X_1195_ d_fabric_in[29] _1195_/Q _1184_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0827__A _0827_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0546__B _0521_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_179 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0562__A _0561_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_393 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_0_0_clk_A clkbuf_3_0_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0979_ _0978_/X _0979_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0746__A2 _0548_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_23 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_143 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0737__A _1126_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_102 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_198 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_146 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_371 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0903__C _0903_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0647__A _0647_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_179 VGND VPWR sky130_fd_sc_hd__fill_2
X_0902_ _1177_/Q _0877_/X _0901_/Y d_sram_in[11] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0976__A2 _0974_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0833_ _0875_/A _0833_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0764_ _0762_/X _1088_/D _0763_/X d_fabric_out[5] VGND VPWR sky130_fd_sc_hd__a21o_4
X_0695_ _1134_/Q _0695_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0900__A2 _0890_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1152__CLK _1152_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0557__A _0556_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_81 VGND VPWR sky130_fd_sc_hd__decap_8
X_1178_ d_fabric_in[12] _1178_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_157 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_108 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_190 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0723__C _0723_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0967__A2 _0966_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_32 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_282 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_116 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0914__B _0913_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1080__A1 _1035_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0958__A2 _0845_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1183__D d_fabric_in[17] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1175__CLK _1188_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1101_ _0594_/A _1101_/Q _1207_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0894__A1 _0891_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1032_ _1031_/X _1032_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_46_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1001__A _1000_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1071__A1 _0984_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0816_ _0813_/X _1109_/Q _0717_/A _0815_/X d_fabric_out[26] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__0840__A _0825_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0747_ _0750_/A _0736_/X _0746_/X _0695_/X _0495_/X _1086_/D VGND VPWR sky130_fd_sc_hd__a32o_4
X_0678_ _1112_/D _0757_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1093__D _0784_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_238 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_249 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0718__C _0501_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_68 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_127 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_149 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1062__A1 _1026_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_89 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0750__A _0750_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1198__CLK _1133_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0573__B1 _0721_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_86 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_271 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0644__B _0644_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_403 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1053__A1 _0974_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_160 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1178__D d_fabric_in[12] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0800__A1 _0714_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0800__B2 _1098_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0601_ _0582_/X _0633_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0532_ _0532_/A _0717_/B _0532_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_21_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0867__A1 _0864_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_260 VGND VPWR sky130_fd_sc_hd__fill_2
X_1015_ _1015_/A _1015_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0835__A _0845_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_263 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1088__D _1088_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_80 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0570__A _0523_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_329 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0729__B _0729_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_34 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_45 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_355 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0745__A _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_22 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0794__B1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_178 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0639__B _0604_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0849__A1 _0830_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1213__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_241 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0655__A _0655_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_263 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_296 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_233 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_255 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0540__D _0540_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0537__B1 _0676_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0515_ _0679_/B _0721_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_66_174 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_314 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0565__A _0584_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_244 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_108 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_347 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_358 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_21 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_204 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_226 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0922__B _0876_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0641__C _0633_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0767__B1 _0709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1191__D d_fabric_in[25] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_130 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_111 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1109__CLK _1096_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0995_ _0995_/A _1026_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0758__B1 _0687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_358 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0726__C _1113_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_328 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0997__B1 _0996_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0742__B _0491_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0749__B1 _0748_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_78 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_43 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0921__B1 _0920_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_358 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0636__C _0635_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_177 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_380 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_350 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_147 VGND VPWR sky130_fd_sc_hd__fill_1
X_0780_ _0779_/X _0778_/X _0762_/X _1091_/Q d_fabric_out[8] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1186__D d_fabric_in[20] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_295 VGND VPWR sky130_fd_sc_hd__decap_8
X_1194_ d_fabric_in[28] _1194_/Q _1184_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1004__A _1031_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0546__C _0537_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0843__A _0843_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_361 VGND VPWR sky130_fd_sc_hd__decap_8
X_0978_ _0973_/A _0952_/B _1021_/C _0982_/D _0978_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__1096__D _0793_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_35 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_280 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0737__B _0720_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_306 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_45 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_361 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_383 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_191 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0903__D _1178_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_217 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_239 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_122 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_111 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0647__B _0647_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_291 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_147 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0663__A _0663_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_361 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_180 VGND VPWR sky130_fd_sc_hd__decap_3
X_0901_ _0854_/A _0901_/B _0901_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_0832_ _0832_/A _0875_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0763_ _0732_/X _0763_/B _0763_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0694_ _0535_/A _0694_/B _0582_/X _1126_/Q _0694_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_51_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0838__A _0838_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_206 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_93 VGND VPWR sky130_fd_sc_hd__decap_4
X_1177_ d_fabric_in[11] _1177_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_24_125 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_109 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_320 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0723__D _0723_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_228 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0748__A _0732_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_66 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_32 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_139 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1080__A2 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_379 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_9_0_clk clkbuf_3_4_0_clk/X _1155_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1100_ _1132_/Q _1100_/Q _1196_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0894__A2 _0877_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1031_ _1007_/A _1021_/B _0999_/X _1031_/D _1031_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_46_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_128 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1071__A2 _1032_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0815_ out_reg _0815_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0746_ _0702_/D _0548_/X _0651_/Y _0745_/X _0746_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_0677_ _0668_/A _0669_/X _0721_/C _0677_/D _0684_/C VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0718__D _0717_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_24 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_46 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1062__A2 _1059_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0573__B2 _0586_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0573__A1 _0540_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_283 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0644__C _0582_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_264 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0941__A _0941_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_132 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1053__A2 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_165 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0800__A2 _1098_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0600_ _0606_/A _0697_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1142__CLK _1096_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0531_ _0530_/X _0717_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1194__D d_fabric_in[28] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0867__A2 _0839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_356 VGND VPWR sky130_fd_sc_hd__decap_12
X_1014_ _0982_/A _1021_/B _1021_/C _1021_/D _1015_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_34_220 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0835__B _0883_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0851__A _0851_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0570__B _1150_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0729_ _0550_/X _0729_/B _0729_/C _0729_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_57_301 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0729__C _0729_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_57 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0745__B _0737_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_223 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_89 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1165__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_289 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0794__A1 _0714_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0794__B2 _1096_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_124 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0849__A2 _0839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_323 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_345 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0655__B _0655_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_245 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1189__D d_fabric_in[23] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0537__A1 _0526_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0514_ _0726_/B _0679_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_39_301 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1007__A _1007_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_367 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0915__B1_N _0914_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0846__A _0846_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1188__CLK _1188_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1099__D _0655_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0581__A _0581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_175 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_197 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_212 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_289 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_278 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0491__A _0491_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0641__D _1117_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0767__A1 _0721_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_182 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_120 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_337 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_189 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_370 VGND VPWR sky130_fd_sc_hd__decap_6
X_0994_ _1010_/A _1010_/B _0999_/A _0972_/A _0995_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_8_260 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0758__A1 _0668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0930__A1 _1189_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_142 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0576__A _0587_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_315 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_134 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_145 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0726__D _0726_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0997__A1 _0968_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0742__C _0726_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0749__A1 _0663_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1203__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_11 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_55 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0921__A1 _0880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_66 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0486__A reb VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0685__B1 _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_87 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_156 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_392 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_230 VGND VPWR sky130_fd_sc_hd__decap_12
X_1193_ d_fabric_in[27] _1193_/Q _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0546__D _0546_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_329 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_159 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1226__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0977_ _1209_/Q _1021_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_10_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_395 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_89 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_229 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_134 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0647__C _0647_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_145 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0658__B1 _0651_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0944__A _0943_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__decap_3
X_0900_ _0851_/A _0890_/X _0899_/X _0901_/B VGND VPWR sky130_fd_sc_hd__a21o_4
X_0831_ _1226_/Q _1156_/D _0831_/C _0832_/A VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__1197__D d_fabric_in[31] VGND VPWR sky130_fd_sc_hd__diode_2
X_0762_ _0663_/A _0762_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0693_ _0676_/D _0627_/Y _0692_/X _0704_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_44_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0838__B _0838_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1015__A _1015_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_251 VGND VPWR sky130_fd_sc_hd__decap_12
X_1176_ d_fabric_in[10] _0895_/D _1188_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0649__B1 _0648_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_115 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0854__A _0854_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_332 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_354 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0821__B1 _1146_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_15 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0748__B _1086_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_148 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_354 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0812__B1 _0656_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_218 VGND VPWR sky130_fd_sc_hd__fill_2
X_1030_ _0944_/X _1025_/X _1029_/Y w_mask[12] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0674__A _0674_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_170 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0803__B1 _0487_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0814_ _0813_/X _1108_/Q _0676_/D _0808_/X d_fabric_out[25] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0745_ _0550_/X _0737_/X _0744_/X _0745_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_0676_ _0676_/A _0492_/C _0676_/C _0676_/D _0676_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0781__A2_N _0496_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1228_ conf[2] _0825_/A _1184_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0584__A _0584_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_295 VGND VPWR sky130_fd_sc_hd__decap_3
X_1159_ _1222_/Q _1159_/Q _1191_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1047__B1 _0958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_298 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_140 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_36 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0573__A2 _0608_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1094__CLK _1096_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0730__C1 _0729_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_99 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0494__A _0493_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_221 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1038__B1 _1037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0644__D _0716_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_100 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_195 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_155 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_188 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_91 VGND VPWR sky130_fd_sc_hd__fill_1
X_0530_ _0529_/Y _0530_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0669__A _0721_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_368 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_284 VGND VPWR sky130_fd_sc_hd__fill_2
X_1013_ _0998_/X _1006_/X _1012_/X w_mask[8] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_34_243 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0835__C _0831_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_93 VGND VPWR sky130_fd_sc_hd__decap_3
X_0728_ _0728_/A _0728_/B _0723_/X _0727_/X _0729_/C VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0579__A _0616_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0659_ _0497_/X _0659_/B _0659_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_57_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_221 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0745__C _0744_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_287 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_213 VGND VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_8_0_clk clkbuf_3_4_0_clk/X _1145_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_43_57 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0794__A2 _0793_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_136 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0489__A _1150_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_331 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_276 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0952__A _1045_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0537__A2 _0532_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0513_ _0616_/B _0726_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_66_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0846__B _0852_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_257 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_268 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_279 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0581__B _1150_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_143 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1132__CLK _1130_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_308 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_239 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_290 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0767__A2 _0497_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_110 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0947__A _0940_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_305 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_382 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0682__A _0722_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0993_ _0968_/X _0992_/X _0989_/X w_mask[5] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_8_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0758__A2 _1128_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1018__A _1018_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0930__A2 _0926_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1155__CLK _1155_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0857__A _1170_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0576__B _0584_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_338 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0592__A _0579_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_37 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_341 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0997__A2 _1026_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_374 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0742__D _0695_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0749__A2 _1086_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0921__A2 _0875_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_78 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_11 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0486__B csb VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0685__A1 _0674_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_113 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_135 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_105 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_396 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_220 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_80 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0929__B1_N _0870_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1178__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0677__A _0668_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1192_ d_fabric_in[26] _1192_/Q _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_36_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_308 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_341 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_190 VGND VPWR sky130_fd_sc_hd__decap_4
X_0976_ _0968_/X _0974_/X _0975_/Y w_mask[2] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0587__A _0587_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0497__A _0497_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0647__D _0646_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0658__A1 _0501_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_157 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0658__B2 _0657_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_127 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_80 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0960__A _0988_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0830_ _0846_/A _0830_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0761_ _0675_/D _0750_/X _0759_/X _0760_/X _1088_/D VGND VPWR sky130_fd_sc_hd__o22a_4
X_0692_ _0739_/D _0558_/X _0692_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_37_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_51 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_clk clkbuf_0_clk/X clkbuf_2_2_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0649__A1 _0626_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_282 VGND VPWR sky130_fd_sc_hd__fill_2
X_1175_ d_fabric_in[9] _0891_/D _1188_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_263 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1031__A _1007_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0821__B2 _0779_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0821__A1 _0663_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0959_ _1065_/B _0838_/B _0958_/X _0959_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_47_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_241 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_116 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_274 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0812__B2 _0808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0812__A1 _0806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_71 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_208 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1216__CLK _1104_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0955__A _1045_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0674__B _0674_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0690__A _0679_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0803__B2 _0801_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0803__A1 _0799_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0813_ _0661_/Y _0813_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0744_ _0738_/X _0739_/X _0740_/X _0744_/D _0744_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_0675_ _0721_/A _0669_/X _0676_/C _0675_/D _0684_/A VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1026__A _0984_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1227_ conf[1] _1156_/D _1133_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0584__B _0584_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_274 VGND VPWR sky130_fd_sc_hd__fill_2
X_1158_ _1158_/D _1150_/D _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_16_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_1089_ _1089_/D _1089_/Q _1155_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1047__A1 _1046_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_307 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_196 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0730__B1 _0719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1038__A1 _0944_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_152 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_112 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_70 VGND VPWR sky130_fd_sc_hd__fill_2
X_1012_ _0985_/X _0983_/X _1011_/Y _1012_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0788__B1 _0739_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0727_ _0508_/A _0724_/X _0725_/X _0726_/X _0727_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0579__B _0530_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0658_ _0501_/X _0551_/Y _0650_/X _0651_/Y _0657_/X _0659_/B VGND VPWR sky130_fd_sc_hd__a32oi_4
X_0589_ _0579_/X _0589_/B _0589_/C _0589_/D _0589_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XANTENNA__0595__A _1132_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0712__B1 _0487_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_37 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_47 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_148 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_288 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0952__B _0952_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_225 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0795__A2_N _0787_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0512_ _0722_/A _0676_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_54_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_28 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_291 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1084__CLK _1155_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_111 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_306 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_391 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_339 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_188 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_350 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_24 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_236 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_328 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0963__A _0950_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0682__B _0679_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_394 VGND VPWR sky130_fd_sc_hd__decap_3
X_0992_ _0992_/A _0992_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_67_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_62 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_7_0_clk clkbuf_4_6_0_clk/A _1152_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__1034__A _1010_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0576__C _0725_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_155 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_125 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_320 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_206 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_353 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_23 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_306 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_328 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0685__A2 _0684_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0783__A _0716_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0677__B _0669_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1191_ d_fabric_in[25] _1191_/Q _1191_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0765__A1_N _0614_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_90 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_331 VGND VPWR sky130_fd_sc_hd__decap_4
X_0975_ _0859_/B _0966_/Y _0960_/X _0975_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__1122__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1029__A _0959_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0587__B _1153_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_37 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_331 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_353 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_183 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0658__A2 _0551_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_117 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_70 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_172 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0960__B _0955_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0760_ _0677_/D _0495_/X _0709_/X _0760_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1145__CLK _1145_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0691_ _0691_/A _0739_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0688__A _0688_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_63 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0649__A2 _0632_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_294 VGND VPWR sky130_fd_sc_hd__decap_4
X_1174_ d_fabric_in[8] _1174_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1031__B _1021_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_161 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0821__A2 _1114_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0958_ _0883_/A _0845_/C _0875_/A _0958_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0889_ _1174_/Q _0877_/X _0888_/Y d_sram_in[8] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0598__A _0579_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_264 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0928__B1_N _0867_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1168__CLK _1133_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0812__A2 _1107_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0955__B _0952_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_161 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_150 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0971__A _1209_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0690__B _0689_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0803__A2 _1100_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0812_ _0806_/X _1107_/Q _0656_/A _0808_/X d_fabric_out[24] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0743_ _0743_/A _0674_/B _0743_/C _0742_/X _0744_/D VGND VPWR sky130_fd_sc_hd__or4_4
X_0674_ _0674_/A _0674_/B _0674_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1026__B _1026_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1226_ conf[0] _1226_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_253 VGND VPWR sky130_fd_sc_hd__fill_2
X_1157_ _0825_/A _1149_/D _1196_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_201 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0584__C _0582_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1042__A _0899_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1088_ _1088_/D _0763_/B _1155_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_267 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1047__A2 _0838_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0881__A _0845_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_16 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_319 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0730__A1 _1117_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1038__A2 _1035_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1102__D _1134_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0_clk clkbuf_0_clk/X clkbuf_1_0_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_11_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_93 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_363 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0966__A _0966_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_264 VGND VPWR sky130_fd_sc_hd__decap_4
X_1011_ _1009_/X _1011_/B _0959_/Y _1011_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_19_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_289 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0788__B2 _0787_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0726_ _0510_/X _0726_/B _1113_/D _0726_/D _0726_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0579__C _0579_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0657_ _0668_/A _0502_/A _0655_/X _0656_/X _0657_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_0588_ _0584_/X _0585_/X _0586_/X _0587_/X _0589_/D VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0712__A1 _0750_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0876__A _0876_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_315 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0595__B _0582_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0712__B2 _0711_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1209_ addr_w[11] _1209_/Q _1196_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_212 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1206__CLK _1188_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_311 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_337 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_267 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0952__C _0878_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_237 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_259 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_92 VGND VPWR sky130_fd_sc_hd__fill_2
X_0511_ _0510_/X _0722_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_3_171 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0696__A _0574_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_3 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_318 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_373 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0933__A1 _1191_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_119 VGND VPWR sky130_fd_sc_hd__decap_3
X_0709_ _0501_/X _0709_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_329 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_226 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_403 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0621__B1 _0620_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0924__A1 _1184_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_145 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0682__C _0682_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0991_ _0982_/A _0952_/B _0982_/C _0982_/D _0992_/A VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0860__B1 _0880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0915__A1 _0912_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_74 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_123 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0576__D _0616_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1034__B _1010_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_137 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_373 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_229 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1200__D addr_w[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_49 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0906__A1 _1178_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_35 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_126 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0783__B _0750_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_118 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_354 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1110__D _0691_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0677__C _0721_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1190_ d_fabric_in[24] _1190_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0974__A _0973_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_321 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_398 VGND VPWR sky130_fd_sc_hd__decap_6
X_0974_ _0973_/X _0974_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1029__B _1026_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0587__C _0586_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1045__A _1045_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0884__A _0903_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_49 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1077__B1 _1076_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_15 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1097__CLK _1207_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_258 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_115 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_126 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1105__D _0723_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0658__A3 _0650_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_295 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1068__B1 _1067_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_71 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_60 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_184 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_93 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0960__C _0959_/Y VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_6_0_clk clkbuf_4_6_0_clk/A _1207_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0690_ _0679_/C _0689_/B _0654_/A _0757_/A _0690_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0969__A _0969_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0688__B _0687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_75 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_97 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0649__A3 _0636_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1173_ d_fabric_in[7] _1173_/Q _1191_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1031__C _0999_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_346 VGND VPWR sky130_fd_sc_hd__fill_2
X_0957_ _1010_/B _1065_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_9_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_0888_ _0880_/X _0888_/B _0905_/A _0888_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0879__A _0878_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_26 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_140 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_162 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_184 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_51 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_62 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0955__C _0982_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_265 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_287 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_140 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1112__CLK _1108_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_257 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0690__C _0654_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0811_ _0806_/X _1106_/Q _1138_/Q _0808_/X d_fabric_out[23] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0742_ _0725_/A _0491_/A _0726_/D _0695_/X _0742_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_6_361 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0699__A _0694_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0673_ _0673_/A _0674_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_42_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1225_ addr_r[13] _1225_/Q _1184_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1156_ _1156_/D _1156_/Q _1155_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0584__D _0677_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1042__B _0899_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_213 VGND VPWR sky130_fd_sc_hd__fill_1
X_1087_ _1087_/D _1087_/Q _1155_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0730__A2 _0548_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1135__CLK _1133_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_265 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_287 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_136 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_61 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_83 VGND VPWR sky130_fd_sc_hd__fill_2
X_1010_ _1010_/A _1010_/B _0878_/Y _1011_/B VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__0982__A _0982_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_224 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_268 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_279 VGND VPWR sky130_fd_sc_hd__decap_3
X_0725_ _0725_/A _0491_/A _0726_/D _0594_/A _0725_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_6_191 VGND VPWR sky130_fd_sc_hd__fill_2
X_0656_ _0656_/A _0717_/B _0656_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0579__D _1130_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0587_ _0587_/A _1153_/Q _0586_/C _0716_/B _0587_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0927__B1_N _0862_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1158__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0712__A2 _0672_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1208_ addr_w[10] _0940_/A _1207_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1203__D addr_w[5] VGND VPWR sky130_fd_sc_hd__diode_2
X_1139_ d_sram_out[24] _0543_/A _1133_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_235 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_323 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_246 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1113__D _1113_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_249 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0510_ _1151_/Q _0510_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0977__A _1209_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0696__B _0701_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_316 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_308 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_360 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_205 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_282 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1048__A _1048_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0933__A2 _0932_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0708_ _0705_/X _0706_/Y _0707_/X _0708_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_0639_ _0723_/D _0604_/Y _0647_/B VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0887__A _0899_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_135 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_146 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_179 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_15 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_396 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0621__A1 _0591_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0924__A2 _0907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1108__D _0602_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0797__A _1146_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_135 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_127 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_60 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0682__D _1128_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0990_ _0968_/X _0983_/X _0989_/X w_mask[4] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_44_81 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0860__A1 _0828_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_91 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0915__A2 _0907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0500__A _0499_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_146 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1034__C _0999_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_396 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0906__A2 _0877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_341 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_333 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_40 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_73 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_267 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1219__CLK _1108_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0677__D _0677_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_396 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_300 VGND VPWR sky130_fd_sc_hd__fill_2
X_0973_ _0973_/A _0982_/B _1045_/C _0982_/D _0973_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__1029__C _1029_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0587__D _0716_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1045__B _1046_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_116 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_403 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1077__A1 _1025_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1211__D addr_w[13] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0760__B1 _0709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_322 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_311 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_160 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1068__A1 _1006_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_50 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1121__D d_sram_out[6] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_72 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_141 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_83 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_152 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_94 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_196 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_7 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0751__B1 _0634_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0985__A _0984_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_241 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1191__CLK _1191_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1172_ d_fabric_in[6] _1172_/Q _1130_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_66_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0649__A4 _0647_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_171 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_193 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1031__D _1031_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_130 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_303 VGND VPWR sky130_fd_sc_hd__decap_3
X_0956_ _1207_/Q _1010_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_20_358 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_19 VGND VPWR sky130_fd_sc_hd__fill_2
X_0887_ _0899_/A _0899_/B _0903_/C _1174_/Q _0888_/B VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0990__B1 _0989_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1056__A _1048_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1206__D addr_w[8] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0895__A _0899_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_222 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_255 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1116__D d_sram_out[1] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0955__D _0859_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_60 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_203 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0690__D _0757_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0810_ _0806_/X _1105_/Q _0723_/D _0808_/X d_fabric_out[22] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0741_ _0510_/X _0726_/B _0741_/C _1130_/Q _0743_/C VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_6_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0699__B _0696_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0672_ _0668_/X _0673_/A _0501_/X _0671_/X _0672_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_35_3 VGND VPWR sky130_fd_sc_hd__decap_4
X_1224_ addr_r[12] _1224_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_266 VGND VPWR sky130_fd_sc_hd__fill_2
X_1155_ _1226_/Q _1155_/Q _1155_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1042__C _0831_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1086_ _1086_/D _1086_/Q _1155_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_247 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_100 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1087__CLK _1155_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0939_ _1197_/Q _0876_/X _0918_/Y d_sram_in[31] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0715__B1 _0714_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_15 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_5_0_clk clkbuf_4_5_0_clk/A _1188_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_57_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_225 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_236 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_104 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_40 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_343 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0706__B1 _0622_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_200 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0982__B _0982_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_247 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_280 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0503__A _1150_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0724_ _0510_/X _0726_/B _0741_/C _0724_/D _0724_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0655_ _0655_/A _0655_/B _0655_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0586_ _0585_/A _0584_/B _0586_/C _1117_/Q _0586_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0712__A3 _0710_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1207_ addr_w[9] _1207_/Q _1207_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1138_ d_sram_out[23] _1138_/Q _1130_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1069_ _1015_/X _1059_/X _1067_/X w_mask[25] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_40_206 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0778__A1_N _0509_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_302 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1102__CLK _1207_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_335 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_368 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_225 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_50 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0696__C _0633_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_306 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_158 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0577__A2_N _0576_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1125__CLK _1131_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1048__B _1048_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0707_ _1116_/Q _0622_/Y _0550_/X _0707_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_0638_ _0717_/A _0558_/X _0647_/A VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0887__B _0899_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0569_ _1153_/Q _0579_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1064__A _1046_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_158 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1214__D addr_r[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_350 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_250 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_283 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0621__A2 _0619_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0909__B1 _0908_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0797__B _0497_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_114 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1124__D d_sram_out[9] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_139 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0911__B1_N _0910_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_342 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0860__A2 _0859_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1148__CLK _1155_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_276 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0988__A _0988_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1034__D _1031_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_117 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_320 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_19 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_209 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1059__A _1042_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1209__D addr_w[11] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_309 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_367 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1119__D d_sram_out[4] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0601__A _0582_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_84 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_401 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_71 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_161 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_345 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_194 VGND VPWR sky130_fd_sc_hd__fill_1
X_0972_ _0972_/A _0982_/D VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_65_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0511__A _0510_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_242 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1045__C _1045_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_106 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_323 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1077__A2 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_142 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0760__A1 _0677_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_109 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_40 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_150 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1068__A2 _1059_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_334 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_51 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_183 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_62 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_389 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_84 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0751__A1 _0668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_7 VGND VPWR sky130_fd_sc_hd__decap_3
X_1171_ d_fabric_in[5] _1171_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0506__A _0505_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_186 VGND VPWR sky130_fd_sc_hd__fill_2
X_0955_ _1045_/A _0952_/B _0982_/C _0859_/A _0955_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0886_ _0908_/C _0903_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0990__A1 _0968_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1056__B _1055_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0895__B _0899_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_245 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_278 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1222__D addr_r[10] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1209__CLK _1196_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_223 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1132__D d_sram_out[17] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_186 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_175 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_93 VGND VPWR sky130_fd_sc_hd__decap_6
X_0740_ _0721_/A _0721_/B _0723_/C _1138_/Q _0740_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_6_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0699__C _0699_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0671_ _0676_/A _0669_/X _0676_/D _0487_/X _0655_/B _0671_/X VGND VPWR sky130_fd_sc_hd__a32o_4
X_1223_ addr_r[11] _1223_/Q _1152_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_28_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_245 VGND VPWR sky130_fd_sc_hd__decap_8
X_1154_ _1162_/Q _1154_/Q _1184_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_278 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1042__D _1042_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_215 VGND VPWR sky130_fd_sc_hd__decap_4
X_1085_ _1085_/D _1085_/Q _1130_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_20_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_178 VGND VPWR sky130_fd_sc_hd__fill_2
X_0938_ _1196_/Q _0876_/X _0914_/Y d_sram_in[30] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0869_ _1172_/Q _0869_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1217__D addr_r[5] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0715__A1 _0663_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_223 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_245 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_112 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_156 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1181__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1127__D d_sram_out[12] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_355 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0706__A1 _0674_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_307 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_215 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0982__C _0982_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_92 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_98 VGND VPWR sky130_fd_sc_hd__fill_2
X_0723_ _0721_/A _0721_/B _0723_/C _0723_/D _0723_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0654_ _0654_/A _0655_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0585_ _0585_/A _0584_/B _0582_/A _1116_/Q _0585_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA_clkbuf_4_7_0_clk_A clkbuf_4_6_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1206_ addr_w[8] baseaddr_w_sync[8] _1188_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_351 VGND VPWR sky130_fd_sc_hd__decap_12
X_1137_ d_sram_out[22] _0723_/D _1108_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_248 VGND VPWR sky130_fd_sc_hd__decap_3
X_1068_ _1006_/X _1059_/X _1067_/X w_mask[24] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0936__A1 _1194_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_215 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_373 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_229 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0604__A _0604_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0927__A1 _1186_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0696__D _0695_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_340 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0863__B1 _0862_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_218 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_229 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0615__B1 _1112_/D VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_4_0_clk clkbuf_4_5_0_clk/A _1133_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0514__A _0726_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1048__C _1048_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0706_ _0674_/A _0703_/A _0622_/Y _0706_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_0637_ _1141_/Q _0717_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0887__C _0903_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0568_ _0560_/Y _0562_/X _0567_/Y _0578_/B VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__1064__B _1046_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0499_ _0620_/A _1147_/Q _0620_/C _0499_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_38_362 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_262 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_295 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0909__A1 _1171_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_340 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1140__D d_sram_out[25] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_251 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0988__B _0988_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_159 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0509__A _0509_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_140 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_195 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1013__B1 _1012_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1075__A _1066_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1225__D addr_r[13] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_49 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_4_0_clk_A clkbuf_3_5_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_313 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_64 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_63 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_15_0_clk_A clkbuf_3_7_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1135__D d_sram_out[20] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_343 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0818__B1 _0532_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1115__CLK _1145_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_335 VGND VPWR sky130_fd_sc_hd__fill_1
X_0971_ _1209_/Q _1045_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0999__A _0999_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1045__D _1045_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0809__B1 _0675_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_357 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_121 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_18 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_187 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0702__A _0741_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_206 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0760__A2 _0495_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1138__CLK _1130_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0925__B1_N _0855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_221 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_265 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_276 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_287 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_30 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_176 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0612__A _0612_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0736__C1 _0735_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0751__A2 _1127_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_254 VGND VPWR sky130_fd_sc_hd__fill_2
X_1170_ d_fabric_in[4] _1170_/Q _1191_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_66_70 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_298 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_198 VGND VPWR sky130_fd_sc_hd__decap_4
X_0954_ _0999_/A _0982_/C VGND VPWR sky130_fd_sc_hd__buf_1
X_0885_ _0845_/C _0908_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0522__A _1151_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0990__A2 _0983_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1056__C _1048_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0895__C _0903_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_73 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_1_0_clk_A clkbuf_1_0_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0607__A _1138_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_132 VGND VPWR sky130_fd_sc_hd__fill_1
X_0670_ _0602_/D _0676_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0699__D _0698_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1222_ addr_r[10] _1222_/Q _1191_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1153_ _1161_/Q _1153_/Q _1130_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1084_ _1084_/D _1084_/Q _1155_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_205 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0517__A _0585_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_290 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_157 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0660__A1 _0487_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0937_ _1195_/Q _0932_/X _0910_/Y d_sram_in[29] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA_clkbuf_4_3_0_clk_A clkbuf_4_2_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0868_ _0864_/Y _0833_/X _0867_/X d_sram_in[5] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0799_ _0661_/Y _0799_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0715__A2 _1084_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_279 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_205 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_293 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0706__A2 _0703_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1143__D d_sram_out[28] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_72 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_268 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0982__D _0982_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_88 VGND VPWR sky130_fd_sc_hd__fill_2
X_0722_ _0722_/A _0492_/C _0723_/C _0717_/A _0728_/B VGND VPWR sky130_fd_sc_hd__and4_4
X_0653_ _0721_/A _0668_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0584_ _0584_/A _0584_/B _0582_/A _0677_/D _0584_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_57_319 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_330 VGND VPWR sky130_fd_sc_hd__fill_2
X_1205_ addr_w[7] baseaddr_w_sync[7] _1145_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_363 VGND VPWR sky130_fd_sc_hd__decap_3
X_1136_ d_sram_out[21] _0675_/D _1104_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_396 VGND VPWR sky130_fd_sc_hd__decap_8
X_1067_ _1044_/X _1025_/X _1066_/Y _1067_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_40_219 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0936__A2 _0932_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1228__D conf[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_75 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_271 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_293 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1138__D d_sram_out[23] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0927__A2 _0926_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0620__A _0620_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_352 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_396 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0863__A1 _0857_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_377 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0615__B2 _0558_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_252 VGND VPWR sky130_fd_sc_hd__fill_2
X_0705_ _0617_/X _0686_/X _0689_/X _0705_/D _0705_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0530__A _0529_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0636_ _0676_/C _0686_/C _0635_/Y _0636_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0887__D _1174_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0567_ _0606_/A _0566_/X _0529_/Y _0702_/D _0567_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__1064__C _1045_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0551__B1 _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0498_ _0498_/A _0620_/C VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1171__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_171 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_374 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_300 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_322 VGND VPWR sky130_fd_sc_hd__fill_2
X_1119_ d_sram_out[4] _0540_/D _1131_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_13_208 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0705__A _0617_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_clk_A clkbuf_3_1_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0909__A2 _0890_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0790__B1 _0532_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_119 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_352 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_322 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_333 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_355 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_366 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_73 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_11_0_clk_A clkbuf_3_5_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_263 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_223 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_83 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0988__C _0959_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0781__B1 _0676_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1194__CLK _1184_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0509__B _0674_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_185 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0525__A _0655_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1013__A1 _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0772__B1 _0668_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0619_ _0597_/X _0612_/Y _0618_/Y _0619_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__1075__B _1075_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_42 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_3_0_clk clkbuf_4_2_0_clk/A _1108_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_39_95 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0818__A1 _0813_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0818__B2 _0815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_193 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1151__D _1159_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_152 VGND VPWR sky130_fd_sc_hd__fill_1
X_0970_ _1207_/Q _0982_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_40_391 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0754__B1 _0752_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_211 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0809__A1 _0806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0809__B2 _0808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0993__B1 _0989_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0702__B _0686_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_255 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_31 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_314 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_42 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_31 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_53 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_53 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_369 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_75 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_75 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_52 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0612__B _0612_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0736__B1 _0501_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1146__D d_sram_out[31] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_222 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_82 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_133 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0672__C1 _0671_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_328 VGND VPWR sky130_fd_sc_hd__fill_2
X_0953_ _1209_/Q _0999_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0975__B1 _0960_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0884_ _0903_/B _0899_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0895__D _0895_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_214 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_225 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_166 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_177 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0713__A out_reg VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1105__CLK _1104_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_99 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0607__B _0529_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_239 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_144 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_7 VGND VPWR sky130_fd_sc_hd__decap_12
X_1221_ addr_r[9] _1158_/D _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_203 VGND VPWR sky130_fd_sc_hd__fill_2
X_1152_ _1160_/Q _1152_/Q _1152_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1083_ _0660_/X _1083_/Q _1145_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_239 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_250 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0660__A2 _0496_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1128__CLK _1130_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0533__A _0584_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0924__B1_N _0849_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0936_ _1194_/Q _0932_/X _0905_/Y d_sram_in[28] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0867_ _0864_/Y _0839_/X _0866_/Y _0867_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0798_ _1130_/Q _0750_/X _0797_/X _1098_/D VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0939__B1_N _0918_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_217 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_272 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_32 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_87 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_62 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0618__A _0552_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_261 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_56 VGND VPWR sky130_fd_sc_hd__decap_12
X_0721_ _0721_/A _0721_/B _0721_/C _0721_/D _0728_/A VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_6_195 VGND VPWR sky130_fd_sc_hd__fill_2
X_0652_ _0681_/A _0721_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0583_ _0606_/A _0579_/C _0582_/X _0673_/A _0589_/C VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_33_3 VGND VPWR sky130_fd_sc_hd__decap_4
X_1204_ addr_w[6] baseaddr_w_sync[6] _1133_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1135_ d_sram_out[20] _0634_/A _1133_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0528__A _0527_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_217 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_239 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_291 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_280 VGND VPWR sky130_fd_sc_hd__fill_2
X_1066_ _1066_/A _1066_/B _1048_/C _1066_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_33_294 VGND VPWR sky130_fd_sc_hd__fill_2
X_0919_ _1181_/Q _0907_/X _0918_/Y d_sram_in[15] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_16_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_54 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_75 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0901__A _0854_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0620__B _1147_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1154__D _1162_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0863__A2 _0833_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_209 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_389 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_264 VGND VPWR sky130_fd_sc_hd__fill_2
X_0704_ _0690_/X _0704_/B _0699_/X _0704_/D _0705_/D VGND VPWR sky130_fd_sc_hd__or4_4
X_0635_ _0526_/X _0635_/B _0634_/X _0635_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_0566_ _0644_/B _0566_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1064__D _0859_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0551__A1 _0509_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0497_ _0497_/A _0497_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_331 VGND VPWR sky130_fd_sc_hd__fill_2
X_1118_ d_sram_out[3] _0702_/D _1152_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1049_ _1044_/X _1006_/X _1048_/Y _1049_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_53_367 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0705__B _0686_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0721__A _0721_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0790__B2 _0787_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_301 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_150 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_378 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_85 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_213 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1149__D _1149_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0631__A _0535_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0781__B2 _0496_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_172 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_345 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0806__A _0661_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0525__B _0608_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0541__A _0535_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1013__A2 _1006_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0772__A1 _0676_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0772__B2 _1130_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_19 VGND VPWR sky130_fd_sc_hd__decap_3
X_0618_ _0552_/Y _0618_/B _0618_/C _0617_/X _0618_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XANTENNA__1075__C _1048_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0549_ _0548_/X _0549_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0716__A _0668_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_44 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_30 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_312 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_301 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0818__A2 _1111_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_367 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0626__A _0682_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_304 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_197 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1161__CLK _1130_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0754__A1 _0634_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0754__B2 _0753_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0809__A2 _1104_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_337 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0536__A _0726_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0790__A2_N _0787_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0993__A1 _0968_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0702__C _0633_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_21 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_164 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_326 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_43 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_197 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_65 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_156 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_87 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1184__CLK _1184_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_75 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0612__C _0612_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0736__A1 _0668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1162__D _1225_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_278 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_289 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_164 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_145 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0672__B1 _0501_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0952_ _1045_/A _0952_/B _0878_/Y _0988_/A VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_9_330 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0975__A1 _0859_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0883_ _0883_/A _0903_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_62_19 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_318 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_2_0_clk clkbuf_4_2_0_clk/A _1104_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_11_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_259 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1157__D _0825_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1220_ addr_r[8] baseaddr_r_sync[8] _1188_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1151_ _1159_/Q _1151_/Q _1130_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_226 VGND VPWR sky130_fd_sc_hd__decap_6
X_1082_ csb web _1163_/D VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_20_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_115 VGND VPWR sky130_fd_sc_hd__fill_2
X_0935_ _1193_/Q _0932_/X _0901_/Y d_sram_in[27] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_9_160 VGND VPWR sky130_fd_sc_hd__fill_1
X_0866_ _0910_/A _0866_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0797_ _1146_/Q _0497_/X _0797_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_28_215 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_104 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0724__A _0510_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_148 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_11 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0939__A1 _1197_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_44 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_55 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_66 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1061__B1 _1056_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_336 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1222__CLK _1191_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_204 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_41 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0618__B _0618_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_96 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_95 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0634__A _0634_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1052__B1 _1048_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0720_ _0716_/B _0720_/B _0729_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_0651_ _0500_/X _0651_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0582_ _0582_/A _0582_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_2_391 VGND VPWR sky130_fd_sc_hd__decap_6
X_1203_ addr_w[5] baseaddr_w_sync[5] _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_26_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1134_ d_sram_out[19] _1134_/Q _1184_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1065_ _1046_/A _1065_/B _0878_/Y _1066_/B VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_33_240 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0544__A _0510_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0918_ _0854_/A _0917_/X _0918_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_0849_ _0830_/Y _0839_/X _0848_/Y _0849_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_0_339 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0719__A _0651_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_310 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_44 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_229 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_398 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_10 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_43 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_54 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_111 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0901__B _0901_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0620__C _0620_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_188 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0605__A1_N _0603_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1118__CLK _1152_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0629__A _0628_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_310 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1170__D d_fabric_in[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_324 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0938__B1_N _0914_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_276 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_287 VGND VPWR sky130_fd_sc_hd__fill_2
X_0703_ _0703_/A _0700_/X _0701_/X _0702_/X _0704_/D VGND VPWR sky130_fd_sc_hd__or4_4
X_0634_ _0634_/A _0654_/A _0634_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0565_ _0584_/B _0644_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0551__A2 _0546_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0496_ _0495_/X _0496_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0539__A _0725_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_398 VGND VPWR sky130_fd_sc_hd__decap_6
X_1117_ d_sram_out[2] _1117_/Q _1130_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_1048_ _1048_/A _1048_/B _1048_/C _1048_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0705__C _0689_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1016__B1 _1012_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0721__B _0721_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_203 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0912__A _0903_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0631__B _0654_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1165__D _1165_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_313 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1090__CLK _1155_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0559__A1_N _0554_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_324 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_305 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_198 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0822__A d_sram_in[0] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0772__A2 _0669_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0617_ _0689_/B _0743_/A _0617_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0548_ _0547_/X _0548_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_368 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0716__B _0716_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_198 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0732__A out_reg VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_22 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_324 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0907__A _0876_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0626__B _0686_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_327 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_360 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0642__A _0587_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0754__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_327 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_371 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0552__A _1154_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0993__A2 _0992_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0702__D _0702_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_235 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0727__A _0508_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_22 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_305 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_44 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_22 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_349 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_66 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0612__D _0611_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0736__A2 _1126_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_110 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0637__A _1141_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_113 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0672__A1 _0668_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0951_ _0950_/Y _0952_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_20_308 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_342 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0975__A2 _0966_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0882_ _0903_/A _0899_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_56_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0547__A _0620_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_282 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_102 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_238 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_43 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1151__CLK _1130_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_124 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_64 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0920__A _1182_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0590__B1 _0578_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1173__D d_fabric_in[7] VGND VPWR sky130_fd_sc_hd__diode_2
X_1150_ _1150_/D _1150_/Q _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_238 VGND VPWR sky130_fd_sc_hd__decap_6
X_1081_ _1040_/X _1042_/Y _1079_/X w_mask[31] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_52_219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_293 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_149 VGND VPWR sky130_fd_sc_hd__fill_2
X_0934_ _1192_/Q _0932_/X _0897_/Y d_sram_in[26] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0865_ _0827_/A _0859_/X _0844_/X _0910_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0830__A _0846_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0796_ _0714_/A _0795_/X _0785_/X _1097_/Q d_fabric_out[14] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1083__D _0660_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_205 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1174__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_249 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_116 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0724__B _0726_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1061__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0939__A2 _0876_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0740__A _0721_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_396 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0618__C _0618_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_282 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_241 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0634__B _0654_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_296 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1168__D d_fabric_in[2] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1052__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0650_ _0621_/Y _0623_/X _0549_/Y _0649_/X _0650_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_0581_ _0581_/A _1150_/Q _0582_/A VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1197__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1202_ addr_w[4] baseaddr_w_sync[4] _1188_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_311 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1133_ d_sram_out[18] _0594_/A _1133_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_1_0_clk clkbuf_3_0_0_clk/X _1096_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_25_208 VGND VPWR sky130_fd_sc_hd__fill_2
X_1064_ _1046_/A _1046_/B _1045_/C _0859_/A _1066_/A VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0825__A _0825_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_403 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0544__B _0491_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_274 VGND VPWR sky130_fd_sc_hd__fill_2
X_0917_ _1173_/Q _0880_/B _0916_/X _0917_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0560__A _1127_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0848_ _0897_/A _0848_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0779_ _0665_/B _0779_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_17_89 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_285 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0793__B1 _0792_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_300 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0645__A _0606_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_274 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0784__B1 _0783_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0702_ _0741_/C _0686_/C _0633_/B _0702_/D _0702_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0633_ _0594_/A _0633_/B _0635_/B VGND VPWR sky130_fd_sc_hd__and2_4
X_0564_ _0555_/Y _0584_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0495_ _0497_/A _0495_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_57_119 VGND VPWR sky130_fd_sc_hd__decap_3
X_1116_ d_sram_out[1] _1116_/Q _1196_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1212__CLK _1188_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0555__A _1153_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1047_ _1046_/B _0838_/B _0958_/X _1048_/C VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0705__D _0705_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_266 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1016__A1 _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_299 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0721__C _0721_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0775__B1 _0773_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_344 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_391 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_266 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_255 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_248 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0912__B _0903_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0631__C _0686_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0766__B1 _0719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1181__D d_fabric_in[15] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_281 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0772__A3 _1146_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0616_ _1151_/Q _0616_/B _1146_/Q _0616_/D _0743_/A VGND VPWR sky130_fd_sc_hd__and4_4
X_0547_ _0620_/A _0488_/Y _0620_/C _0547_/X VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__1091__D _0778_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_325 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_185 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_155 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_317 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_339 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0996__B1 _0988_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1108__CLK _1108_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_56 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_89 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0937__B1_N _0910_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_163 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_347 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_144 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0626__C _0626_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_372 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0642__B _0644_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1176__D d_fabric_in[10] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_295 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_391 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_125 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0833__A _0875_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_158 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1086__D _1086_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0727__B _0724_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_12 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_114 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_67 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0743__A _0743_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_203 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_206 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0918__A _0854_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_144 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0657__C1 _0656_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0672__A2 _0673_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0950_ _1207_/Q _0950_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_32_169 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0653__A _0721_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_372 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0829__B1_N _0828_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_354 VGND VPWR sky130_fd_sc_hd__decap_12
X_0881_ _0845_/A _0903_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_49_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0828__A _0828_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0547__B _0488_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_294 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0563__A _0587_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_169 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0738__A _0681_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_11 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_22 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_21 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_324 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0920__B _0876_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0590__B2 _0589_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0590__A1 _0682_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1080_ _1035_/X _1070_/X _1079_/X w_mask[30] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_52_209 VGND VPWR sky130_fd_sc_hd__decap_4
X_0933_ _1191_/Q _0932_/X _0893_/Y d_sram_in[25] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_9_184 VGND VPWR sky130_fd_sc_hd__fill_2
X_0864_ _1171_/Q _0864_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0795_ _0575_/Y _0787_/X _1113_/D _0711_/X _0795_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__0558__A _0584_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_209 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_272 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_128 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0724__C _0741_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1061__A2 _1022_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0740__B _0721_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_76 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0618__D _0617_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_86 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1052__A2 _1015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_154 VGND VPWR sky130_fd_sc_hd__decap_4
X_0580_ _0616_/D _0566_/X _0530_/X _1122_/Q _0589_/B VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1184__D d_fabric_in[18] VGND VPWR sky130_fd_sc_hd__diode_2
X_1201_ addr_w[3] baseaddr_w_sync[3] _1096_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_334 VGND VPWR sky130_fd_sc_hd__fill_2
X_1132_ d_sram_out[17] _1132_/Q _1130_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_367 VGND VPWR sky130_fd_sc_hd__decap_8
X_1063_ _1001_/X _1059_/X _1061_/X w_mask[23] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_33_253 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0544__C _0679_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0841__A _1226_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0916_ _0903_/A _0903_/B _0908_/C _1181_/Q _0916_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0847_ _0880_/A _0859_/B _0844_/X _0846_/X _0897_/A VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__1141__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0778_ _0509_/A _0496_/X _0656_/A _0496_/X _0778_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_308 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1094__D _0788_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_79 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0793__A1 _0757_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_109 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_334 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_356 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0926__A _0876_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_367 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_253 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0645__B _0644_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1179__D d_fabric_in[13] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0661__A out_reg VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_256 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1164__CLK _1145_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0701_ _0741_/C _0701_/B _0553_/X _1132_/Q _0701_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0784__A1 _0717_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0632_ _0656_/A _0627_/Y _0703_/A _0631_/X _0632_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_0563_ _0587_/A _0606_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_31_3 VGND VPWR sky130_fd_sc_hd__decap_4
X_0494_ _0493_/X _0497_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0836__A _0845_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1115_ d_sram_out[0] _1115_/Q _1145_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_53_315 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82 VGND VPWR sky130_fd_sc_hd__decap_4
X_1046_ _1046_/A _1046_/B _0880_/B _1048_/B VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_21_245 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1089__D _1089_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0571__A _0570_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1016__A2 _1015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0775__A1 _1138_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0721__D _0721_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0775__B2 _0774_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_23 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_56 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_323 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_67 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_356 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_337 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_186 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_77 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1187__CLK _1184_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0912__C _0908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0766__A1 _0609_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_0_0_clk clkbuf_3_0_0_clk/X _1131_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_5_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0631__D _1127_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0656__A _0656_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_189 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0615_ _0614_/Y _0576_/X _1112_/D _0558_/X _0618_/C VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_0546_ _0674_/B _0521_/X _0537_/X _0546_/D _0546_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_38_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0566__A _0644_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_337 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_123 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0693__B1 _0692_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_359 VGND VPWR sky130_fd_sc_hd__decap_3
X_1029_ _0959_/Y _1026_/Y _1029_/C _1029_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_14_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_69 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0996__A1 _0985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_46 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_99 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_197 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_359 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0788__A1_N _0554_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_370 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_167 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_98 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_340 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0642__C _0586_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1202__CLK _1188_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_263 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1192__D d_fabric_in[26] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0911__A1 _0908_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_123 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_178 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_362 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1010__A _1010_/A VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_7_0_clk clkbuf_3_7_0_clk/A clkbuf_3_7_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_58_215 VGND VPWR sky130_fd_sc_hd__decap_6
X_0529_ _0528_/X _0529_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0902__A1 _1177_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_101 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_13 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0727__C _0725_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0666__B1 _0665_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_35 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_318 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_24 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_35 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_79 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_57 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_148 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_340 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0743__B _0674_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_23 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_56 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1225__CLK _1184_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_226 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_237 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0918__B _0917_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_97 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0657__B1 _0655_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_126 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_137 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_170 VGND VPWR sky130_fd_sc_hd__fill_2
X_0880_ _0880_/A _0880_/B _0880_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1187__D d_fabric_in[21] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0896__B1 _0895_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0828__B _0828_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_229 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1005__A _0982_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0648__B1 _0622_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0547__C _0620_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0844__A d_sram_in[0] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0936__B1_N _0905_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1073__B1 _1071_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_192 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0820__B1 _1113_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1097__D _0795_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0738__B _0679_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_56 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_251 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_192 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_99 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0811__B1 _1138_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_398 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0590__A2 _0553_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_262 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0664__A out_reg VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_152 VGND VPWR sky130_fd_sc_hd__fill_2
X_0932_ _0876_/A _0932_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_9_163 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0802__B1 _0655_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0863_ _0857_/Y _0833_/X _0862_/X d_sram_in[4] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_61_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_0794_ _0714_/A _0793_/X _0785_/X _1096_/Q d_fabric_out[13] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_5_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0839__A _0839_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0558__B _1153_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_229 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0574__A _0574_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0724__D _0724_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0740__C _0723_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_339 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_10 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1037__B1 _1036_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_140 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_173 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_177 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_7 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0659__A _0497_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1200_ addr_w[2] baseaddr_w_sync[2] _1131_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1093__CLK _1096_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1131_ d_sram_out[16] _0655_/A _1131_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1062_ _1026_/B _1059_/X _1061_/X w_mask[22] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_18_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_232 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0544__D _0656_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_298 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0841__B _1156_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0915_ _0912_/D _0907_/X _0914_/Y d_sram_in[14] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0846_ _0846_/A _0852_/B _0846_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0777_ _0762_/X _1090_/D _0776_/X d_fabric_out[7] VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0569__A _1153_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_210 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_243 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1019__B1 _1011_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_79 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0793__A2 _0711_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_243 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0645__C _0529_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0942__A _0942_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_235 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_268 VGND VPWR sky130_fd_sc_hd__fill_2
X_0700_ _0535_/A _0694_/B _0717_/B _1130_/Q _0700_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0784__A2 _0711_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0631_ _0535_/A _0654_/A _0686_/C _1127_/Q _0631_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1195__D d_fabric_in[29] VGND VPWR sky130_fd_sc_hd__diode_2
X_0562_ _0561_/X _0562_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0493_ _0493_/A _0493_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_24_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_1114_ _1146_/Q _1114_/Q _1130_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_53_338 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_94 VGND VPWR sky130_fd_sc_hd__decap_3
X_1045_ _1045_/A _1046_/B _1045_/C _1045_/D _1048_/A VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_21_235 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0852__A _0851_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_279 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_92 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0775__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0829_ _0880_/A _0828_/B _0828_/X d_sram_in[1] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_29_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_313 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_121 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_23 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_56 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_89 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0762__A _0663_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0912__D _0912_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_290 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0766__A2 _0765_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0923__C1 _0922_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0656__B _0717_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_176 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1131__CLK _1131_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_349 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0614_ _1113_/D _0614_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1008__A _0950_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0545_ _0540_/X _0545_/B _0545_/C _0546_/D VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_38_154 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0693__A1 _0676_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1028_ _1011_/B _1028_/B _1029_/C VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_53_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0582__A _0582_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0996__A2 _0979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_34 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0757__A _0757_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_154 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1154__CLK _1184_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_113 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_157 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0492__A _0620_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0642__D _0540_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_249 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0667__A _0493_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0911__A2 _0907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_400 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_146 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1010__B _1010_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1177__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0528_ _0527_/X _0528_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_58_205 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0902__A2 _0877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_146 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0727__D _0726_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0666__A1 _0663_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_36 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_179 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_58 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0743__C _0743_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_35 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_79 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_223 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0487__A _1132_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0657__A1 _0668_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_168 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0950__A _1207_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0896__A1 _0846_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1005__B _0982_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0648__A1 _0509_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0844__B _0828_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1021__A _0973_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1073__A1 _1022_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0820__A1 _0663_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0820__B2 _0815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0738__C _0721_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_285 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_56 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0811__A1 _0806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0811__B2 _0808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0590__A3 _0509_/A VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_6_0_clk clkbuf_3_7_0_clk/A clkbuf_3_6_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0945__A _0944_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_403 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_241 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_119 VGND VPWR sky130_fd_sc_hd__fill_2
X_0931_ _1190_/Q _0926_/X _0888_/Y d_sram_in[24] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_60_288 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1198__D addr_w[0] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0680__A _0679_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0802__A1 _0799_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0802__B2 _0801_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0862_ _0857_/Y _0839_/X _0861_/Y _0862_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0793_ _0757_/A _0711_/X _0792_/X _0793_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_54_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0558__C _0725_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1215__CLK _1133_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_252 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0574__B _0579_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_222 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0740__D _1138_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_23 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_403 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_55 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_99 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1037__A1 _0985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0796__B1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_145 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0659__B _0659_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0935__B1_N _0901_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_7 VGND VPWR sky130_fd_sc_hd__fill_2
X_1130_ d_sram_out[15] _1130_/Q _1130_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1061_ _1044_/X _1022_/X _1056_/Y _1061_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0675__A _0721_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_296 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0841__C _0845_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0914_ _0897_/A _0913_/X _0914_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_0845_ _0845_/A _0845_/B _0845_/C _0852_/B VGND VPWR sky130_fd_sc_hd__and3_4
X_0776_ _0665_/B _1090_/Q _0776_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0585__A _0585_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_391 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1019__A1 _0985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_58 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0778__B1 _0656_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_104 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_196 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0495__A _0497_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_211 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_200 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0645__D _0721_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_0630_ _0594_/B _0654_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0561_ _0585_/A _0555_/Y _1151_/Q _1150_/Q _0561_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_0492_ _0620_/A _0488_/Y _0492_/C _0498_/A _0493_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_17_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_314 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0889__B1_N _0888_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1113_ _1113_/D _1113_/Q _1130_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_177 VGND VPWR sky130_fd_sc_hd__fill_2
X_1044_ _0843_/A _1044_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_21_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_214 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0852__B _0852_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0828_ _0828_/A _0828_/B _0828_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_0759_ _0757_/X _0758_/X _0719_/X _0759_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_28_36 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_144 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_361 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1083__CLK _1145_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_56 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0923__B1 _0844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_80 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_188 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0953__A _1209_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_309 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_284 VGND VPWR sky130_fd_sc_hd__fill_2
X_0613_ _0697_/A _0701_/B _0594_/B _1141_/Q _0618_/B VGND VPWR sky130_fd_sc_hd__and4_4
X_0544_ _0510_/X _0491_/A _0679_/C _0656_/A _0545_/C VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_38_100 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1024__A _0982_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_103 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0693__A2 _0627_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_147 VGND VPWR sky130_fd_sc_hd__decap_8
X_1027_ _1007_/A _1010_/B _0999_/A _0859_/A _1028_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_41_309 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_180 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_57 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0757__B _0717_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_306 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_339 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0492__B _0488_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0948__A _0969_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0683__A _0674_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_375 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1010__C _0878_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0596__D1 _0595_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0527_ _0581_/A _0489_/Y _0527_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0858__A _0852_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0666__A2 _0660_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_37 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0593__A _0586_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_26 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_106 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0743__D _0742_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_364 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1121__CLK _1196_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_235 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_44 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0657__A2 _0502_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0678__A _1112_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0896__A2 _0890_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1005__C _1021_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0648__A2 _0703_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_272 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_191 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1021__B _1021_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1073__A2 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0820__A2 _1113_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1144__CLK _1207_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0588__A _0584_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0738__D _1122_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_24 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0811__A2 _1106_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0498__A _0498_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_286 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1167__CLK _1152_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0930_ _1189_/Q _0926_/X _0873_/X d_sram_in[23] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0802__A2 _1099_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0861_ _0905_/A _0861_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0792_ _1128_/Q _0493_/X _0792_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_47_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0558__D _0616_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_209 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_231 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0574__C _0573_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1032__A _1031_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_35 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_367 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_79 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_201 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1037__A2 _1001_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_267 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0796__A1 _0714_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0796__B2 _1097_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0956__A _1207_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_315 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_7 VGND VPWR sky130_fd_sc_hd__fill_2
X_1060_ _0992_/X _1059_/X _1057_/X w_mask[21] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0675__B _0669_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_245 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0691__A _0691_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_278 VGND VPWR sky130_fd_sc_hd__fill_2
X_0913_ _1172_/Q _0880_/B _0912_/X _0913_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_0844_ d_sram_in[0] _0828_/B _0844_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0775_ _1138_/Q _0750_/X _0773_/X _0774_/X _1090_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1027__A _1007_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0866__A _0910_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0585__B _0584_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1189_ d_fabric_in[23] _1189_/Q _1184_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_289 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1019__A2 _0992_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0778__B2 _0496_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_5_0_clk clkbuf_3_5_0_clk/A clkbuf_3_5_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_58_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_142 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0776__A _0665_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_326 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_223 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_204 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_81 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1205__CLK _1145_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0560_ _1127_/Q _0560_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0491_ _0491_/A _0492_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_2_193 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0686__A _0676_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1112_ _1112_/D _1112_/Q _1108_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1043_ _1042_/Y _1043_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_46_370 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63 VGND VPWR sky130_fd_sc_hd__decap_12
X_0827_ _0827_/A _0828_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_0758_ _0668_/X _1128_/Q _0687_/X _0758_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_0689_ _0721_/C _0689_/B _0688_/X _0689_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_29_348 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_318 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_329 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_178 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_36 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_373 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1228__CLK _1184_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0934__B1_N _0897_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_219 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0923__A1 _1183_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_112 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_104 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_362 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0612_ _0612_/A _0612_/B _0612_/C _0611_/Y _0612_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
X_0543_ _0543_/A _0656_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_145 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1024__B _0982_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_318 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_329 VGND VPWR sky130_fd_sc_hd__fill_2
X_1026_ _0984_/X _1026_/B _1026_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_34_351 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1040__A _1039_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0850__B1 _0849_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_137 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_351 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_332 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0492__C _0492_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_376 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_398 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1100__D _1132_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_218 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_80 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0964__A _1007_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0683__B _0679_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_373 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0596__C1 _0526_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0526_ _0526_/A _0526_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1035__A _1034_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_295 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_38 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_310 VGND VPWR sky130_fd_sc_hd__fill_2
X_1009_ _1046_/A _1046_/B _0982_/C _1045_/D _1009_/X VGND VPWR sky130_fd_sc_hd__and4_4
XPHY_49 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1076__B1 _1075_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_332 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_376 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_15 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_229 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_402 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1067__B1 _1066_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_60 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0814__B1 _0676_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_376 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1096__CLK _1096_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_280 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_251 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0694__A _0535_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1005__D _1021_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1058__B1 _1057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_170 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0805__B1 _0695_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1021__C _1021_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0869__A _1172_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0588__B _0585_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0509_ _0509_/A _0674_/B _0509_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_39_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_15 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_284 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1049__B1 _1048_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_7_0_clk_A clkbuf_3_7_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_324 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0779__A _0665_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_81 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_184 VGND VPWR sky130_fd_sc_hd__fill_2
X_0860_ _0828_/B _0859_/X _0880_/A _0905_/A VGND VPWR sky130_fd_sc_hd__o21a_4
X_0791_ _0714_/A _1095_/D _0785_/X _1095_/Q d_fabric_out[12] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_9_188 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0689__A _0721_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_74 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1111__CLK _1207_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0989_ _0985_/X _0974_/X _0988_/Y _0989_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0599__A _0574_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_302 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_254 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_46 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_132 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0796__A2 _0795_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_125 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_327 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_210 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1134__CLK _1184_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0675__C _0676_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_80 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0972__A _0972_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_257 VGND VPWR sky130_fd_sc_hd__fill_2
X_0912_ _0903_/A _0903_/B _0908_/C _0912_/D _0912_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0843_ _0843_/A _0859_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_0774_ _1122_/Q _0497_/X _0709_/X _0774_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1027__B _1010_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_305 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0585__C _0582_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1043__A _1042_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_1188_ d_fabric_in[22] _1188_/Q _1188_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_24_202 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0882__A _0903_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1157__CLK _1196_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0776__B _1090_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_235 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0792__A _1128_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1103__D _0634_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_268 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_257 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_227 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_290 VGND VPWR sky130_fd_sc_hd__decap_4
X_0490_ _0489_/Y _0491_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0686__B _0655_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_327 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_1111_ _0532_/A _1111_/Q _1207_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1042_ _0899_/A _0899_/B _0831_/C _1042_/D _1042_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_53_319 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_396 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_51 VGND VPWR sky130_fd_sc_hd__decap_8
X_0826_ _0845_/A _0845_/B _0831_/C _0828_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA_clkbuf_4_6_0_clk_A clkbuf_4_6_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0757_ _0757_/A _0717_/B _0757_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0688_ _0688_/A _0687_/X _0688_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0877__A _0876_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_15_0_clk clkbuf_3_7_0_clk/X _1191_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_44_26 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_209 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0923__A2 _0876_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0787__A _0495_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_146 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_116 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_352 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_396 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_231 VGND VPWR sky130_fd_sc_hd__fill_2
X_0611_ _0741_/C _0689_/B _0610_/Y _0611_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_50_91 VGND VPWR sky130_fd_sc_hd__fill_1
X_0542_ _0681_/A _0726_/B _0679_/C _0634_/A _0545_/B VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0697__A _0697_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_124 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1024__C _0999_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_4_0_clk clkbuf_3_5_0_clk/A clkbuf_3_4_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1025_ _1025_/A _1025_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_34_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_363 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0850__A1 _0830_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0809_ _0806_/X _1104_/Q _0675_/D _0808_/X d_fabric_out[21] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_39_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_26 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_374 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_311 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_344 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0492__D _0498_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_212 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0964__B _1021_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_190 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0683__C _0681_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_91 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_108 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_171 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_182 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_1_1_0_clk_A clkbuf_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0596__B1 _0718_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0525_ _0655_/A _0608_/B _0526_/A VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0933__B1_N _0893_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0615__A1_N _0614_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1218__CLK _1131_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_274 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_28 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VPWR sky130_fd_sc_hd__decap_3
X_1008_ _0950_/Y _1046_/B VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_39 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1076__A1 _0984_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_182 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0890__A _0880_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1201__D addr_w[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_344 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_388 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_3_0_clk_A clkbuf_3_3_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_230 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1067__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_193 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0814__A1 _0813_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0814__B2 _0808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1111__D _0532_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_388 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_174 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_14_0_clk_A clkbuf_3_7_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_71 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0694__B _0694_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_285 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1058__A1 _0983_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0805__B2 _0801_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1021__D _1021_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0805__A1 _0799_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0588__C _0586_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1046__A _1046_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0508_ _0508_/A _0674_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0885__A _0845_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1190__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_403 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_263 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1049__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_15 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_174 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0980__B1 _0975_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1106__D _1138_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_71 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_93 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_247 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_258 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_167 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_156 VGND VPWR sky130_fd_sc_hd__decap_4
X_0790_ _0560_/Y _0787_/X _0532_/A _0787_/X _1095_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__0689__B _0689_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_236 VGND VPWR sky130_fd_sc_hd__decap_6
X_0988_ _0988_/A _0988_/B _0959_/Y _0988_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0599__B _0701_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_325 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_14 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_247 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1086__CLK _1155_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0650__C1 _0649_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_0_0_clk_A clkbuf_1_0_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_376 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_306 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_200 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_222 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0675__D _0675_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_391 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_236 VGND VPWR sky130_fd_sc_hd__fill_2
X_0911_ _0908_/D _0907_/X _0910_/Y d_sram_in[13] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0842_ _0841_/X _0843_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0773_ _0771_/X _0772_/X _0719_/X _0773_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_52_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1027__C _0999_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_328 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0585__D _1116_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1187_ d_fabric_in[21] _1187_/Q _1184_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA_clkbuf_4_2_0_clk_A clkbuf_4_2_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_28 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_280 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0632__C1 _0631_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0792__B _0493_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_94 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1101__CLK _1207_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_173 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_7 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_114 VGND VPWR sky130_fd_sc_hd__fill_2
X_1110_ _0691_/A _1110_/Q _1108_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0686__C _0686_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_32 VGND VPWR sky130_fd_sc_hd__decap_3
X_1041_ _0944_/X _1040_/X _1037_/X w_mask[15] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0983__A _0983_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_350 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_96 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_85 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_74 VGND VPWR sky130_fd_sc_hd__decap_6
X_0825_ _0825_/A _0831_/C VGND VPWR sky130_fd_sc_hd__buf_1
X_0756_ _0663_/X _1087_/D _0755_/X d_fabric_out[4] VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0917__B1 _0916_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0687_ _0675_/D _0654_/A _0687_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_28_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_317 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1204__D addr_w[6] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0893__A _0910_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_206 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0853__C1 _0852_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_283 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1124__CLK _1104_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_309 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1114__D _1146_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_128 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_191 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_82 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_272 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_243 VGND VPWR sky130_fd_sc_hd__fill_1
X_0610_ _0675_/D _0582_/X _0688_/A _0608_/X _0609_/X _0610_/Y VGND VPWR sky130_fd_sc_hd__a2111oi_4
XANTENNA__0978__A _0973_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0541_ _0535_/A _0679_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0697__B _0694_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1024__D _1021_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_169 VGND VPWR sky130_fd_sc_hd__fill_2
X_1024_ _0982_/A _0982_/B _0999_/X _1021_/D _1025_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_34_320 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_386 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0850__A2 _0833_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_172 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1147__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0808_ _0665_/B _0808_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0888__A _0880_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0739_ _0722_/A _0492_/C _0723_/C _0739_/D _0739_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_39_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_386 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_323 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_183 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1109__D _1141_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_10_0_clk_A clkbuf_3_5_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_93 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0964__C _1209_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_301 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0683__D _0683_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_367 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_14_0_clk clkbuf_3_7_0_clk/X _1171_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0596__A1 _1134_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0524_ _0581_/A _0491_/A _0608_/B VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0501__A _0500_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_29 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VPWR sky130_fd_sc_hd__decap_3
X_1007_ _1007_/A _1046_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1076__A2 _1035_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_39 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_249 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_253 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1067__A2 _1025_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_109 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_62 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_367 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0814__A2 _1108_/Q VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_3_0_clk clkbuf_3_3_0_clk/A clkbuf_4_6_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_31_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_271 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0694__C _0582_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_150 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0991__A _0982_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1058__A2 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0805__A2 _1102_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_153 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0588__D _0587_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1046__B _1046_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0507_ _0720_/B _0508_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_36_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_267 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1212__D addr_r[0] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1049__A2 _1006_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_289 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_120 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0980__A1 _0968_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_267 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1122__D d_sram_out[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_153 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1208__CLK _1207_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_60 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_330 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0689__C _0688_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0986__A _0859_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_98 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_201 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_19 VGND VPWR sky130_fd_sc_hd__fill_2
X_0987_ _1045_/A _1065_/B _0982_/C _1045_/D _0988_/B VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0599__C _0553_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1207__D addr_w[9] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_26 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_278 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_112 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_105 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0650__B1 _0549_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_149 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1117__D d_sram_out[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_267 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_215 VGND VPWR sky130_fd_sc_hd__fill_2
X_0910_ _0910_/A _0909_/X _0910_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_0841_ _1226_/Q _1156_/D _0845_/C _0841_/X VGND VPWR sky130_fd_sc_hd__or3_4
X_0772_ _0676_/A _0669_/X _1146_/Q _0668_/A _1130_/Q _0772_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__1180__CLK _1145_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1027__D _0859_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1186_ d_fabric_in[20] _1186_/Q _1130_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_24_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0632__B1 _0703_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0935__A1 _1193_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_167 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0871__B1 _0870_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_403 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_62 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0623__B1 _0622_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_9 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_185 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0686__D _1128_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_159 VGND VPWR sky130_fd_sc_hd__decap_12
X_1040_ _1039_/X _1040_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_64_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0862__B1 _0861_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_218 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0504__A _1152_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0824_ _1156_/D _0845_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0755_ _0732_/X _1087_/Q _0755_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0917__A1 _1173_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0686_ _0676_/C _0655_/B _0686_/C _1128_/Q _0686_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0893__B _0892_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1169_ d_fabric_in[3] _0851_/A _1188_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1070__A _1042_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_332 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0853__B1 _0844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1220__D addr_r[8] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_398 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0605__B1 _0691_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1030__B1 _1029_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_40 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_332 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_365 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1130__D d_sram_out[15] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_61 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_284 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_93 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0978__B _0952_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0540_ _0681_/A _0679_/B _0682_/C _0540_/D _0540_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1099__CLK _1196_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0697__C _0530_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0994__A _1010_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_310 VGND VPWR sky130_fd_sc_hd__decap_4
X_1023_ _0998_/X _1022_/X _1019_/X w_mask[11] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_53_107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_398 VGND VPWR sky130_fd_sc_hd__decap_6
X_0807_ _0806_/X _1103_/Q _0634_/A _0801_/X d_fabric_out[20] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1012__B1 _1011_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0738_ _0681_/A _0679_/B _0721_/C _1122_/Q _0738_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0888__B _0888_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1065__A _1046_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0669_ _0721_/B _0669_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1215__D addr_r[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_159 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1079__B1 _1075_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_321 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_365 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0826__B1 _0831_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1125__D d_sram_out[10] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0964__D _0972_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0817__B1 _0739_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_184 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_379 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0596__A2 _0530_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0523_ _0523_/A _0581_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_26_118 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_170 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1114__CLK _1130_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1006_ _1005_/X _1006_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0899__A _0899_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_41 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_30 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_198 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_40 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0602__A _0697_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1137__CLK _1108_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0694__D _1126_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_257 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0991__B _0952_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_361 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0512__A _0722_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1046__C _0880_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0506_ _0505_/X _0720_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_36_18 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0980__A2 _0979_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_13_0_clk clkbuf_3_6_0_clk/X _1184_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_60_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_147 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_268 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0507__A _0720_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_249 VGND VPWR sky130_fd_sc_hd__fill_1
X_0986_ _0859_/A _1045_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0599__D _0543_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_213 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1223__D addr_r[11] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_38 VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_2_0_clk clkbuf_3_3_0_clk/A clkbuf_4_5_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0650__A1 _0621_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_117 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_356 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_257 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1133__D d_sram_out[18] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_227 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_290 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_282 VGND VPWR sky130_fd_sc_hd__fill_2
X_0840_ _0825_/A _0845_/C VGND VPWR sky130_fd_sc_hd__inv_8
X_0771_ _1138_/Q _0655_/B _0771_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_38_3 VGND VPWR sky130_fd_sc_hd__fill_1
X_1185_ d_fabric_in[19] _1185_/Q _1191_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_374 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_260 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_271 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0632__A1 _0656_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0969_ _0969_/A _0973_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0935__A2 _0932_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1218__D addr_r[6] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0700__A _0535_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_135 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0931__B1_N _0888_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_249 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0871__A1 _0869_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0623__A1 _1115_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1128__D d_sram_out[13] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_319 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0862__A1 _0857_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_282 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_293 VGND VPWR sky130_fd_sc_hd__decap_12
X_0823_ _1226_/Q _0845_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0754_ _0634_/A _0750_/X _0752_/X _0753_/X _1087_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__0917__A2 _0880_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0685_ _0674_/X _0684_/Y _0550_/X _0685_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0520__A _0682_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_105 VGND VPWR sky130_fd_sc_hd__fill_1
X_1168_ d_fabric_in[2] _0846_/A _1133_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_396 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0853__A1 _0827_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1099_ _0655_/A _1099_/Q _1196_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0605__B2 _0604_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_241 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1030__A1 _0944_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_127 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1170__CLK _1191_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_96 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_171 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_296 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_83 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0978__C _1021_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0697__D _1122_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0780__B1 _0762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_70 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0994__B _1010_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_149 VGND VPWR sky130_fd_sc_hd__fill_2
X_1022_ _1021_/X _1022_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_53_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_396 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0515__A _0679_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0806_ _0661_/Y _0806_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1012__A1 _0985_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0737_ _1126_/Q _0720_/B _0737_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0888__C _0905_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1065__B _1065_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0668_ _0668_/A _0668_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1193__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0599_ _0574_/A _0701_/B _0553_/X _0543_/A _0612_/A VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_57_403 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_116 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1079__A1 _0984_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_355 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0826__A1 _0845_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_196 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_182 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1141__D d_sram_out[26] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0817__A1 _0813_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0817__B2 _0815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_358 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_44 VGND VPWR sky130_fd_sc_hd__decap_12
X_0522_ _1151_/Q _0523_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0753__B1 _0709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_200 VGND VPWR sky130_fd_sc_hd__decap_12
X_1005_ _0982_/A _0982_/B _1021_/C _1021_/D _1005_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_22_314 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0899__B _0899_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1226__D conf[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_174 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1089__CLK _1155_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0602__B _0701_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0735__B1 _0695_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1136__D d_sram_out[21] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_240 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_200 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_244 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_266 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_174 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0991__C _0982_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_100 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_373 VGND VPWR sky130_fd_sc_hd__decap_12
X_0505_ _0616_/B _0584_/A _0505_/X VGND VPWR sky130_fd_sc_hd__or2_4
.ends

