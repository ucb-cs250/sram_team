* NGSPICE file created from sram_ifc.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 D Q CLK VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 X VGND VPWR
.ends

.subckt sram_ifc addr_r[0] addr_r[10] addr_r[11] addr_r[12] addr_r[13] addr_r[1] addr_r[2]
+ addr_r[3] addr_r[4] addr_r[5] addr_r[6] addr_r[7] addr_r[8] addr_r[9] addr_w[0]
+ addr_w[10] addr_w[11] addr_w[12] addr_w[13] addr_w[1] addr_w[2] addr_w[3] addr_w[4]
+ addr_w[5] addr_w[6] addr_w[7] addr_w[8] addr_w[9] baseaddr_r_sync[0] baseaddr_r_sync[1]
+ baseaddr_r_sync[2] baseaddr_r_sync[3] baseaddr_r_sync[4] baseaddr_r_sync[5] baseaddr_r_sync[6]
+ baseaddr_r_sync[7] baseaddr_r_sync[8] baseaddr_w_sync[0] baseaddr_w_sync[1] baseaddr_w_sync[2]
+ baseaddr_w_sync[3] baseaddr_w_sync[4] baseaddr_w_sync[5] baseaddr_w_sync[6] baseaddr_w_sync[7]
+ baseaddr_w_sync[8] clk conf[0] conf[1] conf[2] csb csb0_sync csb1_sync d_fabric_in[0]
+ d_fabric_in[10] d_fabric_in[11] d_fabric_in[12] d_fabric_in[13] d_fabric_in[14]
+ d_fabric_in[15] d_fabric_in[16] d_fabric_in[17] d_fabric_in[18] d_fabric_in[19]
+ d_fabric_in[1] d_fabric_in[20] d_fabric_in[21] d_fabric_in[22] d_fabric_in[23] d_fabric_in[24]
+ d_fabric_in[25] d_fabric_in[26] d_fabric_in[27] d_fabric_in[28] d_fabric_in[29]
+ d_fabric_in[2] d_fabric_in[30] d_fabric_in[31] d_fabric_in[3] d_fabric_in[4] d_fabric_in[5]
+ d_fabric_in[6] d_fabric_in[7] d_fabric_in[8] d_fabric_in[9] d_fabric_out[0] d_fabric_out[10]
+ d_fabric_out[11] d_fabric_out[12] d_fabric_out[13] d_fabric_out[14] d_fabric_out[15]
+ d_fabric_out[16] d_fabric_out[17] d_fabric_out[18] d_fabric_out[19] d_fabric_out[1]
+ d_fabric_out[20] d_fabric_out[21] d_fabric_out[22] d_fabric_out[23] d_fabric_out[24]
+ d_fabric_out[25] d_fabric_out[26] d_fabric_out[27] d_fabric_out[28] d_fabric_out[29]
+ d_fabric_out[2] d_fabric_out[30] d_fabric_out[31] d_fabric_out[3] d_fabric_out[4]
+ d_fabric_out[5] d_fabric_out[6] d_fabric_out[7] d_fabric_out[8] d_fabric_out[9]
+ d_sram_in[0] d_sram_in[10] d_sram_in[11] d_sram_in[12] d_sram_in[13] d_sram_in[14]
+ d_sram_in[15] d_sram_in[16] d_sram_in[17] d_sram_in[18] d_sram_in[19] d_sram_in[1]
+ d_sram_in[20] d_sram_in[21] d_sram_in[22] d_sram_in[23] d_sram_in[24] d_sram_in[25]
+ d_sram_in[26] d_sram_in[27] d_sram_in[28] d_sram_in[29] d_sram_in[2] d_sram_in[30]
+ d_sram_in[31] d_sram_in[3] d_sram_in[4] d_sram_in[5] d_sram_in[6] d_sram_in[7] d_sram_in[8]
+ d_sram_in[9] d_sram_out[0] d_sram_out[10] d_sram_out[11] d_sram_out[12] d_sram_out[13]
+ d_sram_out[14] d_sram_out[15] d_sram_out[16] d_sram_out[17] d_sram_out[18] d_sram_out[19]
+ d_sram_out[1] d_sram_out[20] d_sram_out[21] d_sram_out[22] d_sram_out[23] d_sram_out[24]
+ d_sram_out[25] d_sram_out[26] d_sram_out[27] d_sram_out[28] d_sram_out[29] d_sram_out[2]
+ d_sram_out[30] d_sram_out[31] d_sram_out[3] d_sram_out[4] d_sram_out[5] d_sram_out[6]
+ d_sram_out[7] d_sram_out[8] d_sram_out[9] out_reg reb w_mask[0] w_mask[10] w_mask[11]
+ w_mask[12] w_mask[13] w_mask[14] w_mask[15] w_mask[16] w_mask[17] w_mask[18] w_mask[19]
+ w_mask[1] w_mask[20] w_mask[21] w_mask[22] w_mask[23] w_mask[24] w_mask[25] w_mask[26]
+ w_mask[27] w_mask[28] w_mask[29] w_mask[2] w_mask[30] w_mask[31] w_mask[3] w_mask[4]
+ w_mask[5] w_mask[6] w_mask[7] w_mask[8] w_mask[9] web web0_sync VPWR VGND
XANTENNA__1231__CLK _1256_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0703__A _0861_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1142__B1 _1141_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_41 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_62 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0986__C _0986_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1254__CLK _1288_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1270_ addr_w[10] _1270_/Q _1166_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1133__B1 _1128_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0985_ _0953_/Y _0966_/X _1242_/Q _0919_/Y _0985_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__0523__A _0546_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1124__B1 _1123_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_35 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_68 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_114 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0650__A2 _0649_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_54 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1277__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1115__B1 _1114_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0608__A _0608_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_83 VGND VPWR sky130_fd_sc_hd__decap_3
X_0770_ _0533_/X _0763_/Y _0765_/Y _0767_/Y _0769_/Y _0770_/X VGND VPWR sky130_fd_sc_hd__o41a_4
XFILLER_68_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_114 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0562__D1 _0561_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_147 VGND VPWR sky130_fd_sc_hd__fill_2
X_1253_ d_fabric_in[25] _1253_/Q _1253_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_83_128 VGND VPWR sky130_fd_sc_hd__fill_2
X_1184_ d_sram_out[7] _1184_/Q _1184_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0518__A _0518_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0880__A2 _1167_/Q VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_12_0_clk clkbuf_3_6_0_clk/X _1184_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0968_ _0994_/A _0966_/X _1237_/Q _0967_/X _0968_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
X_0899_ _0899_/A _0994_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_59_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_147 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1234__D d_fabric_in[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_180 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0610__B _0547_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0720__A1_N _0889_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_109 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0862__A2 _1160_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_44 VGND VPWR sky130_fd_sc_hd__decap_3
X_0822_ _0822_/A _0822_/B _0786_/A _0822_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_0753_ _0752_/Y _0753_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0684_ _0600_/X _1161_/D _0683_/Y _0684_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_50_3 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_1_0_clk clkbuf_3_1_0_clk/A clkbuf_4_2_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_56_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_139 VGND VPWR sky130_fd_sc_hd__fill_1
X_1236_ d_fabric_in[8] _0963_/D _1256_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1167_ _0607_/C _1167_/Q _1172_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0853__A2 _1158_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1098_ _1071_/Y _1106_/A _1098_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1079__A _1030_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_174 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1229__D d_fabric_in[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_89 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_27 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1030__A2 _0919_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0711__A _0709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_150 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_120 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_40 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_73 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_185 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0621__A _0621_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0978__D _1240_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0780__A1 _0822_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_106 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0994__C _0960_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_70 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_150 VGND VPWR sky130_fd_sc_hd__decap_4
X_1021_ _1020_/Y _1074_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_61_120 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_80 VGND VPWR sky130_fd_sc_hd__fill_1
X_0805_ _1190_/Q _0805_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1049__D _1083_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0736_ _0736_/A _0736_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_115_111 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0531__A _0528_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0667_ _0606_/B _0667_/B _1173_/D _0667_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__0771__A1 _1179_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1065__C _1102_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0598_ _0635_/A _0621_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_130_147 VGND VPWR sky130_fd_sc_hd__decap_12
X_1219_ _0919_/B _1219_/Q _1177_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_24 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0706__A _1145_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_43 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1003__A2 _1000_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_177 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_172 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_186 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0616__A _0588_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_90 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0521_ _0520_/X _0521_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_158 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_169 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_80 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0808__A2 _0807_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1004_ _1252_/Q _0960_/X _0964_/X d_sram_in[24] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_34_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0526__A _0729_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1160__CLK _1173_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0719_ _0666_/Y _0716_/X _0719_/C _0719_/D _0719_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_106_13 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1092__A _1088_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1242__D d_fabric_in[14] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_54 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0983__A1 _1241_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0602__C _0595_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1152__D _0825_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_101 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1183__CLK _1180_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_192 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0974__B2 _0967_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0726__A1 _0654_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0965__A1 _0963_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_12 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_23 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1237__D d_fabric_in[9] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_55 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1142__A1 _1097_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_86 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1147__D _0772_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0986__D _0930_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_148 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_93 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1133__A1 _1024_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0892__B1 _0891_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0804__A _0608_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0984_ _0960_/A _0984_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0947__A1 _0977_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_115 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_159 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1124__A1 _1067_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0714__A _0576_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_159 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1115__A1 _1049_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_63 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0608__B _0608_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0624__A _0621_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1221__CLK _1218_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_174 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_92 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0562__C1 _0553_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1252_ d_fabric_in[24] _1252_/Q _1252_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1183_ d_sram_out[6] _0628_/C _1180_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0865__B1 _0864_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_173 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0534__A _0542_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0967_ _0919_/Y _0967_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0898_ _0874_/X _1176_/Q _0897_/Y d_fabric_out[31] VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_114_13 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1250__D d_fabric_in[22] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_78 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_56 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1244__CLK _1253_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_95 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_73 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_62 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0619__A _0604_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0847__B1 _0846_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_50 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1160__D _1160_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_60 VGND VPWR sky130_fd_sc_hd__fill_1
X_0821_ _0807_/A _0819_/Y _0897_/A _0763_/C _0821_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_9_89 VGND VPWR sky130_fd_sc_hd__decap_3
X_0752_ _0743_/Y _0751_/Y _0699_/X _0752_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_127_120 VGND VPWR sky130_fd_sc_hd__decap_6
X_0683_ _0682_/X _0683_/B _0683_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_89_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0529__A _0542_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1235_ d_fabric_in[7] _0988_/D _1253_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0838__B1 _0837_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1166_ _0608_/C _0877_/A _1166_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_184 VGND VPWR sky130_fd_sc_hd__decap_6
X_1097_ _1136_/A _1097_/B _1102_/C _1097_/D _1097_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__1267__CLK _1274_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1079__B _1077_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1095__A _1095_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0711__B _0595_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_23 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1245__D d_fabric_in[17] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_49 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_107 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0829__B1 _0828_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_98 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_53 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_75 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0902__A _0902_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1006__B1 _0972_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0621__B _0621_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1155__D _0839_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0780__A2 _0779_/Y VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_clk clkbuf_3_5_0_clk/X _1173_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1020_ _1058_/A _1020_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_46_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_154 VGND VPWR sky130_fd_sc_hd__fill_1
X_0804_ _0608_/C _0804_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0735_ _0667_/B _0520_/X _0729_/B _1174_/D _0736_/A VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__0531__B _0763_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0666_ _0667_/B _0520_/X _0594_/X _0666_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_130_104 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1065__D _1097_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0771__A2 _0566_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0597_ _0588_/C _0597_/B _0635_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_130_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_107 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0781__A1_N _0889_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1218_ _0902_/A _1218_/Q _1218_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_111_47 VGND VPWR sky130_fd_sc_hd__decap_6
X_1149_ _0802_/A _1149_/Q _1159_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_111_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_176 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0706__B _0705_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0722__A _0721_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_85 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0616__B _0587_/A VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_0_0_clk clkbuf_3_1_0_clk/A clkbuf_3_0_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_80 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_51 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_40 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0632__A _0544_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0520_ _0588_/B _0520_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_126 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_92 VGND VPWR sky130_fd_sc_hd__fill_2
X_1003_ _1251_/Q _1000_/X _0958_/X d_sram_in[23] VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0807__A _0807_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_143 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0542__A _0542_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0718_ _0718_/A _0544_/X _0550_/X _0624_/B _0719_/D VGND VPWR sky130_fd_sc_hd__and4_4
X_0649_ _0574_/X _0683_/B _0551_/B _0649_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_106_58 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1092__B _1136_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_121 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0717__A _0612_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_66 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_32 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0983__A2 _0957_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0602__D _0601_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0627__A _0608_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_72 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_135 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_7 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_193 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0726__A2 _1178_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_135 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_80 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0537__A _0518_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_157 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0965__A2 _0960_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1142__A2 _1132_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1253__D d_fabric_in[25] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_42 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0910__A _0922_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1163__D _1195_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1133__A2 _1095_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0892__A1 _0874_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1150__CLK _1166_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0983_ _1241_/Q _0957_/X _0982_/Y d_sram_in[13] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_73_3 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_161 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0947__A2 _0941_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0820__A _1208_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1124__A2 _1121_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_19 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0714__B _0612_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1098__A _1071_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_23 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1248__D d_fabric_in[20] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0730__A _0729_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_49 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1173__CLK _1173_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1115__A2 _1105_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_182 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0608__C _0608_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_63 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_52 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0905__A _0919_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0624__B _0624_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1158__D _1158_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0640__A _0640_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_186 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_82 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0562__B1 _0533_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1251_ d_fabric_in[23] _1251_/Q _1288_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1182_ d_sram_out[5] _1182_/Q _1180_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0865__A1 _0843_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_92 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_185 VGND VPWR sky130_fd_sc_hd__decap_4
X_0966_ _1060_/B _0966_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0550__A _0608_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0897_ _0897_/A _0893_/B _0897_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__1196__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_101 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0792__B1 _0782_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0619__B _0613_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_152 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0847__A1 _0672_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_185 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_73 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0635__A _0635_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_68 VGND VPWR sky130_fd_sc_hd__decap_12
X_0820_ _1208_/Q _0897_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_0751_ _0746_/X _0748_/Y _0750_/X _0751_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_127_154 VGND VPWR sky130_fd_sc_hd__decap_6
X_0682_ _0558_/X _0682_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_36_3 VGND VPWR sky130_fd_sc_hd__decap_4
X_1234_ d_fabric_in[6] _1234_/Q _1252_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_49_182 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0529__B _0573_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0838__A1 _0768_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1165_ _0606_/C _0875_/A _1159_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1096_ _1043_/X _1095_/Y _1093_/X w_mask[13] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0545__A _0544_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1079__C _1093_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0949_ _0949_/A _0949_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1095__B _1102_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0711__C _0711_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_22 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0829__A1 _0683_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1261__D addr_w[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_133 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1211__CLK _1177_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_43 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_110 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1006__A1 _1254_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_53 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0621__C _0621_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0765__B1 _0764_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1171__D _1203_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_166 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_93 VGND VPWR sky130_fd_sc_hd__decap_3
X_0803_ _0704_/X _1149_/Q _0802_/Y d_fabric_out[4] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0734_ _0822_/A _0536_/X _0730_/X _0747_/A _0734_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_115_124 VGND VPWR sky130_fd_sc_hd__decap_6
X_0665_ _0660_/X _0661_/Y _0664_/X _0677_/A VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_115_135 VGND VPWR sky130_fd_sc_hd__fill_2
X_0596_ _0587_/A _0597_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1234__CLK _1252_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1217_ _0914_/A _1217_/Q _1253_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_1_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_1148_ _1148_/D _0795_/B _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1079_ _1030_/Y _1077_/Y _1093_/B _1079_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__1256__D d_fabric_in[28] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_89 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_32 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_122 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_63 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0632__B _0606_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1166__D _0608_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_116 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1257__CLK _1177_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_174 VGND VPWR sky130_fd_sc_hd__fill_2
X_1002_ _1250_/Q _1000_/X _0954_/Y d_sram_in[22] VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0807__B _0807_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0717_ _0612_/A _0621_/B _0637_/B _0719_/C VGND VPWR sky130_fd_sc_hd__and3_4
X_0648_ _1185_/Q _0683_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_103_149 VGND VPWR sky130_fd_sc_hd__decap_4
X_0579_ _0607_/A _0609_/A _1195_/Q _0579_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__1092__C _1102_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0717__B _0621_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_166 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0733__A _0539_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0968__B1 _1237_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_22 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_10_0_clk clkbuf_3_5_0_clk/X _1172_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_103_3 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0908__A d_sram_in[0] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0627__B _0628_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_62 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_161 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0959__B1 _0958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0643__A _0623_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_194 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_114 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0553__A _0541_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0748__A1_N _0747_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0728__A _0807_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_87 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0910__B _0910_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_117 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0638__A _0637_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0892__A2 _1173_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0982_ _0950_/X _0981_/Y _0982_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_66_3 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_150 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0548__A _0615_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_139 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0714__C _0621_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1098__B _1106_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_35 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_68 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_128 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1264__D addr_w[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_43 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0624__C _0624_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_121 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0921__A _0921_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_132 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0640__B _0636_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_8 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1174__D _1174_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0562__A1 _1189_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1250_ d_fabric_in[22] _1250_/Q _1253_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_76_150 VGND VPWR sky130_fd_sc_hd__fill_2
X_1181_ d_sram_out[4] _0627_/C _1180_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0865__A2 _1161_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0965_ _0963_/D _0960_/X _0964_/X d_sram_in[8] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0831__A _0883_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0896_ _0589_/Y _0775_/X _0895_/Y d_fabric_out[30] VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_59_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_139 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_37 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_175 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_23 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1259__D d_fabric_in[31] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_113 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0792__B2 _0791_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1290__CLK _1274_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0619__C _0619_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_131 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0847__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0916__A _0915_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0635__B _0623_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1169__D _1169_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0750_ _0749_/X _0750_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0651__A _0698_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0681_ _0652_/Y _0655_/X _0680_/Y _0681_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_89_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_150 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1233_ d_fabric_in[5] _0949_/A _1288_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_49_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0838__A2 _0760_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1164_ _1196_/Q _1164_/Q _1172_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0826__A _0826_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1095_ _1095_/A _1102_/B _1102_/C _1097_/D _1095_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_100_28 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1163__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0948_ _0977_/D _0916_/X _0947_/X d_sram_in[4] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_109_26 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1095__C _1102_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0879_ _0663_/Y _0889_/B _0879_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_125_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_120 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0829__A2 _0760_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0736__A _0736_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_123 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_22 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_33 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_3 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1006__A2 _1000_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_144 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_65 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0765__A1 _0551_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_80 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0646__A _0640_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_72 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1186__CLK _1184_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0802_ _0802_/A _0893_/B _0802_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_0733_ _0539_/X _0822_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0664_ _0662_/Y _0588_/Y _0663_/Y _0615_/Y _0664_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_0595_ _0528_/X _0621_/B _0594_/X _1208_/Q _0595_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_1216_ _1216_/D _0602_/A _1256_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_101 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0556__A _0555_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1147_ _0772_/X _1147_/Q _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_111_16 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_156 VGND VPWR sky130_fd_sc_hd__decap_4
X_1078_ _1075_/A _1127_/B _1127_/C _1093_/B VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_106_114 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_7 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1272__D addr_w[12] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_164 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_93 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_86 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0632__C _0615_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_7 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1182__D d_sram_out[5] VGND VPWR sky130_fd_sc_hd__diode_2
X_1001_ _1249_/Q _1000_/X _0951_/Y d_sram_in[21] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_34_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0807__C _1174_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0674__B1 _0576_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1000__A _0960_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0716_ _0574_/X _0615_/B _0594_/X _0577_/X _0716_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_103_106 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1201__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0647_ _0634_/Y _0646_/Y _0647_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_103_117 VGND VPWR sky130_fd_sc_hd__fill_2
X_0578_ _0574_/X _1161_/D _0576_/X _0577_/X _0578_/Y VGND VPWR sky130_fd_sc_hd__a22oi_4
XANTENNA__1092__D _1083_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_101 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0717__C _0637_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_115 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0968__B2 _0967_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_67 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1267__D addr_w[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_78 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_86 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0627__C _0627_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0924__A _0920_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_148 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_151 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0643__B _1178_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0959__A1 _0988_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_184 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1081__B1 _1080_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_195 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1224__CLK _1253_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1177__D d_sram_out[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_115 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_126 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_60 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_104 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_137 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0553__B _0551_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1072__B1 _1068_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_37 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_19 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_181 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0886__B1 _0885_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0728__B _0763_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0744__A _0682_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_126 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1247__CLK _1288_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1063__B1 _1062_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0810__B1 _0808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0910__C _0909_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0919__A _0922_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_80 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0654__A _0653_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0981_ _0949_/Y _0966_/X _1241_/Q _0967_/X _0981_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_12_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_152 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0801__B1 _0798_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_39 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0564__A _0691_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_47 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_140 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1280__D addr_r[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0640__C _0639_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_166 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0562__A2 _0531_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0649__A _0574_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1180_ d_sram_out[3] _0624_/B _1180_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_76_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_50 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1190__D d_sram_out[13] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_154 VGND VPWR sky130_fd_sc_hd__fill_2
X_0964_ _0964_/A _0962_/Y _0963_/Y _0964_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__0831__B _0831_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0895_ _1175_/Q _0895_/B _0895_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_59_129 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0559__A _1161_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_15 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_19 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1275__D addr_r[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_43 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_10 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_87 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0635__C _1186_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_92 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1009__B1 _0982_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0651__B _0570_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0680_ _0679_/Y _0566_/A _0680_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_50_7 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_83 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1185__D d_sram_out[8] VGND VPWR sky130_fd_sc_hd__diode_2
X_1232_ d_fabric_in[4] _0977_/D _1288_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1163_ _1195_/Q _1163_/Q _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0826__B _0826_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1094_ _1043_/X _1090_/Y _1093_/X w_mask[12] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0947_ _0977_/D _0941_/Y _0964_/A _0947_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_109_16 VGND VPWR sky130_fd_sc_hd__decap_4
X_0878_ _0804_/Y _0775_/X _0877_/Y d_fabric_out[21] VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__1095__D _1097_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_48 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_132 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_165 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_189 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0765__A2 _0668_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_41 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0927__A _1104_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_74 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0646__B _0646_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_7 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0662__A _1203_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0801_ _0797_/Y _0692_/X _0798_/Y _0800_/Y _0802_/A VGND VPWR sky130_fd_sc_hd__a22oi_4
X_0732_ _0731_/Y _0732_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0663_ _0607_/C _0663_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0594_ _0588_/D _0594_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_130_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_110 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0837__A _0859_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1215_ _1215_/D _0587_/A _1252_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_165 VGND VPWR sky130_fd_sc_hd__fill_2
X_1146_ _0753_/Y _0754_/B _1177_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_111_28 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_113 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_39 VGND VPWR sky130_fd_sc_hd__fill_2
X_1077_ _1136_/A _1136_/B _1097_/B _1074_/C _1077_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__0572__A _0567_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1280__CLK _1159_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_104 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_56 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0747__A _0747_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_113 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_99 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_77 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_72 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_43 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_32 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_121 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0657__A _0611_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_143 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1153__CLK _1173_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1000_ _0960_/A _1000_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0674__A1 _0573_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_135 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0674__B2 _1195_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_3 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_clk_A clk VGND VPWR sky130_fd_sc_hd__diode_2
X_0715_ _0603_/X _1196_/Q _0712_/X _0713_/X _0714_/X _0715_/Y VGND VPWR sky130_fd_sc_hd__a2111oi_4
X_0646_ _0640_/Y _0646_/B _0646_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_106_17 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_9_0_clk_A clkbuf_3_4_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0577_ _0737_/D _0577_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_122_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_49 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_146 VGND VPWR sky130_fd_sc_hd__decap_4
X_1129_ _1106_/X _1090_/Y _1128_/X _1129_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1176__CLK _1172_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1283__D addr_r[9] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_53 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_71 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0924__B _1060_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_152 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_97 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1101__A _1058_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0959__A2 _0957_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0643__C _0624_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_185 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1081__A1 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_196 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1193__D d_sram_out[16] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_127 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0553__C _0552_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_171 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1072__A1 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0850__A _0859_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_16 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1199__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_127 VGND VPWR sky130_fd_sc_hd__fill_2
X_0629_ _0627_/Y _0628_/Y _0629_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_89_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0886__A1 _0870_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0728__C _1186_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_78 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1063__A1 _1050_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1278__D addr_r[4] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0810__B2 _0809_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0810__A1 _0804_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0760__A _0749_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_71 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0919__B _0919_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0935__A _1026_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0980_ _1240_/Q _0960_/X _0979_/X d_sram_in[12] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_80_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_160 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1188__D d_sram_out[11] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0670__A _1189_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0801__B2 _0800_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0801__A1 _0797_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_182 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_141 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0564__B _0568_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0580__A _0667_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_19 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_6_0_clk_A clkbuf_3_7_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_67 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1214__CLK _1252_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_44 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_101 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0649__B _0683_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_73 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0665__A _0660_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_177 VGND VPWR sky130_fd_sc_hd__fill_2
X_0963_ _1104_/A _1026_/A _0961_/X _0963_/D _0963_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_71_3 VGND VPWR sky130_fd_sc_hd__fill_1
X_0894_ _0874_/X _1174_/Q _0893_/Y d_fabric_out[29] VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1237__CLK _1252_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_17 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0575__A _0542_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_36 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_66 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_122 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_72 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_54 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_65 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_71 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1009__A1 _1257_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_86 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0651__C _0570_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_51 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0940__B1 _0939_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1231_ d_fabric_in[3] _0936_/D _1256_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_133 VGND VPWR sky130_fd_sc_hd__decap_3
X_1162_ _0737_/D _0866_/A _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1093_ _1030_/Y _1093_/B _1091_/X _1092_/Y _1093_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0946_ _0994_/B _0945_/Y d_sram_in[0] _0964_/A VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0877_ _0877_/A _0895_/B _0877_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_133_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_114 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_79 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_57 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0998__B1 _0939_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_45 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1286__D addr_r[12] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_3 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_171 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_3_0_clk_A clkbuf_2_3_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_93 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_133 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0927__B _0936_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_103 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1104__A _1104_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0943__A _0942_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0800_ _0556_/Y _0799_/Y _0745_/X _0800_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0731_ _0764_/A _0521_/X _0730_/X _0608_/C _0731_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__1196__D d_sram_out[19] VGND VPWR sky130_fd_sc_hd__diode_2
X_0662_ _1203_/Q _0662_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0593_ _0636_/B _0621_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_130_119 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0913__B1 _0986_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0837__B _0859_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1214_ _1214_/D _0546_/A _1252_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1145_ _0701_/Y _1145_/Q _1274_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1014__A _1057_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1076_ _1126_/B _1136_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_4_5_0_clk_A clkbuf_3_2_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0572__B _0742_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0929_ _0928_/Y _1026_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_136_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_119 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_79 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_147 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_40 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0763__A _0763_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_160 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_41 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0938__A _0937_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0657__B _0636_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0674__A2 _1161_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0714_ _0576_/X _0612_/A _0621_/C _0714_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_0645_ _0645_/A _0645_/B _0643_/Y _0644_/Y _0646_/B VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__1139__B1 _1138_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0576_ _0623_/A _0576_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0848__A _1157_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_174 VGND VPWR sky130_fd_sc_hd__decap_12
X_1128_ _1118_/A _1126_/Y _1137_/B _1128_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_15_26 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0583__A _0583_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1059_ _1057_/X _1059_/B _1018_/X _1097_/D _1059_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_40_139 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_163 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0758__A _0807_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_22 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_169 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_139 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_117 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_142 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1081__A2 _1074_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_197 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0668__A _0607_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1270__CLK _1166_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_1_0_0_clk_A clkbuf_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1072__A2 _1071_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0850__B _0859_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_93 VGND VPWR sky130_fd_sc_hd__fill_2
X_0628_ _0628_/A _0535_/A _0628_/C _0628_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_0559_ _1161_/D _0559_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_133_27 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0886__A2 _1170_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0740__D1 _0739_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_clk_A clkbuf_2_1_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_150 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1063__A2 _1049_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0810__A2 _0692_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_54 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0919__C _0921_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_76 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_13_0_clk_A clkbuf_3_6_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_93 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0935__B _0903_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0801__A2 _0692_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_175 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0564__C _0653_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1022__A _1095_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1166__CLK _1166_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0861__A _0861_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0580__B _0608_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_109 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0725__B1_N _0653_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1289__D conf[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_113 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_31 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0649__C _0551_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0665__B _0661_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_189 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1189__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1199__D d_sram_out[22] VGND VPWR sky130_fd_sc_hd__diode_2
X_0962_ _0921_/X _0961_/X _0988_/C d_sram_in[0] _0962_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_0893_ _0893_/A _0893_/B _0893_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_64_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1017__A _1102_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0856__A _0793_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_156 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0575__B _0628_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_15 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0777__A1 _0772_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_145 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_77 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1009__A2 _0915_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_65 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_7 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0940__A1 _0936_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1230_ d_fabric_in[2] _0927_/D _1256_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1161_ _1161_/D _1161_/Q _1173_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_123 VGND VPWR sky130_fd_sc_hd__fill_1
X_1092_ _1088_/A _1136_/B _1102_/B _1083_/B _1092_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_0945_ _0944_/Y _0945_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0876_ _0797_/Y _0775_/X _0875_/Y d_fabric_out[20] VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__1204__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_117 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_1_0_clk_A clkbuf_3_0_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0586__A _1174_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_104 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_137 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0998__A1 _1247_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_72 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_123 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0927__C _0988_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_156 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_126 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1104__B _1026_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1227__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0730_ _0729_/B _0730_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0661_ _0576_/X _1179_/Q _0718_/A _0661_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_115_139 VGND VPWR sky130_fd_sc_hd__fill_2
X_0592_ _0530_/A _0636_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0913__A1 _0994_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_3 VGND VPWR sky130_fd_sc_hd__fill_1
X_1213_ _1213_/D _0542_/A _1256_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0837__C _0859_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_145 VGND VPWR sky130_fd_sc_hd__fill_2
X_1144_ csb web _1144_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_1075_ _1075_/A _1136_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0928_ _0922_/C _0928_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0859_ _0859_/A _0859_/B _0859_/C _1208_/Q _0859_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_20_49 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_123 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0763__B _0762_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_23 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_3 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_67 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0840__B1 _0839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_82 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_71 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_175 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0657__C _1191_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_104 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1084__B1 _1080_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0792__A1_N _0872_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0713_ _0718_/A _0536_/X _0539_/X _1182_/Q _0713_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0644_ _0599_/Y _1179_/Q _0624_/C _0644_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__1139__A1 _1090_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0575_ _0542_/A _0628_/A _0623_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__0898__B1 _0897_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0848__B _0870_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_186 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_18 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1025__A _1022_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_104 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0864__A _0559_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1127_ _1057_/A _1127_/B _1127_/C _1137_/B VGND VPWR sky130_fd_sc_hd__or3_4
X_1058_ _1058_/A _1097_/D VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_31_26 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_175 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0774__A _0793_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_33 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1066__B1 _1063_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_143 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0813__B1 _0742_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_176 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_81 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_41 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_107 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0949__A _0949_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0668__B _0588_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_118 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0850__C _0859_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_29 VGND VPWR sky130_fd_sc_hd__fill_2
X_0627_ _0608_/A _0628_/A _0627_/C _0627_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__0859__A _0859_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0558_ _0607_/B _0558_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_173 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0740__C1 _0734_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_15 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_37 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0594__A _0588_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_22 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_11 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0935__C _0922_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_65 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_3_0_clk clkbuf_2_3_0_clk/A clkbuf_3_7_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_12_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_173 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0679__A _0677_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1022__B _1097_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0861__B _1160_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0580__C _1196_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0589__A _0589_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_165 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_79 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1008__B1_N _0979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_125 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1260__CLK _1274_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_72 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_83 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_54 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_110 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_102 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_31 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0665__C _0664_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0962__A _0921_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0961_ _0936_/A _0961_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0892_ _0874_/X _1173_/Q _0891_/X d_fabric_out[28] VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_57_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_154 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_113 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_168 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_18 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1033__A _1030_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0872__A _0872_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1283__CLK _1288_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0777__A2 _0775_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_24 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_82 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1118__A _1118_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_121 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_7 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0957__A _0960_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0940__A2 _0916_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_143 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1156__CLK _1173_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1160_ _1160_/D _1160_/Q _1173_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_113 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_102 VGND VPWR sky130_fd_sc_hd__fill_2
X_1091_ _1067_/Y _1106_/A _1091_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_64_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0692__A _0749_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0944_ _1023_/A _1126_/B _0944_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_0875_ _0875_/A _0874_/X _0875_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_118_115 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_129 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1028__A _1031_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_146 VGND VPWR sky130_fd_sc_hd__decap_4
X_1289_ conf[1] _0902_/A _1274_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_34_37 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0998__A2 _0984_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1179__CLK _1180_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0927__D _0927_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_179 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1104__C _1026_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_98 VGND VPWR sky130_fd_sc_hd__fill_2
X_0660_ _0656_/Y _0657_/Y _0660_/C _0659_/Y _0660_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_115_107 VGND VPWR sky130_fd_sc_hd__fill_2
X_0591_ _0893_/A _0588_/Y _0589_/Y _0590_/Y _0591_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__0913__A2 _0994_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0687__A _0698_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1212_ _1212_/D _0518_/A _1252_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0837__D _1203_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1143_ _1102_/Y _1132_/A _1141_/X w_mask[31] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_52_105 VGND VPWR sky130_fd_sc_hd__decap_8
X_1074_ _1057_/X _1059_/B _1074_/C _1073_/X _1074_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_52_127 VGND VPWR sky130_fd_sc_hd__decap_12
X_0927_ _1104_/A _0936_/A _0988_/C _0927_/D _0986_/C VGND VPWR sky130_fd_sc_hd__nand4_4
X_0858_ _0705_/X _1159_/D _0857_/X d_fabric_out[14] VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_20_39 VGND VPWR sky130_fd_sc_hd__fill_2
X_0789_ _0779_/Y _0533_/X _0564_/Y _0789_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_136_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0678__B1_N _0653_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0597__A _0588_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_168 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0763__C _0763_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_182 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_86 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0840__A1 _0794_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_3 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_87 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_102 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_127 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_116 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_80 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1084__A1 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0712_ _0718_/A _0536_/X _0550_/X _1184_/Q _0712_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0643_ _0623_/A _1178_/Q _0624_/C _0643_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__1139__A2 _1132_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0574_ _0573_/Y _0574_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0898__A1 _0874_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_154 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1025__B _1024_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1126_ _1136_/A _1126_/B _1097_/B _1136_/D _1126_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_25_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0864__B _0895_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1057_ _1057_/A _1057_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_33_182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_38 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1217__CLK _1253_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_23 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1066__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_133 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0813__A1 _0628_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_166 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_93 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_64 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0668__C _0589_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1126__A _1136_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_130 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_clk clk clkbuf_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_87_3 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0850__D _1174_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0626_ _0626_/A _0623_/Y _0626_/C _0625_/Y _0634_/A VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__0859__B _0859_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0557_ _0535_/A _0607_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1036__A _1025_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0875__A _0875_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0740__B1 _0732_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1109_ _1057_/A _1109_/B _1060_/B _1118_/B VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_21_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_45 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_71 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0798__B1 _0742_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0970__B1 _0969_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0679__B _0679_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_100 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0695__A _0695_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1022__C _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0789__B1 _0564_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0609_ _0609_/A _0608_/B _0786_/A _0609_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_85_111 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_122 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_40 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0952__B1 _0951_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_125 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0962__B _0961_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0960_ _0960_/A _0960_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0891_ _1173_/D _0883_/B _0891_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_4_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_111 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_188 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1033__B _1033_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1120__B1 _1119_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_180 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0872__B _0889_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_14 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_2_0_clk clkbuf_2_3_0_clk/A clkbuf_3_5_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_48_36 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_20 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_31 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_46 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1111__B1 _1110_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_180 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_30 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_23 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_96 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_43 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_87 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1118__B _1118_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_158 VGND VPWR sky130_fd_sc_hd__fill_2
X_1090_ _1057_/X _1059_/B _1073_/X _1097_/D _1090_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_118_105 VGND VPWR sky130_fd_sc_hd__fill_2
X_0943_ _0942_/X _1126_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0874_ _0871_/A _0874_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_118_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1044__A _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1250__CLK _1253_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1288_ conf[0] _0914_/A _1288_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0883__A _0883_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_41 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_45 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_103 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1104__D _1037_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0793__A _0793_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_88 VGND VPWR sky130_fd_sc_hd__fill_2
X_0590_ _0607_/B _0607_/A _0590_/C _0588_/D _0590_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__1273__CLK _1274_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1211_ _1219_/Q _0570_/A _1177_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_114 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_125 VGND VPWR sky130_fd_sc_hd__fill_2
X_1142_ _1097_/Y _1132_/X _1141_/X w_mask[30] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_1073_ _1102_/C _1073_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_52_139 VGND VPWR sky130_fd_sc_hd__decap_12
X_0926_ _0922_/B _0936_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0857_ _0857_/A _0871_/A _0857_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_106_119 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1039__A _1057_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0788_ _0682_/X _0822_/A _0551_/B _0786_/Y _0787_/Y _0788_/Y VGND VPWR sky130_fd_sc_hd__o41ai_4
XANTENNA__0597__B _0597_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_43 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_161 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0840__A2 _1155_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1146__CLK _1177_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_155 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_147 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_93 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_139 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1084__A2 _1083_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0711_ _0709_/X _0595_/Y _0711_/C _0711_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_0642_ _0635_/A _0599_/Y _1187_/Q _0645_/B VGND VPWR sky130_fd_sc_hd__nand3_4
X_0573_ _0535_/A _0573_/B _0573_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__0698__A _0698_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_122 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0898__A2 _1176_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1125_ _1071_/Y _1121_/X _1123_/X w_mask[23] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_1056_ _1044_/X _1055_/Y _1052_/X w_mask[3] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_33_161 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1169__CLK _1172_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0909_ _0914_/A _0903_/X _0909_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_102_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_31 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_68 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1066__A2 _1065_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_134 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0813__A2 _0692_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_167 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_32 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1126__B _1126_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_80 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0974__A1_N _0934_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_183 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_153 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0625_ _0622_/Y _1189_/Q _0573_/Y _0625_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__0859__C _0859_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0556_ _0555_/Y _0556_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1036__B _1027_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0740__A1 _1182_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0875__B _0874_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1108_ _1095_/A _1136_/B _1097_/B _1136_/D _1108_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__0891__A _1173_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1202__D d_sram_out[25] VGND VPWR sky130_fd_sc_hd__diode_2
X_1039_ _1057_/A _1018_/A _1020_/Y _1109_/B _1039_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_21_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_153 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_97 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_63 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0798__A1 _0627_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0970__A1 _1237_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1137__A _1118_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_186 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1022__D _1074_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0789__A1 _0779_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1207__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1047__A _1127_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0608_ _0608_/A _0608_/B _0608_/C _0608_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_0539_ _0607_/A _0539_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_134 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_27 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_59 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_30 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_23 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0952__A1 _0949_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_78 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_11 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_73 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0962__C _0988_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0890_ _0874_/X _1172_/Q _0889_/Y d_fabric_out[27] VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_138_180 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_31 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_148 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1120__A1 _1059_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0618__A2_N _0615_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_126 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_69 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1111__A1 _1106_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_55 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1118__C _1117_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_91 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0613__B1 _0612_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0942_ _0922_/B _0914_/A _0902_/A _0942_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_0873_ _0870_/X _1164_/Q _0872_/Y d_fabric_out[19] VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_62_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1287_ addr_r[13] _1224_/D _1253_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0883__B _0883_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1060__A _1060_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1210__D _1218_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_49 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0604__B1 _0603_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1096__B1 _1093_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_71 VGND VPWR sky130_fd_sc_hd__fill_2
X_1210_ _1218_/Q _0653_/B _1218_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_1_32 VGND VPWR sky130_fd_sc_hd__decap_12
X_1141_ _1024_/X _1102_/Y _1137_/X _1141_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0984__A _0960_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1072_ _1070_/X _1071_/Y _1068_/X w_mask[7] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_52_118 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1087__B1 _1086_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_140 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0834__B1 _0833_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_151 VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_1_0_clk clkbuf_1_0_0_clk/X clkbuf_2_1_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_60_184 VGND VPWR sky130_fd_sc_hd__decap_6
X_0925_ _0924_/X _0925_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0856_ _0793_/A _0871_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_20_19 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1039__B _1018_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0787_ _0889_/A _0671_/Y _1184_/Q _0729_/Y _0787_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__1011__B1 _0990_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_175 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1055__A _1088_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_104 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1205__D d_sram_out[28] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0825__B1 _0823_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_142 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1002__B1 _0954_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_74 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_45 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_72 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1069__B1 _1068_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0816__B1 _0813_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_140 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_184 VGND VPWR sky130_fd_sc_hd__decap_6
X_0710_ _0763_/A _0600_/X _0597_/B _1190_/Q _0711_/C VGND VPWR sky130_fd_sc_hd__nand4_4
X_0641_ _0576_/X _0611_/A _1182_/Q _0645_/A VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__1240__CLK _1252_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0979__A _0964_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0572_ _0567_/Y _0742_/A _0572_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_111_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_3 VGND VPWR sky130_fd_sc_hd__fill_1
X_1124_ _1067_/Y _1121_/X _1123_/X w_mask[22] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_1055_ _1088_/A _1018_/X _1083_/B _1102_/B _1055_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_0908_ d_sram_in[0] _0910_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_0839_ _0883_/B _0839_/B _0839_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0889__A _0889_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_145 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_36 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_124 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_173 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_157 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1263__CLK _1166_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1126__C _1097_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_4 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_97 VGND VPWR sky130_fd_sc_hd__fill_2
X_0624_ _0621_/B _0624_/B _0624_/C _0626_/C VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__0859__D _1208_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0555_ _0667_/B _0520_/X _1173_/D _0555_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__1036__C _1036_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0740__A2 _0729_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1107_ _1136_/C _0919_/Y _1029_/X _1118_/A VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__1286__CLK _1253_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0891__B _0883_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1038_ _1082_/A _1109_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_21_187 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_14 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_87 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_58 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_62 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_110 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0798__A2 _0749_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_114 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1137__B _1137_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0970__A2 _0957_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1159__CLK _1159_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_146 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_80 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_91 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0992__A _0909_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0789__A2 _0533_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0607_ _0607_/A _0607_/B _0607_/C _0607_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_0538_ _0628_/A _0607_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_157 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1213__D _1213_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0937__C1 _0911_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_46 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0952__A2 _0916_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0676__B1_N _0621_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_85 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_67 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0962__D d_sram_in[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_93 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_172 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_116 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1120__A2 _1105_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0772__A2_N _0693_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1058__A _1058_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0897__A _0897_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1208__D d_sram_out[31] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0787__A2_N _0671_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_135 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_149 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_66 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_15 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1111__A2 _1074_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_87 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_69 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_85 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1032__D1 _1060_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0600__A _0599_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_146 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_138 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_182 VGND VPWR sky130_fd_sc_hd__fill_1
X_0941_ _0920_/Y _1060_/B _0941_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__0613__A1 _0606_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0872_ _0872_/A _0889_/B _0872_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_118_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_3 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_138 VGND VPWR sky130_fd_sc_hd__fill_2
X_1286_ addr_r[12] _1286_/Q _1253_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_63_182 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1060__B _1060_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0604__A1 _1169_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0604__B2 _0747_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_173 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_76 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1096__A1 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_68 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_94 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_1140_ _1095_/Y _1132_/X _1138_/X w_mask[29] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_1_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_149 VGND VPWR sky130_fd_sc_hd__fill_2
X_1071_ _1075_/A _1018_/A _1109_/B _1058_/A _1071_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__1087__A1 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_182 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0834__A1 _0724_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0924_ _0920_/Y _1060_/B _0924_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0855_ _0762_/Y _0750_/X _0854_/Y _1159_/D VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__1039__C _1020_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0786_ _0786_/A _0786_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1011__A1 _1259_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1055__B _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0770__B1 _0769_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1071__A _1075_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1269_ addr_w[9] _1082_/A _1274_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_43_108 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1221__D _1284_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0825__A1 _0786_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0825__B2 _0824_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_31 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1002__A1 _1250_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_13 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_154 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_75 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0761__B1 _0760_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_57 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1192__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_51 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1069__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0816__B2 _0815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_60 VGND VPWR sky130_fd_sc_hd__fill_2
X_0640_ _0640_/A _0636_/Y _0639_/Y _0640_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__0979__B _0977_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0571_ _0745_/A _0742_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_111_113 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0995__A _0909_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0752__B1 _0699_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1123_ _1106_/X _1088_/Y _1118_/X _1123_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_1054_ _1109_/B _1102_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0907_ _0919_/B _0922_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_0838_ _0768_/Y _0760_/X _0837_/Y _0839_/B VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0991__B1 _0990_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0889__B _0889_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0769_ _0768_/Y _0533_/X _0566_/A _0769_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_102_113 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0743__B1 _0742_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_157 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1216__D _1216_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_152 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_125 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1126__D _1136_/D VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_0_0_clk clkbuf_1_0_0_clk/X clkbuf_3_1_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_5 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_7 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_32 VGND VPWR sky130_fd_sc_hd__decap_12
X_0623_ _0623_/A _0622_/Y _1190_/Q _0623_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__0973__B1 _0972_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_100 VGND VPWR sky130_fd_sc_hd__fill_2
X_0554_ _0535_/A _0667_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_177 VGND VPWR sky130_fd_sc_hd__fill_2
X_1106_ _1106_/A _1106_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_1037_ _1037_/A _1037_/B _1037_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_21_111 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1141__B1 _1137_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_69 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1230__CLK _1256_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_52 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_73 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0603__A _0608_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0955__B1 _0954_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1137__C _1136_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0707__B1 _0706_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_114 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0992__B _0961_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_3 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0946__B1 d_sram_in[0] VGND VPWR sky130_fd_sc_hd__diode_2
X_0606_ _0544_/X _0606_/B _0606_/C _0606_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_0537_ _0518_/A _0628_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1253__CLK _1253_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1123__B1 _1118_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_180 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_129 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0937__B1 _0936_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_43 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_58 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_97 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1114__B1 _1110_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_73 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_151 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_55 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1276__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_128 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_172 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1041__C1 _1036_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0897__B _0893_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_103 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_39 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_28 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1074__A _1057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1224__D _1224_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_48 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1149__CLK _1159_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_35 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_97 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1032__C1 _1026_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_50 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_117 VGND VPWR sky130_fd_sc_hd__fill_1
X_0940_ _0936_/D _0916_/X _0939_/Y d_sram_in[3] VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0613__A2 _0607_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0871_ _0871_/A _0889_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_1285_ addr_r[11] _1222_/D _1253_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_63_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_29 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0604__A2 _0621_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1219__D _0919_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_185 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_111 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0701__A _0701_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_172 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1096__A2 _1095_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_111 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0611__A _0611_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_133 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_56 VGND VPWR sky130_fd_sc_hd__decap_12
X_1070_ _1043_/A _1070_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_45_161 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1087__A2 _1085_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0834__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_91 VGND VPWR sky130_fd_sc_hd__fill_1
X_0923_ _1127_/C _1060_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0854_ _0846_/A _0846_/B _0846_/C _0589_/A _0854_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_0785_ _0730_/X _0574_/X _1196_/Q _0531_/Y _0637_/B _0785_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__1039__D _1109_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0521__A _0520_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1011__A2 _0915_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0770__A1 _0533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_19 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1055__C _1083_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1071__B _1018_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1268_ addr_w[8] baseaddr_w_sync[8] _1274_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1199_ d_sram_out[22] _0607_/C _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0825__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_186 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1002__A2 _1000_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0761__A1 _0579_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_114 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_63 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_139 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1069__A2 _1067_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_84 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0606__A _0544_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0979__C _0979_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0570_ _0570_/A _0570_/B _0698_/A _0745_/A VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0752__A1 _0743_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0995__B _0961_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_80 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_91 VGND VPWR sky130_fd_sc_hd__fill_2
X_1122_ _1065_/Y _1121_/X _1119_/X w_mask[21] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_1053_ _1044_/X _1049_/Y _1052_/X w_mask[2] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_33_131 VGND VPWR sky130_fd_sc_hd__fill_2
X_0906_ _1104_/A _0988_/C _1026_/C _0994_/B VGND VPWR sky130_fd_sc_hd__o21a_4
X_0837_ _0859_/A _0859_/B _0859_/C _1203_/Q _0837_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__0991__A1 _1243_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0768_ _1187_/Q _0768_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0699_ _0846_/B _0846_/A _0846_/C _0577_/X _0699_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0743__A1 _0727_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1082__A _1082_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1232__D d_fabric_in[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_27 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_115 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_180 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_6 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_134 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_156 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0973__A1 _1238_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0622_ _0617_/C _0622_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0553_ _0541_/Y _0551_/Y _0552_/Y _0553_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__0725__A1 _0724_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_189 VGND VPWR sky130_fd_sc_hd__fill_1
X_1105_ _1132_/A _1105_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_1036_ _1025_/Y _1027_/Y _1036_/C w_mask[0] VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_42_19 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1182__CLK _1180_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1077__A _1136_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_123 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1227__D _1227_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_49 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_22 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1141__A1 _1024_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0652__B1 _0651_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_41 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_85 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0603__B _0615_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0955__A1 _1234_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0707__A1 _0704_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_167 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0992__C _0992_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_3 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_182 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0946__A1 _0994_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0605_ _0628_/A _0606_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0536_ _0609_/A _0536_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_115 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_126 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_148 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1123__A1 _1106_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0882__B1 _0881_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1019_ _1019_/A _1058_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0704__A _0826_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_11 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0937__A1 _0899_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_66 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_14 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_36 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1114__A1 _1106_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_85 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0873__B1 _0872_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0614__A _1172_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_80 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_91 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0524__A _0588_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1041__B1 _1025_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1004__B1_N _0964_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1220__CLK _1253_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_115 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_18 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1074__B _1059_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0519_ _0573_/B _0588_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_73_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_57 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1090__A _1057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0855__B1 _0854_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_34 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1240__D d_fabric_in[12] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_76 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_87 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_58 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1032__B1 _0928_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0791__C1 _0790_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0609__A _0609_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_83 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1150__D _0811_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0870_ _0870_/A _0870_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_118_109 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_71 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0613__A3 _0608_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1243__CLK _1288_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1284_ addr_r[10] _1284_/Q _1253_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0519__A _0573_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0604__A3 _0574_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0999_ _1248_/Q _0984_/X _0947_/X d_sram_in[20] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_117_142 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1085__A _1088_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1235__D d_fabric_in[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_77 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_20 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1266__CLK _1274_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_86 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1005__B1 _0969_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_145 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1145__D _0701_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_81 VGND VPWR sky130_fd_sc_hd__fill_2
X_0922_ _0921_/X _0922_/B _0922_/C _1127_/C VGND VPWR sky130_fd_sc_hd__nand3_4
X_0853_ _0843_/X _1158_/Q _0852_/X d_fabric_out[13] VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_60_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0802__A _0802_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0784_ _0783_/Y _0784_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_114_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_123 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1055__D _1102_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0770__A2 _0763_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_107 VGND VPWR sky130_fd_sc_hd__decap_4
X_1267_ addr_w[7] baseaddr_w_sync[7] _1274_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1289__CLK _1274_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1071__C _1109_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1198_ d_sram_out[21] _0608_/C _1208_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_51_121 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_36 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_154 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_9 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0712__A _0718_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_112 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_137 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0761__A2 _0745_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_52 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_165 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0606__B _0606_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0622__A _0617_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_7 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0971__A1_N _0917_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0752__A2 _0751_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0995__C _1245_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1121_ _1132_/A _1121_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_1052_ _1050_/X _1051_/Y _1034_/X _1052_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_18_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_165 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0673__D1 _0672_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0905_ _0919_/B _1026_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0532__A _0520_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0836_ _0705_/X _1154_/D _0835_/X d_fabric_out[9] VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0991__A2 _0984_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0767_ _0682_/X _0822_/A _0551_/B _0663_/Y _0766_/Y _0767_/Y VGND VPWR sky130_fd_sc_hd__o41ai_4
X_0698_ _0698_/A _0846_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0743__A2 _0741_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_79 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_121 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_84 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_121 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0617__A _0609_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_50 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_56 VGND VPWR sky130_fd_sc_hd__decap_12
X_0621_ _0621_/A _0621_/B _0621_/C _0626_/A VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__0973__A2 _0957_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0552_ _0764_/A _0550_/X _0528_/X _0606_/C _0552_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__0725__A2 _0666_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_1104_ _1104_/A _1026_/A _1026_/C _1037_/A _1132_/A VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__0527__A _0807_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1035_ _1034_/X _1036_/C VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_21_102 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_179 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_157 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_146 VGND VPWR sky130_fd_sc_hd__decap_4
X_0819_ _0637_/B _0819_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1077__B _1136_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1093__A _1030_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1243__D d_fabric_in[15] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_45 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1141__A2 _1102_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0816__A1_N _0607_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0652__A1 _0620_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_97 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0603__C _0588_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0955__A2 _0916_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0900__A _0914_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0707__A2 _0701_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1153__D _0831_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_161 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0946__A2 _0945_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0604_ _1169_/D _0621_/A _0574_/X _0603_/X _0747_/A _0604_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
X_0535_ _0535_/A _0609_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1123__A2 _1088_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0882__A1 _0870_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1018_ _1018_/A _1018_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1088__A _1088_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0937__A2 _1023_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1238__D d_fabric_in[10] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_127 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1114__A2 _1083_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_171 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0873__A1 _0870_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_41 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1148__D _1148_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0630__A _0629_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_116 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0561__B1 _0763_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1172__CLK _1172_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0805__A _1190_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1041__A1 _1037_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0540__A _1169_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0518_ _0518_/A _0573_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1074__C _1074_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1090__B _1059_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0855__A1 _0762_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_79 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_99 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1032__A1 _1026_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0791__B1 _0745_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1195__CLK _1208_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_85 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0609__B _0608_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_182 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_62 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0625__A _0622_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0613__A4 _0609_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_7 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_165 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0965__B1_N _0964_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0782__B1 _0692_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1283_ addr_r[9] _1220_/D _1288_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0535__A _0535_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0998_ _1247_/Q _0984_/X _0939_/Y d_sram_in[19] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_117_121 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1085__B _1059_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_24 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_46 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_68 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_12 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_182 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1251__D d_fabric_in[23] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_89 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1005__A1 _1253_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_83 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_72 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1161__D _1161_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1210__CLK _1218_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_144 VGND VPWR sky130_fd_sc_hd__fill_2
X_0921_ _0921_/A _0921_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0852_ _0861_/A _1158_/D _0852_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_0783_ _0536_/X _0521_/X _0730_/X _1208_/Q _0783_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__0802__B _0893_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0755__B1 _0754_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0770__A3 _0765_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1266_ addr_w[6] baseaddr_w_sync[6] _1274_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_36_141 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1071__D _1058_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1197_ d_sram_out[20] _0606_/C _1208_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0712__B _0536_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_8 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0746__B1 _0745_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_146 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_45 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1246__D d_fabric_in[18] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_16 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_78 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0761__A3 _0757_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_49 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_149 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_76 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1233__CLK _1288_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_97 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0606__C _0606_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_30 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0903__A _0922_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0985__B1 _1242_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1156__D _1156_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_149 VGND VPWR sky130_fd_sc_hd__fill_2
X_1120_ _1059_/Y _1105_/X _1119_/X w_mask[20] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_18_152 VGND VPWR sky130_fd_sc_hd__decap_4
X_1051_ _1051_/A _1051_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0968__A2_N _0966_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0673__C1 _0669_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_92 VGND VPWR sky130_fd_sc_hd__fill_2
X_0904_ _0903_/X _0988_/C VGND VPWR sky130_fd_sc_hd__buf_1
X_0835_ _1154_/Q _0870_/A _0835_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0976__B1 _0975_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0532__B _0528_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0766_ _0662_/Y _0671_/Y _0628_/C _0729_/Y _0766_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
X_0697_ _0807_/B _0846_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1256__CLK _1256_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_182 VGND VPWR sky130_fd_sc_hd__fill_1
X_1249_ d_fabric_in[21] _1249_/Q _1253_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0796__B1_N _0795_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_106 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0723__A _0711_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_44 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_37 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_99 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_96 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0617__B _0608_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_8 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_114 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0633__A _0630_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0958__B1 _0937_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_68 VGND VPWR sky130_fd_sc_hd__decap_12
X_0620_ _0585_/Y _0602_/Y _0619_/Y _0620_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_0551_ _0764_/A _0551_/B _0550_/X _0627_/C _0551_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__1279__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_125 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1135__B1 _1133_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_3 VGND VPWR sky130_fd_sc_hd__fill_1
X_1103_ _1043_/X _1102_/Y _1099_/X w_mask[15] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_1034_ _1033_/X _1034_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0527__B _1185_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_136 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_8_0_clk_A clkbuf_3_4_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0543__A _0543_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0818_ _0816_/Y _0794_/X _0817_/Y d_fabric_out[6] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__1077__C _1097_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0749_ _0749_/A _0749_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_88_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_47 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_18 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1093__B _1093_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0718__A _0718_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_77 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0652__A2 _0650_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_54 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0985__A1_N _0953_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0603__D _0594_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_84 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0628__A _0628_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_7 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0603_ _0608_/A _0615_/B _0588_/B _0594_/X _0603_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0534_ _0542_/A _0535_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_93_172 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0538__A _0628_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0882__A2 _1168_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1017_ _1102_/C _1018_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1088__B _1083_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_57 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1254__D d_fabric_in[26] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_32 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0873__A2 _1164_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0911__A _0911_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0630__B _0612_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_50 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1164__D _1196_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0561__A1 _0556_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_109 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_183 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_3 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1041__A2 _1051_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0517_ reb csb _1227_/D VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1074__D _1073_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1090__C _1073_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0855__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1099__A _1030_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1249__D d_fabric_in[21] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_78 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_5_0_clk_A clkbuf_3_5_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0731__A _0764_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_89 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1032__A2 _1019_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0791__A1 _0624_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_139 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_75 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0609__C _0786_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0625__B _1189_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1159__D _1159_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0641__A _0576_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_177 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0782__A1 _0780_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_93 VGND VPWR sky130_fd_sc_hd__fill_2
X_1282_ addr_r[8] baseaddr_r_sync[8] _1159_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_48_161 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_186 VGND VPWR sky130_fd_sc_hd__decap_4
X_0997_ _1246_/Q _0984_/X _0932_/Y d_sram_in[18] VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0551__A _0764_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_19 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1085__C _1074_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_11 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_111 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1162__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1005__A2 _1000_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_112 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_186 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0636__A _0612_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_0920_ _0919_/Y _0920_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0851_ _0805_/Y _0749_/X _0850_/Y _1158_/D VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0782_ _0780_/X _0781_/Y _0692_/X _0782_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__0755__A1 _0704_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_3 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0770__A4 _0767_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1265_ addr_w[5] baseaddr_w_sync[5] _1166_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_36_131 VGND VPWR sky130_fd_sc_hd__fill_2
X_1196_ d_sram_out[19] _1196_/Q _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_36_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0546__A _0546_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_145 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1185__CLK _1184_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0712__C _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0746__A1 _0822_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0761__A4 _0759_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_11 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1262__D addr_w[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_32 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_10 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_86 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_75 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_64 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0985__B2 _0919_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_2_0_clk_A clkbuf_2_3_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1172__D _1172_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1050_ _1024_/X _1050_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_18_175 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_145 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0673__B1 _0666_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0903_ _0922_/C _0903_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0834_ _0724_/Y _0750_/X _0833_/Y _1154_/D VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0976__A1 _1239_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0765_ _0551_/B _0668_/Y _0764_/Y _0765_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0696_ _0859_/B _0846_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_102_117 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_4_0_clk_A clkbuf_3_2_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1248_ d_fabric_in[20] _1248_/Q _1253_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_24_123 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0664__B1 _0663_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_107 VGND VPWR sky130_fd_sc_hd__decap_3
X_1179_ d_sram_out[2] _1179_/Q _1180_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_24_156 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_129 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0723__B _0715_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_89 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1257__D d_fabric_in[29] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_27 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1200__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_112 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0655__B1 _0654_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0617__C _0617_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_126 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_104 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_189 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0914__A _0914_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0633__B _0633_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0958__A1 _0988_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1080__B1 _1079_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1167__D _0607_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0550_ _0608_/B _0550_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_104 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1135__A1 _1088_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0894__B1 _0893_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1102_ _1136_/A _1102_/B _1102_/C _1136_/D _1102_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_1033_ _1030_/Y _1033_/B _1033_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0527__C _0763_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_115 VGND VPWR sky130_fd_sc_hd__fill_2
X_0817_ _0826_/A _1151_/Q _0817_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__1223__CLK _1253_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1077__D _1074_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0748_ _0747_/Y _0763_/C _0577_/X _0600_/X _0748_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
X_0679_ _0677_/Y _0679_/B _0679_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_107_59 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1093__C _1091_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0718__B _0544_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_89 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0734__A _0822_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_126 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_159 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0909__A _0914_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0876__B1 _0875_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0628__B _0535_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0644__A _0599_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1246__CLK _1288_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_170 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1053__B1 _1052_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0800__B1 _0745_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0602_ _0602_/A _0591_/X _0595_/Y _0601_/Y _0602_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_0533_ _0533_/A _0533_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0819__A _0637_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0867__B1 _0866_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_184 VGND VPWR sky130_fd_sc_hd__decap_6
X_1016_ _1031_/B _1097_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0554__A _0535_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1088__C _1136_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_36 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_13 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0729__A _0558_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_clk_A clkbuf_3_1_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0858__B1 _0857_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_66 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1270__D addr_w[10] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1269__CLK _1274_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12_0_clk_A clkbuf_3_6_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_91 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_62 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0639__A _0621_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0561__A2 _0560_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0849__B1 _0848_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1180__D d_sram_out[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_176 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_3 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0549__A _0573_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_16 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1090__D _1097_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_154 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_176 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1099__B _1093_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_68 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_39 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0731__B _0521_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0791__A2 _0566_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1265__D addr_w[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_21 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_54 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_97 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0625__C _0573_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0922__A _0921_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_96 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0641__B _0611_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1175__D _0589_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0782__A2 _0781_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180 VGND VPWR sky130_fd_sc_hd__decap_6
X_1281_ addr_r[7] baseaddr_r_sync[7] _1159_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_48_140 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_121 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_101 VGND VPWR sky130_fd_sc_hd__fill_2
X_0996_ _0996_/A _0986_/A _0996_/C d_sram_in[17] VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_117_134 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0551__B _0551_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_189 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1085__D _1073_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_176 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_45 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0742__A _0742_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_167 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_115 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_64 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0917__A _0927_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_102 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_165 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0636__B _0636_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_73 VGND VPWR sky130_fd_sc_hd__fill_2
X_0850_ _0859_/A _0859_/B _0859_/C _1174_/D _0850_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_0781_ _0889_/A _0763_/C _1196_/Q _0600_/X _0781_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__0755__A2 _0752_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_148 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_3 VGND VPWR sky130_fd_sc_hd__fill_1
X_1264_ addr_w[4] baseaddr_w_sync[4] _1166_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_36_121 VGND VPWR sky130_fd_sc_hd__fill_1
X_1195_ d_sram_out[18] _1195_/Q _1208_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_51_102 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_0_0_clk_A clkbuf_3_0_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0979_ _0964_/A _0977_/Y _0979_/C _0979_/X VGND VPWR sky130_fd_sc_hd__and3_4
XANTENNA__0712__D _1184_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0746__A2 _0724_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0737__A _0544_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_113 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_51 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_62 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_95 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0647__A _0634_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_135 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0673__A1 _0617_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_83 VGND VPWR sky130_fd_sc_hd__decap_3
X_0902_ _0902_/A _0922_/C VGND VPWR sky130_fd_sc_hd__buf_1
X_0833_ _0846_/A _0846_/B _0846_/C _0747_/A _0833_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__0976__A2 _0957_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0764_ _0764_/A _0822_/A _0730_/X _1195_/Q _0764_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_0695_ _0695_/A _0859_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_110_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1152__CLK _1173_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0557__A _0535_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1247_ d_fabric_in[19] _1247_/Q _1288_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_112_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_1178_ d_sram_out[1] _1178_/Q _1180_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_24_113 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0664__A1 _0662_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0664__B2 _0615_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_119 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0723__C _0719_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1273__D addr_w[13] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_76 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0655__A1 _1177_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_82 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_31 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0914__B _0922_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_149 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1080__A1 _1050_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0958__A2 _0941_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0633__C _0632_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0930__A _0921_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_7 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0591__B1 _0589_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1183__D d_sram_out[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_83 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1175__CLK _1173_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1135__A2 _1132_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0894__A1 _0874_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1101_ _1058_/A _1136_/D VGND VPWR sky130_fd_sc_hd__buf_1
X_1032_ _1026_/B _1019_/A _0928_/Y _1026_/C _1060_/A _1033_/B VGND VPWR sky130_fd_sc_hd__a2111o_4
X_0816_ _0607_/C _0693_/Y _0813_/Y _0815_/X _0816_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
X_0747_ _0747_/A _0747_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_107_27 VGND VPWR sky130_fd_sc_hd__fill_2
X_0678_ _0683_/B _0666_/Y _0653_/Y _0679_/B VGND VPWR sky130_fd_sc_hd__a21boi_4
XFILLER_88_127 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1093__D _1092_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_26 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0718__C _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0734__B _0536_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1268__D addr_w[8] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0750__A _0749_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1198__CLK _1208_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0909__B _0903_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_182 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0876__A1 _0797_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0628__C _0628_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_63 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0925__A _0924_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0644__B _1179_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1053__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1178__D d_sram_out[1] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0660__A _0656_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0800__A1 _0556_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0601_ _0621_/A _0600_/X _1203_/Q _0601_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_0532_ _0520_/X _0528_/X _0533_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_21_3 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0867__A1 _0577_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0835__A _1154_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1015_ _1082_/A _1031_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1088__D _1073_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0570__A _0570_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_25 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_47 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0729__B _0729_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0858__A1 _0705_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_89 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0745__A _0745_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_66 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_187 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_74 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0849__A1 _0705_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0639__B _0638_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1213__CLK _1256_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_95 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0785__B1 _0531_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_174 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0565__A _0564_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_188 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1099__C _1098_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0731__C _0730_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_108 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_11 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1236__CLK _1256_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_130 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1281__D addr_r[7] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0700__B1 _0699_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_82 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_31 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1008__A1 _1256_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0922__B _0922_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0641__C _1182_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0767__B1 _0766_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_40 VGND VPWR sky130_fd_sc_hd__fill_2
X_1280_ addr_r[6] baseaddr_r_sync[6] _1159_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1191__D d_sram_out[14] VGND VPWR sky130_fd_sc_hd__diode_2
X_0995_ _0909_/Y _0961_/X _1245_/Q _0996_/C VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__0551__C _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1259__CLK _1177_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_19 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_155 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_57 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0997__B1 _0932_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_45 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1276__D addr_r[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_93 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_111 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0636__C _1184_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_85 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_96 VGND VPWR sky130_fd_sc_hd__fill_2
X_0780_ _0822_/B _0779_/Y _0745_/A _0780_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_60_7 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1186__D d_sram_out[9] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_116 VGND VPWR sky130_fd_sc_hd__decap_6
X_1263_ addr_w[3] baseaddr_w_sync[3] _1166_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1194_ d_sram_out[17] _0737_/D _1184_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_51_114 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0843__A _0870_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0978_ _1104_/A _1026_/A _0936_/A _1240_/Q _0979_/C VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_10_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_182 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0737__B _0606_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0753__A _0752_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_119 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0928__A _0922_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0720__A2_N _0588_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_85 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0647__B _0646_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0673__A2 _0883_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0663__A _0607_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0901_ _1026_/B _1104_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0832_ _0794_/X _1153_/Q _0831_/X d_fabric_out[8] VGND VPWR sky130_fd_sc_hd__o21a_4
X_0763_ _0763_/A _0762_/Y _0763_/C _0763_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_0694_ _0691_/A _0568_/A _0695_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_51_3 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1138__B1 _1137_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_130 VGND VPWR sky130_fd_sc_hd__decap_4
X_1246_ d_fabric_in[18] _1246_/Q _1288_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1177_ d_sram_out[0] _1177_/Q _1177_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0664__A2 _0588_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0573__A _0535_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_109 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_180 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0723__D _0722_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_8 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_69 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1129__B1 _1128_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_55 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_125 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0655__A2 _0651_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_54 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0914__C _0919_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_76 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1080__A2 _1059_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0930__B _1026_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_80 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0591__B2 _0590_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0591__A1 _0893_/A VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_9_0_clk clkbuf_3_4_0_clk/X _1163_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_87_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0658__A _0599_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1100_ _1043_/X _1097_/Y _1099_/X w_mask[14] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0894__A2 _1174_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1031_ _1013_/A _1031_/B _1060_/A VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_99_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_180 VGND VPWR sky130_fd_sc_hd__decap_3
X_0815_ _0814_/X _0607_/Y _0742_/X _0815_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_0746_ _0822_/B _0724_/Y _0745_/X _0746_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_107_39 VGND VPWR sky130_fd_sc_hd__fill_2
X_0677_ _0677_/A _0673_/Y _0677_/C _0677_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__0568__A _0568_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0718__D _0624_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1229_ d_fabric_in[1] _0899_/A _1256_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0734__C _0730_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_46 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1284__D addr_r[10] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_21 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_87 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_76 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0876__A2 _0775_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_98 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1102__A _1136_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0644__C _0624_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_150 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0941__A _0920_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1053__A2 _1049_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_165 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_154 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0800__A2 _0799_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0660__B _0657_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0600_ _0599_/Y _0600_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0531_ _0528_/X _0763_/C _0531_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__1194__D d_sram_out[17] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_83 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_150 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0867__A2 _0704_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0835__B _0870_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1014_ _1057_/A _1095_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1012__A _1270_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0570__B _0570_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0729_ _0558_/X _0729_/B _0606_/B _0729_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_134_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_183 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0858__A2 _1159_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0729__C _0606_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_45 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1279__D addr_r[5] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1165__CLK _1159_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_135 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_168 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0849__A2 _1157_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0639__C _0590_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_123 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0936__A _0936_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_7 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1189__D d_sram_out[12] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_270 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0671__A _0607_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0785__B2 _0637_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0785__A1 _0730_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_142 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0846__A _0846_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_123 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_145 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1188__CLK _1184_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1099__D _1092_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_15 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0581__A _0579_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_26 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0731__D _0608_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_186 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0756__A _1195_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0700__A1 _0690_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_55 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_44 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1008__A2 _0960_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0922__C _0922_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0767__A1 _0682_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_153 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0666__A _0667_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_3 VGND VPWR sky130_fd_sc_hd__fill_1
X_0994_ _0994_/A _0994_/B _0960_/A _0996_/A VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_117_114 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0551__D _0627_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_28 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_186 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0576__A _0623_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_27 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0997__A1 _1246_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_147 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_57 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1203__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_61 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_93 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_159 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1110__A _1118_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_7 VGND VPWR sky130_fd_sc_hd__fill_2
X_1262_ addr_w[2] baseaddr_w_sync[2] _1274_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_36_123 VGND VPWR sky130_fd_sc_hd__decap_4
X_1193_ d_sram_out[16] _1161_/D _1184_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_51_137 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1020__A _1058_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1226__CLK _1208_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0977_ _0921_/X _0961_/X _0988_/C _0977_/D _0977_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_105_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_49 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_69 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_112 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0737__C _0729_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_46 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_12 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1287__D addr_r[13] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_109 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1105__A _1132_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_70 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_156 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_41 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_92 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0944__A _1023_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1249__CLK _1253_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__decap_3
X_0900_ _0914_/A _1026_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0831_ _0883_/B _0831_/B _0831_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__1197__D d_sram_out[20] VGND VPWR sky130_fd_sc_hd__diode_2
X_0762_ _1191_/Q _0762_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0693_ _0692_/X _0693_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_44_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1138__A1 _1024_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_164 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1015__A _1082_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1245_ d_fabric_in[17] _1245_/Q _1288_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1176_ _1208_/Q _1176_/Q _1172_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0854__A _0846_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0573__B _0573_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0821__B1 _0897_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_15 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_19 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1129__A1 _1106_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_131 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0888__B1 _0887_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0764__A _0764_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_118 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0930__C _1026_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_129 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0591__A2 _0588_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0658__B _0627_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1030_ _1127_/B _0919_/Y _1029_/X _1030_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_21_107 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1056__B1 _1052_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0814_ _0807_/A _0762_/Y _0668_/Y _0814_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0745_ _0745_/A _0745_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0676_ _0674_/Y _0675_/Y _0621_/A _0677_/C VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_88_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_151 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0781__A2_N _0763_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1228_ d_fabric_in[0] d_sram_in[0] _1256_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0584__A _0624_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1159_ _1159_/D _0857_/A _1159_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_12_118 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0734__D _0747_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_173 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_162 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0759__A _0822_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_11 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_32 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1102__B _1102_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0941__B _1060_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0660__C _0660_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0530_ _0530_/A _0763_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_154 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_176 VGND VPWR sky130_fd_sc_hd__fill_2
X_1013_ _1013_/A _1057_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1029__B1 _0914_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0570__C _0698_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0728_ _0807_/B _0763_/A _1186_/Q _0728_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_0659_ _0636_/B _0628_/C _0583_/A _0659_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__0579__A _0607_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_36 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_58 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_24 VGND VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_8_0_clk clkbuf_3_4_0_clk/X _1159_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_138_156 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_54 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_31 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0936__B _1026_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_101 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_260 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0671__B _0609_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0785__A2 _0574_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0846__B _0846_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1023__A _1023_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0581__B _0580_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_49 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0766__A1_N _0662_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0700__A2 _0693_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_23 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_40 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_11 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1282__CLK _1159_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_115 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0767__A2 _0822_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_159 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_86 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1108__A _1095_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_63 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0688__D1 _0859_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0666__B _0520_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_157 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0682__A _0558_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0993_ _0910_/B _0960_/X _0992_/Y d_sram_in[16] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_74_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1018__A _1018_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1155__CLK _1172_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0857__A _0857_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_154 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0592__A _0530_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0997__A2 _0984_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_56 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_124 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_77 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_65 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_81 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_70 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1110__B _1108_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1178__CLK _1180_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0677__A _0677_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1261_ addr_w[1] baseaddr_w_sync[1] _1166_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1192_ d_sram_out[15] _0637_/B _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_36_135 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0676__A1 _0674_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_149 VGND VPWR sky130_fd_sc_hd__fill_2
X_0976_ _1239_/Q _0957_/X _0975_/Y d_sram_in[11] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_10_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_26 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_15 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0587__A _0587_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0737__D _0737_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_14 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_24 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_94 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_60 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0944__B _1126_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1121__A _1132_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_91 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_91 VGND VPWR sky130_fd_sc_hd__fill_1
X_0830_ _0861_/A _0883_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0960__A _0960_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0761_ _0579_/Y _0745_/X _0757_/Y _0759_/Y _0760_/X _0761_/Y VGND VPWR sky130_fd_sc_hd__a41oi_4
X_0692_ _0749_/A _0692_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1138__A2 _1097_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_62 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_clk clkbuf_0_clk/X clkbuf_2_3_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1244_ d_fabric_in[16] _0992_/C _1253_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_110_176 VGND VPWR sky130_fd_sc_hd__decap_6
X_1175_ _0589_/A _1175_/Q _1173_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0854__B _0846_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1031__A _1013_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0870__A _0870_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0821__A1 _0807_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0821__B2 _0763_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_0959_ _0988_/D _0957_/X _0958_/X d_sram_in[7] VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1129__A2 _1090_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_182 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0888__A1 _0662_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_46 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_116 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0764__B _0822_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_149 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_96 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0812__A1 _0704_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0930__D d_sram_in[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_93 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0658__C _0624_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1216__CLK _1256_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_160 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1056__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0803__A1 _0704_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0813_ _0628_/C _0692_/X _0742_/X _0813_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0744_ _0682_/X _0822_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0567__B1 _0566_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0675_ _0539_/X _0558_/X _0606_/C _0675_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__1026__A _1026_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_18 VGND VPWR sky130_fd_sc_hd__fill_2
X_1227_ _1227_/D csb1_sync _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1158_ _1158_/D _1158_/Q _1173_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1089_ _1070_/X _1088_/Y _1086_/X w_mask[11] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_113_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_108 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1239__CLK _1252_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0759__B _0859_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0775__A _0870_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_51 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1102__C _1102_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_141 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_174 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_101 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_145 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0660__D _0659_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_30 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0721__B1 _0720_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0685__A _0682_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1012_ _1270_/Q _1013_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1029__A1 _0903_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0788__B1 _0787_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_94 VGND VPWR sky130_fd_sc_hd__fill_1
X_0727_ _0723_/Y _0725_/Y _0726_/X _0727_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_0658_ _0599_/Y _0627_/C _0624_/C _0660_/C VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__0981__A1_N _0949_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0579__B _0609_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0589_ _0589_/A _0589_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0595__A _0528_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_168 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_19 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_95 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_33 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0951__B1 _0950_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_111 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_50 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0936__C _0903_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_147 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_261 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0671__C _0590_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0785__A3 _1196_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_100 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0846__C _0846_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_19 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_105 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0748__A2_N _0763_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_129 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0933__B1 _0932_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_114 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_35 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_52 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_74 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_105 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0767__A3 _0551_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_83 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_65 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_171 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1108__B _1136_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_20 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0666__C _0594_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0688__C1 _0570_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0963__A _1104_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0992_ _0909_/Y _0961_/X _0992_/C _0992_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_117_105 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_138 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_73 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_19 VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_7_0_clk clkbuf_4_6_0_clk/A _1218_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_39_133 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0857__B _0871_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_166 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1034__A _1033_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_114 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0906__B1 _1026_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_68 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0783__A _0536_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_77 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1110__C _1118_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_130 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0677__B _0673_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1260_ addr_w[0] baseaddr_w_sync[0] _1274_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1191_ d_sram_out[14] _1191_/Q _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0676__A2 _0675_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0693__A _0692_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0975_ _0938_/Y _0974_/Y _0975_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__0868__A _0868_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1272__CLK _1180_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_26 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_36 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_172 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0778__A _1196_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_44 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_21 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_139 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_161 VGND VPWR sky130_fd_sc_hd__fill_2
X_0760_ _0749_/A _0760_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1145__CLK _1274_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0691_ _0691_/A _0698_/A _0521_/X _0570_/B _0749_/A VGND VPWR sky130_fd_sc_hd__and4_4
X_1243_ d_fabric_in[15] _1243_/Q _1288_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_2_74 VGND VPWR sky130_fd_sc_hd__decap_12
X_1174_ _1174_/D _1174_/Q _1173_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_24_117 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0854__C _0846_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1031__B _1031_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_172 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0821__A2 _0819_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0958_ _0988_/D _0941_/Y _0937_/X _0958_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0585__A1 _0578_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0889_ _0889_/A _0889_/B _0889_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__0598__A _0635_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0888__A2 _0775_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_20 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0764__C _0730_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_53 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_57 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1168__CLK _1172_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_3 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0812__A2 _1150_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_87 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1132__A _1132_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_172 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1056__A2 _1055_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0803__A2 _1149_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0812_ _0704_/X _1150_/Q _0811_/Y d_fabric_out[5] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0743_ _0727_/Y _0741_/X _0742_/X _0743_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0567__A1 _0527_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0674_ _0573_/Y _1161_/D _0576_/X _1195_/Q _0674_/Y VGND VPWR sky130_fd_sc_hd__a22oi_4
XANTENNA__1026__B _1026_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_175 VGND VPWR sky130_fd_sc_hd__decap_8
X_1226_ web web0_sync _1208_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1157_ _1157_/D _1157_/Q _1173_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1042__A _1037_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1088_ _1088_/A _1083_/B _1136_/C _1073_/X _1088_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__0881__A _0786_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_7 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0759__C _1203_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0715__D1 _0714_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_67 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1102__D _1136_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_186 VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_clk clkbuf_0_clk/X clkbuf_1_0_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_98_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_86 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1127__A _1057_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0966__A _1060_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0721__A1 _0893_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1011_ _1259_/Q _0915_/X _0990_/X d_sram_in[31] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_97_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1029__A2 _0919_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0788__A1 _0682_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_19 VGND VPWR sky130_fd_sc_hd__decap_8
X_0726_ _0654_/Y _1178_/Q _0566_/Y _0726_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_0657_ _0611_/A _0636_/B _1191_/Q _0657_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__0579__C _1195_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1037__A _1037_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0588_ _0608_/A _0588_/B _0588_/C _0588_/D _0588_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_69_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0595__B _0621_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_167 VGND VPWR sky130_fd_sc_hd__fill_2
X_1209_ _1217_/Q _0568_/A _1218_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_138_125 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1206__CLK _1208_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_74 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0951__A1 _0949_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0786__A _0786_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0936__D _0936_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_93 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_251 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0696__A _0859_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_104 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_167 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0846__D _1173_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_115 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1229__CLK _1256_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_18 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_0709_ _0609_/Y _0708_/Y _0621_/A _0709_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0933__A1 _0927_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_57 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0767__A4 _0663_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_44 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1108__C _1097_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_43 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0688__B1 _0570_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0963__B _1026_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0860__B1 _0859_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0991_ _1243_/Q _0984_/X _0990_/X d_sram_in[15] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_125_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_85 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_126 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_17 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1050__A _1024_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0851__B1 _0850_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1200__D d_sram_out[23] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_49 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_38 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0906__A1 _1104_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_36 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0783__B _0521_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0842__B1 _0841_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_60 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0677__C _0677_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_80 VGND VPWR sky130_fd_sc_hd__fill_2
X_1190_ d_sram_out[13] _1190_/Q _1208_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_51_118 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1086__B1 _1079_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0974_ _0934_/Y _0966_/X _1239_/Q _0967_/X _0974_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_113_131 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1010__B1 _0986_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0868__B _0895_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1045__A _1270_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_137 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0824__B1 _0742_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1001__B1 _0951_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_153 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_52 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0794__A _0893_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_11 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_51 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_148 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1068__B1 _1062_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0815__B1 _0742_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_82 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_93 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_93 VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_6_0_clk clkbuf_4_6_0_clk/A _1177_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0690_ _0572_/Y _0681_/Y _0689_/Y _0690_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0969__A _0950_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_134 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_156 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_31 VGND VPWR sky130_fd_sc_hd__decap_12
X_1242_ d_fabric_in[14] _1242_/Q _1253_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_2_86 VGND VPWR sky130_fd_sc_hd__decap_12
X_1173_ _1173_/D _1173_/Q _1173_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_17_170 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0854__D _0589_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_140 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0806__B1 _0708_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_184 VGND VPWR sky130_fd_sc_hd__decap_6
X_0957_ _0960_/A _0957_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0585__A2 _0581_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0888_ _0662_/Y _0775_/X _0887_/Y d_fabric_out[26] VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__0990__C1 _0937_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0879__A _0663_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_43 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0764__D _1195_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_76 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_162 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_11 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_81 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_7 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_184 VGND VPWR sky130_fd_sc_hd__decap_6
X_0811_ _0811_/A _0893_/B _0811_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__1262__CLK _1274_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0742_ _0742_/A _0742_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0567__A2 _0562_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0673_ _0617_/Y _0883_/A _0666_/Y _0669_/Y _0672_/Y _0673_/Y VGND VPWR sky130_fd_sc_hd__a2111oi_4
XANTENNA__0699__A _0846_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1026__C _1026_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1225_ _1144_/X csb0_sync _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1156_ _1156_/D _1156_/Q _1173_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1087_ _1070_/X _1085_/Y _1086_/X w_mask[10] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0881__B _0889_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_25 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0715__C1 _0713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_165 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1285__CLK _1253_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_94 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1127__B _1127_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0721__A2 _0590_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1010_ _1258_/Q _0915_/X _0986_/Y d_sram_in[30] VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0982__A _0950_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0788__A2 _0822_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_74 VGND VPWR sky130_fd_sc_hd__decap_12
X_0725_ _0724_/Y _0666_/Y _0653_/Y _0725_/Y VGND VPWR sky130_fd_sc_hd__a21boi_4
X_0656_ _0623_/A _0611_/A _1187_/Q _0656_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__1037__B _1037_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0587_ _0587_/A _0588_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1158__CLK _1173_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_113 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0595__C _0594_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1208_ d_sram_out[31] _1208_/Q _1208_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1203__D d_sram_out[26] VGND VPWR sky130_fd_sc_hd__diode_2
X_1139_ _1090_/Y _1132_/X _1138_/X w_mask[28] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_43_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_16 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_42 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0951__A2 _0925_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_46 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_79 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_85 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_61 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_252 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_93 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_161 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0977__A _0921_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_129 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1048__A _1020_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0708_ _0539_/X _0558_/X _0608_/C _0708_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__0933__A2 _0916_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0639_ _0621_/B _0638_/Y _0590_/C _0639_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__0887__A _1171_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_27 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_48 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_23 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0797__A _0606_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1108__D _1136_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0688__A1 _0684_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_116 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0963__C _0961_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0860__A1 _0819_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0990_ _1243_/Q _0967_/X _0989_/Y _0937_/X _0990_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_117_118 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_64 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_138 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0851__A1 _0805_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_162 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0906__A2 _0988_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_21 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_149 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0783__C _0730_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_97 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0842__A1 _0779_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_62 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_165 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1219__CLK _1177_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_127 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_80 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1086__A1 _1050_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_91 VGND VPWR sky130_fd_sc_hd__fill_1
X_0973_ _1238_/Q _0957_/X _0972_/Y d_sram_in[10] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_72_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_110 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1010__A1 _1258_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_119 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_182 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0824__A1 _1184_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1211__D _1219_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1001__A1 _1249_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_165 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_45 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_96 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_56 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1068__A1 _1050_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0815__A1 _0814_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_83 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_8 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0969__B _0968_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0751__B1 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_43 VGND VPWR sky130_fd_sc_hd__decap_12
X_1241_ d_fabric_in[13] _1241_/Q _1256_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1191__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1172_ _1172_/D _1172_/Q _1172_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_2_98 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0806__A1 _0807_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_19 VGND VPWR sky130_fd_sc_hd__decap_12
X_0956_ _0914_/Y _0960_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0887_ _1171_/Q _0895_/B _0887_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__0990__B1 _0989_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0879__B _0889_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0895__A _1175_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1206__D d_sram_out[29] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0981__B1 _1241_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_63 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_60 VGND VPWR sky130_fd_sc_hd__fill_1
X_0810_ _0804_/Y _0692_/X _0808_/X _0809_/Y _0811_/A VGND VPWR sky130_fd_sc_hd__a22oi_4
X_0741_ _0728_/Y _0740_/Y _0566_/Y _0741_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0672_ _0672_/A _0594_/X _0671_/Y _0672_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0699__B _0846_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_3 VGND VPWR sky130_fd_sc_hd__decap_4
X_1224_ _1224_/D _1216_/D _1253_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1155_ _0839_/B _1155_/Q _1172_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1086_ _1050_/X _1065_/Y _1079_/X _1086_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_20_166 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_133 VGND VPWR sky130_fd_sc_hd__fill_2
X_0939_ _0934_/Y _0925_/X _0938_/Y _0939_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0715__B1 _0712_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_5_0_clk clkbuf_3_2_0_clk/X _1256_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_113_32 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1140__B1 _1138_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_58 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_133 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_40 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_11 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0954__B1 _0931_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_55 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1127__C _1127_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_147 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1131__B1 _1129_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0982__B _0981_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0788__A3 _0551_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_86 VGND VPWR sky130_fd_sc_hd__decap_8
X_0724_ _1186_/Q _0724_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0655_ _1177_/Q _0651_/X _0654_/Y _0655_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0586_ _1174_/D _0893_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_69_111 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0595__D _1208_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1207_ d_sram_out[30] _0589_/A _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1122__B1 _1119_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1138_ _1024_/X _1097_/Y _1137_/X _1138_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_1069_ _1044_/X _1067_/Y _1068_/X w_mask[6] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_138_149 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_54 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_36 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_31 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_53 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_42 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_147 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1252__CLK _1252_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_57 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1113__B1 _1111_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_84 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_242 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_127 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_173 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0977__B _0961_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_171 VGND VPWR sky130_fd_sc_hd__decap_12
X_0707_ _0704_/X _0701_/A _0706_/Y d_fabric_out[0] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0638_ _0637_/Y _0638_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0887__B _0895_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0569_ _0653_/B _0698_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_38_17 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1275__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_147 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1214__D _1214_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_38 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0688__A2 _0686_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_128 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0963__D _0963_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0860__A2 _0749_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1148__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0988__A _0921_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_158 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0851__A2 _0749_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_119 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1059__A _1057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_152 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1209__D _1217_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_128 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0783__D _1208_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_161 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0842__A2 _0760_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_41 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_111 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0601__A _0621_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_177 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_117 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1086__A2 _1065_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0972_ _0986_/A _0971_/Y _0986_/C _0930_/Y _0972_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_65_3 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1010__A2 _0915_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0803__B1_N _0802_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_19 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0818__B1_N _0817_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0824__A2 _0760_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_153 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_7 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1001__A2 _1000_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_177 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1068__A2 _1055_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_40 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0815__A2 _0607_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_73 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_83 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_114 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0751__A1 _0746_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1240_ d_fabric_in[12] _1240_/Q _1252_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_2_55 VGND VPWR sky130_fd_sc_hd__decap_6
X_1171_ _1203_/Q _1171_/Q _1173_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0806__A2 _0805_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0955_ _1234_/Q _0916_/X _0954_/Y d_sram_in[6] VGND VPWR sky130_fd_sc_hd__a21o_4
X_0886_ _0870_/X _1170_/Q _0885_/Y d_fabric_out[25] VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0990__A1 _1243_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_147 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0895__B _0895_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_158 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1222__D _1222_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_131 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1209__CLK _1218_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0981__B2 _0967_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_164 VGND VPWR sky130_fd_sc_hd__fill_2
X_0740_ _1182_/Q _0729_/Y _0732_/Y _0734_/X _0739_/X _0740_/Y VGND VPWR sky130_fd_sc_hd__a2111oi_4
X_0671_ _0607_/A _0609_/A _0590_/C _0671_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__0699__C _0846_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0996__A _0996_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_3 VGND VPWR sky130_fd_sc_hd__fill_1
X_1223_ _1286_/Q _1215_/D _1253_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1154_ _1154_/D _1154_/Q _1172_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1085_ _1088_/A _1059_/B _1074_/C _1073_/X _1085_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_32_19 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_123 VGND VPWR sky130_fd_sc_hd__fill_1
X_0938_ _0937_/X _0938_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0869_ _0843_/X _1163_/Q _0868_/Y d_fabric_out[18] VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1067__A _1075_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1217__D _0914_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0715__A1 _0603_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_55 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1140__A1 _1095_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_37 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_88 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_105 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1181__CLK _1180_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_63 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0954__A1 _0953_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1131__A1 _1083_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_93 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0890__B1 _0889_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0788__A4 _0786_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0792__A2_N _0693_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0723_ _0711_/X _0715_/Y _0719_/Y _0722_/Y _0723_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_0654_ _0653_/Y _0654_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0585_ _0578_/Y _0581_/X _0718_/A _0585_/Y VGND VPWR sky130_fd_sc_hd__a21boi_4
XFILLER_69_189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_148 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_7_0_clk_A clkbuf_4_6_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1206_ d_sram_out[29] _1174_/D _1208_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1122__A1 _1065_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1137_ _1118_/A _1137_/B _1136_/Y _1137_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_1068_ _1050_/X _1055_/Y _1062_/X _1068_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_138_106 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_99 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_115 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1113__A1 _1051_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_210 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_51 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_276 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_139 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_73 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_185 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0977__C _0988_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_104 VGND VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_4_0_clk clkbuf_3_2_0_clk/X _1252_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0706_ _1145_/Q _0705_/X _0706_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_0637_ _0588_/D _0637_/B _0637_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_0568_ _0568_/A _0570_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_80_140 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_12 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1230__D d_fabric_in[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_49 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_21 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_109 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_36 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_62 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0845__B1 _0844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_94 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_142 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0988__B _0936_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1089__B1 _1086_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0836__B1 _0835_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1242__CLK _1253_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1059__B _1059_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1075__A _1075_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1225__D _1144_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_78 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_107 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_4_0_clk_A clkbuf_3_5_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0601__B _0600_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_145 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_134 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_50 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_15_0_clk_A clkbuf_3_7_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_71 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1265__CLK _1166_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0971_ _0917_/Y _0966_/X _1238_/Q _0967_/X _0971_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_58_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0809__B1 _0742_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_176 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0702__A out_reg VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_101 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_11 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_48 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1288__CLK _1288_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_30 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_63 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_74 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_154 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_96 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_51 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0612__A _0612_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0751__A2 _0748_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_126 VGND VPWR sky130_fd_sc_hd__fill_2
X_1170_ _0747_/A _1170_/Q _1172_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_66_92 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_176 VGND VPWR sky130_fd_sc_hd__fill_2
X_0954_ _0953_/Y _0925_/X _0931_/X _0954_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0885_ _0747_/Y _0889_/B _0885_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__0522__A _0521_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0990__A2 _0967_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_24 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_154 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_187 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_58 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_1_0_clk_A clkbuf_1_0_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0607__A _0607_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_94 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_72 VGND VPWR sky130_fd_sc_hd__fill_2
X_0670_ _1189_/Q _0672_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0699__D _0577_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0996__B _0986_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_80 VGND VPWR sky130_fd_sc_hd__decap_3
X_1222_ _1222_/D _1214_/D _1253_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1153_ _0831_/B _1153_/Q _1173_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1084_ _1070_/X _1083_/Y _1080_/X w_mask[9] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0517__A reb VGND VPWR sky130_fd_sc_hd__diode_2
X_0937_ _0899_/A _1023_/A _0936_/X _0911_/A _0937_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_9_180 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_3_0_clk_A clkbuf_4_2_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0868_ _0868_/A _0895_/B _0868_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__1067__B _1127_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0799_ _0822_/B _0672_/A _0675_/Y _0799_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0715__A2 _1196_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_157 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1083__A _1057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1233__D d_fabric_in[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_27 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1140__A2 _1132_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_146 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0954__A2 _0925_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_79 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1131__A2 _1121_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0890__A1 _0874_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_7 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_82 VGND VPWR sky130_fd_sc_hd__fill_2
X_0722_ _0721_/Y _0722_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0653_ _0570_/B _0653_/B _0691_/A _0653_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_0584_ _0624_/C _0718_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_40_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_102 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_146 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_179 VGND VPWR sky130_fd_sc_hd__fill_2
X_1205_ d_sram_out[28] _1173_/D _1208_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1122__A2 _1121_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1136_ _1136_/A _1136_/B _1136_/C _1136_/D _1136_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__0709__B1_N _0621_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1067_ _1075_/A _1127_/B _1018_/A _1058_/A _1067_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_138_118 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1078__A _1075_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1228__D d_fabric_in[0] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0710__A _0763_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1113__A2 _1105_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_171 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_200 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_233 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0620__A _0585_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0977__D _0977_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_119 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_70 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_0705_ _0861_/A _0705_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_128_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0530__A _0530_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0636_ _0612_/A _0636_/B _1184_/Q _0636_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_0567_ _0527_/Y _0562_/Y _0566_/Y _0567_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_57_138 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1171__CLK _1173_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1119_ _1106_/X _1085_/Y _1118_/X _1119_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0705__A _0861_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_0_0_clk_A clkbuf_3_1_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0790__B1 _0789_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_105 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_58 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0845__A1 _0843_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_185 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_73 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_11_0_clk_A clkbuf_3_5_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0615__A _0607_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_94 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0988__C _0988_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_56 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0781__B1 _1196_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_81 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1194__CLK _1184_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_182 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1089__A1 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0836__A1 _0705_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_163 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0525__A _0590_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1059__C _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_165 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0772__B1 _0761_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0619_ _0604_/Y _0613_/X _0619_/C _0619_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_131_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_57 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1091__A _1067_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_141 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0827__A1 _0825_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1241__D d_fabric_in[13] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_31 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1004__A1 _1252_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0601__C _1203_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_157 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_84 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_3_0_clk clkbuf_4_2_0_clk/A _1274_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0818__A1 _0816_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1151__D _0816_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0970_ _1237_/Q _0957_/X _0969_/Y d_sram_in[9] VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0809__A1 _1182_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0993__B1 _0992_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_113 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1236__D d_fabric_in[8] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_56 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_66 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_99 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_31 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_122 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_64 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_133 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_75 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_97 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1146__D _0753_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_71 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1232__CLK _1288_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_92 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_144 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_166 VGND VPWR sky130_fd_sc_hd__decap_4
X_0953_ _1234_/Q _0953_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_70_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_0884_ _0870_/X _1169_/Q _0883_/X d_fabric_out[24] VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_99_111 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_144 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0727__B1 _0726_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_127 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0713__A _0718_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1255__CLK _1288_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1143__B1 _1141_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0607__B _0607_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_62 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0623__A _0623_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_103 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_7 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0996__C _0996_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1221_ _1284_/Q _1213_/D _1218_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1134__B1 _1133_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1152_ _0825_/Y _0826_/B _1173_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1083_ _1057_/X _1083_/B _1136_/C _1073_/X _1083_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__0517__B csb VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_114 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_169 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0533__A _0533_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0936_ _0936_/A _1026_/B _0903_/X _0936_/D _0936_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0948__B1 _0947_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0867_ _0577_/X _0704_/X _0866_/X d_fabric_out[17] VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1067__C _1018_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0798_ _0627_/C _0749_/X _0742_/A _0798_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__1278__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1083__B _1083_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1125__B1 _1123_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0708__A _0539_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_32 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0939__B1 _0938_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_14 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_98 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_47 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_87 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1116__B1 _1114_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0890__A2 _1172_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0721_ _0893_/A _0590_/Y _0720_/Y _0721_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_10_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_140 VGND VPWR sky130_fd_sc_hd__fill_2
X_0652_ _0620_/Y _0650_/Y _0651_/X _0652_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_6_184 VGND VPWR sky130_fd_sc_hd__decap_6
X_0583_ _0583_/A _0624_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_33_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1107__B1 _1029_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_180 VGND VPWR sky130_fd_sc_hd__fill_2
X_1204_ d_sram_out[27] _1172_/D _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0528__A _0590_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1135_ _1088_/Y _1132_/X _1133_/X w_mask[27] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_92_161 VGND VPWR sky130_fd_sc_hd__fill_2
X_1066_ _1044_/X _1065_/Y _1063_/X w_mask[5] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__1078__B _1127_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0919_ _0922_/C _0919_/B _0921_/A _0919_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0710__B _0600_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_34 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_23 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1244__D d_fabric_in[16] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_183 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_54 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_201 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0901__A _1026_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_154 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0620__B _0602_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_50 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1154__D _1154_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0974__A2_N _0966_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0704_ _0826_/A _0704_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0811__A _0811_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0635_ _0635_/A _0623_/A _1186_/Q _0640_/A VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_99_90 VGND VPWR sky130_fd_sc_hd__fill_2
X_0566_ _0566_/A _0566_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_57_106 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_183 VGND VPWR sky130_fd_sc_hd__decap_6
X_1118_ _1118_/A _1118_/B _1117_/Y _1118_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_80_175 VGND VPWR sky130_fd_sc_hd__fill_2
X_1049_ _1088_/A _1059_/B _1018_/X _1083_/B _1049_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_110_36 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1239__D d_fabric_in[11] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0790__A1 _0784_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_113 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_31 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0845__A2 _1156_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0615__B _0615_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1149__D _0802_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_13 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0631__A _0599_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0988__D _0988_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0781__B2 _0600_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_161 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1089__A2 _1088_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_142 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0836__A2 _1154_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1059__D _1097_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_100 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0541__A _0536_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_177 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0772__B2 _0771_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0618_ _0889_/A _0615_/Y _1173_/D _0617_/Y _0619_/C VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_131_147 VGND VPWR sky130_fd_sc_hd__decap_6
X_0549_ _0573_/B _0608_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_105_25 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1091__B _1106_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0827__A2 _0794_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0716__A _0574_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_79 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_33 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1004__A2 _0960_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_98 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0818__A2 _0794_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_84 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0626__A _0626_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1161__CLK _1173_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0739__D1 _0738_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_158 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_80 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0809__A2 _0749_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_186 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0536__A _0609_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_156 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0690__B1 _0689_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0993__A1 _0910_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1252__D d_fabric_in[24] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_56 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_131 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_21 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_87 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0681__B1 _0680_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_98 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1184__CLK _1184_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_50 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1162__D _0737_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0952_ _0949_/A _0916_/X _0951_/Y d_sram_in[5] VGND VPWR sky130_fd_sc_hd__a21o_4
X_0883_ _0883_/A _0883_/B _0883_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_63_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0727__A1 _0723_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_19 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_101 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_145 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1097__A _1136_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0713__B _0536_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_2_0_clk clkbuf_4_2_0_clk/A _1166_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_11_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1247__D d_fabric_in[19] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_7 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1143__A1 _1102_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_53 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_112 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0607__C _0607_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0904__A _0903_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0623__B _0622_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1157__D _1157_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0709__A1 _0609_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_7 VGND VPWR sky130_fd_sc_hd__fill_1
X_1220_ _1220_/D _1212_/D _1253_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1134__A1 _1085_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1151_ _0816_/Y _1151_/Q _1173_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1082_ _1082_/A _1136_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_20_137 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0948__A1 _0977_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0935_ _1026_/B _0903_/X _0922_/B _1023_/A VGND VPWR sky130_fd_sc_hd__nor3_4
X_0866_ _0866_/A _0871_/A _0866_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_0797_ _0606_/C _0797_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1067__D _1058_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1083__C _1136_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1125__A1 _1071_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_58 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0884__B1 _0883_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0708__B _0558_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_104 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_137 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0724__A _1186_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_108 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0939__A1 _0934_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_55 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1061__B1 _1060_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_26 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1222__CLK _1253_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1116__A1 _1055_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_41 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0634__A _0634_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0720_ _0889_/A _0588_/Y _0747_/A _0617_/Y _0720_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__1052__B1 _1034_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0651_ _0698_/A _0570_/A _0570_/B _0651_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_0582_ _0588_/C _0587_/A _0583_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_88_70 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1107__A1 _1136_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1203_ d_sram_out[26] _1203_/Q _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_92_140 VGND VPWR sky130_fd_sc_hd__fill_2
X_1134_ _1085_/Y _1132_/X _1133_/X w_mask[26] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_92_184 VGND VPWR sky130_fd_sc_hd__decap_6
X_1065_ _1057_/X _1018_/X _1102_/B _1097_/D _1065_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__0618__B1 _1173_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0544__A _0608_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1245__CLK _1288_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1078__C _1127_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0918_ _0914_/A _0921_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_0849_ _0705_/X _1157_/D _0848_/X d_fabric_out[12] VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0710__C _0597_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_29 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_46 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0719__A _0666_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_140 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_39 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_22 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1260__D addr_w[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_99 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_224 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_144 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0620__C _0619_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0629__A _0627_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1170__D _0747_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1268__CLK _1274_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0703_ _0861_/A _0826_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0811__B _0893_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0634_ _0634_/A _0633_/Y _0634_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_0565_ _0564_/Y _0566_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_57_118 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0539__A _0607_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_140 VGND VPWR sky130_fd_sc_hd__fill_2
X_1117_ _1095_/A _1136_/B _1136_/C _1136_/D _1117_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_80_132 VGND VPWR sky130_fd_sc_hd__fill_2
X_1048_ _1020_/Y _1083_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_119_13 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_79 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0790__A2 _0533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_125 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1255__D d_fabric_in[27] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_16 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_98 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_143 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0615__C _0588_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_41 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1007__B1 _0975_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0912__A _0911_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0631__B _0622_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_69 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1165__D _0606_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_129 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_93 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_3 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0822__A _0822_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0541__B _0539_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_156 VGND VPWR sky130_fd_sc_hd__decap_6
X_0617_ _0609_/A _0608_/B _0617_/C _0617_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_0548_ _0615_/B _0551_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_105_37 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_151 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_165 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0716__B _0615_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_23 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0732__A _0731_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_55 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_126 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_115 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0907__A _0919_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0626__B _0623_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0642__A _0635_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0739__C1 _0736_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_148 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_121 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0817__A _0826_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_154 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_132 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0690__A1 _0572_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_168 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0552__A _0764_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0993__A2 _0960_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_14 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_13 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_110 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_22 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0681__A1 _0652_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_88 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_80 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_91 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0637__A _0588_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_154 VGND VPWR sky130_fd_sc_hd__decap_3
X_0951_ _0949_/Y _0925_/X _0950_/X _0951_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0882_ _0870_/X _1168_/Q _0881_/Y d_fabric_out[23] VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0727__A2 _0725_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0547__A _0547_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_16 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_49 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_135 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_124 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_179 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1097__B _1097_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0713__C _0539_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1263__D addr_w[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_140 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1143__A2 _1132_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_173 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1151__CLK _1173_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_97 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0623__C _1190_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0920__A _0919_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0709__A2 _0708_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_127 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1173__D _1173_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1134__A2 _1132_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1150_ _0811_/A _1150_/Q _1166_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1081_ _1070_/X _1074_/Y _1080_/X w_mask[8] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_93_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_150 VGND VPWR sky130_fd_sc_hd__fill_1
X_0934_ _0936_/D _0934_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0865_ _0843_/X _1161_/Q _0864_/Y d_fabric_out[16] VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0948__A2 _0916_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0830__A _0861_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0796_ _1148_/D _0794_/X _0795_/Y d_fabric_out[3] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_87_127 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1083__D _1073_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1174__CLK _1173_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1125__A2 _1121_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_171 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0708__C _0608_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0884__A1 _0870_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1279_ addr_r[5] baseaddr_r_sync[5] _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1061__A1 _1095_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0939__A2 _0925_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1258__D d_fabric_in[30] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_56 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_127 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1116__A2 _1105_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0585__B1_N _0718_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_97 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0915__A _0914_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0634__B _0633_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_47 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1168__D _0786_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1052__A1 _1050_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0650_ _0647_/Y _0649_/Y _0602_/A _0650_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_6_175 VGND VPWR sky130_fd_sc_hd__fill_2
X_0581_ _0579_/Y _0580_/Y _0581_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1197__CLK _1208_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1107__A2 _0919_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1202_ d_sram_out[25] _0747_/A _1208_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_19_3 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_1_0_clk clkbuf_3_0_0_clk/X _1253_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1133_ _1024_/X _1095_/Y _1128_/X _1133_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_1064_ _1044_/X _1059_/Y _1063_/X w_mask[4] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0618__B2 _0617_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0917_ _0927_/D _0917_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0560__A _0558_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0848_ _1157_/Q _0870_/A _0848_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_0779_ _0621_/C _0779_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_68_19 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0710__D _1190_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_119 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0719__B _0716_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0735__A _0667_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_225 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_11 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_258 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_55 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_269 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_182 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0629__B _0628_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_91 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_73 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0645__A _0645_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_72 VGND VPWR sky130_fd_sc_hd__fill_2
X_0702_ out_reg _0861_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0633_ _0630_/Y _0633_/B _0632_/Y _0633_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_0564_ _0691_/A _0568_/A _0653_/B _0564_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_1116_ _1055_/Y _1105_/X _1114_/X w_mask[19] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__1212__CLK _1252_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_155 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_16 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0555__A _0667_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1047_ _1127_/B _1059_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_119_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_58 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0790__A3 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_28 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_66 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1271__D addr_w[11] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_98 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0615__D _0588_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1007__A1 _1255_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_86 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0631__C _1191_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0766__B1 _0628_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_51 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_108 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1235__CLK _1253_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1181__D d_sram_out[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_83 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0822__B _0822_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0541__C _0883_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0616_ _0588_/C _0587_/A _0617_/C VGND VPWR sky130_fd_sc_hd__nand2_4
X_0547_ _0547_/A _0615_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_144 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0716__C _0594_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_135 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0748__B1 _0577_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1266__D addr_w[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_32 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1258__CLK _1177_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_54 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0626__C _0626_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_52 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0987__B1 _0986_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0923__A _1127_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0642__B _0599_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0739__B1 _0533_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1176__D _1208_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_160 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_182 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0817__B _1151_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_147 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_136 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0690__A2 _0681_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0833__A _0846_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0552__B _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_36 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_23 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_56 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0681__A2 _0655_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_89 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_22 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_55 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0918__A _0914_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0637__B _0637_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0653__A _0570_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0950_ _0994_/A _0944_/Y _0986_/A _0950_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0881_ _0786_/Y _0889_/B _0881_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_99_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_158 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_3 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0828__A _0846_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_28 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0563__A _0570_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0713__D _1182_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1097__C _1102_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_36 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_152 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0738__A _0737_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_33 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_117 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1119__B1 _1118_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0648__A _1185_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1080_ _1050_/X _1059_/Y _1079_/X _1080_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0933_ _0927_/D _0916_/X _0932_/Y d_sram_in[2] VGND VPWR sky130_fd_sc_hd__a21o_4
X_0864_ _0559_/Y _0895_/B _0864_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_0795_ _0826_/A _0795_/B _0795_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__0558__A _0607_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_183 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_38 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0884__A2 _1169_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1278_ addr_r[4] baseaddr_r_sync[4] _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1061__A2 _1126_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1274__D addr_r[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1052__A2 _1051_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0931__A _0911_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_90 VGND VPWR sky130_fd_sc_hd__fill_1
X_0580_ _0667_/B _0608_/B _1196_/Q _0580_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_40_7 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1184__D d_sram_out[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_109 VGND VPWR sky130_fd_sc_hd__decap_4
X_1201_ d_sram_out[24] _1169_/D _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_92_120 VGND VPWR sky130_fd_sc_hd__fill_2
X_1132_ _1132_/A _1132_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_92_175 VGND VPWR sky130_fd_sc_hd__decap_8
X_1063_ _1050_/X _1049_/Y _1062_/X _1063_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0841__A _0859_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0916_ _0915_/X _0916_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0847_ _0672_/A _0750_/X _0846_/Y _1157_/D VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0560__B _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0778_ _1196_/Q _0872_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_108_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_19 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0719__C _0719_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0735__B _0520_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_215 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1269__D addr_w[9] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_42 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0926__A _0922_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_96 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0645__B _0645_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_7 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_62 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1179__D d_sram_out[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_111 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1164__CLK _1172_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0661__A _0576_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0701_ _0701_/A _0701_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0632_ _0544_/X _0606_/B _0615_/B _0632_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_0563_ _0570_/A _0691_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_99_93 VGND VPWR sky130_fd_sc_hd__fill_2
X_1115_ _1049_/Y _1105_/X _1114_/X w_mask[18] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0555__B _0520_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1046_ _1075_/A _1088_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_119_111 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_80 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0571__A _0745_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_37 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_147 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0790__A4 _0788_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_153 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_77 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1187__CLK _1180_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_83 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_54 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_32 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1007__A2 _0915_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_98 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0766__B2 _0729_/Y VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_0_0_clk clkbuf_3_0_0_clk/X _1288_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_109_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_85 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_186 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0656__A _0623_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_3 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0822__C _0786_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0541__D _0528_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0615_ _0607_/B _0615_/B _0588_/B _0588_/D _0615_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_0546_ _0546_/A _0547_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_38_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0566__A _0566_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_27 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0716__D _0577_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1029_ _0903_/X _0919_/B _0914_/Y _1029_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0748__B2 _0600_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_147 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_158 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1282__D addr_r[8] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_175 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_87 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_145 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_123 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0684__B1 _0683_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0626__D _0625_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0987__A1 _1242_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0642__C _1187_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0739__A1 _0531_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_106 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1202__CLK _1208_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1192__D d_sram_out[15] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_101 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_145 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0833__B _0846_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0552__C _0528_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_7_0_clk clkbuf_3_7_0_clk/A clkbuf_3_7_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_104_128 VGND VPWR sky130_fd_sc_hd__decap_3
X_0529_ _0542_/A _0573_/B _0530_/A VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_26_123 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_13 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_156 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_46 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1225__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1277__D addr_r[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0934__A _0936_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0653__B _0653_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_7 VGND VPWR sky130_fd_sc_hd__fill_2
X_0880_ _0870_/X _1167_/Q _0879_/Y d_fabric_out[22] VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1187__D d_sram_out[10] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_115 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0896__B1 _0895_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0828__B _0846_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0844__A _0883_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1248__CLK _1253_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0618__A1_N _0889_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1097__D _1097_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_15 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_89 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0754__A _0705_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1064__B1 _1063_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_88 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1119__A1 _1106_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_63 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0929__A _0928_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_85 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0878__B1 _0877_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_118 VGND VPWR sky130_fd_sc_hd__fill_1
X_0932_ _0917_/Y _0925_/X _0931_/X _0932_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0863_ _0871_/A _0895_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_61_3 VGND VPWR sky130_fd_sc_hd__fill_1
X_0794_ _0893_/B _0794_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0839__A _0883_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0869__B1 _0868_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_93 VGND VPWR sky130_fd_sc_hd__decap_4
X_1277_ addr_r[3] baseaddr_r_sync[3] _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0574__A _0573_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_129 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1061__A3 _1109_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0749__A _0749_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1290__D conf[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0931__B _0986_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_155 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0971__A2_N _0966_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0659__A _0636_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1200_ d_sram_out[23] _0786_/A _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_77_184 VGND VPWR sky130_fd_sc_hd__decap_6
X_1131_ _1083_/Y _1121_/X _1129_/X w_mask[25] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_92_165 VGND VPWR sky130_fd_sc_hd__fill_2
X_1062_ _1030_/Y _1061_/Y _1062_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0841__B _0859_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0915_ _0914_/Y _0915_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0846_ _0846_/A _0846_/B _0846_/C _1173_/D _0846_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__0560__C _0559_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0777_ _0772_/X _0775_/X _0776_/Y d_fabric_out[2] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0569__A _0653_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_151 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0719__D _0719_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_58 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0735__C _0729_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_216 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_24 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_249 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_3 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1285__D addr_r[11] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_54 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_87 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0645__C _0643_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_52 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0942__A _0922_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0661__B _1179_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0700_ _0690_/Y _0693_/Y _0699_/X _0701_/A VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_128_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_0631_ _0599_/Y _0622_/Y _1191_/Q _0633_/B VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_99_72 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1195__D d_sram_out[18] VGND VPWR sky130_fd_sc_hd__diode_2
X_0562_ _1189_/Q _0531_/Y _0533_/X _0553_/Y _0561_/X _0562_/Y VGND VPWR sky130_fd_sc_hd__a2111oi_4
XFILLER_24_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_154 VGND VPWR sky130_fd_sc_hd__fill_2
X_1114_ _1106_/X _1083_/Y _1110_/X _1114_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0555__C _1173_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1013__A _1013_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1045_ _1270_/Q _1075_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_80_179 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0852__A _0861_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_134 VGND VPWR sky130_fd_sc_hd__fill_2
X_0829_ _0683_/B _0760_/X _0828_/Y _0831_/B VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_134_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_35 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0816__A2_N _0693_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_45 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0762__A _1191_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_17 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_165 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0656__B _0611_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0672__A _0672_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1281__CLK _1159_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_104 VGND VPWR sky130_fd_sc_hd__fill_1
X_0614_ _1172_/D _0889_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_0545_ _0544_/X _0764_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_105_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_1028_ _1031_/B _1127_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0582__A _0588_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_37 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_47 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0757__A _0764_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1154__CLK _1172_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_187 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0684__A1 _0600_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_157 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_32 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0987__A2 _0984_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0739__A2 _1190_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_40 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_62 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_140 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0667__A _0606_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_113 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0833__C _0846_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0552__D _0606_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_107 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_118 VGND VPWR sky130_fd_sc_hd__fill_2
X_0528_ _0590_/C _0528_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1177__CLK _1177_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0577__A _0737_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_135 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_47 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_50 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_54 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_65 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_124 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0653__C _0691_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_7 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0896__A1 _0589_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0828__C _0883_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0844__B _1156_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1021__A _1020_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_182 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0772__A1_N _0868_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0787__A1_N _0889_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_57 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_127 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0754__B _0754_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1064__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1288__D conf[0] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1119__A2 _1085_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_42 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_182 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0878__A1 _0804_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1106__A _1106_/A VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_6_0_clk clkbuf_3_7_0_clk/A clkbuf_3_6_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_93_74 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0945__A _0944_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0931_ _0911_/Y _0986_/C _0930_/Y _0931_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_13_182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_142 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0680__A _0679_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1198__D d_sram_out[21] VGND VPWR sky130_fd_sc_hd__diode_2
X_0862_ _0843_/X _1160_/Q _0861_/X d_fabric_out[15] VGND VPWR sky130_fd_sc_hd__o21a_4
X_0793_ _0793_/A _0893_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_54_3 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0839__B _0839_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0869__A1 _0843_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1016__A _1031_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1215__CLK _1252_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1276_ addr_r[2] baseaddr_r_sync[2] _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1061__A4 _1074_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0590__A _0607_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_39 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0931__C _0930_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0659__B _0628_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1238__CLK _1256_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1130_ _1074_/Y _1121_/X _1129_/X w_mask[24] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0720__B1 _0747_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0675__A _0539_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1061_ _1095_/A _1126_/B _1109_/B _1074_/C _1060_/Y _1061_/Y VGND VPWR sky130_fd_sc_hd__a41oi_4
XANTENNA__0841__C _0859_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0914_ _0914_/A _0922_/C _0919_/B _0914_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_0845_ _0843_/X _1156_/Q _0844_/X d_fabric_out[11] VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0787__B1 _1184_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0776_ _0826_/A _1147_/Q _0776_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_68_174 VGND VPWR sky130_fd_sc_hd__fill_2
X_1259_ d_fabric_in[31] _1259_/Q _1177_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0735__D _1174_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_206 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_148 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0950__B1 _0986_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0645__D _0644_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_71 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0942__B _0914_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_91 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0661__C _0718_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0769__B1 _0566_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0630_ _0629_/Y _0612_/A _0630_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_99_51 VGND VPWR sky130_fd_sc_hd__fill_2
X_0561_ _0556_/Y _0560_/Y _0763_/A _0561_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_99_84 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_111 VGND VPWR sky130_fd_sc_hd__decap_4
X_1113_ _1051_/Y _1105_/X _1111_/X w_mask[17] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_80_114 VGND VPWR sky130_fd_sc_hd__fill_2
X_1044_ _1043_/X _1044_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_80_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0812__B1_N _0811_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0852__B _1158_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_17 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_93 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0827__B1_N _0826_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0828_ _0846_/A _0846_/B _0883_/A _0846_/C _0828_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_0759_ _0822_/B _0859_/A _1203_/Q _0759_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_135_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0932__B1 _0931_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_47 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_24 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0999__B1 _0947_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_3 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0985__A2_N _0966_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_60 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_93 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_100 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_86 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_114 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0656__C _1187_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0953__A _1234_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1100__B1 _1099_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0672__B _0594_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_127 VGND VPWR sky130_fd_sc_hd__fill_2
X_0613_ _0606_/Y _0607_/Y _0608_/Y _0609_/Y _0612_/Y _0613_/X VGND VPWR sky130_fd_sc_hd__a41o_4
X_0544_ _0608_/A _0544_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_124_171 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1024__A _1106_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_125 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0863__A _0871_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1027_ _1037_/A _1037_/B _1022_/Y _1027_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0582__B _0587_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_160 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_182 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0757__B _1187_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0684__A2 _1161_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0773__A out_reg VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1109__A _1057_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_152 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0667__B _0667_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0683__A _0682_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0833__D _0747_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1019__A _1019_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_18 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_29 VGND VPWR sky130_fd_sc_hd__fill_2
X_0527_ _0807_/B _1185_/Q _0763_/A _0527_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_112_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_169 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0593__A _0636_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_37 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0768__A _1187_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_19 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1271__CLK _1166_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_32 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_117 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_128 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0896__A2 _0775_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0828__D _0846_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_128 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_161 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_39 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0588__A _0608_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_111 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_47 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1064__A2 _1059_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_161 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0878__A2 _0775_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_86 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1167__CLK _1172_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0961__A _0936_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0930_ _0921_/X _1026_/A _1026_/C d_sram_in[0] _0930_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_9_121 VGND VPWR sky130_fd_sc_hd__fill_2
X_0861_ _0861_/A _1160_/D _0861_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_9_154 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0680__B _0566_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0792_ _0872_/A _0693_/Y _0782_/Y _0791_/X _1148_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0869__A2 _1163_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_175 VGND VPWR sky130_fd_sc_hd__fill_2
X_1275_ addr_r[1] baseaddr_r_sync[1] _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0871__A _0871_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0590__B _0607_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_46 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_68 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_78 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0796__A1 _1148_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_75 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0659__C _0583_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1117__A _1095_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0956__A _0914_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0720__B2 _0617_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0675__B _0558_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1060_ _1060_/A _1060_/B _1060_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__0691__A _0691_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0913_ _0994_/A _0994_/B _0986_/A d_sram_in[1] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0844_ _0883_/B _1156_/D _0844_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0841__D _1172_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0787__B2 _0729_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0775_ _0870_/A _0775_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1027__A _1037_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0866__A _0866_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_27 VGND VPWR sky130_fd_sc_hd__fill_2
X_1258_ d_fabric_in[30] _1258_/Q _1177_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_83_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_189 VGND VPWR sky130_fd_sc_hd__fill_1
X_1189_ d_sram_out[12] _1189_/Q _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_207 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_229 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_clk clkbuf_3_5_0_clk/A clkbuf_3_5_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0950__A1 _0994_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_186 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0776__A _0826_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_11 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_44 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_55 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_66 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_167 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0942__C _0902_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_76 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0769__A1 _0768_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_147 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1205__CLK _1208_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0560_ _0558_/X _0550_/X _0559_/Y _0560_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_2_171 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0686__A _0807_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_145 VGND VPWR sky130_fd_sc_hd__fill_2
X_1112_ _1022_/Y _1105_/X _1111_/X w_mask[16] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_65_189 VGND VPWR sky130_fd_sc_hd__fill_1
X_1043_ _1043_/A _1043_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_63 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_158 VGND VPWR sky130_fd_sc_hd__decap_3
X_0827_ _0825_/Y _0794_/X _0826_/Y d_fabric_out[7] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0758_ _0807_/B _0859_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0689_ _0689_/A _0689_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0932__A1 _0917_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0596__A _0587_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0999__A1 _1248_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1228__CLK _1256_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_51 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_32 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_81 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1100__A1 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0672__C _0671_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_7 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0612_ _0612_/A _0612_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0543_ _0543_/A _0608_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_148 VGND VPWR sky130_fd_sc_hd__fill_2
X_1026_ _1026_/A _1026_/B _1026_/C _1037_/B VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__1040__A _1039_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_139 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0669__B1 _0617_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1094__B1 _1093_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_23 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_56 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_60 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1109__B _1109_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_93 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_53 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0667__C _1173_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_91 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0964__A _0964_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0683__B _0683_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0832__B1 _0831_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_3 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_62 VGND VPWR sky130_fd_sc_hd__decap_4
X_0526_ _0729_/B _0763_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1035__A _1034_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0874__A _0871_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_148 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_27 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_38 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_118 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VPWR sky130_fd_sc_hd__decap_3
X_1009_ _1257_/Q _0915_/X _0982_/Y d_sram_in[29] VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0823__B1 _0742_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0784__A _0783_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_170 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_71 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0814__B1 _0668_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0694__A _0691_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_29 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0588__B _0588_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_7_0_clk_A clkbuf_3_7_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_25 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_173 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0779__A _0621_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_72 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_92 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_162 VGND VPWR sky130_fd_sc_hd__fill_2
X_0860_ _0819_/Y _0749_/X _0859_/Y _1160_/D VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0791_ _0624_/B _0566_/A _0745_/X _0790_/X _0791_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_9_188 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0689__A _0689_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_110 VGND VPWR sky130_fd_sc_hd__fill_2
X_1274_ addr_r[0] baseaddr_r_sync[0] _1274_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0590__C _0590_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1261__CLK _1166_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0989_ _0988_/Y _0989_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0599__A _0573_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_132 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_64 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_110 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0796__A2 _0794_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_50 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1117__B _1136_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_154 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0675__C _0606_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0972__A _0986_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1284__CLK _1253_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0691__B _0698_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0912_ _0911_/Y _0986_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0843_ _0870_/A _0843_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0774_ _0793_/A _0870_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1027__B _1037_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_102 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0866__B _0871_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1043__A _1043_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1257_ d_fabric_in[29] _1257_/Q _1177_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1188_ d_sram_out[11] _0621_/C _1184_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_219 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_8 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0950__A2 _0944_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_154 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1157__CLK _1173_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_41 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_52 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0776__B _1147_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_146 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_60 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0769__A2 _0533_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_97 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1128__A _1118_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0967__A _0919_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_102 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0686__B _0521_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1111_ _1106_/X _1074_/Y _1110_/X _1111_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_65_179 VGND VPWR sky130_fd_sc_hd__fill_2
X_1042_ _1037_/Y _1043_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_0_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_115 VGND VPWR sky130_fd_sc_hd__decap_3
X_0826_ _0826_/A _0826_/B _0826_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_0757_ _0764_/A _1187_/Q _0757_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA_clkbuf_4_6_0_clk_A clkbuf_4_6_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1038__A _1082_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0688_ _0684_/Y _0686_/Y _0570_/A _0570_/B _0859_/C _0689_/A VGND VPWR sky130_fd_sc_hd__a2111oi_4
XANTENNA__0877__A _0877_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0932__A2 _0925_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_15_0_clk clkbuf_3_7_0_clk/X _1201_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_56_135 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_157 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0999__A2 _0984_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_63 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_85 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_89 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_40 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_124 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_93 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1100__A2 _1097_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_182 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_92 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_118 VGND VPWR sky130_fd_sc_hd__decap_4
X_0611_ _0611_/A _0612_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_50_91 VGND VPWR sky130_fd_sc_hd__decap_8
X_0542_ _0542_/A _0543_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_124_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0697__A _0807_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_3 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0678__A1 _0683_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_179 VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_clk clkbuf_3_5_0_clk/A clkbuf_3_4_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1025_ _1022_/Y _1024_/X _1025_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_61_182 VGND VPWR sky130_fd_sc_hd__fill_2
X_0809_ _1182_/Q _0749_/X _0742_/A _0809_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_30_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_37 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0669__A1 _0667_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_20 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_53 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_160 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1094__A1 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1109__C _1060_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_21 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_154 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_98 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0964__B _0962_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_108 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_91 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0980__B1_N _0979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_182 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0832__A1 _0794_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_1_1_0_clk_A clkbuf_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_30 VGND VPWR sky130_fd_sc_hd__decap_12
X_0525_ _0590_/C _0729_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_165 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1218__CLK _1218_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_127 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1051__A _1051_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_28 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VPWR sky130_fd_sc_hd__decap_3
X_1008_ _1256_/Q _0960_/X _0979_/X d_sram_in[28] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0823__A1 _0821_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1201__D d_sram_out[24] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_27 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_3_0_clk_A clkbuf_2_1_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_42 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_97 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_152 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0814__A1 _0807_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_14_0_clk_A clkbuf_3_7_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0578__B1 _0576_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_93 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1136__A _1136_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1290_ conf[2] _0919_/B _1274_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0975__A _0938_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0694__B _0568_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_130 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1046__A _1075_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0588__C _0588_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0741__B1 _0566_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1190__CLK _1208_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0885__A _0747_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_37 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_152 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_89 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0795__A _0826_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_84 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_101 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0799__B1 _0675_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0790_ _0784_/Y _0533_/X _0785_/X _0788_/Y _0789_/Y _0790_/X VGND VPWR sky130_fd_sc_hd__o41a_4
XFILLER_42_92 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0971__B1 _1238_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_144 VGND VPWR sky130_fd_sc_hd__fill_2
X_1273_ addr_w[13] _1037_/A _1274_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0590__D _0588_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0988_ _0921_/X _0936_/A _0988_/C _0988_/D _0988_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__0599__B _0543_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_111 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_155 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_15 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_58 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_25 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_73 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_62 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_44 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_99 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_0_0_clk_A clkbuf_1_0_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1117__C _1136_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_133 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_114 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_169 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1130__B1 _1129_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0972__B _0971_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0691__C _0521_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0911_ _0911_/A _0911_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0842_ _0779_/Y _0760_/X _0841_/Y _1156_/D VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0773_ out_reg _0793_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_52_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_170 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1027__C _1022_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_136 VGND VPWR sky130_fd_sc_hd__fill_2
X_1256_ d_fabric_in[28] _1256_/Q _1256_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1187_ d_sram_out[10] _1187_/Q _1180_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA_clkbuf_4_2_0_clk_A clkbuf_4_2_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_209 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_118 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_166 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1112__B1 _1111_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_52 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_34 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_56 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_21 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_76 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_171 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1128__B _1126_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0686__C _0883_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1144__A csb VGND VPWR sky130_fd_sc_hd__diode_2
X_1110_ _1118_/A _1108_/Y _1118_/B _1110_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_65_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1251__CLK _1288_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1103__B1 _1099_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1041_ _1037_/Y _1051_/A _1025_/Y _1036_/C w_mask[1] VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__0968__A1_N _0994_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_85 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_138 VGND VPWR sky130_fd_sc_hd__fill_2
X_0825_ _0786_/Y _0750_/X _0823_/X _0824_/Y _0825_/Y VGND VPWR sky130_fd_sc_hd__a22oi_4
XFILLER_127_160 VGND VPWR sky130_fd_sc_hd__fill_1
X_0756_ _1195_/Q _0868_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_127_182 VGND VPWR sky130_fd_sc_hd__decap_8
X_0687_ _0698_/A _0859_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0877__B _0895_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1054__A _1109_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_114 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0893__A _0893_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1204__D d_sram_out[27] VGND VPWR sky130_fd_sc_hd__diode_2
X_1239_ d_fabric_in[11] _1239_/Q _1252_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_71_139 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_33 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_37 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_108 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_75 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1274__CLK _1274_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_23 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0610_ _0587_/A _0547_/A _0611_/A VGND VPWR sky130_fd_sc_hd__nor2_4
X_0541_ _0536_/X _0539_/X _0883_/A _0528_/X _0541_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__0978__A _1104_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0678__A2 _0666_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1024_ _1106_/A _1024_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1147__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1049__A _1088_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0808_ _0806_/X _0807_/Y _0742_/A _0808_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_0739_ _0531_/Y _1190_/Q _0533_/A _0736_/Y _0738_/Y _0739_/X VGND VPWR sky130_fd_sc_hd__a2111o_4
XFILLER_130_100 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_111 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_103 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0669__A2 _0668_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_59 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_128 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_106 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_43 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_65 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1094__A2 _1090_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_36 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_11 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_62 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_33 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_144 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_10_0_clk_A clkbuf_3_5_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_117 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0964__C _0963_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_161 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0832__A2 _1153_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_14_0_clk clkbuf_3_7_0_clk/X _1208_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_42 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_86 VGND VPWR sky130_fd_sc_hd__decap_8
X_0524_ _0588_/C _0590_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_111 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VPWR sky130_fd_sc_hd__decap_3
X_1007_ _1255_/Q _0915_/X _0975_/Y d_sram_in[27] VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0823__A2 _0822_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_21 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_53 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_42 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_109 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_150 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_84 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0814__A2 _0762_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_164 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0578__B2 _0577_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0578__A1 _0574_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_3_0_clk clkbuf_2_1_0_clk/X clkbuf_4_6_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__1136__B _1136_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0975__B _0974_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0588__D _0588_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_175 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0741__A1 _0728_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0885__B _0889_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1062__A _1030_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1212__D _1212_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_131 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_131 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0980__A1 _1240_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_97 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_186 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0795__B _0795_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_78 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0799__A1 _0822_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_146 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1208__CLK _1208_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_168 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0971__B2 _0967_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0947__B1_N _0964_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0986__A _0986_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1272_ addr_w[12] _1102_/C _1180_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_95_189 VGND VPWR sky130_fd_sc_hd__fill_1
X_0987_ _1242_/Q _0984_/X _0986_/Y d_sram_in[14] VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1057__A _1057_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1207__D d_sram_out[30] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_37 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0650__B1 _0602_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1117__D _1136_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_71 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1130__A1 _1074_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0972__C _0986_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0691__D _0570_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0910_ _0922_/B _0910_/B _0909_/Y _0911_/A VGND VPWR sky130_fd_sc_hd__nor3_4
X_0841_ _0859_/A _0859_/B _0859_/C _1172_/D _0841_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_0772_ _0868_/A _0693_/Y _0761_/Y _0771_/X _0772_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1180__CLK _1180_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_123 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_148 VGND VPWR sky130_fd_sc_hd__decap_3
X_1255_ d_fabric_in[27] _1255_/Q _1288_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1186_ d_sram_out[9] _1186_/Q _1184_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_91_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0880__B1 _0879_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_15 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_87 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1112__A1 _1022_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_24 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_75 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_73 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_55 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1128__C _1137_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_70 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1144__B web VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_115 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1103__A1 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1040_ _1039_/X _1051_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_80_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0862__B1 _0861_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0824_ _1184_/Q _0760_/X _0742_/X _0824_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_134_109 VGND VPWR sky130_fd_sc_hd__decap_12
X_0755_ _0704_/X _0752_/Y _0754_/Y d_fabric_out[1] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0686_ _0807_/A _0521_/X _0883_/A _0686_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__0893__B _0893_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1238_ d_fabric_in[10] _1238_/Q _1256_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_44_28 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1070__A _1043_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1169_ _1169_/D _1169_/Q _1172_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0853__B1 _0852_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1220__D _1220_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_49 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_47 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1030__B1 _1029_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_104 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_79 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_184 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0540_ _1169_/D _0883_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0978__B _1026_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_126 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0994__A _0994_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_1023_ _1023_/A _1106_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_61_162 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_109 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_19 VGND VPWR sky130_fd_sc_hd__decap_12
X_0807_ _0807_/A _0807_/B _1174_/D _0807_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XANTENNA__1049__B _1059_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0738_ _0737_/Y _0738_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0669_ _0667_/Y _0668_/Y _0617_/C _0669_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_130_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1065__A _1057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0771__C1 _0770_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1215__D _1215_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_151 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_3 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1241__CLK _1256_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_52 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1003__B1 _0958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_153 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_96 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_93 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_7 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0989__A _0988_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_54 VGND VPWR sky130_fd_sc_hd__decap_6
X_0523_ _0546_/A _0588_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_134 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_107 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_170 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0808__B1 _0742_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1006_ _1254_/Q _1000_/X _0972_/Y d_sram_in[26] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_34_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1264__CLK _1166_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0766__A2_N _0671_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0899__A _0899_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_112 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_66 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_69 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_121 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0578__A2 _1161_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0602__A _0602_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1136__C _1136_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_70 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1287__CLK _1253_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_143 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_190 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0741__A2 _0740_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1062__B _1061_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_54 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0980__A2 _0960_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_36 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_165 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_13_0_clk clkbuf_3_6_0_clk/X _1180_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_93_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_95 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_125 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0799__A2 _0672_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_22 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0986__B _0985_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1271_ addr_w[11] _1019_/A _1166_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_95_179 VGND VPWR sky130_fd_sc_hd__fill_2
X_0986_ _0986_/A _0985_/Y _0986_/C _0930_/Y _0986_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__1073__A _1102_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_23 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1223__D _1286_/Q VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_2_0_clk clkbuf_2_1_0_clk/X clkbuf_3_2_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_10_102 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0650__A1 _0647_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_168 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_117 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_86 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_35 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_97 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_3 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1130__A2 _1121_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0972__D _0930_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_93 VGND VPWR sky130_fd_sc_hd__fill_2
X_0840_ _0794_/X _1155_/Q _0839_/X d_fabric_out[10] VGND VPWR sky130_fd_sc_hd__o21a_4
X_0771_ _1179_/Q _0566_/A _0745_/X _0770_/X _0771_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_38_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1254_ d_fabric_in[26] _1254_/Q _1288_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1185_ d_sram_out[8] _1185_/Q _1184_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0880__A1 _0870_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_19 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_0969_ _0950_/X _0968_/Y _0969_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XANTENNA__1218__D _0902_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_15 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_44 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_48 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1112__A2 _1105_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_85 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_184 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0610__A _0587_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1103__A2 _1102_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0862__A1 _0843_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_107 VGND VPWR sky130_fd_sc_hd__fill_2
X_0823_ _0821_/X _0822_/Y _0742_/X _0823_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_0754_ _0705_/X _0754_/B _0754_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_0685_ _0682_/X _0807_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0520__A _0588_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1237_ d_fabric_in[9] _1237_/Q _1252_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1168_ _0786_/A _1168_/Q _1172_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0853__A1 _0843_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1099_ _1030_/Y _1093_/B _1098_/X _1092_/Y _1099_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_100_24 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_79 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_7 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_15 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1030__A1 _1127_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_30 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1170__CLK _1172_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_182 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_174 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0605__A _0628_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_173 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_110 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0978__C _0936_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0780__B1 _0745_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_81 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0994__B _0994_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_138 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_108 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_160 VGND VPWR sky130_fd_sc_hd__fill_1
X_1022_ _1095_/A _1097_/B _1018_/X _1074_/C _1022_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
X_0806_ _0807_/A _0805_/Y _0708_/Y _0806_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1049__C _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0737_ _0544_/X _0606_/B _0729_/B _0737_/D _0737_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_115_143 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_154 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0981__A2_N _0966_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0668_ _0607_/B _0588_/B _0589_/A _0668_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_130_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1065__B _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0771__B1 _0745_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0599_ _0573_/B _0543_/A _0599_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__1193__CLK _1184_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_127 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_182 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1231__D d_fabric_in[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1003__A1 _1251_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_165 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_160 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_7 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_93 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_66 VGND VPWR sky130_fd_sc_hd__fill_1
X_0522_ _0521_/X _0807_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0777__B1_N _0776_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0808__A1 _0806_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1005_ _1253_/Q _1000_/X _0969_/Y d_sram_in[25] VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__1076__A _1126_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_124 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1226__D web VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_22 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_111 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_63 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0983__B1 _0982_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0602__B _0591_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1136__D _1136_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_82 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_166 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0974__B1 _1239_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_111 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0726__B1 _0566_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_155 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_105 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_116 VGND VPWR sky130_fd_sc_hd__decap_3
.ends

