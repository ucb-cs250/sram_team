VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sram_ifc
  CLASS BLOCK ;
  FOREIGN sram_ifc ;
  ORIGIN 0.000 0.000 ;
  SIZE 198.260 BY 208.980 ;
  PIN addr_r[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END addr_r[0]
  PIN addr_r[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 194.260 180.240 198.260 180.840 ;
    END
  END addr_r[10]
  PIN addr_r[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 194.260 47.640 198.260 48.240 ;
    END
  END addr_r[11]
  PIN addr_r[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.990 204.980 122.270 208.980 ;
    END
  END addr_r[12]
  PIN addr_r[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 194.260 142.840 198.260 143.440 ;
    END
  END addr_r[13]
  PIN addr_r[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END addr_r[1]
  PIN addr_r[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 204.980 115.370 208.980 ;
    END
  END addr_r[2]
  PIN addr_r[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END addr_r[3]
  PIN addr_r[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END addr_r[4]
  PIN addr_r[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.190 204.980 39.470 208.980 ;
    END
  END addr_r[5]
  PIN addr_r[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END addr_r[6]
  PIN addr_r[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END addr_r[7]
  PIN addr_r[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END addr_r[8]
  PIN addr_r[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.790 204.980 21.070 208.980 ;
    END
  END addr_r[9]
  PIN addr_w[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END addr_w[0]
  PIN addr_w[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END addr_w[10]
  PIN addr_w[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END addr_w[11]
  PIN addr_w[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END addr_w[12]
  PIN addr_w[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END addr_w[13]
  PIN addr_w[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END addr_w[1]
  PIN addr_w[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 194.260 23.840 198.260 24.440 ;
    END
  END addr_w[2]
  PIN addr_w[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END addr_w[3]
  PIN addr_w[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END addr_w[4]
  PIN addr_w[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.390 204.980 48.670 208.980 ;
    END
  END addr_w[5]
  PIN addr_w[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END addr_w[6]
  PIN addr_w[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END addr_w[7]
  PIN addr_w[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 204.980 4.970 208.980 ;
    END
  END addr_w[8]
  PIN addr_w[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END addr_w[9]
  PIN baseaddr_r_sync[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 85.040 198.260 85.640 ;
    END
  END baseaddr_r_sync[0]
  PIN baseaddr_r_sync[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 138.090 204.980 138.370 208.980 ;
    END
  END baseaddr_r_sync[1]
  PIN baseaddr_r_sync[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END baseaddr_r_sync[2]
  PIN baseaddr_r_sync[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END baseaddr_r_sync[3]
  PIN baseaddr_r_sync[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 10.240 198.260 10.840 ;
    END
  END baseaddr_r_sync[4]
  PIN baseaddr_r_sync[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END baseaddr_r_sync[5]
  PIN baseaddr_r_sync[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END baseaddr_r_sync[6]
  PIN baseaddr_r_sync[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.690 204.980 27.970 208.980 ;
    END
  END baseaddr_r_sync[7]
  PIN baseaddr_r_sync[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 142.690 204.980 142.970 208.980 ;
    END
  END baseaddr_r_sync[8]
  PIN baseaddr_w_sync[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.090 204.980 69.370 208.980 ;
    END
  END baseaddr_w_sync[0]
  PIN baseaddr_w_sync[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 183.640 198.260 184.240 ;
    END
  END baseaddr_w_sync[1]
  PIN baseaddr_w_sync[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END baseaddr_w_sync[2]
  PIN baseaddr_w_sync[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 52.990 204.980 53.270 208.980 ;
    END
  END baseaddr_w_sync[3]
  PIN baseaddr_w_sync[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.590 204.980 80.870 208.980 ;
    END
  END baseaddr_w_sync[4]
  PIN baseaddr_w_sync[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 172.590 204.980 172.870 208.980 ;
    END
  END baseaddr_w_sync[5]
  PIN baseaddr_w_sync[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END baseaddr_w_sync[6]
  PIN baseaddr_w_sync[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END baseaddr_w_sync[7]
  PIN baseaddr_w_sync[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END baseaddr_w_sync[8]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END clk
  PIN conf[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.490 204.980 133.770 208.980 ;
    END
  END conf[0]
  PIN conf[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END conf[1]
  PIN conf[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 194.260 71.440 198.260 72.040 ;
    END
  END conf[2]
  PIN csb
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END csb
  PIN csb0_sync
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 188.690 204.980 188.970 208.980 ;
    END
  END csb0_sync
  PIN csb1_sync
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.490 204.980 18.770 208.980 ;
    END
  END csb1_sync
  PIN d_fabric_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END d_fabric_in[0]
  PIN d_fabric_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END d_fabric_in[10]
  PIN d_fabric_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.390 204.980 117.670 208.980 ;
    END
  END d_fabric_in[11]
  PIN d_fabric_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 194.260 200.640 198.260 201.240 ;
    END
  END d_fabric_in[12]
  PIN d_fabric_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END d_fabric_in[13]
  PIN d_fabric_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END d_fabric_in[14]
  PIN d_fabric_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.290 204.980 32.570 208.980 ;
    END
  END d_fabric_in[15]
  PIN d_fabric_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 147.290 204.980 147.570 208.980 ;
    END
  END d_fabric_in[16]
  PIN d_fabric_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 194.260 197.240 198.260 197.840 ;
    END
  END d_fabric_in[17]
  PIN d_fabric_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 194.260 156.440 198.260 157.040 ;
    END
  END d_fabric_in[18]
  PIN d_fabric_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.990 204.980 191.270 208.980 ;
    END
  END d_fabric_in[19]
  PIN d_fabric_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END d_fabric_in[1]
  PIN d_fabric_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END d_fabric_in[20]
  PIN d_fabric_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 194.260 146.240 198.260 146.840 ;
    END
  END d_fabric_in[21]
  PIN d_fabric_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END d_fabric_in[22]
  PIN d_fabric_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 194.260 112.240 198.260 112.840 ;
    END
  END d_fabric_in[23]
  PIN d_fabric_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END d_fabric_in[24]
  PIN d_fabric_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 158.790 204.980 159.070 208.980 ;
    END
  END d_fabric_in[25]
  PIN d_fabric_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.290 204.980 55.570 208.980 ;
    END
  END d_fabric_in[26]
  PIN d_fabric_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 204.980 14.170 208.980 ;
    END
  END d_fabric_in[27]
  PIN d_fabric_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 194.260 98.640 198.260 99.240 ;
    END
  END d_fabric_in[28]
  PIN d_fabric_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 194.260 125.840 198.260 126.440 ;
    END
  END d_fabric_in[29]
  PIN d_fabric_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END d_fabric_in[2]
  PIN d_fabric_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END d_fabric_in[30]
  PIN d_fabric_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END d_fabric_in[31]
  PIN d_fabric_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END d_fabric_in[3]
  PIN d_fabric_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 149.590 204.980 149.870 208.980 ;
    END
  END d_fabric_in[4]
  PIN d_fabric_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 131.190 204.980 131.470 208.980 ;
    END
  END d_fabric_in[5]
  PIN d_fabric_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END d_fabric_in[6]
  PIN d_fabric_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 194.260 207.440 198.260 208.040 ;
    END
  END d_fabric_in[7]
  PIN d_fabric_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END d_fabric_in[8]
  PIN d_fabric_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END d_fabric_in[9]
  PIN d_fabric_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END d_fabric_out[0]
  PIN d_fabric_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END d_fabric_out[10]
  PIN d_fabric_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END d_fabric_out[11]
  PIN d_fabric_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 170.040 198.260 170.640 ;
    END
  END d_fabric_out[12]
  PIN d_fabric_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END d_fabric_out[13]
  PIN d_fabric_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END d_fabric_out[14]
  PIN d_fabric_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.890 204.980 83.170 208.980 ;
    END
  END d_fabric_out[15]
  PIN d_fabric_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 122.440 198.260 123.040 ;
    END
  END d_fabric_out[16]
  PIN d_fabric_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 128.890 204.980 129.170 208.980 ;
    END
  END d_fabric_out[17]
  PIN d_fabric_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END d_fabric_out[18]
  PIN d_fabric_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 17.040 198.260 17.640 ;
    END
  END d_fabric_out[19]
  PIN d_fabric_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END d_fabric_out[1]
  PIN d_fabric_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END d_fabric_out[20]
  PIN d_fabric_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END d_fabric_out[21]
  PIN d_fabric_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END d_fabric_out[22]
  PIN d_fabric_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END d_fabric_out[23]
  PIN d_fabric_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 74.840 198.260 75.440 ;
    END
  END d_fabric_out[24]
  PIN d_fabric_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END d_fabric_out[25]
  PIN d_fabric_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END d_fabric_out[26]
  PIN d_fabric_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END d_fabric_out[27]
  PIN d_fabric_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.490 204.980 87.770 208.980 ;
    END
  END d_fabric_out[28]
  PIN d_fabric_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END d_fabric_out[29]
  PIN d_fabric_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.390 204.980 71.670 208.980 ;
    END
  END d_fabric_out[2]
  PIN d_fabric_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.990 204.980 99.270 208.980 ;
    END
  END d_fabric_out[30]
  PIN d_fabric_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 197.890 204.980 198.170 208.980 ;
    END
  END d_fabric_out[31]
  PIN d_fabric_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.390 204.980 163.670 208.980 ;
    END
  END d_fabric_out[3]
  PIN d_fabric_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END d_fabric_out[4]
  PIN d_fabric_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 163.240 198.260 163.840 ;
    END
  END d_fabric_out[5]
  PIN d_fabric_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 149.640 198.260 150.240 ;
    END
  END d_fabric_out[6]
  PIN d_fabric_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 105.440 198.260 106.040 ;
    END
  END d_fabric_out[7]
  PIN d_fabric_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END d_fabric_out[8]
  PIN d_fabric_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END d_fabric_out[9]
  PIN d_sram_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END d_sram_in[0]
  PIN d_sram_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 61.240 198.260 61.840 ;
    END
  END d_sram_in[10]
  PIN d_sram_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 57.840 198.260 58.440 ;
    END
  END d_sram_in[11]
  PIN d_sram_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.590 204.980 103.870 208.980 ;
    END
  END d_sram_in[12]
  PIN d_sram_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.990 204.980 7.270 208.980 ;
    END
  END d_sram_in[13]
  PIN d_sram_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END d_sram_in[14]
  PIN d_sram_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END d_sram_in[15]
  PIN d_sram_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 37.440 198.260 38.040 ;
    END
  END d_sram_in[16]
  PIN d_sram_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 0.040 198.260 0.640 ;
    END
  END d_sram_in[17]
  PIN d_sram_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END d_sram_in[18]
  PIN d_sram_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 187.040 198.260 187.640 ;
    END
  END d_sram_in[19]
  PIN d_sram_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 204.980 73.970 208.980 ;
    END
  END d_sram_in[1]
  PIN d_sram_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.790 204.980 44.070 208.980 ;
    END
  END d_sram_in[20]
  PIN d_sram_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 136.040 198.260 136.640 ;
    END
  END d_sram_in[21]
  PIN d_sram_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END d_sram_in[22]
  PIN d_sram_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END d_sram_in[23]
  PIN d_sram_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END d_sram_in[24]
  PIN d_sram_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 181.790 204.980 182.070 208.980 ;
    END
  END d_sram_in[25]
  PIN d_sram_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END d_sram_in[26]
  PIN d_sram_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.490 204.980 64.770 208.980 ;
    END
  END d_sram_in[27]
  PIN d_sram_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END d_sram_in[28]
  PIN d_sram_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END d_sram_in[29]
  PIN d_sram_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END d_sram_in[2]
  PIN d_sram_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.890 204.980 106.170 208.980 ;
    END
  END d_sram_in[30]
  PIN d_sram_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 30.640 198.260 31.240 ;
    END
  END d_sram_in[31]
  PIN d_sram_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.390 204.980 2.670 208.980 ;
    END
  END d_sram_in[3]
  PIN d_sram_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 204.980 90.070 208.980 ;
    END
  END d_sram_in[4]
  PIN d_sram_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 51.040 198.260 51.640 ;
    END
  END d_sram_in[5]
  PIN d_sram_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.890 204.980 37.170 208.980 ;
    END
  END d_sram_in[6]
  PIN d_sram_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END d_sram_in[7]
  PIN d_sram_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END d_sram_in[8]
  PIN d_sram_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 68.040 198.260 68.640 ;
    END
  END d_sram_in[9]
  PIN d_sram_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END d_sram_out[0]
  PIN d_sram_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END d_sram_out[10]
  PIN d_sram_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END d_sram_out[11]
  PIN d_sram_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.990 204.980 30.270 208.980 ;
    END
  END d_sram_out[12]
  PIN d_sram_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.790 204.980 113.070 208.980 ;
    END
  END d_sram_out[13]
  PIN d_sram_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END d_sram_out[14]
  PIN d_sram_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 174.890 204.980 175.170 208.980 ;
    END
  END d_sram_out[15]
  PIN d_sram_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END d_sram_out[16]
  PIN d_sram_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 194.260 193.840 198.260 194.440 ;
    END
  END d_sram_out[17]
  PIN d_sram_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END d_sram_out[18]
  PIN d_sram_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 165.690 204.980 165.970 208.980 ;
    END
  END d_sram_out[19]
  PIN d_sram_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 194.260 132.640 198.260 133.240 ;
    END
  END d_sram_out[1]
  PIN d_sram_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END d_sram_out[20]
  PIN d_sram_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END d_sram_out[21]
  PIN d_sram_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END d_sram_out[22]
  PIN d_sram_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 167.990 204.980 168.270 208.980 ;
    END
  END d_sram_out[23]
  PIN d_sram_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END d_sram_out[24]
  PIN d_sram_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END d_sram_out[25]
  PIN d_sram_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 179.490 204.980 179.770 208.980 ;
    END
  END d_sram_out[26]
  PIN d_sram_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END d_sram_out[27]
  PIN d_sram_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END d_sram_out[28]
  PIN d_sram_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END d_sram_out[29]
  PIN d_sram_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 194.260 173.440 198.260 174.040 ;
    END
  END d_sram_out[2]
  PIN d_sram_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END d_sram_out[30]
  PIN d_sram_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END d_sram_out[31]
  PIN d_sram_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 194.260 44.240 198.260 44.840 ;
    END
  END d_sram_out[3]
  PIN d_sram_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END d_sram_out[4]
  PIN d_sram_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END d_sram_out[5]
  PIN d_sram_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 194.260 108.840 198.260 109.440 ;
    END
  END d_sram_out[6]
  PIN d_sram_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 204.980 23.370 208.980 ;
    END
  END d_sram_out[7]
  PIN d_sram_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END d_sram_out[8]
  PIN d_sram_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END d_sram_out[9]
  PIN out_reg
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 154.190 204.980 154.470 208.980 ;
    END
  END out_reg
  PIN reb
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END reb
  PIN w_mask[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END w_mask[0]
  PIN w_mask[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 96.690 204.980 96.970 208.980 ;
    END
  END w_mask[10]
  PIN w_mask[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 159.840 198.260 160.440 ;
    END
  END w_mask[11]
  PIN w_mask[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END w_mask[12]
  PIN w_mask[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END w_mask[13]
  PIN w_mask[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END w_mask[14]
  PIN w_mask[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END w_mask[15]
  PIN w_mask[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 156.490 204.980 156.770 208.980 ;
    END
  END w_mask[16]
  PIN w_mask[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 193.290 204.980 193.570 208.980 ;
    END
  END w_mask[17]
  PIN w_mask[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 119.040 198.260 119.640 ;
    END
  END w_mask[18]
  PIN w_mask[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END w_mask[19]
  PIN w_mask[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END w_mask[1]
  PIN w_mask[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 62.190 204.980 62.470 208.980 ;
    END
  END w_mask[20]
  PIN w_mask[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 11.590 204.980 11.870 208.980 ;
    END
  END w_mask[21]
  PIN w_mask[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 140.390 204.980 140.670 208.980 ;
    END
  END w_mask[22]
  PIN w_mask[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END w_mask[23]
  PIN w_mask[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END w_mask[24]
  PIN w_mask[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END w_mask[25]
  PIN w_mask[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.290 204.980 124.570 208.980 ;
    END
  END w_mask[26]
  PIN w_mask[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 57.590 204.980 57.870 208.980 ;
    END
  END w_mask[27]
  PIN w_mask[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.190 204.980 108.470 208.980 ;
    END
  END w_mask[28]
  PIN w_mask[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 184.090 204.980 184.370 208.980 ;
    END
  END w_mask[29]
  PIN w_mask[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.290 204.980 78.570 208.980 ;
    END
  END w_mask[2]
  PIN w_mask[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END w_mask[30]
  PIN w_mask[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END w_mask[31]
  PIN w_mask[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 95.240 198.260 95.840 ;
    END
  END w_mask[3]
  PIN w_mask[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 81.640 198.260 82.240 ;
    END
  END w_mask[4]
  PIN w_mask[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.090 204.980 92.370 208.980 ;
    END
  END w_mask[5]
  PIN w_mask[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 34.040 198.260 34.640 ;
    END
  END w_mask[6]
  PIN w_mask[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 6.840 198.260 7.440 ;
    END
  END w_mask[7]
  PIN w_mask[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 88.440 198.260 89.040 ;
    END
  END w_mask[8]
  PIN w_mask[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 194.260 20.440 198.260 21.040 ;
    END
  END w_mask[9]
  PIN web
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.090 204.980 46.370 208.980 ;
    END
  END web
  PIN web0_sync
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END web0_sync
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 192.740 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 192.740 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 192.740 195.925 ;
      LAYER met1 ;
        RECT 0.070 5.820 193.590 201.240 ;
      LAYER met2 ;
        RECT 0.090 204.700 2.110 207.925 ;
        RECT 2.950 204.700 4.410 207.925 ;
        RECT 5.250 204.700 6.710 207.925 ;
        RECT 7.550 204.700 11.310 207.925 ;
        RECT 12.150 204.700 13.610 207.925 ;
        RECT 14.450 204.700 18.210 207.925 ;
        RECT 19.050 204.700 20.510 207.925 ;
        RECT 21.350 204.700 22.810 207.925 ;
        RECT 23.650 204.700 27.410 207.925 ;
        RECT 28.250 204.700 29.710 207.925 ;
        RECT 30.550 204.700 32.010 207.925 ;
        RECT 32.850 204.700 36.610 207.925 ;
        RECT 37.450 204.700 38.910 207.925 ;
        RECT 39.750 204.700 43.510 207.925 ;
        RECT 44.350 204.700 45.810 207.925 ;
        RECT 46.650 204.700 48.110 207.925 ;
        RECT 48.950 204.700 52.710 207.925 ;
        RECT 53.550 204.700 55.010 207.925 ;
        RECT 55.850 204.700 57.310 207.925 ;
        RECT 58.150 204.700 61.910 207.925 ;
        RECT 62.750 204.700 64.210 207.925 ;
        RECT 65.050 204.700 68.810 207.925 ;
        RECT 69.650 204.700 71.110 207.925 ;
        RECT 71.950 204.700 73.410 207.925 ;
        RECT 74.250 204.700 78.010 207.925 ;
        RECT 78.850 204.700 80.310 207.925 ;
        RECT 81.150 204.700 82.610 207.925 ;
        RECT 83.450 204.700 87.210 207.925 ;
        RECT 88.050 204.700 89.510 207.925 ;
        RECT 90.350 204.700 91.810 207.925 ;
        RECT 92.650 204.700 96.410 207.925 ;
        RECT 97.250 204.700 98.710 207.925 ;
        RECT 99.550 204.700 103.310 207.925 ;
        RECT 104.150 204.700 105.610 207.925 ;
        RECT 106.450 204.700 107.910 207.925 ;
        RECT 108.750 204.700 112.510 207.925 ;
        RECT 113.350 204.700 114.810 207.925 ;
        RECT 115.650 204.700 117.110 207.925 ;
        RECT 117.950 204.700 121.710 207.925 ;
        RECT 122.550 204.700 124.010 207.925 ;
        RECT 124.850 204.700 128.610 207.925 ;
        RECT 129.450 204.700 130.910 207.925 ;
        RECT 131.750 204.700 133.210 207.925 ;
        RECT 134.050 204.700 137.810 207.925 ;
        RECT 138.650 204.700 140.110 207.925 ;
        RECT 140.950 204.700 142.410 207.925 ;
        RECT 143.250 204.700 147.010 207.925 ;
        RECT 147.850 204.700 149.310 207.925 ;
        RECT 150.150 204.700 153.910 207.925 ;
        RECT 154.750 204.700 156.210 207.925 ;
        RECT 157.050 204.700 158.510 207.925 ;
        RECT 159.350 204.700 163.110 207.925 ;
        RECT 163.950 204.700 165.410 207.925 ;
        RECT 166.250 204.700 167.710 207.925 ;
        RECT 168.550 204.700 172.310 207.925 ;
        RECT 173.150 204.700 174.610 207.925 ;
        RECT 175.450 204.700 179.210 207.925 ;
        RECT 180.050 204.700 181.510 207.925 ;
        RECT 182.350 204.700 183.810 207.925 ;
        RECT 184.650 204.700 188.410 207.925 ;
        RECT 189.250 204.700 190.710 207.925 ;
        RECT 191.550 204.700 193.010 207.925 ;
        RECT 193.850 204.700 197.610 207.925 ;
        RECT 0.090 4.280 198.170 204.700 ;
        RECT 0.650 0.155 2.110 4.280 ;
        RECT 2.950 0.155 4.410 4.280 ;
        RECT 5.250 0.155 9.010 4.280 ;
        RECT 9.850 0.155 11.310 4.280 ;
        RECT 12.150 0.155 13.610 4.280 ;
        RECT 14.450 0.155 18.210 4.280 ;
        RECT 19.050 0.155 20.510 4.280 ;
        RECT 21.350 0.155 22.810 4.280 ;
        RECT 23.650 0.155 27.410 4.280 ;
        RECT 28.250 0.155 29.710 4.280 ;
        RECT 30.550 0.155 34.310 4.280 ;
        RECT 35.150 0.155 36.610 4.280 ;
        RECT 37.450 0.155 38.910 4.280 ;
        RECT 39.750 0.155 43.510 4.280 ;
        RECT 44.350 0.155 45.810 4.280 ;
        RECT 46.650 0.155 48.110 4.280 ;
        RECT 48.950 0.155 52.710 4.280 ;
        RECT 53.550 0.155 55.010 4.280 ;
        RECT 55.850 0.155 59.610 4.280 ;
        RECT 60.450 0.155 61.910 4.280 ;
        RECT 62.750 0.155 64.210 4.280 ;
        RECT 65.050 0.155 68.810 4.280 ;
        RECT 69.650 0.155 71.110 4.280 ;
        RECT 71.950 0.155 73.410 4.280 ;
        RECT 74.250 0.155 78.010 4.280 ;
        RECT 78.850 0.155 80.310 4.280 ;
        RECT 81.150 0.155 84.910 4.280 ;
        RECT 85.750 0.155 87.210 4.280 ;
        RECT 88.050 0.155 89.510 4.280 ;
        RECT 90.350 0.155 94.110 4.280 ;
        RECT 94.950 0.155 96.410 4.280 ;
        RECT 97.250 0.155 98.710 4.280 ;
        RECT 99.550 0.155 103.310 4.280 ;
        RECT 104.150 0.155 105.610 4.280 ;
        RECT 106.450 0.155 110.210 4.280 ;
        RECT 111.050 0.155 112.510 4.280 ;
        RECT 113.350 0.155 114.810 4.280 ;
        RECT 115.650 0.155 119.410 4.280 ;
        RECT 120.250 0.155 121.710 4.280 ;
        RECT 122.550 0.155 124.010 4.280 ;
        RECT 124.850 0.155 128.610 4.280 ;
        RECT 129.450 0.155 130.910 4.280 ;
        RECT 131.750 0.155 135.510 4.280 ;
        RECT 136.350 0.155 137.810 4.280 ;
        RECT 138.650 0.155 140.110 4.280 ;
        RECT 140.950 0.155 144.710 4.280 ;
        RECT 145.550 0.155 147.010 4.280 ;
        RECT 147.850 0.155 149.310 4.280 ;
        RECT 150.150 0.155 153.910 4.280 ;
        RECT 154.750 0.155 156.210 4.280 ;
        RECT 157.050 0.155 160.810 4.280 ;
        RECT 161.650 0.155 163.110 4.280 ;
        RECT 163.950 0.155 165.410 4.280 ;
        RECT 166.250 0.155 170.010 4.280 ;
        RECT 170.850 0.155 172.310 4.280 ;
        RECT 173.150 0.155 174.610 4.280 ;
        RECT 175.450 0.155 179.210 4.280 ;
        RECT 180.050 0.155 181.510 4.280 ;
        RECT 182.350 0.155 186.110 4.280 ;
        RECT 186.950 0.155 188.410 4.280 ;
        RECT 189.250 0.155 190.710 4.280 ;
        RECT 191.550 0.155 195.310 4.280 ;
        RECT 196.150 0.155 197.610 4.280 ;
      LAYER met3 ;
        RECT 4.400 207.040 193.860 207.905 ;
        RECT 0.065 205.040 198.195 207.040 ;
        RECT 4.400 203.640 198.195 205.040 ;
        RECT 0.065 201.640 198.195 203.640 ;
        RECT 4.400 200.240 193.860 201.640 ;
        RECT 0.065 198.240 198.195 200.240 ;
        RECT 0.065 196.840 193.860 198.240 ;
        RECT 0.065 194.840 198.195 196.840 ;
        RECT 4.400 193.440 193.860 194.840 ;
        RECT 0.065 191.440 198.195 193.440 ;
        RECT 4.400 190.040 198.195 191.440 ;
        RECT 0.065 188.040 198.195 190.040 ;
        RECT 0.065 186.640 193.860 188.040 ;
        RECT 0.065 184.640 198.195 186.640 ;
        RECT 4.400 183.240 193.860 184.640 ;
        RECT 0.065 181.240 198.195 183.240 ;
        RECT 4.400 179.840 193.860 181.240 ;
        RECT 0.065 177.840 198.195 179.840 ;
        RECT 4.400 176.440 198.195 177.840 ;
        RECT 0.065 174.440 198.195 176.440 ;
        RECT 0.065 173.040 193.860 174.440 ;
        RECT 0.065 171.040 198.195 173.040 ;
        RECT 4.400 169.640 193.860 171.040 ;
        RECT 0.065 167.640 198.195 169.640 ;
        RECT 4.400 166.240 198.195 167.640 ;
        RECT 0.065 164.240 198.195 166.240 ;
        RECT 4.400 162.840 193.860 164.240 ;
        RECT 0.065 160.840 198.195 162.840 ;
        RECT 0.065 159.440 193.860 160.840 ;
        RECT 0.065 157.440 198.195 159.440 ;
        RECT 4.400 156.040 193.860 157.440 ;
        RECT 0.065 154.040 198.195 156.040 ;
        RECT 4.400 152.640 198.195 154.040 ;
        RECT 0.065 150.640 198.195 152.640 ;
        RECT 0.065 149.240 193.860 150.640 ;
        RECT 0.065 147.240 198.195 149.240 ;
        RECT 4.400 145.840 193.860 147.240 ;
        RECT 0.065 143.840 198.195 145.840 ;
        RECT 4.400 142.440 193.860 143.840 ;
        RECT 0.065 140.440 198.195 142.440 ;
        RECT 4.400 139.040 198.195 140.440 ;
        RECT 0.065 137.040 198.195 139.040 ;
        RECT 0.065 135.640 193.860 137.040 ;
        RECT 0.065 133.640 198.195 135.640 ;
        RECT 4.400 132.240 193.860 133.640 ;
        RECT 0.065 130.240 198.195 132.240 ;
        RECT 4.400 128.840 198.195 130.240 ;
        RECT 0.065 126.840 198.195 128.840 ;
        RECT 4.400 125.440 193.860 126.840 ;
        RECT 0.065 123.440 198.195 125.440 ;
        RECT 0.065 122.040 193.860 123.440 ;
        RECT 0.065 120.040 198.195 122.040 ;
        RECT 4.400 118.640 193.860 120.040 ;
        RECT 0.065 116.640 198.195 118.640 ;
        RECT 4.400 115.240 198.195 116.640 ;
        RECT 0.065 113.240 198.195 115.240 ;
        RECT 0.065 111.840 193.860 113.240 ;
        RECT 0.065 109.840 198.195 111.840 ;
        RECT 4.400 108.440 193.860 109.840 ;
        RECT 0.065 106.440 198.195 108.440 ;
        RECT 4.400 105.040 193.860 106.440 ;
        RECT 0.065 103.040 198.195 105.040 ;
        RECT 4.400 101.640 198.195 103.040 ;
        RECT 0.065 99.640 198.195 101.640 ;
        RECT 0.065 98.240 193.860 99.640 ;
        RECT 0.065 96.240 198.195 98.240 ;
        RECT 4.400 94.840 193.860 96.240 ;
        RECT 0.065 92.840 198.195 94.840 ;
        RECT 4.400 91.440 198.195 92.840 ;
        RECT 0.065 89.440 198.195 91.440 ;
        RECT 4.400 88.040 193.860 89.440 ;
        RECT 0.065 86.040 198.195 88.040 ;
        RECT 0.065 84.640 193.860 86.040 ;
        RECT 0.065 82.640 198.195 84.640 ;
        RECT 4.400 81.240 193.860 82.640 ;
        RECT 0.065 79.240 198.195 81.240 ;
        RECT 4.400 77.840 198.195 79.240 ;
        RECT 0.065 75.840 198.195 77.840 ;
        RECT 0.065 74.440 193.860 75.840 ;
        RECT 0.065 72.440 198.195 74.440 ;
        RECT 4.400 71.040 193.860 72.440 ;
        RECT 0.065 69.040 198.195 71.040 ;
        RECT 4.400 67.640 193.860 69.040 ;
        RECT 0.065 65.640 198.195 67.640 ;
        RECT 4.400 64.240 198.195 65.640 ;
        RECT 0.065 62.240 198.195 64.240 ;
        RECT 0.065 60.840 193.860 62.240 ;
        RECT 0.065 58.840 198.195 60.840 ;
        RECT 4.400 57.440 193.860 58.840 ;
        RECT 0.065 55.440 198.195 57.440 ;
        RECT 4.400 54.040 198.195 55.440 ;
        RECT 0.065 52.040 198.195 54.040 ;
        RECT 4.400 50.640 193.860 52.040 ;
        RECT 0.065 48.640 198.195 50.640 ;
        RECT 0.065 47.240 193.860 48.640 ;
        RECT 0.065 45.240 198.195 47.240 ;
        RECT 4.400 43.840 193.860 45.240 ;
        RECT 0.065 41.840 198.195 43.840 ;
        RECT 4.400 40.440 198.195 41.840 ;
        RECT 0.065 38.440 198.195 40.440 ;
        RECT 0.065 37.040 193.860 38.440 ;
        RECT 0.065 35.040 198.195 37.040 ;
        RECT 4.400 33.640 193.860 35.040 ;
        RECT 0.065 31.640 198.195 33.640 ;
        RECT 4.400 30.240 193.860 31.640 ;
        RECT 0.065 28.240 198.195 30.240 ;
        RECT 4.400 26.840 198.195 28.240 ;
        RECT 0.065 24.840 198.195 26.840 ;
        RECT 0.065 23.440 193.860 24.840 ;
        RECT 0.065 21.440 198.195 23.440 ;
        RECT 4.400 20.040 193.860 21.440 ;
        RECT 0.065 18.040 198.195 20.040 ;
        RECT 4.400 16.640 193.860 18.040 ;
        RECT 0.065 14.640 198.195 16.640 ;
        RECT 4.400 13.240 198.195 14.640 ;
        RECT 0.065 11.240 198.195 13.240 ;
        RECT 0.065 9.840 193.860 11.240 ;
        RECT 0.065 7.840 198.195 9.840 ;
        RECT 4.400 6.440 193.860 7.840 ;
        RECT 0.065 4.440 198.195 6.440 ;
        RECT 4.400 3.040 198.195 4.440 ;
        RECT 0.065 1.040 198.195 3.040 ;
        RECT 0.065 0.175 193.860 1.040 ;
      LAYER met4 ;
        RECT 19.190 6.295 178.610 196.080 ;
      LAYER met5 ;
        RECT 5.520 106.280 192.740 181.270 ;
        RECT 5.520 72.300 192.740 101.480 ;
  END
END sram_ifc
END LIBRARY

